/* modified netlist. Source: module Keccak in file /mnt/c/Users/amirm/Desktop/Papers_in_progress/SAUBER/Design for our FPGA/8-Keccak-200_RoundBased_PortSerial/4-AGEMA/Keccak.v */
/* 0 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 1 register stage(s) in total */

module Keccak_SAUBER_Pipeline_d1 (InData_s0_t, Reset_t, Reset_f, InData_s0_f, InData_s1_t, InData_s1_f, OutData_s0_t, Ready_t, OutData_s0_f, OutData_s1_t, OutData_s1_f, Ready_f);
    input [7:0] InData_s0_t ;
    input Reset_t ;
    input Reset_f ;
    input [7:0] InData_s0_f ;
    input [7:0] InData_s1_t ;
    input [7:0] InData_s1_f ;
    output [7:0] OutData_s0_t ;
    output Ready_t ;
    output [7:0] OutData_s0_f ;
    output [7:0] OutData_s1_t ;
    output [7:0] OutData_s1_f ;
    output Ready_f ;
    wire IotaRC_7 ;
    wire IotaRC_3 ;
    wire n9 ;
    wire THETA_n200 ;
    wire THETA_n199 ;
    wire THETA_n198 ;
    wire THETA_n197 ;
    wire THETA_n196 ;
    wire THETA_n195 ;
    wire THETA_n194 ;
    wire THETA_n193 ;
    wire THETA_n192 ;
    wire THETA_n191 ;
    wire THETA_n190 ;
    wire THETA_n189 ;
    wire THETA_n188 ;
    wire THETA_n187 ;
    wire THETA_n186 ;
    wire THETA_n185 ;
    wire THETA_n184 ;
    wire THETA_n183 ;
    wire THETA_n182 ;
    wire THETA_n181 ;
    wire THETA_n180 ;
    wire THETA_n179 ;
    wire THETA_n178 ;
    wire THETA_n177 ;
    wire THETA_n176 ;
    wire THETA_n175 ;
    wire THETA_n174 ;
    wire THETA_n173 ;
    wire THETA_n172 ;
    wire THETA_n171 ;
    wire THETA_n170 ;
    wire THETA_n169 ;
    wire THETA_n168 ;
    wire THETA_n167 ;
    wire THETA_n166 ;
    wire THETA_n165 ;
    wire THETA_n164 ;
    wire THETA_n163 ;
    wire THETA_n162 ;
    wire THETA_n161 ;
    wire THETA_n160 ;
    wire THETA_n159 ;
    wire THETA_n158 ;
    wire THETA_n157 ;
    wire THETA_n156 ;
    wire THETA_n155 ;
    wire THETA_n154 ;
    wire THETA_n153 ;
    wire THETA_n152 ;
    wire THETA_n151 ;
    wire THETA_n150 ;
    wire THETA_n149 ;
    wire THETA_n148 ;
    wire THETA_n147 ;
    wire THETA_n146 ;
    wire THETA_n145 ;
    wire THETA_n144 ;
    wire THETA_n143 ;
    wire THETA_n142 ;
    wire THETA_n141 ;
    wire THETA_n140 ;
    wire THETA_n139 ;
    wire THETA_n138 ;
    wire THETA_n137 ;
    wire THETA_n136 ;
    wire THETA_n135 ;
    wire THETA_n134 ;
    wire THETA_n133 ;
    wire THETA_n132 ;
    wire THETA_n131 ;
    wire THETA_n130 ;
    wire THETA_n129 ;
    wire THETA_n128 ;
    wire THETA_n127 ;
    wire THETA_n126 ;
    wire THETA_n125 ;
    wire THETA_n124 ;
    wire THETA_n123 ;
    wire THETA_n122 ;
    wire THETA_n121 ;
    wire THETA_n120 ;
    wire THETA_n119 ;
    wire THETA_n118 ;
    wire THETA_n117 ;
    wire THETA_n116 ;
    wire THETA_n115 ;
    wire THETA_n114 ;
    wire THETA_n113 ;
    wire THETA_n112 ;
    wire THETA_n111 ;
    wire THETA_n110 ;
    wire THETA_n109 ;
    wire THETA_n108 ;
    wire THETA_n107 ;
    wire THETA_n106 ;
    wire THETA_n105 ;
    wire THETA_n104 ;
    wire THETA_n103 ;
    wire THETA_n102 ;
    wire THETA_n101 ;
    wire THETA_n100 ;
    wire THETA_n99 ;
    wire THETA_n98 ;
    wire THETA_n97 ;
    wire THETA_n96 ;
    wire THETA_n95 ;
    wire THETA_n94 ;
    wire THETA_n93 ;
    wire THETA_n92 ;
    wire THETA_n91 ;
    wire THETA_n90 ;
    wire THETA_n89 ;
    wire THETA_n88 ;
    wire THETA_n87 ;
    wire THETA_n86 ;
    wire THETA_n85 ;
    wire THETA_n84 ;
    wire THETA_n83 ;
    wire THETA_n82 ;
    wire THETA_n81 ;
    wire THETA_n80 ;
    wire THETA_n79 ;
    wire THETA_n78 ;
    wire THETA_n77 ;
    wire THETA_n76 ;
    wire THETA_n75 ;
    wire THETA_n74 ;
    wire THETA_n73 ;
    wire THETA_n72 ;
    wire THETA_n71 ;
    wire THETA_n70 ;
    wire THETA_n69 ;
    wire THETA_n68 ;
    wire THETA_n67 ;
    wire THETA_n66 ;
    wire THETA_n65 ;
    wire THETA_n64 ;
    wire THETA_n63 ;
    wire THETA_n62 ;
    wire THETA_n61 ;
    wire THETA_n60 ;
    wire THETA_n59 ;
    wire THETA_n58 ;
    wire THETA_n57 ;
    wire THETA_n56 ;
    wire THETA_n55 ;
    wire THETA_n54 ;
    wire THETA_n53 ;
    wire THETA_n52 ;
    wire THETA_n51 ;
    wire THETA_n50 ;
    wire THETA_n49 ;
    wire THETA_n48 ;
    wire THETA_n47 ;
    wire THETA_n46 ;
    wire THETA_n45 ;
    wire THETA_n44 ;
    wire THETA_n43 ;
    wire THETA_n42 ;
    wire THETA_n41 ;
    wire THETA_n40 ;
    wire THETA_n39 ;
    wire THETA_n38 ;
    wire THETA_n37 ;
    wire THETA_n36 ;
    wire THETA_n35 ;
    wire THETA_n34 ;
    wire THETA_n33 ;
    wire THETA_n32 ;
    wire THETA_n31 ;
    wire THETA_n30 ;
    wire THETA_n29 ;
    wire THETA_n28 ;
    wire THETA_n27 ;
    wire THETA_n26 ;
    wire THETA_n25 ;
    wire THETA_n24 ;
    wire THETA_n23 ;
    wire THETA_n22 ;
    wire THETA_n21 ;
    wire THETA_n20 ;
    wire THETA_n19 ;
    wire THETA_n18 ;
    wire THETA_n17 ;
    wire THETA_n16 ;
    wire THETA_n15 ;
    wire THETA_n14 ;
    wire THETA_n13 ;
    wire THETA_n12 ;
    wire THETA_n11 ;
    wire THETA_n10 ;
    wire THETA_n9 ;
    wire THETA_n8 ;
    wire THETA_n7 ;
    wire THETA_n6 ;
    wire THETA_n5 ;
    wire THETA_n4 ;
    wire THETA_n3 ;
    wire THETA_n2 ;
    wire THETA_n1 ;
    wire CHI_ChiOut_3 ;
    wire CHI_ChiOut_7 ;
    wire CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_1__GEN_ROWS_0__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_1__GEN_ROWS_0__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_1__GEN_ROWS_0__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_1__GEN_ROWS_0__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_1__GEN_ROWS_0__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_1__GEN_ROWS_1__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_1__GEN_ROWS_1__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_1__GEN_ROWS_1__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_1__GEN_ROWS_1__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_1__GEN_ROWS_1__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_1__GEN_ROWS_2__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_1__GEN_ROWS_2__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_1__GEN_ROWS_2__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_1__GEN_ROWS_2__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_1__GEN_ROWS_2__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_1__GEN_ROWS_3__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_1__GEN_ROWS_3__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_1__GEN_ROWS_3__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_1__GEN_ROWS_3__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_1__GEN_ROWS_3__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_1__GEN_ROWS_4__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_1__GEN_ROWS_4__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_1__GEN_ROWS_4__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_1__GEN_ROWS_4__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_1__GEN_ROWS_4__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_2__GEN_ROWS_0__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_2__GEN_ROWS_0__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_2__GEN_ROWS_0__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_2__GEN_ROWS_0__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_2__GEN_ROWS_0__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_2__GEN_ROWS_1__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_2__GEN_ROWS_1__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_2__GEN_ROWS_1__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_2__GEN_ROWS_1__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_2__GEN_ROWS_1__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_2__GEN_ROWS_2__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_2__GEN_ROWS_2__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_2__GEN_ROWS_2__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_2__GEN_ROWS_2__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_2__GEN_ROWS_2__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_2__GEN_ROWS_3__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_2__GEN_ROWS_3__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_2__GEN_ROWS_3__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_2__GEN_ROWS_3__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_2__GEN_ROWS_3__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_2__GEN_ROWS_4__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_2__GEN_ROWS_4__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_2__GEN_ROWS_4__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_2__GEN_ROWS_4__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_2__GEN_ROWS_4__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_3__GEN_ROWS_0__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_3__GEN_ROWS_0__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_3__GEN_ROWS_0__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_3__GEN_ROWS_0__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_3__GEN_ROWS_0__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_3__GEN_ROWS_1__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_3__GEN_ROWS_1__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_3__GEN_ROWS_1__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_3__GEN_ROWS_1__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_3__GEN_ROWS_1__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_3__GEN_ROWS_2__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_3__GEN_ROWS_2__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_3__GEN_ROWS_2__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_3__GEN_ROWS_2__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_3__GEN_ROWS_2__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_3__GEN_ROWS_3__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_3__GEN_ROWS_3__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_3__GEN_ROWS_3__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_3__GEN_ROWS_3__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_3__GEN_ROWS_3__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_3__GEN_ROWS_4__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_3__GEN_ROWS_4__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_3__GEN_ROWS_4__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_3__GEN_ROWS_4__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_3__GEN_ROWS_4__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_4__GEN_ROWS_0__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_4__GEN_ROWS_0__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_4__GEN_ROWS_0__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_4__GEN_ROWS_0__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_4__GEN_ROWS_0__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_4__GEN_ROWS_1__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_4__GEN_ROWS_1__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_4__GEN_ROWS_1__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_4__GEN_ROWS_1__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_4__GEN_ROWS_1__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_4__GEN_ROWS_2__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_4__GEN_ROWS_2__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_4__GEN_ROWS_2__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_4__GEN_ROWS_2__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_4__GEN_ROWS_2__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_4__GEN_ROWS_3__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_4__GEN_ROWS_3__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_4__GEN_ROWS_3__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_4__GEN_ROWS_3__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_4__GEN_ROWS_3__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_4__GEN_ROWS_4__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_4__GEN_ROWS_4__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_4__GEN_ROWS_4__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_4__GEN_ROWS_4__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_4__GEN_ROWS_4__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_5__GEN_ROWS_0__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_5__GEN_ROWS_0__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_5__GEN_ROWS_0__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_5__GEN_ROWS_0__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_5__GEN_ROWS_0__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_5__GEN_ROWS_1__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_5__GEN_ROWS_1__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_5__GEN_ROWS_1__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_5__GEN_ROWS_1__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_5__GEN_ROWS_1__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_5__GEN_ROWS_2__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_5__GEN_ROWS_2__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_5__GEN_ROWS_2__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_5__GEN_ROWS_2__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_5__GEN_ROWS_2__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_5__GEN_ROWS_3__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_5__GEN_ROWS_3__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_5__GEN_ROWS_3__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_5__GEN_ROWS_3__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_5__GEN_ROWS_3__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_5__GEN_ROWS_4__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_5__GEN_ROWS_4__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_5__GEN_ROWS_4__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_5__GEN_ROWS_4__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_5__GEN_ROWS_4__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_6__GEN_ROWS_0__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_6__GEN_ROWS_0__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_6__GEN_ROWS_0__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_6__GEN_ROWS_0__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_6__GEN_ROWS_0__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_6__GEN_ROWS_1__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_6__GEN_ROWS_1__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_6__GEN_ROWS_1__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_6__GEN_ROWS_1__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_6__GEN_ROWS_1__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_6__GEN_ROWS_2__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_6__GEN_ROWS_2__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_6__GEN_ROWS_2__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_6__GEN_ROWS_2__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_6__GEN_ROWS_2__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_6__GEN_ROWS_3__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_6__GEN_ROWS_3__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_6__GEN_ROWS_3__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_6__GEN_ROWS_3__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_6__GEN_ROWS_3__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_6__GEN_ROWS_4__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_6__GEN_ROWS_4__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_6__GEN_ROWS_4__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_6__GEN_ROWS_4__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_6__GEN_ROWS_4__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_7__GEN_ROWS_0__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_7__GEN_ROWS_0__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_7__GEN_ROWS_0__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_7__GEN_ROWS_0__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_7__GEN_ROWS_0__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_7__GEN_ROWS_1__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_7__GEN_ROWS_1__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_7__GEN_ROWS_1__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_7__GEN_ROWS_1__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_7__GEN_ROWS_1__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_7__GEN_ROWS_2__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_7__GEN_ROWS_2__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_7__GEN_ROWS_2__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_7__GEN_ROWS_2__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_7__GEN_ROWS_2__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_7__GEN_ROWS_3__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_7__GEN_ROWS_3__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_7__GEN_ROWS_3__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_7__GEN_ROWS_3__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_7__GEN_ROWS_3__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_7__GEN_ROWS_4__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_7__GEN_ROWS_4__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_7__GEN_ROWS_4__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_7__GEN_ROWS_4__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_7__GEN_ROWS_4__sbox_and_xor_inst_e_nxy ;
    wire KECCAK_CONTROL_n47 ;
    wire KECCAK_CONTROL_n45 ;
    wire KECCAK_CONTROL_n44 ;
    wire KECCAK_CONTROL_n43 ;
    wire KECCAK_CONTROL_n34 ;
    wire KECCAK_CONTROL_n33 ;
    wire KECCAK_CONTROL_n32 ;
    wire KECCAK_CONTROL_n30 ;
    wire KECCAK_CONTROL_n29 ;
    wire KECCAK_CONTROL_n28 ;
    wire KECCAK_CONTROL_n27 ;
    wire KECCAK_CONTROL_n25 ;
    wire KECCAK_CONTROL_n23 ;
    wire KECCAK_CONTROL_n22 ;
    wire KECCAK_CONTROL_n21 ;
    wire KECCAK_CONTROL_n20 ;
    wire KECCAK_CONTROL_n19 ;
    wire KECCAK_CONTROL_n18 ;
    wire KECCAK_CONTROL_n17 ;
    wire KECCAK_CONTROL_n16 ;
    wire KECCAK_CONTROL_n15 ;
    wire KECCAK_CONTROL_n14 ;
    wire KECCAK_CONTROL_n13 ;
    wire KECCAK_CONTROL_n11 ;
    wire KECCAK_CONTROL_n10 ;
    wire KECCAK_CONTROL_n8 ;
    wire KECCAK_CONTROL_CtrlStatexDP_reg_1__Q ;
    wire KECCAK_CONTROL_RoundCountLastxDP_reg_Q ;
    wire KECCAK_CONTROL_RC_GEN_n28 ;
    wire KECCAK_CONTROL_RC_GEN_n27 ;
    wire KECCAK_CONTROL_RC_GEN_n26 ;
    wire KECCAK_CONTROL_RC_GEN_n25 ;
    wire KECCAK_CONTROL_RC_GEN_n22 ;
    wire KECCAK_CONTROL_RC_GEN_n19 ;
    wire KECCAK_CONTROL_RC_GEN_n18 ;
    wire KECCAK_CONTROL_RC_GEN_n17 ;
    wire KECCAK_CONTROL_RC_GEN_n15 ;
    wire KECCAK_CONTROL_RC_GEN_n14 ;
    wire KECCAK_CONTROL_RC_GEN_n13 ;
    wire KECCAK_CONTROL_RC_GEN_n12 ;
    wire KECCAK_CONTROL_RC_GEN_n11 ;
    wire KECCAK_CONTROL_RC_GEN_n9 ;
    wire KECCAK_CONTROL_RC_GEN_n8 ;
    wire KECCAK_CONTROL_RC_GEN_n6 ;
    wire KECCAK_CONTROL_RC_GEN_n5 ;
    wire KECCAK_CONTROL_RC_GEN_n4 ;
    wire KECCAK_CONTROL_RC_GEN_n3 ;
    wire KECCAK_CONTROL_RC_GEN_n2 ;
    wire KECCAK_CONTROL_RC_GEN_n30 ;
    wire KECCAK_CONTROL_RC_GEN_n31 ;
    wire KECCAK_CONTROL_RC_GEN_n23 ;
    wire KECCAK_CONTROL_RC_GEN_n24 ;
    wire KECCAK_CONTROL_RC_GEN_n20 ;
    wire KECCAK_CONTROL_RC_GEN_n21 ;
    wire KECCAK_CONTROL_RC_GEN_U25_Y ;
    wire KECCAK_CONTROL_RC_GEN_U25_X ;
    wire KECCAK_CONTROL_RC_GEN_U28_Y ;
    wire KECCAK_CONTROL_RC_GEN_U28_X ;
    wire KECCAK_CONTROL_RC_GEN_U32_Y ;
    wire KECCAK_CONTROL_RC_GEN_U32_X ;
    wire U810_Y ;
    wire U810_X ;
    wire U812_Y ;
    wire U812_X ;
    wire U814_Y ;
    wire U814_X ;
    wire U816_Y ;
    wire U816_X ;
    wire U817_Y ;
    wire U817_X ;
    wire U818_Y ;
    wire U818_X ;
    wire U820_Y ;
    wire U820_X ;
    wire U821_Y ;
    wire U821_X ;
    wire U822_Y ;
    wire U822_X ;
    wire U823_Y ;
    wire U823_X ;
    wire U824_Y ;
    wire U824_X ;
    wire U825_Y ;
    wire U825_X ;
    wire U827_Y ;
    wire U827_X ;
    wire U828_Y ;
    wire U828_X ;
    wire U830_Y ;
    wire U830_X ;
    wire U831_Y ;
    wire U831_X ;
    wire U832_Y ;
    wire U832_X ;
    wire U833_Y ;
    wire U833_X ;
    wire U834_Y ;
    wire U834_X ;
    wire U835_Y ;
    wire U835_X ;
    wire U836_Y ;
    wire U836_X ;
    wire U837_Y ;
    wire U837_X ;
    wire U838_Y ;
    wire U838_X ;
    wire U839_Y ;
    wire U839_X ;
    wire U841_Y ;
    wire U841_X ;
    wire U842_Y ;
    wire U842_X ;
    wire U843_Y ;
    wire U843_X ;
    wire U844_Y ;
    wire U844_X ;
    wire U845_Y ;
    wire U845_X ;
    wire U846_Y ;
    wire U846_X ;
    wire U847_Y ;
    wire U847_X ;
    wire U848_Y ;
    wire U848_X ;
    wire U849_Y ;
    wire U849_X ;
    wire U850_Y ;
    wire U850_X ;
    wire U851_Y ;
    wire U851_X ;
    wire U852_Y ;
    wire U852_X ;
    wire U853_Y ;
    wire U853_X ;
    wire U854_Y ;
    wire U854_X ;
    wire U855_Y ;
    wire U855_X ;
    wire U856_Y ;
    wire U856_X ;
    wire U857_Y ;
    wire U857_X ;
    wire U858_Y ;
    wire U858_X ;
    wire U859_Y ;
    wire U859_X ;
    wire U860_Y ;
    wire U860_X ;
    wire U861_Y ;
    wire U861_X ;
    wire U862_Y ;
    wire U862_X ;
    wire U863_Y ;
    wire U863_X ;
    wire U864_Y ;
    wire U864_X ;
    wire U865_Y ;
    wire U865_X ;
    wire U866_Y ;
    wire U866_X ;
    wire U867_Y ;
    wire U867_X ;
    wire U868_Y ;
    wire U868_X ;
    wire U869_Y ;
    wire U869_X ;
    wire U870_Y ;
    wire U870_X ;
    wire U871_Y ;
    wire U871_X ;
    wire U872_Y ;
    wire U872_X ;
    wire U873_Y ;
    wire U873_X ;
    wire U874_Y ;
    wire U874_X ;
    wire U875_Y ;
    wire U875_X ;
    wire U876_Y ;
    wire U876_X ;
    wire U877_Y ;
    wire U877_X ;
    wire U878_Y ;
    wire U878_X ;
    wire U879_Y ;
    wire U879_X ;
    wire U880_Y ;
    wire U880_X ;
    wire U881_Y ;
    wire U881_X ;
    wire U882_Y ;
    wire U882_X ;
    wire U883_Y ;
    wire U883_X ;
    wire U884_Y ;
    wire U884_X ;
    wire U885_Y ;
    wire U885_X ;
    wire U886_Y ;
    wire U886_X ;
    wire U887_Y ;
    wire U887_X ;
    wire U888_Y ;
    wire U888_X ;
    wire U889_Y ;
    wire U889_X ;
    wire U890_Y ;
    wire U890_X ;
    wire U891_Y ;
    wire U891_X ;
    wire U892_Y ;
    wire U892_X ;
    wire U893_Y ;
    wire U893_X ;
    wire U894_Y ;
    wire U894_X ;
    wire U895_Y ;
    wire U895_X ;
    wire U896_Y ;
    wire U896_X ;
    wire U897_Y ;
    wire U897_X ;
    wire U898_Y ;
    wire U898_X ;
    wire U899_Y ;
    wire U899_X ;
    wire U900_Y ;
    wire U900_X ;
    wire U901_Y ;
    wire U901_X ;
    wire U902_Y ;
    wire U902_X ;
    wire U903_Y ;
    wire U903_X ;
    wire U904_Y ;
    wire U904_X ;
    wire U905_Y ;
    wire U905_X ;
    wire U906_Y ;
    wire U906_X ;
    wire U907_Y ;
    wire U907_X ;
    wire U908_Y ;
    wire U908_X ;
    wire U909_Y ;
    wire U909_X ;
    wire U910_Y ;
    wire U910_X ;
    wire U911_Y ;
    wire U911_X ;
    wire U912_Y ;
    wire U912_X ;
    wire U913_Y ;
    wire U913_X ;
    wire U914_Y ;
    wire U914_X ;
    wire U915_Y ;
    wire U915_X ;
    wire U916_Y ;
    wire U916_X ;
    wire U917_Y ;
    wire U917_X ;
    wire U918_Y ;
    wire U918_X ;
    wire U919_Y ;
    wire U919_X ;
    wire U920_Y ;
    wire U920_X ;
    wire U921_Y ;
    wire U921_X ;
    wire U922_Y ;
    wire U922_X ;
    wire U923_Y ;
    wire U923_X ;
    wire U924_Y ;
    wire U924_X ;
    wire U925_Y ;
    wire U925_X ;
    wire U926_Y ;
    wire U926_X ;
    wire U927_Y ;
    wire U927_X ;
    wire U928_Y ;
    wire U928_X ;
    wire U929_Y ;
    wire U929_X ;
    wire U930_Y ;
    wire U930_X ;
    wire U931_Y ;
    wire U931_X ;
    wire U932_Y ;
    wire U932_X ;
    wire U933_Y ;
    wire U933_X ;
    wire U934_Y ;
    wire U934_X ;
    wire U935_Y ;
    wire U935_X ;
    wire U936_Y ;
    wire U936_X ;
    wire U937_Y ;
    wire U937_X ;
    wire U938_Y ;
    wire U938_X ;
    wire U939_Y ;
    wire U939_X ;
    wire U940_Y ;
    wire U940_X ;
    wire U941_Y ;
    wire U941_X ;
    wire U942_Y ;
    wire U942_X ;
    wire U943_Y ;
    wire U943_X ;
    wire U944_Y ;
    wire U944_X ;
    wire U945_Y ;
    wire U945_X ;
    wire U946_Y ;
    wire U946_X ;
    wire U947_Y ;
    wire U947_X ;
    wire U948_Y ;
    wire U948_X ;
    wire U949_Y ;
    wire U949_X ;
    wire U950_Y ;
    wire U950_X ;
    wire U951_Y ;
    wire U951_X ;
    wire U952_Y ;
    wire U952_X ;
    wire U953_Y ;
    wire U953_X ;
    wire U954_Y ;
    wire U954_X ;
    wire U955_Y ;
    wire U955_X ;
    wire U956_Y ;
    wire U956_X ;
    wire U957_Y ;
    wire U957_X ;
    wire U958_Y ;
    wire U958_X ;
    wire U959_Y ;
    wire U959_X ;
    wire U960_Y ;
    wire U960_X ;
    wire U961_Y ;
    wire U961_X ;
    wire U962_Y ;
    wire U962_X ;
    wire U963_Y ;
    wire U963_X ;
    wire U964_Y ;
    wire U964_X ;
    wire U965_Y ;
    wire U965_X ;
    wire U966_Y ;
    wire U966_X ;
    wire U967_Y ;
    wire U967_X ;
    wire U968_Y ;
    wire U968_X ;
    wire U969_Y ;
    wire U969_X ;
    wire U970_Y ;
    wire U970_X ;
    wire U971_Y ;
    wire U971_X ;
    wire U972_Y ;
    wire U972_X ;
    wire U973_Y ;
    wire U973_X ;
    wire U974_Y ;
    wire U974_X ;
    wire U975_Y ;
    wire U975_X ;
    wire U976_Y ;
    wire U976_X ;
    wire U977_Y ;
    wire U977_X ;
    wire U978_Y ;
    wire U978_X ;
    wire U979_Y ;
    wire U979_X ;
    wire U980_Y ;
    wire U980_X ;
    wire U981_Y ;
    wire U981_X ;
    wire U982_Y ;
    wire U982_X ;
    wire U983_Y ;
    wire U983_X ;
    wire U984_Y ;
    wire U984_X ;
    wire U985_Y ;
    wire U985_X ;
    wire U986_Y ;
    wire U986_X ;
    wire U987_Y ;
    wire U987_X ;
    wire U988_Y ;
    wire U988_X ;
    wire U989_Y ;
    wire U989_X ;
    wire U990_Y ;
    wire U990_X ;
    wire U991_Y ;
    wire U991_X ;
    wire U992_Y ;
    wire U992_X ;
    wire U993_Y ;
    wire U993_X ;
    wire U994_Y ;
    wire U994_X ;
    wire U995_Y ;
    wire U995_X ;
    wire U996_Y ;
    wire U996_X ;
    wire U997_Y ;
    wire U997_X ;
    wire U998_Y ;
    wire U998_X ;
    wire U999_Y ;
    wire U999_X ;
    wire U1000_Y ;
    wire U1000_X ;
    wire U1001_Y ;
    wire U1001_X ;
    wire U1002_Y ;
    wire U1002_X ;
    wire U1003_Y ;
    wire U1003_X ;
    wire U1004_Y ;
    wire U1004_X ;
    wire U1005_Y ;
    wire U1005_X ;
    wire U1006_Y ;
    wire U1006_X ;
    wire U1007_Y ;
    wire U1007_X ;
    wire U1008_Y ;
    wire U1008_X ;
    wire U1009_Y ;
    wire U1009_X ;
    wire U1010_Y ;
    wire U1010_X ;
    wire U1011_Y ;
    wire U1011_X ;
    wire U1012_Y ;
    wire U1012_X ;
    wire U1013_Y ;
    wire U1013_X ;
    wire U1014_Y ;
    wire U1014_X ;
    wire U1015_Y ;
    wire U1015_X ;
    wire U1016_Y ;
    wire U1016_X ;
    wire [199:8] StateOut ;
    wire [199:0] StateFromRhoPi ;
    wire [199:0] StateFromChi ;
    wire [1:0] IotaRC ;
    wire [1:0] CHI_ChiOut ;
    wire [4:0] KECCAK_CONTROL_RoundCountxDP ;
    wire [2:0] KECCAK_CONTROL_CtrlStatexDP ;
    wire new_AGEMA_signal_2130 ;
    wire new_AGEMA_signal_2131 ;
    wire new_AGEMA_signal_2132 ;
    wire new_AGEMA_signal_2133 ;
    wire new_AGEMA_signal_2134 ;
    wire new_AGEMA_signal_2135 ;
    wire new_AGEMA_signal_2136 ;
    wire new_AGEMA_signal_2137 ;
    wire new_AGEMA_signal_2138 ;
    wire new_AGEMA_signal_2139 ;
    wire new_AGEMA_signal_2140 ;
    wire new_AGEMA_signal_2141 ;
    wire new_AGEMA_signal_2142 ;
    wire new_AGEMA_signal_2143 ;
    wire new_AGEMA_signal_2144 ;
    wire new_AGEMA_signal_2145 ;
    wire new_AGEMA_signal_2146 ;
    wire new_AGEMA_signal_2147 ;
    wire new_AGEMA_signal_2148 ;
    wire new_AGEMA_signal_2149 ;
    wire new_AGEMA_signal_2150 ;
    wire new_AGEMA_signal_2151 ;
    wire new_AGEMA_signal_2152 ;
    wire new_AGEMA_signal_2153 ;
    wire new_AGEMA_signal_2154 ;
    wire new_AGEMA_signal_2155 ;
    wire new_AGEMA_signal_2156 ;
    wire new_AGEMA_signal_2157 ;
    wire new_AGEMA_signal_2158 ;
    wire new_AGEMA_signal_2159 ;
    wire new_AGEMA_signal_2160 ;
    wire new_AGEMA_signal_2161 ;
    wire new_AGEMA_signal_2162 ;
    wire new_AGEMA_signal_2163 ;
    wire new_AGEMA_signal_2164 ;
    wire new_AGEMA_signal_2165 ;
    wire new_AGEMA_signal_2166 ;
    wire new_AGEMA_signal_2167 ;
    wire new_AGEMA_signal_2168 ;
    wire new_AGEMA_signal_2169 ;
    wire new_AGEMA_signal_2170 ;
    wire new_AGEMA_signal_2171 ;
    wire new_AGEMA_signal_2172 ;
    wire new_AGEMA_signal_2173 ;
    wire new_AGEMA_signal_2174 ;
    wire new_AGEMA_signal_2175 ;
    wire new_AGEMA_signal_2176 ;
    wire new_AGEMA_signal_2177 ;
    wire new_AGEMA_signal_2178 ;
    wire new_AGEMA_signal_2179 ;
    wire new_AGEMA_signal_2180 ;
    wire new_AGEMA_signal_2181 ;
    wire new_AGEMA_signal_2182 ;
    wire new_AGEMA_signal_2183 ;
    wire new_AGEMA_signal_2184 ;
    wire new_AGEMA_signal_2185 ;
    wire new_AGEMA_signal_2186 ;
    wire new_AGEMA_signal_2187 ;
    wire new_AGEMA_signal_2188 ;
    wire new_AGEMA_signal_2189 ;
    wire new_AGEMA_signal_2190 ;
    wire new_AGEMA_signal_2191 ;
    wire new_AGEMA_signal_2192 ;
    wire new_AGEMA_signal_2193 ;
    wire new_AGEMA_signal_2194 ;
    wire new_AGEMA_signal_2195 ;
    wire new_AGEMA_signal_2196 ;
    wire new_AGEMA_signal_2197 ;
    wire new_AGEMA_signal_2198 ;
    wire new_AGEMA_signal_2199 ;
    wire new_AGEMA_signal_2200 ;
    wire new_AGEMA_signal_2201 ;
    wire new_AGEMA_signal_2202 ;
    wire new_AGEMA_signal_2203 ;
    wire new_AGEMA_signal_2204 ;
    wire new_AGEMA_signal_2205 ;
    wire new_AGEMA_signal_2206 ;
    wire new_AGEMA_signal_2207 ;
    wire new_AGEMA_signal_2208 ;
    wire new_AGEMA_signal_2209 ;
    wire new_AGEMA_signal_2210 ;
    wire new_AGEMA_signal_2211 ;
    wire new_AGEMA_signal_2212 ;
    wire new_AGEMA_signal_2213 ;
    wire new_AGEMA_signal_2214 ;
    wire new_AGEMA_signal_2215 ;
    wire new_AGEMA_signal_2216 ;
    wire new_AGEMA_signal_2217 ;
    wire new_AGEMA_signal_2218 ;
    wire new_AGEMA_signal_2219 ;
    wire new_AGEMA_signal_2220 ;
    wire new_AGEMA_signal_2221 ;
    wire new_AGEMA_signal_2222 ;
    wire new_AGEMA_signal_2223 ;
    wire new_AGEMA_signal_2224 ;
    wire new_AGEMA_signal_2225 ;
    wire new_AGEMA_signal_2226 ;
    wire new_AGEMA_signal_2227 ;
    wire new_AGEMA_signal_2228 ;
    wire new_AGEMA_signal_2229 ;
    wire new_AGEMA_signal_2230 ;
    wire new_AGEMA_signal_2231 ;
    wire new_AGEMA_signal_2232 ;
    wire new_AGEMA_signal_2233 ;
    wire new_AGEMA_signal_2234 ;
    wire new_AGEMA_signal_2235 ;
    wire new_AGEMA_signal_2236 ;
    wire new_AGEMA_signal_2237 ;
    wire new_AGEMA_signal_2238 ;
    wire new_AGEMA_signal_2239 ;
    wire new_AGEMA_signal_2240 ;
    wire new_AGEMA_signal_2241 ;
    wire new_AGEMA_signal_2242 ;
    wire new_AGEMA_signal_2243 ;
    wire new_AGEMA_signal_2244 ;
    wire new_AGEMA_signal_2245 ;
    wire new_AGEMA_signal_2246 ;
    wire new_AGEMA_signal_2247 ;
    wire new_AGEMA_signal_2248 ;
    wire new_AGEMA_signal_2249 ;
    wire new_AGEMA_signal_2250 ;
    wire new_AGEMA_signal_2251 ;
    wire new_AGEMA_signal_2252 ;
    wire new_AGEMA_signal_2253 ;
    wire new_AGEMA_signal_2254 ;
    wire new_AGEMA_signal_2255 ;
    wire new_AGEMA_signal_2256 ;
    wire new_AGEMA_signal_2257 ;
    wire new_AGEMA_signal_2258 ;
    wire new_AGEMA_signal_2259 ;
    wire new_AGEMA_signal_2260 ;
    wire new_AGEMA_signal_2261 ;
    wire new_AGEMA_signal_2262 ;
    wire new_AGEMA_signal_2263 ;
    wire new_AGEMA_signal_2264 ;
    wire new_AGEMA_signal_2265 ;
    wire new_AGEMA_signal_2266 ;
    wire new_AGEMA_signal_2267 ;
    wire new_AGEMA_signal_2268 ;
    wire new_AGEMA_signal_2269 ;
    wire new_AGEMA_signal_2270 ;
    wire new_AGEMA_signal_2271 ;
    wire new_AGEMA_signal_2272 ;
    wire new_AGEMA_signal_2273 ;
    wire new_AGEMA_signal_2274 ;
    wire new_AGEMA_signal_2275 ;
    wire new_AGEMA_signal_2276 ;
    wire new_AGEMA_signal_2277 ;
    wire new_AGEMA_signal_2278 ;
    wire new_AGEMA_signal_2279 ;
    wire new_AGEMA_signal_2280 ;
    wire new_AGEMA_signal_2281 ;
    wire new_AGEMA_signal_2282 ;
    wire new_AGEMA_signal_2283 ;
    wire new_AGEMA_signal_2284 ;
    wire new_AGEMA_signal_2285 ;
    wire new_AGEMA_signal_2286 ;
    wire new_AGEMA_signal_2287 ;
    wire new_AGEMA_signal_2288 ;
    wire new_AGEMA_signal_2289 ;
    wire new_AGEMA_signal_2290 ;
    wire new_AGEMA_signal_2291 ;
    wire new_AGEMA_signal_2292 ;
    wire new_AGEMA_signal_2293 ;
    wire new_AGEMA_signal_2294 ;
    wire new_AGEMA_signal_2295 ;
    wire new_AGEMA_signal_2296 ;
    wire new_AGEMA_signal_2297 ;
    wire new_AGEMA_signal_2298 ;
    wire new_AGEMA_signal_2299 ;
    wire new_AGEMA_signal_2300 ;
    wire new_AGEMA_signal_2301 ;
    wire new_AGEMA_signal_2302 ;
    wire new_AGEMA_signal_2303 ;
    wire new_AGEMA_signal_2304 ;
    wire new_AGEMA_signal_2305 ;
    wire new_AGEMA_signal_2306 ;
    wire new_AGEMA_signal_2307 ;
    wire new_AGEMA_signal_2308 ;
    wire new_AGEMA_signal_2309 ;
    wire new_AGEMA_signal_2310 ;
    wire new_AGEMA_signal_2311 ;
    wire new_AGEMA_signal_2312 ;
    wire new_AGEMA_signal_2313 ;
    wire new_AGEMA_signal_2314 ;
    wire new_AGEMA_signal_2315 ;
    wire new_AGEMA_signal_2316 ;
    wire new_AGEMA_signal_2317 ;
    wire new_AGEMA_signal_2318 ;
    wire new_AGEMA_signal_2319 ;
    wire new_AGEMA_signal_2320 ;
    wire new_AGEMA_signal_2321 ;
    wire new_AGEMA_signal_2322 ;
    wire new_AGEMA_signal_2323 ;
    wire new_AGEMA_signal_2324 ;
    wire new_AGEMA_signal_2325 ;
    wire new_AGEMA_signal_2326 ;
    wire new_AGEMA_signal_2327 ;
    wire new_AGEMA_signal_2328 ;
    wire new_AGEMA_signal_2329 ;
    wire new_AGEMA_signal_2330 ;
    wire new_AGEMA_signal_2331 ;
    wire new_AGEMA_signal_2332 ;
    wire new_AGEMA_signal_2333 ;
    wire new_AGEMA_signal_2334 ;
    wire new_AGEMA_signal_2335 ;
    wire new_AGEMA_signal_2336 ;
    wire new_AGEMA_signal_2337 ;
    wire new_AGEMA_signal_2338 ;
    wire new_AGEMA_signal_2339 ;
    wire new_AGEMA_signal_2340 ;
    wire new_AGEMA_signal_2341 ;
    wire new_AGEMA_signal_2342 ;
    wire new_AGEMA_signal_2343 ;
    wire new_AGEMA_signal_2344 ;
    wire new_AGEMA_signal_2345 ;
    wire new_AGEMA_signal_2346 ;
    wire new_AGEMA_signal_2347 ;
    wire new_AGEMA_signal_2348 ;
    wire new_AGEMA_signal_2349 ;
    wire new_AGEMA_signal_2350 ;
    wire new_AGEMA_signal_2351 ;
    wire new_AGEMA_signal_2352 ;
    wire new_AGEMA_signal_2353 ;
    wire new_AGEMA_signal_2354 ;
    wire new_AGEMA_signal_2355 ;
    wire new_AGEMA_signal_2356 ;
    wire new_AGEMA_signal_2357 ;
    wire new_AGEMA_signal_2358 ;
    wire new_AGEMA_signal_2359 ;
    wire new_AGEMA_signal_2360 ;
    wire new_AGEMA_signal_2361 ;
    wire new_AGEMA_signal_2362 ;
    wire new_AGEMA_signal_2363 ;
    wire new_AGEMA_signal_2364 ;
    wire new_AGEMA_signal_2365 ;
    wire new_AGEMA_signal_2366 ;
    wire new_AGEMA_signal_2367 ;
    wire new_AGEMA_signal_2368 ;
    wire new_AGEMA_signal_2369 ;
    wire new_AGEMA_signal_2370 ;
    wire new_AGEMA_signal_2371 ;
    wire new_AGEMA_signal_2372 ;
    wire new_AGEMA_signal_2373 ;
    wire new_AGEMA_signal_2374 ;
    wire new_AGEMA_signal_2375 ;
    wire new_AGEMA_signal_2376 ;
    wire new_AGEMA_signal_2377 ;
    wire new_AGEMA_signal_2378 ;
    wire new_AGEMA_signal_2379 ;
    wire new_AGEMA_signal_2380 ;
    wire new_AGEMA_signal_2381 ;
    wire new_AGEMA_signal_2382 ;
    wire new_AGEMA_signal_2383 ;
    wire new_AGEMA_signal_2384 ;
    wire new_AGEMA_signal_2385 ;
    wire new_AGEMA_signal_2386 ;
    wire new_AGEMA_signal_2387 ;
    wire new_AGEMA_signal_2388 ;
    wire new_AGEMA_signal_2389 ;
    wire new_AGEMA_signal_2390 ;
    wire new_AGEMA_signal_2391 ;
    wire new_AGEMA_signal_2392 ;
    wire new_AGEMA_signal_2393 ;
    wire new_AGEMA_signal_2394 ;
    wire new_AGEMA_signal_2395 ;
    wire new_AGEMA_signal_2396 ;
    wire new_AGEMA_signal_2397 ;
    wire new_AGEMA_signal_2398 ;
    wire new_AGEMA_signal_2399 ;
    wire new_AGEMA_signal_2400 ;
    wire new_AGEMA_signal_2401 ;
    wire new_AGEMA_signal_2402 ;
    wire new_AGEMA_signal_2403 ;
    wire new_AGEMA_signal_2404 ;
    wire new_AGEMA_signal_2405 ;
    wire new_AGEMA_signal_2406 ;
    wire new_AGEMA_signal_2407 ;
    wire new_AGEMA_signal_2408 ;
    wire new_AGEMA_signal_2409 ;
    wire new_AGEMA_signal_2410 ;
    wire new_AGEMA_signal_2411 ;
    wire new_AGEMA_signal_2412 ;
    wire new_AGEMA_signal_2413 ;
    wire new_AGEMA_signal_2414 ;
    wire new_AGEMA_signal_2415 ;
    wire new_AGEMA_signal_2416 ;
    wire new_AGEMA_signal_2417 ;
    wire new_AGEMA_signal_2418 ;
    wire new_AGEMA_signal_2419 ;
    wire new_AGEMA_signal_2420 ;
    wire new_AGEMA_signal_2421 ;
    wire new_AGEMA_signal_2422 ;
    wire new_AGEMA_signal_2423 ;
    wire new_AGEMA_signal_2424 ;
    wire new_AGEMA_signal_2425 ;
    wire new_AGEMA_signal_2426 ;
    wire new_AGEMA_signal_2427 ;
    wire new_AGEMA_signal_2428 ;
    wire new_AGEMA_signal_2429 ;
    wire new_AGEMA_signal_2430 ;
    wire new_AGEMA_signal_2431 ;
    wire new_AGEMA_signal_2432 ;
    wire new_AGEMA_signal_2433 ;
    wire new_AGEMA_signal_2434 ;
    wire new_AGEMA_signal_2435 ;
    wire new_AGEMA_signal_2436 ;
    wire new_AGEMA_signal_2437 ;
    wire new_AGEMA_signal_2438 ;
    wire new_AGEMA_signal_2439 ;
    wire new_AGEMA_signal_2440 ;
    wire new_AGEMA_signal_2441 ;
    wire new_AGEMA_signal_2442 ;
    wire new_AGEMA_signal_2443 ;
    wire new_AGEMA_signal_2444 ;
    wire new_AGEMA_signal_2445 ;
    wire new_AGEMA_signal_2446 ;
    wire new_AGEMA_signal_2447 ;
    wire new_AGEMA_signal_2448 ;
    wire new_AGEMA_signal_2449 ;
    wire new_AGEMA_signal_2450 ;
    wire new_AGEMA_signal_2451 ;
    wire new_AGEMA_signal_2452 ;
    wire new_AGEMA_signal_2453 ;
    wire new_AGEMA_signal_2454 ;
    wire new_AGEMA_signal_2455 ;
    wire new_AGEMA_signal_2456 ;
    wire new_AGEMA_signal_2457 ;
    wire new_AGEMA_signal_2458 ;
    wire new_AGEMA_signal_2459 ;
    wire new_AGEMA_signal_2460 ;
    wire new_AGEMA_signal_2461 ;
    wire new_AGEMA_signal_2462 ;
    wire new_AGEMA_signal_2463 ;
    wire new_AGEMA_signal_2464 ;
    wire new_AGEMA_signal_2465 ;
    wire new_AGEMA_signal_2466 ;
    wire new_AGEMA_signal_2467 ;
    wire new_AGEMA_signal_2468 ;
    wire new_AGEMA_signal_2469 ;
    wire new_AGEMA_signal_2470 ;
    wire new_AGEMA_signal_2471 ;
    wire new_AGEMA_signal_2472 ;
    wire new_AGEMA_signal_2473 ;
    wire new_AGEMA_signal_2474 ;
    wire new_AGEMA_signal_2475 ;
    wire new_AGEMA_signal_2476 ;
    wire new_AGEMA_signal_2477 ;
    wire new_AGEMA_signal_2478 ;
    wire new_AGEMA_signal_2479 ;
    wire new_AGEMA_signal_2480 ;
    wire new_AGEMA_signal_2481 ;
    wire new_AGEMA_signal_2482 ;
    wire new_AGEMA_signal_2483 ;
    wire new_AGEMA_signal_2484 ;
    wire new_AGEMA_signal_2485 ;
    wire new_AGEMA_signal_2486 ;
    wire new_AGEMA_signal_2487 ;
    wire new_AGEMA_signal_2488 ;
    wire new_AGEMA_signal_2489 ;
    wire new_AGEMA_signal_2490 ;
    wire new_AGEMA_signal_2491 ;
    wire new_AGEMA_signal_2492 ;
    wire new_AGEMA_signal_2493 ;
    wire new_AGEMA_signal_2494 ;
    wire new_AGEMA_signal_2495 ;
    wire new_AGEMA_signal_2496 ;
    wire new_AGEMA_signal_2497 ;
    wire new_AGEMA_signal_2498 ;
    wire new_AGEMA_signal_2499 ;
    wire new_AGEMA_signal_2500 ;
    wire new_AGEMA_signal_2501 ;
    wire new_AGEMA_signal_2502 ;
    wire new_AGEMA_signal_2503 ;
    wire new_AGEMA_signal_2504 ;
    wire new_AGEMA_signal_2505 ;
    wire new_AGEMA_signal_2506 ;
    wire new_AGEMA_signal_2507 ;
    wire new_AGEMA_signal_2508 ;
    wire new_AGEMA_signal_2509 ;
    wire new_AGEMA_signal_2510 ;
    wire new_AGEMA_signal_2511 ;
    wire new_AGEMA_signal_2512 ;
    wire new_AGEMA_signal_2513 ;
    wire new_AGEMA_signal_2514 ;
    wire new_AGEMA_signal_2515 ;
    wire new_AGEMA_signal_2516 ;
    wire new_AGEMA_signal_2517 ;
    wire new_AGEMA_signal_2518 ;
    wire new_AGEMA_signal_2519 ;
    wire new_AGEMA_signal_2520 ;
    wire new_AGEMA_signal_2521 ;
    wire new_AGEMA_signal_2522 ;
    wire new_AGEMA_signal_2523 ;
    wire new_AGEMA_signal_2524 ;
    wire new_AGEMA_signal_2525 ;
    wire new_AGEMA_signal_2526 ;
    wire new_AGEMA_signal_2527 ;
    wire new_AGEMA_signal_2528 ;
    wire new_AGEMA_signal_2532 ;
    wire new_AGEMA_signal_2533 ;
    wire new_AGEMA_signal_2534 ;
    wire new_AGEMA_signal_2535 ;
    wire new_AGEMA_signal_2536 ;
    wire new_AGEMA_signal_2537 ;
    wire new_AGEMA_signal_2538 ;
    wire new_AGEMA_signal_2539 ;
    wire new_AGEMA_signal_2540 ;
    wire new_AGEMA_signal_2541 ;
    wire new_AGEMA_signal_2542 ;
    wire new_AGEMA_signal_2543 ;
    wire new_AGEMA_signal_2544 ;
    wire new_AGEMA_signal_2545 ;
    wire new_AGEMA_signal_2546 ;
    wire new_AGEMA_signal_2547 ;
    wire new_AGEMA_signal_2548 ;
    wire new_AGEMA_signal_2549 ;
    wire new_AGEMA_signal_2550 ;
    wire new_AGEMA_signal_2551 ;
    wire new_AGEMA_signal_2552 ;
    wire new_AGEMA_signal_2553 ;
    wire new_AGEMA_signal_2554 ;
    wire new_AGEMA_signal_2555 ;
    wire new_AGEMA_signal_2556 ;
    wire new_AGEMA_signal_2557 ;
    wire new_AGEMA_signal_2558 ;
    wire new_AGEMA_signal_2559 ;
    wire new_AGEMA_signal_2560 ;
    wire new_AGEMA_signal_2561 ;
    wire new_AGEMA_signal_2562 ;
    wire new_AGEMA_signal_2563 ;
    wire new_AGEMA_signal_2564 ;
    wire new_AGEMA_signal_2565 ;
    wire new_AGEMA_signal_2566 ;
    wire new_AGEMA_signal_2567 ;
    wire new_AGEMA_signal_2568 ;
    wire new_AGEMA_signal_2569 ;
    wire new_AGEMA_signal_2570 ;
    wire new_AGEMA_signal_2571 ;
    wire new_AGEMA_signal_2572 ;
    wire new_AGEMA_signal_2573 ;
    wire new_AGEMA_signal_2574 ;
    wire new_AGEMA_signal_2575 ;
    wire new_AGEMA_signal_2576 ;
    wire new_AGEMA_signal_2577 ;
    wire new_AGEMA_signal_2578 ;
    wire new_AGEMA_signal_2579 ;
    wire new_AGEMA_signal_2580 ;
    wire new_AGEMA_signal_2581 ;
    wire new_AGEMA_signal_2582 ;
    wire new_AGEMA_signal_2583 ;
    wire new_AGEMA_signal_2584 ;
    wire new_AGEMA_signal_2585 ;
    wire new_AGEMA_signal_2586 ;
    wire new_AGEMA_signal_2587 ;
    wire new_AGEMA_signal_2588 ;
    wire new_AGEMA_signal_2589 ;
    wire new_AGEMA_signal_2590 ;
    wire new_AGEMA_signal_2591 ;
    wire new_AGEMA_signal_2592 ;
    wire new_AGEMA_signal_2593 ;
    wire new_AGEMA_signal_2594 ;
    wire new_AGEMA_signal_2595 ;
    wire new_AGEMA_signal_2596 ;
    wire new_AGEMA_signal_2597 ;
    wire new_AGEMA_signal_2598 ;
    wire new_AGEMA_signal_2599 ;
    wire new_AGEMA_signal_2600 ;
    wire new_AGEMA_signal_2601 ;
    wire new_AGEMA_signal_2602 ;
    wire new_AGEMA_signal_2603 ;
    wire new_AGEMA_signal_2604 ;
    wire new_AGEMA_signal_2605 ;
    wire new_AGEMA_signal_2606 ;
    wire new_AGEMA_signal_2607 ;
    wire new_AGEMA_signal_2608 ;
    wire new_AGEMA_signal_2609 ;
    wire new_AGEMA_signal_2610 ;
    wire new_AGEMA_signal_2611 ;
    wire new_AGEMA_signal_2612 ;
    wire new_AGEMA_signal_2613 ;
    wire new_AGEMA_signal_2614 ;
    wire new_AGEMA_signal_2615 ;
    wire new_AGEMA_signal_2616 ;
    wire new_AGEMA_signal_2617 ;
    wire new_AGEMA_signal_2618 ;
    wire new_AGEMA_signal_2619 ;
    wire new_AGEMA_signal_2620 ;
    wire new_AGEMA_signal_2621 ;
    wire new_AGEMA_signal_2622 ;
    wire new_AGEMA_signal_2623 ;
    wire new_AGEMA_signal_2624 ;
    wire new_AGEMA_signal_2625 ;
    wire new_AGEMA_signal_2626 ;
    wire new_AGEMA_signal_2627 ;
    wire new_AGEMA_signal_2628 ;
    wire new_AGEMA_signal_2629 ;
    wire new_AGEMA_signal_2630 ;
    wire new_AGEMA_signal_2631 ;
    wire new_AGEMA_signal_2632 ;
    wire new_AGEMA_signal_2633 ;
    wire new_AGEMA_signal_2634 ;
    wire new_AGEMA_signal_2635 ;
    wire new_AGEMA_signal_2636 ;
    wire new_AGEMA_signal_2640 ;
    wire new_AGEMA_signal_2641 ;
    wire new_AGEMA_signal_2642 ;
    wire new_AGEMA_signal_2643 ;
    wire new_AGEMA_signal_2644 ;
    wire new_AGEMA_signal_2645 ;
    wire new_AGEMA_signal_2646 ;
    wire new_AGEMA_signal_2647 ;
    wire new_AGEMA_signal_2648 ;
    wire new_AGEMA_signal_2649 ;
    wire new_AGEMA_signal_2650 ;
    wire new_AGEMA_signal_2651 ;
    wire new_AGEMA_signal_2652 ;
    wire new_AGEMA_signal_2653 ;
    wire new_AGEMA_signal_2654 ;
    wire new_AGEMA_signal_2655 ;
    wire new_AGEMA_signal_2656 ;
    wire new_AGEMA_signal_2657 ;
    wire new_AGEMA_signal_2658 ;
    wire new_AGEMA_signal_2659 ;
    wire new_AGEMA_signal_2660 ;
    wire new_AGEMA_signal_2661 ;
    wire new_AGEMA_signal_2662 ;
    wire new_AGEMA_signal_2663 ;
    wire new_AGEMA_signal_2664 ;
    wire new_AGEMA_signal_2665 ;
    wire new_AGEMA_signal_2666 ;
    wire new_AGEMA_signal_2667 ;
    wire new_AGEMA_signal_2668 ;
    wire new_AGEMA_signal_2669 ;
    wire new_AGEMA_signal_2670 ;
    wire new_AGEMA_signal_2671 ;
    wire new_AGEMA_signal_2672 ;
    wire new_AGEMA_signal_2673 ;
    wire new_AGEMA_signal_2674 ;
    wire new_AGEMA_signal_2675 ;
    wire new_AGEMA_signal_2676 ;
    wire new_AGEMA_signal_2677 ;
    wire new_AGEMA_signal_2678 ;
    wire new_AGEMA_signal_2679 ;
    wire new_AGEMA_signal_2680 ;
    wire new_AGEMA_signal_2681 ;
    wire new_AGEMA_signal_2682 ;
    wire new_AGEMA_signal_2683 ;
    wire new_AGEMA_signal_2684 ;
    wire new_AGEMA_signal_2685 ;
    wire new_AGEMA_signal_2686 ;
    wire new_AGEMA_signal_2687 ;
    wire new_AGEMA_signal_2688 ;
    wire new_AGEMA_signal_2689 ;
    wire new_AGEMA_signal_2690 ;
    wire new_AGEMA_signal_2691 ;
    wire new_AGEMA_signal_2692 ;
    wire new_AGEMA_signal_2693 ;
    wire new_AGEMA_signal_2694 ;
    wire new_AGEMA_signal_2695 ;
    wire new_AGEMA_signal_2696 ;
    wire new_AGEMA_signal_2697 ;
    wire new_AGEMA_signal_2698 ;
    wire new_AGEMA_signal_2699 ;
    wire new_AGEMA_signal_2700 ;
    wire new_AGEMA_signal_2701 ;
    wire new_AGEMA_signal_2702 ;
    wire new_AGEMA_signal_2703 ;
    wire new_AGEMA_signal_2704 ;
    wire new_AGEMA_signal_2705 ;
    wire new_AGEMA_signal_2706 ;
    wire new_AGEMA_signal_2707 ;
    wire new_AGEMA_signal_2708 ;
    wire new_AGEMA_signal_2709 ;
    wire new_AGEMA_signal_2710 ;
    wire new_AGEMA_signal_2711 ;
    wire new_AGEMA_signal_2712 ;
    wire new_AGEMA_signal_2713 ;
    wire new_AGEMA_signal_2714 ;
    wire new_AGEMA_signal_2715 ;
    wire new_AGEMA_signal_2716 ;
    wire new_AGEMA_signal_2717 ;
    wire new_AGEMA_signal_2718 ;
    wire new_AGEMA_signal_2719 ;
    wire new_AGEMA_signal_2720 ;
    wire new_AGEMA_signal_2721 ;
    wire new_AGEMA_signal_2722 ;
    wire new_AGEMA_signal_2723 ;
    wire new_AGEMA_signal_2724 ;
    wire new_AGEMA_signal_2725 ;
    wire new_AGEMA_signal_2726 ;
    wire new_AGEMA_signal_2727 ;
    wire new_AGEMA_signal_2728 ;
    wire new_AGEMA_signal_2729 ;
    wire new_AGEMA_signal_2730 ;
    wire new_AGEMA_signal_2731 ;
    wire new_AGEMA_signal_2732 ;
    wire new_AGEMA_signal_2733 ;
    wire new_AGEMA_signal_2734 ;
    wire new_AGEMA_signal_2735 ;
    wire new_AGEMA_signal_2736 ;
    wire new_AGEMA_signal_2737 ;
    wire new_AGEMA_signal_2738 ;
    wire new_AGEMA_signal_2739 ;
    wire new_AGEMA_signal_2740 ;
    wire new_AGEMA_signal_2741 ;
    wire new_AGEMA_signal_2742 ;
    wire new_AGEMA_signal_2743 ;
    wire new_AGEMA_signal_2744 ;
    wire new_AGEMA_signal_2745 ;
    wire new_AGEMA_signal_2746 ;
    wire new_AGEMA_signal_2747 ;
    wire new_AGEMA_signal_2748 ;
    wire new_AGEMA_signal_2749 ;
    wire new_AGEMA_signal_2750 ;
    wire new_AGEMA_signal_2751 ;
    wire new_AGEMA_signal_2752 ;
    wire new_AGEMA_signal_2753 ;
    wire new_AGEMA_signal_2754 ;
    wire new_AGEMA_signal_2755 ;
    wire new_AGEMA_signal_2756 ;
    wire new_AGEMA_signal_2757 ;
    wire new_AGEMA_signal_2758 ;
    wire new_AGEMA_signal_2759 ;
    wire new_AGEMA_signal_2760 ;
    wire new_AGEMA_signal_2761 ;
    wire new_AGEMA_signal_2762 ;
    wire new_AGEMA_signal_2766 ;
    wire new_AGEMA_signal_2767 ;
    wire new_AGEMA_signal_2768 ;
    wire new_AGEMA_signal_2769 ;
    wire new_AGEMA_signal_2770 ;
    wire new_AGEMA_signal_2771 ;
    wire new_AGEMA_signal_2772 ;
    wire new_AGEMA_signal_2773 ;
    wire new_AGEMA_signal_2774 ;
    wire new_AGEMA_signal_2775 ;
    wire new_AGEMA_signal_2776 ;
    wire new_AGEMA_signal_2777 ;
    wire new_AGEMA_signal_2778 ;
    wire new_AGEMA_signal_2779 ;
    wire new_AGEMA_signal_2780 ;
    wire new_AGEMA_signal_2781 ;
    wire new_AGEMA_signal_2782 ;
    wire new_AGEMA_signal_2783 ;
    wire new_AGEMA_signal_2784 ;
    wire new_AGEMA_signal_2785 ;
    wire new_AGEMA_signal_2786 ;
    wire new_AGEMA_signal_2787 ;
    wire new_AGEMA_signal_2788 ;
    wire new_AGEMA_signal_2789 ;
    wire new_AGEMA_signal_2790 ;
    wire new_AGEMA_signal_2791 ;
    wire new_AGEMA_signal_2792 ;
    wire new_AGEMA_signal_2793 ;
    wire new_AGEMA_signal_2794 ;
    wire new_AGEMA_signal_2795 ;
    wire new_AGEMA_signal_2796 ;
    wire new_AGEMA_signal_2797 ;
    wire new_AGEMA_signal_2798 ;
    wire new_AGEMA_signal_2799 ;
    wire new_AGEMA_signal_2800 ;
    wire new_AGEMA_signal_2801 ;
    wire new_AGEMA_signal_2802 ;
    wire new_AGEMA_signal_2803 ;
    wire new_AGEMA_signal_2804 ;
    wire new_AGEMA_signal_2805 ;
    wire new_AGEMA_signal_2806 ;
    wire new_AGEMA_signal_2807 ;
    wire new_AGEMA_signal_2808 ;
    wire new_AGEMA_signal_2809 ;
    wire new_AGEMA_signal_2810 ;
    wire new_AGEMA_signal_2811 ;
    wire new_AGEMA_signal_2812 ;
    wire new_AGEMA_signal_2813 ;
    wire new_AGEMA_signal_2814 ;
    wire new_AGEMA_signal_2815 ;
    wire new_AGEMA_signal_2816 ;
    wire new_AGEMA_signal_2817 ;
    wire new_AGEMA_signal_2818 ;
    wire new_AGEMA_signal_2819 ;
    wire new_AGEMA_signal_2820 ;
    wire new_AGEMA_signal_2821 ;
    wire new_AGEMA_signal_2822 ;
    wire new_AGEMA_signal_2823 ;
    wire new_AGEMA_signal_2824 ;
    wire new_AGEMA_signal_2825 ;
    wire new_AGEMA_signal_2826 ;
    wire new_AGEMA_signal_2827 ;
    wire new_AGEMA_signal_2828 ;
    wire new_AGEMA_signal_2829 ;
    wire new_AGEMA_signal_2830 ;
    wire new_AGEMA_signal_2831 ;
    wire new_AGEMA_signal_2832 ;
    wire new_AGEMA_signal_2833 ;
    wire new_AGEMA_signal_2834 ;
    wire new_AGEMA_signal_2835 ;
    wire new_AGEMA_signal_2836 ;
    wire new_AGEMA_signal_2837 ;
    wire new_AGEMA_signal_2838 ;
    wire new_AGEMA_signal_2839 ;
    wire new_AGEMA_signal_2840 ;
    wire new_AGEMA_signal_2841 ;
    wire new_AGEMA_signal_2842 ;
    wire new_AGEMA_signal_2843 ;
    wire new_AGEMA_signal_2844 ;
    wire new_AGEMA_signal_2845 ;
    wire new_AGEMA_signal_2846 ;
    wire new_AGEMA_signal_2847 ;
    wire new_AGEMA_signal_2848 ;
    wire new_AGEMA_signal_2849 ;
    wire new_AGEMA_signal_2850 ;
    wire new_AGEMA_signal_2851 ;
    wire new_AGEMA_signal_2852 ;
    wire new_AGEMA_signal_2853 ;
    wire new_AGEMA_signal_2854 ;
    wire new_AGEMA_signal_2855 ;
    wire new_AGEMA_signal_2856 ;
    wire new_AGEMA_signal_2857 ;
    wire new_AGEMA_signal_2858 ;
    wire new_AGEMA_signal_2859 ;
    wire new_AGEMA_signal_2860 ;
    wire new_AGEMA_signal_2861 ;
    wire new_AGEMA_signal_2862 ;
    wire new_AGEMA_signal_2863 ;
    wire new_AGEMA_signal_2864 ;
    wire new_AGEMA_signal_2865 ;
    wire new_AGEMA_signal_2866 ;
    wire new_AGEMA_signal_2867 ;
    wire new_AGEMA_signal_2868 ;
    wire new_AGEMA_signal_2869 ;
    wire new_AGEMA_signal_2870 ;
    wire new_AGEMA_signal_2871 ;
    wire new_AGEMA_signal_2872 ;
    wire new_AGEMA_signal_2873 ;
    wire new_AGEMA_signal_2874 ;
    wire new_AGEMA_signal_2875 ;
    wire new_AGEMA_signal_2876 ;
    wire new_AGEMA_signal_2877 ;
    wire new_AGEMA_signal_2878 ;
    wire new_AGEMA_signal_2879 ;
    wire new_AGEMA_signal_2880 ;
    wire new_AGEMA_signal_2881 ;
    wire new_AGEMA_signal_2882 ;
    wire new_AGEMA_signal_2883 ;
    wire new_AGEMA_signal_2884 ;
    wire new_AGEMA_signal_2885 ;
    wire new_AGEMA_signal_2886 ;
    wire new_AGEMA_signal_2887 ;
    wire new_AGEMA_signal_2888 ;
    wire new_AGEMA_signal_2889 ;
    wire new_AGEMA_signal_2890 ;
    wire new_AGEMA_signal_2891 ;
    wire new_AGEMA_signal_2892 ;
    wire new_AGEMA_signal_2893 ;
    wire new_AGEMA_signal_2894 ;
    wire new_AGEMA_signal_2895 ;
    wire new_AGEMA_signal_2896 ;
    wire new_AGEMA_signal_2897 ;
    wire new_AGEMA_signal_2898 ;
    wire new_AGEMA_signal_2899 ;
    wire new_AGEMA_signal_2900 ;
    wire new_AGEMA_signal_2901 ;
    wire new_AGEMA_signal_2902 ;
    wire new_AGEMA_signal_2903 ;
    wire new_AGEMA_signal_2904 ;
    wire new_AGEMA_signal_2905 ;
    wire new_AGEMA_signal_2906 ;
    wire new_AGEMA_signal_2907 ;
    wire new_AGEMA_signal_2908 ;
    wire new_AGEMA_signal_2909 ;
    wire new_AGEMA_signal_2910 ;
    wire new_AGEMA_signal_2911 ;
    wire new_AGEMA_signal_2912 ;
    wire new_AGEMA_signal_2913 ;
    wire new_AGEMA_signal_2914 ;
    wire new_AGEMA_signal_2915 ;
    wire new_AGEMA_signal_2916 ;
    wire new_AGEMA_signal_2917 ;
    wire new_AGEMA_signal_2918 ;
    wire new_AGEMA_signal_2919 ;
    wire new_AGEMA_signal_2920 ;
    wire new_AGEMA_signal_2921 ;
    wire new_AGEMA_signal_2922 ;
    wire new_AGEMA_signal_2923 ;
    wire new_AGEMA_signal_2924 ;
    wire new_AGEMA_signal_2925 ;
    wire new_AGEMA_signal_2926 ;
    wire new_AGEMA_signal_2927 ;
    wire new_AGEMA_signal_2928 ;
    wire new_AGEMA_signal_2929 ;
    wire new_AGEMA_signal_2930 ;
    wire new_AGEMA_signal_2931 ;
    wire new_AGEMA_signal_2932 ;
    wire new_AGEMA_signal_2933 ;
    wire new_AGEMA_signal_2934 ;
    wire new_AGEMA_signal_2935 ;
    wire new_AGEMA_signal_2936 ;
    wire new_AGEMA_signal_2937 ;
    wire new_AGEMA_signal_2938 ;
    wire new_AGEMA_signal_2939 ;
    wire new_AGEMA_signal_2940 ;
    wire new_AGEMA_signal_2941 ;
    wire new_AGEMA_signal_2942 ;
    wire new_AGEMA_signal_2943 ;
    wire new_AGEMA_signal_2944 ;
    wire new_AGEMA_signal_2945 ;
    wire new_AGEMA_signal_2946 ;
    wire new_AGEMA_signal_2947 ;
    wire new_AGEMA_signal_2948 ;
    wire new_AGEMA_signal_2949 ;
    wire new_AGEMA_signal_2950 ;
    wire new_AGEMA_signal_2951 ;
    wire new_AGEMA_signal_2952 ;
    wire new_AGEMA_signal_2953 ;
    wire new_AGEMA_signal_2954 ;
    wire new_AGEMA_signal_2955 ;
    wire new_AGEMA_signal_2956 ;
    wire new_AGEMA_signal_2957 ;
    wire new_AGEMA_signal_2958 ;
    wire new_AGEMA_signal_2959 ;
    wire new_AGEMA_signal_2960 ;
    wire new_AGEMA_signal_2961 ;
    wire new_AGEMA_signal_2962 ;
    wire new_AGEMA_signal_2963 ;
    wire new_AGEMA_signal_2964 ;
    wire new_AGEMA_signal_2965 ;
    wire new_AGEMA_signal_2966 ;
    wire new_AGEMA_signal_2967 ;
    wire new_AGEMA_signal_2968 ;
    wire new_AGEMA_signal_2969 ;
    wire new_AGEMA_signal_2970 ;
    wire new_AGEMA_signal_2971 ;
    wire new_AGEMA_signal_2972 ;
    wire new_AGEMA_signal_2973 ;
    wire new_AGEMA_signal_2974 ;
    wire new_AGEMA_signal_2975 ;
    wire new_AGEMA_signal_2976 ;
    wire new_AGEMA_signal_2977 ;
    wire new_AGEMA_signal_2978 ;
    wire new_AGEMA_signal_2979 ;
    wire new_AGEMA_signal_2980 ;
    wire new_AGEMA_signal_2981 ;
    wire new_AGEMA_signal_2982 ;
    wire new_AGEMA_signal_2983 ;
    wire new_AGEMA_signal_2984 ;
    wire new_AGEMA_signal_2985 ;
    wire new_AGEMA_signal_2986 ;
    wire new_AGEMA_signal_2987 ;
    wire new_AGEMA_signal_2988 ;
    wire new_AGEMA_signal_2989 ;
    wire new_AGEMA_signal_2990 ;
    wire new_AGEMA_signal_2991 ;
    wire new_AGEMA_signal_2992 ;
    wire new_AGEMA_signal_2993 ;
    wire new_AGEMA_signal_2995 ;
    wire new_AGEMA_signal_2996 ;
    wire new_AGEMA_signal_2997 ;
    wire new_AGEMA_signal_2998 ;
    wire new_AGEMA_signal_2999 ;
    wire new_AGEMA_signal_3000 ;
    wire new_AGEMA_signal_3001 ;
    wire new_AGEMA_signal_3002 ;
    wire new_AGEMA_signal_3003 ;
    wire new_AGEMA_signal_3005 ;
    wire new_AGEMA_signal_3009 ;
    wire new_AGEMA_signal_3010 ;
    wire new_AGEMA_signal_3011 ;
    wire new_AGEMA_signal_3012 ;
    wire new_AGEMA_signal_3013 ;
    wire new_AGEMA_signal_3014 ;
    wire new_AGEMA_signal_3015 ;
    wire new_AGEMA_signal_3016 ;
    wire new_AGEMA_signal_3017 ;
    wire new_AGEMA_signal_3018 ;
    wire new_AGEMA_signal_3019 ;
    wire new_AGEMA_signal_3020 ;
    wire new_AGEMA_signal_3021 ;
    wire new_AGEMA_signal_3022 ;
    wire new_AGEMA_signal_3023 ;
    wire new_AGEMA_signal_3027 ;
    wire new_AGEMA_signal_3028 ;
    wire new_AGEMA_signal_3029 ;
    wire new_AGEMA_signal_3033 ;
    wire new_AGEMA_signal_3034 ;
    wire new_AGEMA_signal_3035 ;
    wire new_AGEMA_signal_3036 ;
    wire new_AGEMA_signal_3037 ;
    wire new_AGEMA_signal_3038 ;
    wire new_AGEMA_signal_3039 ;
    wire new_AGEMA_signal_3040 ;
    wire new_AGEMA_signal_3041 ;
    wire new_AGEMA_signal_3042 ;
    wire new_AGEMA_signal_3043 ;
    wire new_AGEMA_signal_3044 ;
    wire new_AGEMA_signal_3045 ;
    wire new_AGEMA_signal_3046 ;
    wire new_AGEMA_signal_3047 ;
    wire new_AGEMA_signal_3048 ;
    wire new_AGEMA_signal_3049 ;
    wire new_AGEMA_signal_3050 ;
    wire new_AGEMA_signal_3051 ;
    wire new_AGEMA_signal_3052 ;
    wire new_AGEMA_signal_3053 ;
    wire new_AGEMA_signal_3054 ;
    wire new_AGEMA_signal_3055 ;
    wire new_AGEMA_signal_3056 ;
    wire new_AGEMA_signal_3057 ;
    wire new_AGEMA_signal_3058 ;
    wire new_AGEMA_signal_3059 ;
    wire new_AGEMA_signal_3060 ;
    wire new_AGEMA_signal_3061 ;
    wire new_AGEMA_signal_3062 ;
    wire new_AGEMA_signal_3063 ;
    wire new_AGEMA_signal_3064 ;
    wire new_AGEMA_signal_3065 ;
    wire new_AGEMA_signal_3066 ;
    wire new_AGEMA_signal_3067 ;
    wire new_AGEMA_signal_3068 ;
    wire new_AGEMA_signal_3069 ;
    wire new_AGEMA_signal_3070 ;
    wire new_AGEMA_signal_3071 ;
    wire new_AGEMA_signal_3072 ;
    wire new_AGEMA_signal_3073 ;
    wire new_AGEMA_signal_3074 ;
    wire new_AGEMA_signal_3075 ;
    wire new_AGEMA_signal_3076 ;
    wire new_AGEMA_signal_3077 ;
    wire new_AGEMA_signal_3081 ;
    wire new_AGEMA_signal_3082 ;
    wire new_AGEMA_signal_3083 ;
    wire new_AGEMA_signal_3084 ;
    wire new_AGEMA_signal_3085 ;
    wire new_AGEMA_signal_3086 ;
    wire new_AGEMA_signal_3087 ;
    wire new_AGEMA_signal_3088 ;
    wire new_AGEMA_signal_3089 ;
    wire new_AGEMA_signal_3090 ;
    wire new_AGEMA_signal_3091 ;
    wire new_AGEMA_signal_3092 ;
    wire new_AGEMA_signal_3093 ;
    wire new_AGEMA_signal_3094 ;
    wire new_AGEMA_signal_3095 ;
    wire new_AGEMA_signal_3096 ;
    wire new_AGEMA_signal_3097 ;
    wire new_AGEMA_signal_3098 ;
    wire new_AGEMA_signal_3099 ;
    wire new_AGEMA_signal_3100 ;
    wire new_AGEMA_signal_3101 ;
    wire new_AGEMA_signal_3102 ;
    wire new_AGEMA_signal_3103 ;
    wire new_AGEMA_signal_3104 ;
    wire new_AGEMA_signal_3105 ;
    wire new_AGEMA_signal_3106 ;
    wire new_AGEMA_signal_3107 ;
    wire new_AGEMA_signal_3108 ;
    wire new_AGEMA_signal_3109 ;
    wire new_AGEMA_signal_3110 ;
    wire new_AGEMA_signal_3111 ;
    wire new_AGEMA_signal_3112 ;
    wire new_AGEMA_signal_3113 ;
    wire new_AGEMA_signal_3114 ;
    wire new_AGEMA_signal_3115 ;
    wire new_AGEMA_signal_3116 ;
    wire new_AGEMA_signal_3117 ;
    wire new_AGEMA_signal_3118 ;
    wire new_AGEMA_signal_3119 ;
    wire new_AGEMA_signal_3120 ;
    wire new_AGEMA_signal_3121 ;
    wire new_AGEMA_signal_3122 ;
    wire new_AGEMA_signal_3123 ;
    wire new_AGEMA_signal_3124 ;
    wire new_AGEMA_signal_3125 ;
    wire new_AGEMA_signal_3126 ;
    wire new_AGEMA_signal_3127 ;
    wire new_AGEMA_signal_3128 ;
    wire new_AGEMA_signal_3129 ;
    wire new_AGEMA_signal_3130 ;
    wire new_AGEMA_signal_3131 ;
    wire new_AGEMA_signal_3132 ;
    wire new_AGEMA_signal_3133 ;
    wire new_AGEMA_signal_3134 ;
    wire new_AGEMA_signal_3135 ;
    wire new_AGEMA_signal_3136 ;
    wire new_AGEMA_signal_3137 ;
    wire new_AGEMA_signal_3138 ;
    wire new_AGEMA_signal_3139 ;
    wire new_AGEMA_signal_3140 ;
    wire new_AGEMA_signal_3141 ;
    wire new_AGEMA_signal_3142 ;
    wire new_AGEMA_signal_3143 ;
    wire new_AGEMA_signal_3144 ;
    wire new_AGEMA_signal_3145 ;
    wire new_AGEMA_signal_3146 ;
    wire new_AGEMA_signal_3147 ;
    wire new_AGEMA_signal_3148 ;
    wire new_AGEMA_signal_3149 ;
    wire new_AGEMA_signal_3153 ;
    wire new_AGEMA_signal_3154 ;
    wire new_AGEMA_signal_3155 ;
    wire new_AGEMA_signal_3156 ;
    wire new_AGEMA_signal_3157 ;
    wire new_AGEMA_signal_3158 ;
    wire new_AGEMA_signal_3159 ;
    wire new_AGEMA_signal_3160 ;
    wire new_AGEMA_signal_3161 ;
    wire new_AGEMA_signal_3162 ;
    wire new_AGEMA_signal_3163 ;
    wire new_AGEMA_signal_3164 ;
    wire new_AGEMA_signal_3165 ;
    wire new_AGEMA_signal_3166 ;
    wire new_AGEMA_signal_3167 ;
    wire new_AGEMA_signal_3168 ;
    wire new_AGEMA_signal_3169 ;
    wire new_AGEMA_signal_3170 ;
    wire new_AGEMA_signal_3171 ;
    wire new_AGEMA_signal_3172 ;
    wire new_AGEMA_signal_3173 ;
    wire new_AGEMA_signal_3174 ;
    wire new_AGEMA_signal_3175 ;
    wire new_AGEMA_signal_3176 ;
    wire new_AGEMA_signal_3177 ;
    wire new_AGEMA_signal_3178 ;
    wire new_AGEMA_signal_3179 ;
    wire new_AGEMA_signal_3180 ;
    wire new_AGEMA_signal_3181 ;
    wire new_AGEMA_signal_3182 ;
    wire new_AGEMA_signal_3183 ;
    wire new_AGEMA_signal_3184 ;
    wire new_AGEMA_signal_3185 ;
    wire new_AGEMA_signal_3186 ;
    wire new_AGEMA_signal_3187 ;
    wire new_AGEMA_signal_3188 ;
    wire new_AGEMA_signal_3189 ;
    wire new_AGEMA_signal_3190 ;
    wire new_AGEMA_signal_3191 ;
    wire new_AGEMA_signal_3192 ;
    wire new_AGEMA_signal_3193 ;
    wire new_AGEMA_signal_3194 ;
    wire new_AGEMA_signal_3195 ;
    wire new_AGEMA_signal_3196 ;
    wire new_AGEMA_signal_3197 ;
    wire new_AGEMA_signal_3198 ;
    wire new_AGEMA_signal_3199 ;
    wire new_AGEMA_signal_3200 ;
    wire new_AGEMA_signal_3201 ;
    wire new_AGEMA_signal_3202 ;
    wire new_AGEMA_signal_3203 ;
    wire new_AGEMA_signal_3204 ;
    wire new_AGEMA_signal_3205 ;
    wire new_AGEMA_signal_3206 ;
    wire new_AGEMA_signal_3207 ;
    wire new_AGEMA_signal_3208 ;
    wire new_AGEMA_signal_3209 ;
    wire new_AGEMA_signal_3210 ;
    wire new_AGEMA_signal_3211 ;
    wire new_AGEMA_signal_3212 ;
    wire new_AGEMA_signal_3213 ;
    wire new_AGEMA_signal_3214 ;
    wire new_AGEMA_signal_3215 ;
    wire new_AGEMA_signal_3216 ;
    wire new_AGEMA_signal_3217 ;
    wire new_AGEMA_signal_3218 ;
    wire new_AGEMA_signal_3219 ;
    wire new_AGEMA_signal_3220 ;
    wire new_AGEMA_signal_3221 ;
    wire new_AGEMA_signal_3222 ;
    wire new_AGEMA_signal_3223 ;
    wire new_AGEMA_signal_3224 ;
    wire new_AGEMA_signal_3225 ;
    wire new_AGEMA_signal_3226 ;
    wire new_AGEMA_signal_3227 ;
    wire new_AGEMA_signal_3228 ;
    wire new_AGEMA_signal_3229 ;
    wire new_AGEMA_signal_3230 ;
    wire new_AGEMA_signal_3231 ;
    wire new_AGEMA_signal_3232 ;
    wire new_AGEMA_signal_3233 ;
    wire new_AGEMA_signal_3234 ;
    wire new_AGEMA_signal_3235 ;
    wire new_AGEMA_signal_3236 ;
    wire new_AGEMA_signal_3237 ;
    wire new_AGEMA_signal_3238 ;
    wire new_AGEMA_signal_3239 ;
    wire new_AGEMA_signal_3240 ;
    wire new_AGEMA_signal_3241 ;
    wire new_AGEMA_signal_3242 ;
    wire new_AGEMA_signal_3243 ;
    wire new_AGEMA_signal_3244 ;
    wire new_AGEMA_signal_3245 ;
    wire new_AGEMA_signal_3246 ;
    wire new_AGEMA_signal_3247 ;
    wire new_AGEMA_signal_3248 ;
    wire new_AGEMA_signal_3249 ;
    wire new_AGEMA_signal_3250 ;
    wire new_AGEMA_signal_3251 ;
    wire new_AGEMA_signal_3252 ;
    wire new_AGEMA_signal_3253 ;
    wire new_AGEMA_signal_3254 ;
    wire new_AGEMA_signal_3255 ;
    wire new_AGEMA_signal_3256 ;
    wire new_AGEMA_signal_3257 ;
    wire new_AGEMA_signal_3258 ;
    wire new_AGEMA_signal_3259 ;
    wire new_AGEMA_signal_3260 ;
    wire new_AGEMA_signal_3261 ;
    wire new_AGEMA_signal_3262 ;
    wire new_AGEMA_signal_3263 ;
    wire new_AGEMA_signal_3264 ;
    wire new_AGEMA_signal_3265 ;
    wire new_AGEMA_signal_3266 ;
    wire new_AGEMA_signal_3267 ;
    wire new_AGEMA_signal_3268 ;
    wire new_AGEMA_signal_3269 ;
    wire new_AGEMA_signal_3270 ;
    wire new_AGEMA_signal_3271 ;
    wire new_AGEMA_signal_3272 ;
    wire new_AGEMA_signal_3273 ;
    wire new_AGEMA_signal_3274 ;
    wire new_AGEMA_signal_3275 ;
    wire new_AGEMA_signal_3276 ;
    wire new_AGEMA_signal_3277 ;
    wire new_AGEMA_signal_3278 ;
    wire new_AGEMA_signal_3279 ;
    wire new_AGEMA_signal_3280 ;
    wire new_AGEMA_signal_3281 ;
    wire new_AGEMA_signal_3282 ;
    wire new_AGEMA_signal_3283 ;
    wire new_AGEMA_signal_3284 ;
    wire new_AGEMA_signal_3285 ;
    wire new_AGEMA_signal_3286 ;
    wire new_AGEMA_signal_3287 ;
    wire new_AGEMA_signal_3288 ;
    wire new_AGEMA_signal_3289 ;
    wire new_AGEMA_signal_3290 ;
    wire new_AGEMA_signal_3291 ;
    wire new_AGEMA_signal_3292 ;
    wire new_AGEMA_signal_3293 ;
    wire new_AGEMA_signal_3294 ;
    wire new_AGEMA_signal_3295 ;
    wire new_AGEMA_signal_3296 ;
    wire new_AGEMA_signal_3297 ;
    wire new_AGEMA_signal_3298 ;
    wire new_AGEMA_signal_3299 ;
    wire new_AGEMA_signal_3300 ;
    wire new_AGEMA_signal_3301 ;
    wire new_AGEMA_signal_3302 ;
    wire new_AGEMA_signal_3303 ;
    wire new_AGEMA_signal_3304 ;
    wire new_AGEMA_signal_3305 ;
    wire new_AGEMA_signal_3306 ;
    wire new_AGEMA_signal_3307 ;
    wire new_AGEMA_signal_3308 ;
    wire new_AGEMA_signal_3309 ;
    wire new_AGEMA_signal_3310 ;
    wire new_AGEMA_signal_3311 ;
    wire new_AGEMA_signal_3312 ;
    wire new_AGEMA_signal_3313 ;
    wire new_AGEMA_signal_3314 ;
    wire new_AGEMA_signal_3315 ;
    wire new_AGEMA_signal_3316 ;
    wire new_AGEMA_signal_3317 ;
    wire new_AGEMA_signal_3318 ;
    wire new_AGEMA_signal_3319 ;
    wire new_AGEMA_signal_3320 ;
    wire new_AGEMA_signal_3321 ;
    wire new_AGEMA_signal_3322 ;
    wire new_AGEMA_signal_3323 ;
    wire new_AGEMA_signal_3324 ;
    wire new_AGEMA_signal_3325 ;
    wire new_AGEMA_signal_3326 ;
    wire new_AGEMA_signal_3327 ;
    wire new_AGEMA_signal_3328 ;
    wire new_AGEMA_signal_3329 ;
    wire new_AGEMA_signal_3330 ;
    wire new_AGEMA_signal_3331 ;
    wire new_AGEMA_signal_3332 ;
    wire new_AGEMA_signal_3333 ;
    wire new_AGEMA_signal_3334 ;
    wire new_AGEMA_signal_3335 ;
    wire new_AGEMA_signal_3336 ;
    wire new_AGEMA_signal_3337 ;
    wire new_AGEMA_signal_3338 ;
    wire new_AGEMA_signal_3339 ;
    wire new_AGEMA_signal_3340 ;
    wire new_AGEMA_signal_3341 ;
    wire new_AGEMA_signal_3342 ;
    wire new_AGEMA_signal_3343 ;
    wire new_AGEMA_signal_3344 ;
    wire new_AGEMA_signal_3345 ;
    wire new_AGEMA_signal_3346 ;
    wire new_AGEMA_signal_3347 ;
    wire new_AGEMA_signal_3348 ;
    wire new_AGEMA_signal_3349 ;
    wire new_AGEMA_signal_3350 ;
    wire new_AGEMA_signal_3351 ;
    wire new_AGEMA_signal_3352 ;
    wire new_AGEMA_signal_3353 ;
    wire new_AGEMA_signal_3354 ;
    wire new_AGEMA_signal_3355 ;
    wire new_AGEMA_signal_3356 ;
    wire new_AGEMA_signal_3357 ;
    wire new_AGEMA_signal_3358 ;
    wire new_AGEMA_signal_3359 ;
    wire new_AGEMA_signal_3360 ;
    wire new_AGEMA_signal_3361 ;
    wire new_AGEMA_signal_3362 ;
    wire new_AGEMA_signal_3363 ;
    wire new_AGEMA_signal_3364 ;
    wire new_AGEMA_signal_3365 ;
    wire new_AGEMA_signal_3366 ;
    wire new_AGEMA_signal_3367 ;
    wire new_AGEMA_signal_3368 ;
    wire new_AGEMA_signal_3369 ;
    wire new_AGEMA_signal_3370 ;
    wire new_AGEMA_signal_3371 ;
    wire new_AGEMA_signal_3372 ;
    wire new_AGEMA_signal_3373 ;
    wire new_AGEMA_signal_3374 ;
    wire new_AGEMA_signal_3375 ;
    wire new_AGEMA_signal_3376 ;
    wire new_AGEMA_signal_3377 ;
    wire new_AGEMA_signal_3378 ;
    wire new_AGEMA_signal_3379 ;
    wire new_AGEMA_signal_3380 ;
    wire new_AGEMA_signal_3381 ;
    wire new_AGEMA_signal_3382 ;
    wire new_AGEMA_signal_3383 ;
    wire new_AGEMA_signal_3384 ;
    wire new_AGEMA_signal_3385 ;
    wire new_AGEMA_signal_3386 ;
    wire new_AGEMA_signal_3387 ;
    wire new_AGEMA_signal_3388 ;
    wire new_AGEMA_signal_3389 ;
    wire new_AGEMA_signal_3390 ;
    wire new_AGEMA_signal_3391 ;
    wire new_AGEMA_signal_3392 ;
    wire new_AGEMA_signal_3393 ;
    wire new_AGEMA_signal_3394 ;
    wire new_AGEMA_signal_3395 ;
    wire new_AGEMA_signal_3396 ;
    wire new_AGEMA_signal_3397 ;
    wire new_AGEMA_signal_3398 ;
    wire new_AGEMA_signal_3399 ;
    wire new_AGEMA_signal_3400 ;
    wire new_AGEMA_signal_3401 ;
    wire new_AGEMA_signal_3402 ;
    wire new_AGEMA_signal_3403 ;
    wire new_AGEMA_signal_3404 ;
    wire new_AGEMA_signal_3405 ;
    wire new_AGEMA_signal_3406 ;
    wire new_AGEMA_signal_3407 ;
    wire new_AGEMA_signal_3408 ;
    wire new_AGEMA_signal_3409 ;
    wire new_AGEMA_signal_3410 ;
    wire new_AGEMA_signal_3411 ;
    wire new_AGEMA_signal_3412 ;
    wire new_AGEMA_signal_3413 ;
    wire new_AGEMA_signal_3414 ;
    wire new_AGEMA_signal_3415 ;
    wire new_AGEMA_signal_3416 ;
    wire new_AGEMA_signal_3417 ;
    wire new_AGEMA_signal_3418 ;
    wire new_AGEMA_signal_3419 ;
    wire new_AGEMA_signal_3420 ;
    wire new_AGEMA_signal_3421 ;
    wire new_AGEMA_signal_3422 ;
    wire new_AGEMA_signal_3423 ;
    wire new_AGEMA_signal_3424 ;
    wire new_AGEMA_signal_3425 ;
    wire new_AGEMA_signal_3426 ;
    wire new_AGEMA_signal_3427 ;
    wire new_AGEMA_signal_3428 ;
    wire new_AGEMA_signal_3429 ;
    wire new_AGEMA_signal_3430 ;
    wire new_AGEMA_signal_3431 ;
    wire new_AGEMA_signal_3432 ;
    wire new_AGEMA_signal_3433 ;
    wire new_AGEMA_signal_3434 ;
    wire new_AGEMA_signal_3435 ;
    wire new_AGEMA_signal_3436 ;
    wire new_AGEMA_signal_3437 ;
    wire new_AGEMA_signal_3438 ;
    wire new_AGEMA_signal_3439 ;
    wire new_AGEMA_signal_3440 ;
    wire new_AGEMA_signal_3441 ;
    wire new_AGEMA_signal_3442 ;
    wire new_AGEMA_signal_3443 ;
    wire new_AGEMA_signal_3444 ;
    wire new_AGEMA_signal_3445 ;
    wire new_AGEMA_signal_3446 ;
    wire new_AGEMA_signal_3447 ;
    wire new_AGEMA_signal_3448 ;
    wire new_AGEMA_signal_3449 ;
    wire new_AGEMA_signal_3450 ;
    wire new_AGEMA_signal_3451 ;
    wire new_AGEMA_signal_3452 ;
    wire new_AGEMA_signal_3453 ;
    wire new_AGEMA_signal_3454 ;
    wire new_AGEMA_signal_3455 ;
    wire new_AGEMA_signal_3456 ;
    wire new_AGEMA_signal_3457 ;
    wire new_AGEMA_signal_3458 ;
    wire new_AGEMA_signal_3459 ;
    wire new_AGEMA_signal_3460 ;
    wire new_AGEMA_signal_3461 ;
    wire new_AGEMA_signal_3462 ;
    wire new_AGEMA_signal_3463 ;
    wire new_AGEMA_signal_3464 ;
    wire new_AGEMA_signal_3465 ;
    wire new_AGEMA_signal_3466 ;
    wire new_AGEMA_signal_3467 ;
    wire new_AGEMA_signal_3468 ;
    wire new_AGEMA_signal_3469 ;
    wire new_AGEMA_signal_3470 ;
    wire new_AGEMA_signal_3471 ;
    wire new_AGEMA_signal_3472 ;
    wire new_AGEMA_signal_3473 ;
    wire new_AGEMA_signal_3474 ;
    wire new_AGEMA_signal_3475 ;
    wire new_AGEMA_signal_3476 ;
    wire new_AGEMA_signal_3477 ;
    wire new_AGEMA_signal_3478 ;
    wire new_AGEMA_signal_3479 ;
    wire new_AGEMA_signal_3480 ;
    wire new_AGEMA_signal_3481 ;
    wire new_AGEMA_signal_3482 ;
    wire new_AGEMA_signal_3483 ;
    wire new_AGEMA_signal_3484 ;
    wire new_AGEMA_signal_3485 ;
    wire new_AGEMA_signal_3486 ;
    wire new_AGEMA_signal_3487 ;
    wire new_AGEMA_signal_3488 ;
    wire new_AGEMA_signal_3489 ;
    wire new_AGEMA_signal_3490 ;
    wire new_AGEMA_signal_3491 ;
    wire new_AGEMA_signal_3492 ;
    wire new_AGEMA_signal_3493 ;
    wire new_AGEMA_signal_3494 ;
    wire new_AGEMA_signal_3495 ;
    wire new_AGEMA_signal_3496 ;
    wire new_AGEMA_signal_3497 ;
    wire new_AGEMA_signal_3498 ;
    wire new_AGEMA_signal_3499 ;
    wire new_AGEMA_signal_3500 ;
    wire new_AGEMA_signal_3501 ;
    wire new_AGEMA_signal_3502 ;
    wire new_AGEMA_signal_3503 ;
    wire new_AGEMA_signal_3504 ;
    wire new_AGEMA_signal_3505 ;
    wire new_AGEMA_signal_3506 ;
    wire new_AGEMA_signal_3507 ;
    wire new_AGEMA_signal_3508 ;
    wire new_AGEMA_signal_3509 ;
    wire new_AGEMA_signal_3510 ;
    wire new_AGEMA_signal_3511 ;
    wire new_AGEMA_signal_3512 ;
    wire new_AGEMA_signal_3513 ;
    wire new_AGEMA_signal_3514 ;
    wire new_AGEMA_signal_3515 ;
    wire new_AGEMA_signal_3516 ;
    wire new_AGEMA_signal_3517 ;
    wire new_AGEMA_signal_3518 ;
    wire new_AGEMA_signal_3519 ;
    wire new_AGEMA_signal_3520 ;
    wire new_AGEMA_signal_3521 ;
    wire new_AGEMA_signal_3522 ;
    wire new_AGEMA_signal_3523 ;
    wire new_AGEMA_signal_3524 ;
    wire new_AGEMA_signal_3525 ;
    wire new_AGEMA_signal_3526 ;
    wire new_AGEMA_signal_3527 ;
    wire new_AGEMA_signal_3528 ;
    wire new_AGEMA_signal_3529 ;
    wire new_AGEMA_signal_3530 ;
    wire new_AGEMA_signal_3531 ;
    wire new_AGEMA_signal_3532 ;
    wire new_AGEMA_signal_3533 ;
    wire new_AGEMA_signal_3534 ;
    wire new_AGEMA_signal_3535 ;
    wire new_AGEMA_signal_3536 ;
    wire new_AGEMA_signal_3537 ;
    wire new_AGEMA_signal_3538 ;
    wire new_AGEMA_signal_3539 ;
    wire new_AGEMA_signal_3540 ;
    wire new_AGEMA_signal_3541 ;
    wire new_AGEMA_signal_3542 ;
    wire new_AGEMA_signal_3543 ;
    wire new_AGEMA_signal_3544 ;
    wire new_AGEMA_signal_3545 ;
    wire new_AGEMA_signal_3546 ;
    wire new_AGEMA_signal_3547 ;
    wire new_AGEMA_signal_3548 ;
    wire new_AGEMA_signal_3549 ;
    wire new_AGEMA_signal_3550 ;
    wire new_AGEMA_signal_3551 ;
    wire new_AGEMA_signal_3552 ;
    wire new_AGEMA_signal_3553 ;
    wire new_AGEMA_signal_3554 ;
    wire new_AGEMA_signal_3555 ;
    wire new_AGEMA_signal_3556 ;
    wire new_AGEMA_signal_3557 ;
    wire new_AGEMA_signal_3558 ;
    wire new_AGEMA_signal_3559 ;
    wire new_AGEMA_signal_3560 ;
    wire new_AGEMA_signal_3561 ;
    wire new_AGEMA_signal_3562 ;
    wire new_AGEMA_signal_3563 ;
    wire new_AGEMA_signal_3564 ;
    wire new_AGEMA_signal_3565 ;
    wire new_AGEMA_signal_3566 ;
    wire new_AGEMA_signal_3567 ;
    wire new_AGEMA_signal_3568 ;
    wire new_AGEMA_signal_3569 ;
    wire new_AGEMA_signal_3570 ;
    wire new_AGEMA_signal_3571 ;
    wire new_AGEMA_signal_3572 ;
    wire new_AGEMA_signal_3573 ;
    wire new_AGEMA_signal_3574 ;
    wire new_AGEMA_signal_3575 ;
    wire new_AGEMA_signal_3576 ;
    wire new_AGEMA_signal_3577 ;
    wire new_AGEMA_signal_3578 ;
    wire new_AGEMA_signal_3579 ;
    wire new_AGEMA_signal_3580 ;
    wire new_AGEMA_signal_3581 ;
    wire new_AGEMA_signal_3582 ;
    wire new_AGEMA_signal_3583 ;
    wire new_AGEMA_signal_3584 ;
    wire new_AGEMA_signal_3585 ;
    wire new_AGEMA_signal_3586 ;
    wire new_AGEMA_signal_3587 ;
    wire new_AGEMA_signal_3588 ;
    wire new_AGEMA_signal_3589 ;
    wire new_AGEMA_signal_3590 ;
    wire new_AGEMA_signal_3591 ;
    wire new_AGEMA_signal_3592 ;
    wire new_AGEMA_signal_3593 ;
    wire new_AGEMA_signal_3594 ;
    wire new_AGEMA_signal_3595 ;
    wire new_AGEMA_signal_3596 ;
    wire new_AGEMA_signal_3597 ;
    wire new_AGEMA_signal_3598 ;
    wire new_AGEMA_signal_3599 ;
    wire new_AGEMA_signal_3600 ;
    wire new_AGEMA_signal_3601 ;
    wire new_AGEMA_signal_3602 ;
    wire new_AGEMA_signal_3603 ;
    wire new_AGEMA_signal_3604 ;
    wire new_AGEMA_signal_3605 ;
    wire new_AGEMA_signal_3606 ;
    wire new_AGEMA_signal_3607 ;
    wire new_AGEMA_signal_3608 ;
    wire new_AGEMA_signal_3609 ;
    wire new_AGEMA_signal_3610 ;
    wire new_AGEMA_signal_3611 ;
    wire new_AGEMA_signal_3612 ;
    wire new_AGEMA_signal_3613 ;
    wire new_AGEMA_signal_3614 ;
    wire new_AGEMA_signal_3615 ;
    wire new_AGEMA_signal_3616 ;
    wire new_AGEMA_signal_3617 ;
    wire new_AGEMA_signal_3618 ;
    wire new_AGEMA_signal_3619 ;
    wire new_AGEMA_signal_3620 ;
    wire new_AGEMA_signal_3621 ;
    wire new_AGEMA_signal_3622 ;
    wire new_AGEMA_signal_3623 ;
    wire new_AGEMA_signal_3624 ;
    wire new_AGEMA_signal_3625 ;
    wire new_AGEMA_signal_3626 ;
    wire new_AGEMA_signal_3627 ;
    wire new_AGEMA_signal_3628 ;
    wire new_AGEMA_signal_3629 ;
    wire new_AGEMA_signal_3630 ;
    wire new_AGEMA_signal_3631 ;
    wire new_AGEMA_signal_3632 ;
    wire new_AGEMA_signal_3633 ;
    wire new_AGEMA_signal_3634 ;
    wire new_AGEMA_signal_3635 ;
    wire new_AGEMA_signal_3636 ;
    wire new_AGEMA_signal_3637 ;
    wire new_AGEMA_signal_3638 ;
    wire new_AGEMA_signal_3639 ;
    wire new_AGEMA_signal_3640 ;
    wire new_AGEMA_signal_3641 ;
    wire new_AGEMA_signal_3642 ;
    wire new_AGEMA_signal_3643 ;
    wire new_AGEMA_signal_3644 ;
    wire new_AGEMA_signal_3645 ;
    wire new_AGEMA_signal_3646 ;
    wire new_AGEMA_signal_3647 ;
    wire new_AGEMA_signal_3648 ;
    wire new_AGEMA_signal_3649 ;
    wire new_AGEMA_signal_3650 ;
    wire new_AGEMA_signal_3651 ;
    wire new_AGEMA_signal_3652 ;
    wire new_AGEMA_signal_3653 ;
    wire new_AGEMA_signal_3654 ;
    wire new_AGEMA_signal_3655 ;
    wire new_AGEMA_signal_3656 ;
    wire new_AGEMA_signal_3657 ;
    wire new_AGEMA_signal_3658 ;
    wire new_AGEMA_signal_3659 ;
    wire new_AGEMA_signal_3660 ;
    wire new_AGEMA_signal_3661 ;
    wire new_AGEMA_signal_3662 ;
    wire new_AGEMA_signal_3663 ;
    wire new_AGEMA_signal_3664 ;
    wire new_AGEMA_signal_3665 ;
    wire new_AGEMA_signal_3666 ;
    wire new_AGEMA_signal_3667 ;
    wire new_AGEMA_signal_3668 ;
    wire new_AGEMA_signal_3669 ;
    wire new_AGEMA_signal_3670 ;
    wire new_AGEMA_signal_3671 ;
    wire new_AGEMA_signal_3672 ;
    wire new_AGEMA_signal_3673 ;
    wire new_AGEMA_signal_3674 ;
    wire new_AGEMA_signal_3675 ;
    wire new_AGEMA_signal_3676 ;
    wire new_AGEMA_signal_3677 ;
    wire new_AGEMA_signal_3678 ;
    wire new_AGEMA_signal_3679 ;
    wire new_AGEMA_signal_3680 ;
    wire new_AGEMA_signal_3681 ;
    wire new_AGEMA_signal_3682 ;
    wire new_AGEMA_signal_3683 ;
    wire new_AGEMA_signal_3684 ;
    wire new_AGEMA_signal_3685 ;
    wire new_AGEMA_signal_3686 ;
    wire new_AGEMA_signal_3687 ;
    wire new_AGEMA_signal_3688 ;
    wire new_AGEMA_signal_3689 ;
    wire new_AGEMA_signal_3690 ;
    wire new_AGEMA_signal_3691 ;
    wire new_AGEMA_signal_3692 ;
    wire new_AGEMA_signal_3693 ;
    wire new_AGEMA_signal_3694 ;
    wire new_AGEMA_signal_3695 ;
    wire new_AGEMA_signal_3696 ;
    wire new_AGEMA_signal_3697 ;
    wire new_AGEMA_signal_3698 ;
    wire new_AGEMA_signal_3699 ;
    wire new_AGEMA_signal_3700 ;
    wire new_AGEMA_signal_3701 ;
    wire new_AGEMA_signal_3702 ;
    wire new_AGEMA_signal_3703 ;
    wire new_AGEMA_signal_3704 ;
    wire new_AGEMA_signal_3705 ;
    wire new_AGEMA_signal_3706 ;
    wire new_AGEMA_signal_3707 ;
    wire new_AGEMA_signal_3708 ;
    wire new_AGEMA_signal_3709 ;
    wire new_AGEMA_signal_3710 ;
    wire new_AGEMA_signal_3711 ;
    wire new_AGEMA_signal_3712 ;
    wire new_AGEMA_signal_3713 ;
    wire new_AGEMA_signal_3714 ;
    wire new_AGEMA_signal_3715 ;
    wire new_AGEMA_signal_3716 ;
    wire new_AGEMA_signal_3717 ;
    wire new_AGEMA_signal_3718 ;
    wire new_AGEMA_signal_3719 ;
    wire new_AGEMA_signal_3720 ;
    wire new_AGEMA_signal_3721 ;
    wire new_AGEMA_signal_3722 ;
    wire new_AGEMA_signal_3723 ;
    wire new_AGEMA_signal_3724 ;
    wire new_AGEMA_signal_3725 ;
    wire new_AGEMA_signal_3726 ;
    wire new_AGEMA_signal_3727 ;
    wire new_AGEMA_signal_3728 ;
    wire new_AGEMA_signal_3729 ;
    wire new_AGEMA_signal_3730 ;
    wire new_AGEMA_signal_3731 ;
    wire new_AGEMA_signal_3732 ;
    wire new_AGEMA_signal_3733 ;
    wire new_AGEMA_signal_3734 ;
    wire new_AGEMA_signal_3735 ;
    wire new_AGEMA_signal_3736 ;
    wire new_AGEMA_signal_3737 ;
    wire new_AGEMA_signal_3738 ;
    wire new_AGEMA_signal_3739 ;
    wire new_AGEMA_signal_3740 ;
    wire new_AGEMA_signal_3741 ;
    wire new_AGEMA_signal_3742 ;
    wire new_AGEMA_signal_3743 ;
    wire new_AGEMA_signal_3744 ;
    wire new_AGEMA_signal_3745 ;
    wire new_AGEMA_signal_3746 ;
    wire new_AGEMA_signal_3747 ;
    wire new_AGEMA_signal_3748 ;
    wire new_AGEMA_signal_3749 ;
    wire new_AGEMA_signal_3750 ;
    wire new_AGEMA_signal_3751 ;
    wire new_AGEMA_signal_3752 ;
    wire new_AGEMA_signal_3753 ;
    wire new_AGEMA_signal_3754 ;
    wire new_AGEMA_signal_3755 ;
    wire new_AGEMA_signal_3756 ;
    wire new_AGEMA_signal_3757 ;
    wire new_AGEMA_signal_3758 ;
    wire new_AGEMA_signal_3759 ;
    wire new_AGEMA_signal_3760 ;
    wire new_AGEMA_signal_3761 ;
    wire new_AGEMA_signal_3762 ;
    wire new_AGEMA_signal_3763 ;
    wire new_AGEMA_signal_3764 ;
    wire new_AGEMA_signal_3765 ;
    wire new_AGEMA_signal_3766 ;
    wire new_AGEMA_signal_3767 ;
    wire new_AGEMA_signal_3768 ;
    wire new_AGEMA_signal_3769 ;
    wire new_AGEMA_signal_3770 ;
    wire new_AGEMA_signal_3771 ;
    wire new_AGEMA_signal_3772 ;
    wire new_AGEMA_signal_3773 ;
    wire new_AGEMA_signal_3774 ;
    wire new_AGEMA_signal_3775 ;
    wire new_AGEMA_signal_3776 ;
    wire new_AGEMA_signal_3777 ;
    wire new_AGEMA_signal_3778 ;
    wire new_AGEMA_signal_3779 ;
    wire new_AGEMA_signal_3780 ;
    wire new_AGEMA_signal_3781 ;
    wire new_AGEMA_signal_3782 ;
    wire new_AGEMA_signal_3783 ;
    wire new_AGEMA_signal_3784 ;
    wire new_AGEMA_signal_3785 ;
    wire new_AGEMA_signal_3786 ;
    wire new_AGEMA_signal_3787 ;
    wire new_AGEMA_signal_3788 ;
    wire new_AGEMA_signal_3789 ;
    wire new_AGEMA_signal_3790 ;
    wire new_AGEMA_signal_3791 ;
    wire new_AGEMA_signal_3792 ;
    wire new_AGEMA_signal_3793 ;
    wire new_AGEMA_signal_3794 ;
    wire new_AGEMA_signal_3795 ;
    wire new_AGEMA_signal_3796 ;
    wire new_AGEMA_signal_3797 ;
    wire new_AGEMA_signal_3798 ;
    wire new_AGEMA_signal_3799 ;
    wire new_AGEMA_signal_3800 ;
    wire new_AGEMA_signal_3801 ;
    wire new_AGEMA_signal_3802 ;
    wire new_AGEMA_signal_3803 ;
    wire new_AGEMA_signal_3804 ;
    wire new_AGEMA_signal_3805 ;
    wire new_AGEMA_signal_3806 ;
    wire new_AGEMA_signal_3807 ;
    wire new_AGEMA_signal_3808 ;
    wire new_AGEMA_signal_3809 ;
    wire new_AGEMA_signal_3810 ;
    wire new_AGEMA_signal_3811 ;
    wire new_AGEMA_signal_3812 ;
    wire new_AGEMA_signal_3813 ;
    wire new_AGEMA_signal_3814 ;
    wire new_AGEMA_signal_3815 ;
    wire new_AGEMA_signal_3816 ;
    wire new_AGEMA_signal_3817 ;
    wire new_AGEMA_signal_3818 ;
    wire new_AGEMA_signal_3819 ;
    wire new_AGEMA_signal_3820 ;
    wire new_AGEMA_signal_3821 ;
    wire new_AGEMA_signal_3822 ;
    wire new_AGEMA_signal_3823 ;
    wire new_AGEMA_signal_3824 ;
    wire new_AGEMA_signal_3825 ;
    wire new_AGEMA_signal_3826 ;
    wire new_AGEMA_signal_3827 ;
    wire new_AGEMA_signal_3828 ;
    wire new_AGEMA_signal_3829 ;
    wire new_AGEMA_signal_3830 ;
    wire new_AGEMA_signal_3831 ;
    wire new_AGEMA_signal_3832 ;
    wire new_AGEMA_signal_3833 ;
    wire new_AGEMA_signal_3834 ;
    wire new_AGEMA_signal_3835 ;
    wire new_AGEMA_signal_3836 ;
    wire new_AGEMA_signal_3837 ;
    wire new_AGEMA_signal_3838 ;
    wire new_AGEMA_signal_3839 ;
    wire new_AGEMA_signal_3840 ;
    wire new_AGEMA_signal_3841 ;
    wire new_AGEMA_signal_3842 ;
    wire new_AGEMA_signal_3843 ;
    wire new_AGEMA_signal_3844 ;
    wire new_AGEMA_signal_3845 ;
    wire new_AGEMA_signal_3846 ;
    wire new_AGEMA_signal_3847 ;
    wire new_AGEMA_signal_3848 ;
    wire new_AGEMA_signal_3849 ;
    wire new_AGEMA_signal_3850 ;
    wire new_AGEMA_signal_3851 ;
    wire new_AGEMA_signal_3852 ;
    wire new_AGEMA_signal_3853 ;
    wire new_AGEMA_signal_3854 ;
    wire new_AGEMA_signal_3855 ;
    wire new_AGEMA_signal_3856 ;
    wire new_AGEMA_signal_3857 ;
    wire new_AGEMA_signal_3858 ;
    wire new_AGEMA_signal_3859 ;
    wire new_AGEMA_signal_3860 ;
    wire new_AGEMA_signal_3861 ;
    wire new_AGEMA_signal_3862 ;
    wire new_AGEMA_signal_3863 ;
    wire new_AGEMA_signal_3864 ;
    wire new_AGEMA_signal_3865 ;
    wire new_AGEMA_signal_3866 ;
    wire new_AGEMA_signal_3867 ;
    wire new_AGEMA_signal_3868 ;
    wire new_AGEMA_signal_3869 ;
    wire new_AGEMA_signal_3870 ;
    wire new_AGEMA_signal_3871 ;
    wire new_AGEMA_signal_3872 ;
    wire new_AGEMA_signal_3873 ;
    wire new_AGEMA_signal_3874 ;
    wire new_AGEMA_signal_3875 ;
    wire new_AGEMA_signal_3876 ;
    wire new_AGEMA_signal_3877 ;
    wire new_AGEMA_signal_3878 ;
    wire new_AGEMA_signal_3879 ;
    wire new_AGEMA_signal_3880 ;
    wire new_AGEMA_signal_3881 ;
    wire new_AGEMA_signal_3882 ;
    wire new_AGEMA_signal_3883 ;
    wire new_AGEMA_signal_3884 ;
    wire new_AGEMA_signal_3885 ;
    wire new_AGEMA_signal_3886 ;
    wire new_AGEMA_signal_3887 ;
    wire new_AGEMA_signal_3888 ;
    wire new_AGEMA_signal_3889 ;
    wire new_AGEMA_signal_3890 ;
    wire new_AGEMA_signal_3891 ;
    wire new_AGEMA_signal_3892 ;
    wire new_AGEMA_signal_3893 ;
    wire new_AGEMA_signal_3894 ;
    wire new_AGEMA_signal_3895 ;
    wire new_AGEMA_signal_3896 ;
    wire new_AGEMA_signal_3897 ;
    wire new_AGEMA_signal_3898 ;
    wire new_AGEMA_signal_3899 ;
    wire new_AGEMA_signal_3900 ;
    wire new_AGEMA_signal_3901 ;
    wire new_AGEMA_signal_3902 ;
    wire new_AGEMA_signal_3903 ;
    wire new_AGEMA_signal_3904 ;
    wire new_AGEMA_signal_3905 ;
    wire new_AGEMA_signal_3906 ;
    wire new_AGEMA_signal_3907 ;
    wire new_AGEMA_signal_3908 ;
    wire new_AGEMA_signal_3909 ;
    wire new_AGEMA_signal_3910 ;
    wire new_AGEMA_signal_3911 ;
    wire new_AGEMA_signal_3912 ;
    wire new_AGEMA_signal_3913 ;
    wire new_AGEMA_signal_3914 ;
    wire new_AGEMA_signal_3915 ;
    wire new_AGEMA_signal_3916 ;
    wire new_AGEMA_signal_3917 ;
    wire new_AGEMA_signal_3918 ;
    wire new_AGEMA_signal_3919 ;
    wire new_AGEMA_signal_3920 ;
    wire new_AGEMA_signal_3921 ;
    wire new_AGEMA_signal_3922 ;
    wire new_AGEMA_signal_3923 ;
    wire new_AGEMA_signal_3924 ;
    wire new_AGEMA_signal_3925 ;
    wire new_AGEMA_signal_3926 ;
    wire new_AGEMA_signal_3927 ;
    wire new_AGEMA_signal_3928 ;
    wire new_AGEMA_signal_3929 ;
    wire new_AGEMA_signal_3930 ;
    wire new_AGEMA_signal_3931 ;
    wire new_AGEMA_signal_3932 ;
    wire new_AGEMA_signal_3933 ;
    wire new_AGEMA_signal_3934 ;
    wire new_AGEMA_signal_3935 ;
    wire new_AGEMA_signal_3936 ;
    wire new_AGEMA_signal_3937 ;
    wire new_AGEMA_signal_3938 ;
    wire new_AGEMA_signal_3939 ;
    wire new_AGEMA_signal_3940 ;
    wire new_AGEMA_signal_3941 ;
    wire new_AGEMA_signal_3942 ;
    wire new_AGEMA_signal_3943 ;
    wire new_AGEMA_signal_3944 ;
    wire new_AGEMA_signal_3945 ;
    wire new_AGEMA_signal_3946 ;
    wire new_AGEMA_signal_3947 ;
    wire new_AGEMA_signal_3948 ;
    wire new_AGEMA_signal_3949 ;
    wire new_AGEMA_signal_3950 ;
    wire new_AGEMA_signal_3951 ;
    wire new_AGEMA_signal_3952 ;
    wire new_AGEMA_signal_3953 ;
    wire new_AGEMA_signal_3954 ;
    wire new_AGEMA_signal_3955 ;
    wire new_AGEMA_signal_3956 ;
    wire new_AGEMA_signal_3957 ;
    wire new_AGEMA_signal_3958 ;
    wire new_AGEMA_signal_3959 ;
    wire new_AGEMA_signal_3960 ;
    wire new_AGEMA_signal_3961 ;
    wire new_AGEMA_signal_3962 ;
    wire new_AGEMA_signal_3963 ;
    wire new_AGEMA_signal_3964 ;
    wire new_AGEMA_signal_3965 ;
    wire new_AGEMA_signal_3966 ;
    wire new_AGEMA_signal_3967 ;
    wire new_AGEMA_signal_3968 ;
    wire new_AGEMA_signal_3969 ;
    wire new_AGEMA_signal_3970 ;
    wire new_AGEMA_signal_3971 ;
    wire new_AGEMA_signal_3972 ;
    wire new_AGEMA_signal_3973 ;
    wire new_AGEMA_signal_3974 ;
    wire new_AGEMA_signal_3975 ;
    wire new_AGEMA_signal_3976 ;
    wire new_AGEMA_signal_3977 ;
    wire new_AGEMA_signal_3978 ;
    wire new_AGEMA_signal_3979 ;
    wire new_AGEMA_signal_3980 ;
    wire new_AGEMA_signal_3981 ;
    wire new_AGEMA_signal_3982 ;
    wire new_AGEMA_signal_3983 ;
    wire new_AGEMA_signal_3984 ;
    wire new_AGEMA_signal_3985 ;
    wire new_AGEMA_signal_3986 ;
    wire new_AGEMA_signal_3987 ;
    wire new_AGEMA_signal_3988 ;
    wire new_AGEMA_signal_3989 ;
    wire new_AGEMA_signal_3990 ;
    wire new_AGEMA_signal_3991 ;
    wire new_AGEMA_signal_3992 ;
    wire new_AGEMA_signal_3993 ;
    wire new_AGEMA_signal_3994 ;
    wire new_AGEMA_signal_3995 ;
    wire new_AGEMA_signal_3996 ;
    wire new_AGEMA_signal_3997 ;
    wire new_AGEMA_signal_3998 ;
    wire new_AGEMA_signal_3999 ;
    wire new_AGEMA_signal_4000 ;
    wire new_AGEMA_signal_4001 ;
    wire new_AGEMA_signal_4002 ;
    wire new_AGEMA_signal_4003 ;
    wire new_AGEMA_signal_4004 ;
    wire new_AGEMA_signal_4005 ;
    wire new_AGEMA_signal_4006 ;
    wire new_AGEMA_signal_4007 ;
    wire new_AGEMA_signal_4008 ;
    wire new_AGEMA_signal_4009 ;
    wire new_AGEMA_signal_4010 ;
    wire new_AGEMA_signal_4011 ;
    wire new_AGEMA_signal_4012 ;
    wire new_AGEMA_signal_4013 ;
    wire new_AGEMA_signal_4014 ;
    wire new_AGEMA_signal_4015 ;
    wire new_AGEMA_signal_4016 ;
    wire new_AGEMA_signal_4017 ;
    wire new_AGEMA_signal_4018 ;
    wire new_AGEMA_signal_4019 ;
    wire new_AGEMA_signal_4020 ;
    wire new_AGEMA_signal_4021 ;
    wire new_AGEMA_signal_4022 ;
    wire new_AGEMA_signal_4023 ;
    wire new_AGEMA_signal_4024 ;
    wire new_AGEMA_signal_4025 ;
    wire new_AGEMA_signal_4026 ;
    wire new_AGEMA_signal_4027 ;
    wire new_AGEMA_signal_4028 ;
    wire new_AGEMA_signal_4029 ;
    wire new_AGEMA_signal_4030 ;
    wire new_AGEMA_signal_4031 ;
    wire new_AGEMA_signal_4032 ;
    wire new_AGEMA_signal_4033 ;
    wire new_AGEMA_signal_4034 ;
    wire new_AGEMA_signal_4035 ;
    wire new_AGEMA_signal_4036 ;
    wire new_AGEMA_signal_4037 ;
    wire new_AGEMA_signal_4038 ;
    wire new_AGEMA_signal_4039 ;
    wire new_AGEMA_signal_4040 ;
    wire new_AGEMA_signal_4041 ;
    wire new_AGEMA_signal_4042 ;
    wire new_AGEMA_signal_4043 ;
    wire new_AGEMA_signal_4044 ;
    wire new_AGEMA_signal_4045 ;
    wire new_AGEMA_signal_4046 ;
    wire new_AGEMA_signal_4047 ;
    wire new_AGEMA_signal_4048 ;
    wire new_AGEMA_signal_4049 ;
    wire new_AGEMA_signal_4050 ;
    wire new_AGEMA_signal_4051 ;
    wire new_AGEMA_signal_4052 ;
    wire new_AGEMA_signal_4053 ;
    wire new_AGEMA_signal_4054 ;
    wire new_AGEMA_signal_4055 ;
    wire new_AGEMA_signal_4056 ;
    wire new_AGEMA_signal_4057 ;
    wire new_AGEMA_signal_4058 ;
    wire new_AGEMA_signal_4059 ;
    wire new_AGEMA_signal_4060 ;
    wire new_AGEMA_signal_4061 ;
    wire new_AGEMA_signal_4062 ;
    wire new_AGEMA_signal_4063 ;
    wire new_AGEMA_signal_4064 ;
    wire new_AGEMA_signal_4065 ;
    wire new_AGEMA_signal_4066 ;
    wire new_AGEMA_signal_4067 ;
    wire new_AGEMA_signal_4068 ;
    wire new_AGEMA_signal_4069 ;
    wire new_AGEMA_signal_4070 ;
    wire new_AGEMA_signal_4071 ;
    wire new_AGEMA_signal_4072 ;
    wire new_AGEMA_signal_4073 ;
    wire new_AGEMA_signal_4074 ;
    wire new_AGEMA_signal_4075 ;
    wire new_AGEMA_signal_4076 ;
    wire new_AGEMA_signal_4077 ;
    wire new_AGEMA_signal_4078 ;
    wire new_AGEMA_signal_4079 ;
    wire new_AGEMA_signal_4080 ;
    wire new_AGEMA_signal_4081 ;
    wire new_AGEMA_signal_4082 ;
    wire new_AGEMA_signal_4083 ;
    wire new_AGEMA_signal_4084 ;
    wire new_AGEMA_signal_4085 ;
    wire new_AGEMA_signal_4086 ;
    wire new_AGEMA_signal_4087 ;
    wire new_AGEMA_signal_4088 ;
    wire new_AGEMA_signal_4089 ;
    wire new_AGEMA_signal_4090 ;
    wire new_AGEMA_signal_4091 ;
    wire new_AGEMA_signal_4092 ;
    wire new_AGEMA_signal_4093 ;
    wire new_AGEMA_signal_4094 ;
    wire new_AGEMA_signal_4095 ;
    wire new_AGEMA_signal_4096 ;
    wire new_AGEMA_signal_4097 ;
    wire new_AGEMA_signal_4098 ;
    wire new_AGEMA_signal_4099 ;
    wire new_AGEMA_signal_4100 ;
    wire new_AGEMA_signal_4101 ;
    wire new_AGEMA_signal_4102 ;
    wire new_AGEMA_signal_4103 ;
    wire new_AGEMA_signal_4104 ;
    wire new_AGEMA_signal_4105 ;
    wire new_AGEMA_signal_4106 ;
    wire new_AGEMA_signal_4107 ;
    wire new_AGEMA_signal_4108 ;
    wire new_AGEMA_signal_4109 ;
    wire new_AGEMA_signal_4110 ;
    wire new_AGEMA_signal_4111 ;
    wire new_AGEMA_signal_4112 ;
    wire new_AGEMA_signal_4113 ;
    wire new_AGEMA_signal_4114 ;
    wire new_AGEMA_signal_4115 ;
    wire new_AGEMA_signal_4116 ;
    wire new_AGEMA_signal_4117 ;
    wire new_AGEMA_signal_4118 ;
    wire new_AGEMA_signal_4119 ;
    wire new_AGEMA_signal_4120 ;
    wire new_AGEMA_signal_4121 ;
    wire new_AGEMA_signal_4122 ;
    wire new_AGEMA_signal_4123 ;
    wire new_AGEMA_signal_4124 ;
    wire new_AGEMA_signal_4125 ;
    wire new_AGEMA_signal_4126 ;
    wire new_AGEMA_signal_4127 ;
    wire new_AGEMA_signal_4128 ;
    wire new_AGEMA_signal_4129 ;
    wire new_AGEMA_signal_4130 ;
    wire new_AGEMA_signal_4131 ;
    wire new_AGEMA_signal_4132 ;
    wire new_AGEMA_signal_4133 ;
    wire new_AGEMA_signal_4134 ;
    wire new_AGEMA_signal_4135 ;
    wire new_AGEMA_signal_4136 ;
    wire new_AGEMA_signal_4137 ;
    wire new_AGEMA_signal_4138 ;
    wire new_AGEMA_signal_4139 ;
    wire new_AGEMA_signal_4140 ;
    wire new_AGEMA_signal_4141 ;
    wire new_AGEMA_signal_4142 ;
    wire new_AGEMA_signal_4143 ;
    wire new_AGEMA_signal_4144 ;
    wire new_AGEMA_signal_4145 ;
    wire new_AGEMA_signal_4146 ;
    wire new_AGEMA_signal_4147 ;
    wire new_AGEMA_signal_4148 ;
    wire new_AGEMA_signal_4149 ;
    wire new_AGEMA_signal_4150 ;
    wire new_AGEMA_signal_4151 ;
    wire new_AGEMA_signal_4152 ;
    wire new_AGEMA_signal_4153 ;
    wire new_AGEMA_signal_4154 ;
    wire new_AGEMA_signal_4155 ;
    wire new_AGEMA_signal_4156 ;
    wire new_AGEMA_signal_4157 ;
    wire new_AGEMA_signal_4158 ;
    wire new_AGEMA_signal_4159 ;
    wire new_AGEMA_signal_4160 ;
    wire new_AGEMA_signal_4161 ;
    wire new_AGEMA_signal_4162 ;
    wire new_AGEMA_signal_4163 ;
    wire new_AGEMA_signal_4164 ;
    wire new_AGEMA_signal_4165 ;
    wire new_AGEMA_signal_4166 ;
    wire new_AGEMA_signal_4167 ;
    wire new_AGEMA_signal_4168 ;
    wire new_AGEMA_signal_4169 ;
    wire new_AGEMA_signal_4170 ;
    wire new_AGEMA_signal_4171 ;
    wire new_AGEMA_signal_4172 ;
    wire new_AGEMA_signal_4173 ;
    wire new_AGEMA_signal_4174 ;
    wire new_AGEMA_signal_4175 ;
    wire new_AGEMA_signal_4176 ;
    wire new_AGEMA_signal_4177 ;
    wire new_AGEMA_signal_4178 ;
    wire new_AGEMA_signal_4179 ;
    wire new_AGEMA_signal_4180 ;
    wire new_AGEMA_signal_4181 ;
    wire new_AGEMA_signal_4182 ;
    wire new_AGEMA_signal_4183 ;
    wire new_AGEMA_signal_4184 ;
    wire new_AGEMA_signal_4185 ;
    wire new_AGEMA_signal_4186 ;
    wire new_AGEMA_signal_4187 ;
    wire new_AGEMA_signal_4188 ;
    wire new_AGEMA_signal_4189 ;
    wire new_AGEMA_signal_4190 ;
    wire new_AGEMA_signal_4191 ;
    wire new_AGEMA_signal_4192 ;
    wire new_AGEMA_signal_4193 ;
    wire new_AGEMA_signal_4194 ;
    wire new_AGEMA_signal_4195 ;
    wire new_AGEMA_signal_4196 ;
    wire new_AGEMA_signal_4197 ;
    wire new_AGEMA_signal_4198 ;
    wire new_AGEMA_signal_4199 ;
    wire new_AGEMA_signal_4200 ;
    wire new_AGEMA_signal_4201 ;
    wire new_AGEMA_signal_4202 ;
    wire new_AGEMA_signal_4203 ;
    wire new_AGEMA_signal_4204 ;
    wire new_AGEMA_signal_4205 ;
    wire new_AGEMA_signal_4206 ;
    wire new_AGEMA_signal_4207 ;
    wire new_AGEMA_signal_4208 ;
    wire new_AGEMA_signal_4209 ;
    wire new_AGEMA_signal_4210 ;
    wire new_AGEMA_signal_4211 ;
    wire new_AGEMA_signal_4212 ;
    wire new_AGEMA_signal_4213 ;
    wire new_AGEMA_signal_4214 ;
    wire new_AGEMA_signal_4215 ;
    wire new_AGEMA_signal_4216 ;
    wire new_AGEMA_signal_4217 ;
    wire new_AGEMA_signal_4218 ;
    wire new_AGEMA_signal_4219 ;
    wire new_AGEMA_signal_4220 ;
    wire new_AGEMA_signal_4221 ;
    wire new_AGEMA_signal_4222 ;
    wire new_AGEMA_signal_4223 ;
    wire new_AGEMA_signal_4224 ;
    wire new_AGEMA_signal_4225 ;
    wire new_AGEMA_signal_4226 ;
    wire new_AGEMA_signal_4227 ;
    wire new_AGEMA_signal_4228 ;
    wire new_AGEMA_signal_4229 ;
    wire new_AGEMA_signal_4230 ;
    wire new_AGEMA_signal_4231 ;
    wire new_AGEMA_signal_4232 ;
    wire new_AGEMA_signal_4233 ;
    wire new_AGEMA_signal_4234 ;
    wire new_AGEMA_signal_4235 ;
    wire new_AGEMA_signal_4236 ;
    wire new_AGEMA_signal_4237 ;
    wire new_AGEMA_signal_4238 ;
    wire new_AGEMA_signal_4239 ;
    wire new_AGEMA_signal_4240 ;
    wire new_AGEMA_signal_4241 ;
    wire new_AGEMA_signal_4242 ;
    wire new_AGEMA_signal_4243 ;
    wire new_AGEMA_signal_4244 ;
    wire new_AGEMA_signal_4245 ;
    wire new_AGEMA_signal_4246 ;
    wire new_AGEMA_signal_4247 ;
    wire new_AGEMA_signal_4248 ;
    wire new_AGEMA_signal_4249 ;
    wire new_AGEMA_signal_4250 ;
    wire new_AGEMA_signal_4251 ;
    wire new_AGEMA_signal_4252 ;
    wire new_AGEMA_signal_4253 ;
    wire new_AGEMA_signal_4254 ;
    wire new_AGEMA_signal_4255 ;
    wire new_AGEMA_signal_4256 ;
    wire new_AGEMA_signal_4257 ;
    wire new_AGEMA_signal_4258 ;
    wire new_AGEMA_signal_4259 ;
    wire new_AGEMA_signal_4260 ;
    wire new_AGEMA_signal_4261 ;
    wire new_AGEMA_signal_4262 ;
    wire new_AGEMA_signal_4263 ;
    wire new_AGEMA_signal_4264 ;
    wire new_AGEMA_signal_4265 ;
    wire new_AGEMA_signal_4266 ;
    wire new_AGEMA_signal_4267 ;
    wire new_AGEMA_signal_4268 ;
    wire new_AGEMA_signal_4269 ;
    wire new_AGEMA_signal_4270 ;
    wire new_AGEMA_signal_4271 ;
    wire new_AGEMA_signal_4272 ;
    wire new_AGEMA_signal_4273 ;
    wire new_AGEMA_signal_4274 ;
    wire new_AGEMA_signal_4275 ;
    wire new_AGEMA_signal_4276 ;
    wire new_AGEMA_signal_4277 ;
    wire new_AGEMA_signal_4278 ;
    wire new_AGEMA_signal_4279 ;
    wire new_AGEMA_signal_4280 ;
    wire new_AGEMA_signal_4281 ;
    wire new_AGEMA_signal_4282 ;
    wire new_AGEMA_signal_4283 ;
    wire new_AGEMA_signal_4284 ;
    wire new_AGEMA_signal_4285 ;
    wire new_AGEMA_signal_4286 ;
    wire new_AGEMA_signal_4287 ;
    wire new_AGEMA_signal_4288 ;
    wire new_AGEMA_signal_4289 ;
    wire new_AGEMA_signal_4290 ;
    wire new_AGEMA_signal_4291 ;
    wire new_AGEMA_signal_4292 ;
    wire new_AGEMA_signal_4293 ;
    wire new_AGEMA_signal_4294 ;
    wire new_AGEMA_signal_4295 ;
    wire new_AGEMA_signal_4296 ;
    wire new_AGEMA_signal_4297 ;
    wire new_AGEMA_signal_4298 ;
    wire new_AGEMA_signal_4299 ;
    wire new_AGEMA_signal_4300 ;
    wire new_AGEMA_signal_4301 ;
    wire new_AGEMA_signal_4302 ;
    wire new_AGEMA_signal_4303 ;
    wire new_AGEMA_signal_4304 ;
    wire new_AGEMA_signal_4305 ;
    wire new_AGEMA_signal_4306 ;
    wire new_AGEMA_signal_4307 ;
    wire new_AGEMA_signal_4308 ;
    wire new_AGEMA_signal_4309 ;
    wire new_AGEMA_signal_4310 ;
    wire new_AGEMA_signal_4311 ;
    wire new_AGEMA_signal_4312 ;
    wire new_AGEMA_signal_4313 ;
    wire new_AGEMA_signal_4314 ;
    wire new_AGEMA_signal_4315 ;
    wire new_AGEMA_signal_4316 ;
    wire new_AGEMA_signal_4317 ;
    wire new_AGEMA_signal_4318 ;
    wire new_AGEMA_signal_4319 ;
    wire new_AGEMA_signal_4320 ;
    wire new_AGEMA_signal_4321 ;
    wire new_AGEMA_signal_4322 ;
    wire new_AGEMA_signal_4323 ;
    wire new_AGEMA_signal_4324 ;
    wire new_AGEMA_signal_4325 ;
    wire new_AGEMA_signal_4326 ;
    wire new_AGEMA_signal_4327 ;
    wire new_AGEMA_signal_4328 ;
    wire new_AGEMA_signal_4329 ;
    wire new_AGEMA_signal_4330 ;
    wire new_AGEMA_signal_4331 ;
    wire new_AGEMA_signal_4332 ;
    wire new_AGEMA_signal_4333 ;
    wire new_AGEMA_signal_4334 ;
    wire new_AGEMA_signal_4335 ;
    wire new_AGEMA_signal_4336 ;
    wire new_AGEMA_signal_4337 ;
    wire new_AGEMA_signal_4338 ;
    wire new_AGEMA_signal_4339 ;
    wire new_AGEMA_signal_4340 ;
    wire new_AGEMA_signal_4341 ;
    wire new_AGEMA_signal_4342 ;
    wire new_AGEMA_signal_4343 ;
    wire new_AGEMA_signal_4344 ;
    wire new_AGEMA_signal_4345 ;
    wire new_AGEMA_signal_4346 ;
    wire new_AGEMA_signal_4347 ;
    wire new_AGEMA_signal_4348 ;
    wire new_AGEMA_signal_4349 ;
    wire new_AGEMA_signal_4350 ;
    wire new_AGEMA_signal_4351 ;
    wire new_AGEMA_signal_4352 ;
    wire new_AGEMA_signal_4353 ;
    wire new_AGEMA_signal_4354 ;
    wire new_AGEMA_signal_4355 ;
    wire new_AGEMA_signal_4356 ;
    wire new_AGEMA_signal_4357 ;
    wire new_AGEMA_signal_4358 ;
    wire new_AGEMA_signal_4359 ;
    wire new_AGEMA_signal_4360 ;
    wire new_AGEMA_signal_4361 ;
    wire new_AGEMA_signal_4362 ;
    wire new_AGEMA_signal_4363 ;
    wire new_AGEMA_signal_4364 ;
    wire new_AGEMA_signal_4365 ;
    wire new_AGEMA_signal_4366 ;
    wire new_AGEMA_signal_4367 ;
    wire new_AGEMA_signal_4368 ;
    wire new_AGEMA_signal_4369 ;
    wire new_AGEMA_signal_4370 ;
    wire new_AGEMA_signal_4371 ;
    wire new_AGEMA_signal_4372 ;
    wire new_AGEMA_signal_4373 ;
    wire new_AGEMA_signal_4374 ;
    wire new_AGEMA_signal_4375 ;
    wire new_AGEMA_signal_4376 ;
    wire new_AGEMA_signal_4377 ;
    wire new_AGEMA_signal_4378 ;
    wire new_AGEMA_signal_4379 ;
    wire new_AGEMA_signal_4380 ;
    wire new_AGEMA_signal_4381 ;
    wire new_AGEMA_signal_4382 ;
    wire new_AGEMA_signal_4383 ;
    wire new_AGEMA_signal_4384 ;
    wire new_AGEMA_signal_4385 ;
    wire new_AGEMA_signal_4386 ;
    wire new_AGEMA_signal_4387 ;
    wire new_AGEMA_signal_4388 ;
    wire new_AGEMA_signal_4389 ;
    wire new_AGEMA_signal_4390 ;
    wire new_AGEMA_signal_4391 ;
    wire new_AGEMA_signal_4392 ;
    wire new_AGEMA_signal_4393 ;
    wire new_AGEMA_signal_4394 ;
    wire new_AGEMA_signal_4395 ;
    wire new_AGEMA_signal_4396 ;
    wire new_AGEMA_signal_4397 ;
    wire new_AGEMA_signal_4398 ;
    wire new_AGEMA_signal_4399 ;
    wire new_AGEMA_signal_4400 ;
    wire new_AGEMA_signal_4401 ;
    wire new_AGEMA_signal_4402 ;
    wire new_AGEMA_signal_4403 ;
    wire new_AGEMA_signal_4404 ;
    wire new_AGEMA_signal_4405 ;
    wire new_AGEMA_signal_4406 ;
    wire new_AGEMA_signal_4407 ;
    wire new_AGEMA_signal_4408 ;
    wire new_AGEMA_signal_4409 ;
    wire new_AGEMA_signal_4410 ;
    wire new_AGEMA_signal_4411 ;
    wire new_AGEMA_signal_4412 ;
    wire new_AGEMA_signal_4413 ;
    wire new_AGEMA_signal_4414 ;
    wire new_AGEMA_signal_4415 ;
    wire new_AGEMA_signal_4416 ;
    wire new_AGEMA_signal_4417 ;
    wire new_AGEMA_signal_4418 ;
    wire new_AGEMA_signal_4419 ;
    wire new_AGEMA_signal_4420 ;
    wire new_AGEMA_signal_4421 ;
    wire new_AGEMA_signal_4422 ;
    wire new_AGEMA_signal_4423 ;
    wire new_AGEMA_signal_4424 ;
    wire new_AGEMA_signal_4425 ;
    wire new_AGEMA_signal_4426 ;
    wire new_AGEMA_signal_4427 ;
    wire new_AGEMA_signal_4428 ;
    wire new_AGEMA_signal_4429 ;
    wire new_AGEMA_signal_4430 ;
    wire new_AGEMA_signal_4431 ;
    wire new_AGEMA_signal_4432 ;
    wire new_AGEMA_signal_4433 ;
    wire new_AGEMA_signal_4434 ;
    wire new_AGEMA_signal_4435 ;
    wire new_AGEMA_signal_4436 ;
    wire new_AGEMA_signal_4437 ;
    wire new_AGEMA_signal_4438 ;
    wire new_AGEMA_signal_4439 ;
    wire new_AGEMA_signal_4440 ;
    wire new_AGEMA_signal_4441 ;
    wire new_AGEMA_signal_4442 ;
    wire new_AGEMA_signal_4443 ;
    wire new_AGEMA_signal_4444 ;
    wire new_AGEMA_signal_4445 ;
    wire new_AGEMA_signal_4446 ;
    wire new_AGEMA_signal_4447 ;
    wire new_AGEMA_signal_4448 ;
    wire new_AGEMA_signal_4449 ;
    wire new_AGEMA_signal_4450 ;
    wire new_AGEMA_signal_4451 ;
    wire new_AGEMA_signal_4452 ;
    wire new_AGEMA_signal_4453 ;
    wire new_AGEMA_signal_4454 ;
    wire new_AGEMA_signal_4455 ;
    wire new_AGEMA_signal_4456 ;
    wire new_AGEMA_signal_4457 ;
    wire new_AGEMA_signal_4458 ;
    wire new_AGEMA_signal_4459 ;
    wire new_AGEMA_signal_4460 ;
    wire new_AGEMA_signal_4461 ;
    wire new_AGEMA_signal_4462 ;
    wire new_AGEMA_signal_4463 ;
    wire new_AGEMA_signal_4464 ;
    wire new_AGEMA_signal_4465 ;
    wire new_AGEMA_signal_4466 ;
    wire new_AGEMA_signal_4467 ;
    wire new_AGEMA_signal_4468 ;
    wire new_AGEMA_signal_4469 ;
    wire new_AGEMA_signal_4470 ;
    wire new_AGEMA_signal_4471 ;
    wire new_AGEMA_signal_4472 ;
    wire new_AGEMA_signal_4473 ;
    wire new_AGEMA_signal_4474 ;
    wire new_AGEMA_signal_4475 ;
    wire new_AGEMA_signal_4476 ;
    wire new_AGEMA_signal_4477 ;
    wire new_AGEMA_signal_4478 ;
    wire new_AGEMA_signal_4479 ;
    wire new_AGEMA_signal_4480 ;
    wire new_AGEMA_signal_4481 ;
    wire new_AGEMA_signal_4482 ;
    wire new_AGEMA_signal_4483 ;
    wire new_AGEMA_signal_4484 ;
    wire new_AGEMA_signal_4485 ;
    wire new_AGEMA_signal_4486 ;
    wire new_AGEMA_signal_4487 ;
    wire new_AGEMA_signal_4488 ;
    wire new_AGEMA_signal_4489 ;
    wire new_AGEMA_signal_4490 ;
    wire new_AGEMA_signal_4491 ;
    wire new_AGEMA_signal_4492 ;
    wire new_AGEMA_signal_4493 ;
    wire new_AGEMA_signal_4494 ;
    wire new_AGEMA_signal_4495 ;
    wire new_AGEMA_signal_4496 ;
    wire new_AGEMA_signal_4497 ;
    wire new_AGEMA_signal_4498 ;
    wire new_AGEMA_signal_4499 ;
    wire new_AGEMA_signal_4500 ;
    wire new_AGEMA_signal_4501 ;
    wire new_AGEMA_signal_4502 ;
    wire new_AGEMA_signal_4503 ;
    wire new_AGEMA_signal_4504 ;
    wire new_AGEMA_signal_4505 ;
    wire new_AGEMA_signal_4506 ;
    wire new_AGEMA_signal_4507 ;
    wire new_AGEMA_signal_4508 ;
    wire new_AGEMA_signal_4509 ;
    wire new_AGEMA_signal_4510 ;
    wire new_AGEMA_signal_4511 ;
    wire new_AGEMA_signal_4512 ;
    wire new_AGEMA_signal_4513 ;
    wire new_AGEMA_signal_4514 ;
    wire new_AGEMA_signal_4515 ;
    wire new_AGEMA_signal_4516 ;
    wire new_AGEMA_signal_4517 ;
    wire new_AGEMA_signal_4518 ;
    wire new_AGEMA_signal_4519 ;
    wire new_AGEMA_signal_4520 ;
    wire new_AGEMA_signal_4521 ;
    wire new_AGEMA_signal_4522 ;
    wire new_AGEMA_signal_4523 ;
    wire new_AGEMA_signal_4524 ;
    wire new_AGEMA_signal_4525 ;
    wire new_AGEMA_signal_4526 ;
    wire new_AGEMA_signal_4527 ;
    wire new_AGEMA_signal_4528 ;
    wire new_AGEMA_signal_4529 ;
    wire new_AGEMA_signal_4530 ;
    wire new_AGEMA_signal_4531 ;
    wire new_AGEMA_signal_4532 ;
    wire new_AGEMA_signal_4533 ;
    wire new_AGEMA_signal_4534 ;
    wire new_AGEMA_signal_4535 ;
    wire new_AGEMA_signal_4536 ;
    wire new_AGEMA_signal_4537 ;
    wire new_AGEMA_signal_4538 ;
    wire new_AGEMA_signal_4539 ;
    wire new_AGEMA_signal_4540 ;
    wire new_AGEMA_signal_4541 ;
    wire new_AGEMA_signal_4542 ;
    wire new_AGEMA_signal_4543 ;
    wire new_AGEMA_signal_4544 ;
    wire new_AGEMA_signal_4545 ;
    wire new_AGEMA_signal_4546 ;
    wire new_AGEMA_signal_4547 ;
    wire new_AGEMA_signal_4548 ;
    wire new_AGEMA_signal_4549 ;
    wire new_AGEMA_signal_4550 ;
    wire new_AGEMA_signal_4551 ;
    wire new_AGEMA_signal_4552 ;
    wire new_AGEMA_signal_4553 ;
    wire new_AGEMA_signal_4554 ;
    wire new_AGEMA_signal_4555 ;
    wire new_AGEMA_signal_4556 ;
    wire new_AGEMA_signal_4557 ;
    wire new_AGEMA_signal_4558 ;
    wire new_AGEMA_signal_4559 ;
    wire new_AGEMA_signal_4560 ;
    wire new_AGEMA_signal_4561 ;
    wire new_AGEMA_signal_4562 ;
    wire new_AGEMA_signal_4563 ;
    wire new_AGEMA_signal_4564 ;
    wire new_AGEMA_signal_4565 ;
    wire new_AGEMA_signal_4566 ;
    wire new_AGEMA_signal_4567 ;
    wire new_AGEMA_signal_4568 ;
    wire new_AGEMA_signal_4569 ;
    wire new_AGEMA_signal_4570 ;
    wire new_AGEMA_signal_4571 ;
    wire new_AGEMA_signal_4572 ;
    wire new_AGEMA_signal_4573 ;
    wire new_AGEMA_signal_4574 ;
    wire new_AGEMA_signal_4575 ;
    wire new_AGEMA_signal_4576 ;
    wire new_AGEMA_signal_4577 ;
    wire new_AGEMA_signal_4578 ;
    wire new_AGEMA_signal_4579 ;
    wire new_AGEMA_signal_4580 ;
    wire new_AGEMA_signal_4581 ;
    wire new_AGEMA_signal_4582 ;
    wire new_AGEMA_signal_4583 ;
    wire new_AGEMA_signal_4584 ;
    wire new_AGEMA_signal_4585 ;
    wire new_AGEMA_signal_4586 ;
    wire new_AGEMA_signal_4587 ;
    wire new_AGEMA_signal_4588 ;
    wire new_AGEMA_signal_4589 ;
    wire new_AGEMA_signal_4590 ;
    wire new_AGEMA_signal_4591 ;
    wire new_AGEMA_signal_4592 ;
    wire new_AGEMA_signal_4593 ;
    wire new_AGEMA_signal_4594 ;
    wire new_AGEMA_signal_4595 ;
    wire new_AGEMA_signal_4596 ;
    wire new_AGEMA_signal_4597 ;
    wire new_AGEMA_signal_4598 ;
    wire new_AGEMA_signal_4599 ;
    wire new_AGEMA_signal_4600 ;
    wire new_AGEMA_signal_4601 ;
    wire new_AGEMA_signal_4602 ;
    wire new_AGEMA_signal_4603 ;
    wire new_AGEMA_signal_4604 ;
    wire new_AGEMA_signal_4605 ;
    wire new_AGEMA_signal_4606 ;
    wire new_AGEMA_signal_4607 ;
    wire new_AGEMA_signal_4608 ;
    wire new_AGEMA_signal_4609 ;
    wire new_AGEMA_signal_4610 ;
    wire new_AGEMA_signal_4611 ;
    wire new_AGEMA_signal_4612 ;
    wire new_AGEMA_signal_4613 ;
    wire new_AGEMA_signal_4614 ;
    wire new_AGEMA_signal_4615 ;
    wire new_AGEMA_signal_4616 ;
    wire new_AGEMA_signal_4617 ;
    wire new_AGEMA_signal_4618 ;
    wire new_AGEMA_signal_4619 ;
    wire new_AGEMA_signal_4620 ;
    wire new_AGEMA_signal_4621 ;
    wire new_AGEMA_signal_4622 ;
    wire new_AGEMA_signal_4623 ;
    wire new_AGEMA_signal_4624 ;
    wire new_AGEMA_signal_4625 ;
    wire new_AGEMA_signal_4626 ;
    wire new_AGEMA_signal_4627 ;
    wire new_AGEMA_signal_4628 ;
    wire new_AGEMA_signal_4629 ;
    wire new_AGEMA_signal_4630 ;
    wire new_AGEMA_signal_4631 ;
    wire new_AGEMA_signal_4632 ;
    wire new_AGEMA_signal_4633 ;
    wire new_AGEMA_signal_4634 ;
    wire new_AGEMA_signal_4635 ;
    wire new_AGEMA_signal_4636 ;
    wire new_AGEMA_signal_4637 ;
    wire new_AGEMA_signal_4638 ;
    wire new_AGEMA_signal_4639 ;
    wire new_AGEMA_signal_4640 ;
    wire new_AGEMA_signal_4641 ;
    wire new_AGEMA_signal_4642 ;
    wire new_AGEMA_signal_4643 ;
    wire new_AGEMA_signal_4644 ;
    wire new_AGEMA_signal_4645 ;
    wire new_AGEMA_signal_4646 ;
    wire new_AGEMA_signal_4647 ;
    wire new_AGEMA_signal_4648 ;
    wire new_AGEMA_signal_4649 ;
    wire new_AGEMA_signal_4650 ;
    wire new_AGEMA_signal_4651 ;
    wire new_AGEMA_signal_4652 ;
    wire new_AGEMA_signal_4653 ;
    wire new_AGEMA_signal_4654 ;
    wire new_AGEMA_signal_4655 ;
    wire new_AGEMA_signal_4656 ;
    wire new_AGEMA_signal_4657 ;
    wire new_AGEMA_signal_4658 ;
    wire new_AGEMA_signal_4659 ;
    wire new_AGEMA_signal_4660 ;
    wire new_AGEMA_signal_4661 ;
    wire new_AGEMA_signal_4662 ;
    wire new_AGEMA_signal_4663 ;
    wire new_AGEMA_signal_4664 ;
    wire new_AGEMA_signal_4665 ;
    wire new_AGEMA_signal_4666 ;
    wire new_AGEMA_signal_4667 ;
    wire new_AGEMA_signal_4668 ;
    wire new_AGEMA_signal_4669 ;
    wire new_AGEMA_signal_4670 ;
    wire new_AGEMA_signal_4671 ;
    wire new_AGEMA_signal_4672 ;
    wire new_AGEMA_signal_4673 ;
    wire new_AGEMA_signal_4674 ;
    wire new_AGEMA_signal_4675 ;
    wire new_AGEMA_signal_4676 ;
    wire new_AGEMA_signal_4677 ;
    wire new_AGEMA_signal_4678 ;
    wire new_AGEMA_signal_4679 ;
    wire new_AGEMA_signal_4680 ;
    wire new_AGEMA_signal_4681 ;
    wire new_AGEMA_signal_4682 ;
    wire new_AGEMA_signal_4683 ;
    wire new_AGEMA_signal_4684 ;
    wire new_AGEMA_signal_4685 ;
    wire new_AGEMA_signal_4686 ;
    wire new_AGEMA_signal_4687 ;
    wire new_AGEMA_signal_4688 ;
    wire new_AGEMA_signal_4689 ;
    wire new_AGEMA_signal_4690 ;
    wire new_AGEMA_signal_4691 ;
    wire new_AGEMA_signal_4692 ;
    wire new_AGEMA_signal_4693 ;
    wire new_AGEMA_signal_4694 ;
    wire new_AGEMA_signal_4695 ;
    wire new_AGEMA_signal_4696 ;
    wire new_AGEMA_signal_4697 ;
    wire new_AGEMA_signal_4698 ;
    wire new_AGEMA_signal_4699 ;
    wire new_AGEMA_signal_4700 ;
    wire new_AGEMA_signal_4701 ;
    wire new_AGEMA_signal_4702 ;
    wire new_AGEMA_signal_4703 ;
    wire new_AGEMA_signal_4704 ;
    wire new_AGEMA_signal_4705 ;
    wire new_AGEMA_signal_4706 ;
    wire new_AGEMA_signal_4707 ;
    wire new_AGEMA_signal_4708 ;
    wire new_AGEMA_signal_4709 ;
    wire new_AGEMA_signal_4710 ;
    wire new_AGEMA_signal_4711 ;
    wire new_AGEMA_signal_4712 ;
    wire new_AGEMA_signal_4713 ;
    wire new_AGEMA_signal_4714 ;
    wire new_AGEMA_signal_4715 ;
    wire new_AGEMA_signal_4716 ;
    wire new_AGEMA_signal_4717 ;
    wire new_AGEMA_signal_4718 ;
    wire new_AGEMA_signal_4719 ;
    wire new_AGEMA_signal_4720 ;
    wire new_AGEMA_signal_4721 ;
    wire new_AGEMA_signal_4722 ;
    wire new_AGEMA_signal_4723 ;
    wire new_AGEMA_signal_4724 ;
    wire new_AGEMA_signal_4725 ;
    wire new_AGEMA_signal_4726 ;
    wire new_AGEMA_signal_4727 ;
    wire new_AGEMA_signal_4728 ;
    wire new_AGEMA_signal_4729 ;
    wire new_AGEMA_signal_4730 ;
    wire new_AGEMA_signal_4731 ;
    wire new_AGEMA_signal_4732 ;
    wire new_AGEMA_signal_4733 ;
    wire new_AGEMA_signal_4734 ;
    wire new_AGEMA_signal_4735 ;
    wire new_AGEMA_signal_4736 ;
    wire new_AGEMA_signal_4737 ;
    wire new_AGEMA_signal_4738 ;
    wire new_AGEMA_signal_4739 ;
    wire new_AGEMA_signal_4740 ;
    wire new_AGEMA_signal_4741 ;
    wire new_AGEMA_signal_4742 ;
    wire new_AGEMA_signal_4743 ;
    wire new_AGEMA_signal_4744 ;
    wire new_AGEMA_signal_4745 ;
    wire new_AGEMA_signal_4746 ;
    wire new_AGEMA_signal_4747 ;
    wire new_AGEMA_signal_4748 ;
    wire new_AGEMA_signal_4749 ;
    wire new_AGEMA_signal_4750 ;
    wire new_AGEMA_signal_4751 ;
    wire new_AGEMA_signal_4752 ;
    wire new_AGEMA_signal_4753 ;
    wire new_AGEMA_signal_4754 ;
    wire new_AGEMA_signal_4755 ;
    wire new_AGEMA_signal_4756 ;
    wire new_AGEMA_signal_4757 ;
    wire new_AGEMA_signal_4758 ;
    wire new_AGEMA_signal_4759 ;
    wire new_AGEMA_signal_4760 ;
    wire new_AGEMA_signal_4761 ;
    wire new_AGEMA_signal_4762 ;
    wire new_AGEMA_signal_4763 ;
    wire new_AGEMA_signal_4764 ;
    wire new_AGEMA_signal_4765 ;
    wire new_AGEMA_signal_4766 ;
    wire new_AGEMA_signal_4767 ;
    wire new_AGEMA_signal_4768 ;
    wire new_AGEMA_signal_4769 ;
    wire new_AGEMA_signal_4770 ;
    wire new_AGEMA_signal_4771 ;
    wire new_AGEMA_signal_4772 ;
    wire new_AGEMA_signal_4773 ;
    wire new_AGEMA_signal_4774 ;
    wire new_AGEMA_signal_4775 ;
    wire new_AGEMA_signal_4776 ;
    wire new_AGEMA_signal_4777 ;
    wire new_AGEMA_signal_4778 ;
    wire new_AGEMA_signal_4779 ;
    wire new_AGEMA_signal_4780 ;
    wire new_AGEMA_signal_4781 ;
    wire new_AGEMA_signal_4782 ;
    wire new_AGEMA_signal_4783 ;
    wire new_AGEMA_signal_4784 ;
    wire new_AGEMA_signal_4785 ;
    wire new_AGEMA_signal_4786 ;
    wire new_AGEMA_signal_4787 ;
    wire new_AGEMA_signal_4788 ;
    wire new_AGEMA_signal_4789 ;
    wire new_AGEMA_signal_4790 ;
    wire new_AGEMA_signal_4791 ;
    wire new_AGEMA_signal_4792 ;
    wire new_AGEMA_signal_4793 ;
    wire new_AGEMA_signal_4794 ;
    wire new_AGEMA_signal_4795 ;
    wire new_AGEMA_signal_4796 ;
    wire new_AGEMA_signal_4797 ;
    wire new_AGEMA_signal_4798 ;
    wire new_AGEMA_signal_4799 ;
    wire new_AGEMA_signal_4800 ;
    wire new_AGEMA_signal_4801 ;
    wire new_AGEMA_signal_4802 ;
    wire new_AGEMA_signal_4803 ;
    wire new_AGEMA_signal_4804 ;
    wire new_AGEMA_signal_4805 ;
    wire new_AGEMA_signal_4806 ;
    wire new_AGEMA_signal_4807 ;
    wire new_AGEMA_signal_4808 ;
    wire new_AGEMA_signal_4809 ;
    wire new_AGEMA_signal_4810 ;
    wire new_AGEMA_signal_4811 ;
    wire new_AGEMA_signal_4812 ;
    wire new_AGEMA_signal_4813 ;
    wire new_AGEMA_signal_4814 ;
    wire new_AGEMA_signal_4815 ;
    wire new_AGEMA_signal_4816 ;
    wire new_AGEMA_signal_4817 ;
    wire new_AGEMA_signal_4818 ;
    wire new_AGEMA_signal_4819 ;
    wire new_AGEMA_signal_4820 ;
    wire new_AGEMA_signal_4821 ;
    wire new_AGEMA_signal_4822 ;
    wire new_AGEMA_signal_4823 ;
    wire new_AGEMA_signal_4824 ;
    wire new_AGEMA_signal_4825 ;
    wire new_AGEMA_signal_4826 ;
    wire new_AGEMA_signal_4827 ;
    wire new_AGEMA_signal_4828 ;
    wire new_AGEMA_signal_4829 ;
    wire new_AGEMA_signal_4830 ;
    wire new_AGEMA_signal_4831 ;
    wire new_AGEMA_signal_4832 ;
    wire new_AGEMA_signal_4833 ;
    wire new_AGEMA_signal_4834 ;
    wire new_AGEMA_signal_4835 ;
    wire new_AGEMA_signal_4836 ;
    wire new_AGEMA_signal_4837 ;
    wire new_AGEMA_signal_4838 ;
    wire new_AGEMA_signal_4839 ;
    wire new_AGEMA_signal_4840 ;
    wire new_AGEMA_signal_4841 ;
    wire new_AGEMA_signal_4842 ;
    wire new_AGEMA_signal_4843 ;
    wire new_AGEMA_signal_4844 ;
    wire new_AGEMA_signal_4845 ;
    wire new_AGEMA_signal_4846 ;
    wire new_AGEMA_signal_4847 ;
    wire new_AGEMA_signal_4848 ;
    wire new_AGEMA_signal_4849 ;
    wire new_AGEMA_signal_4850 ;
    wire new_AGEMA_signal_4851 ;
    wire new_AGEMA_signal_4852 ;
    wire new_AGEMA_signal_4853 ;
    wire new_AGEMA_signal_4854 ;
    wire new_AGEMA_signal_4855 ;
    wire new_AGEMA_signal_4856 ;
    wire new_AGEMA_signal_4857 ;
    wire new_AGEMA_signal_4858 ;
    wire new_AGEMA_signal_4859 ;
    wire new_AGEMA_signal_4860 ;
    wire new_AGEMA_signal_4861 ;
    wire new_AGEMA_signal_4862 ;
    wire new_AGEMA_signal_4863 ;
    wire new_AGEMA_signal_4864 ;
    wire new_AGEMA_signal_4865 ;
    wire new_AGEMA_signal_4866 ;
    wire new_AGEMA_signal_4867 ;
    wire new_AGEMA_signal_4868 ;
    wire new_AGEMA_signal_4869 ;
    wire new_AGEMA_signal_4870 ;
    wire new_AGEMA_signal_4871 ;
    wire new_AGEMA_signal_4872 ;
    wire new_AGEMA_signal_4873 ;
    wire new_AGEMA_signal_4874 ;
    wire new_AGEMA_signal_4875 ;
    wire new_AGEMA_signal_4876 ;
    wire new_AGEMA_signal_4877 ;
    wire new_AGEMA_signal_4878 ;
    wire new_AGEMA_signal_4879 ;
    wire new_AGEMA_signal_4880 ;
    wire new_AGEMA_signal_4881 ;
    wire new_AGEMA_signal_4882 ;
    wire new_AGEMA_signal_4883 ;
    wire new_AGEMA_signal_4884 ;
    wire new_AGEMA_signal_4885 ;
    wire new_AGEMA_signal_4886 ;
    wire new_AGEMA_signal_4887 ;
    wire new_AGEMA_signal_4888 ;
    wire new_AGEMA_signal_4889 ;
    wire new_AGEMA_signal_4890 ;
    wire new_AGEMA_signal_4891 ;
    wire new_AGEMA_signal_4892 ;
    wire new_AGEMA_signal_4893 ;
    wire new_AGEMA_signal_4894 ;
    wire new_AGEMA_signal_4895 ;
    wire new_AGEMA_signal_4896 ;
    wire new_AGEMA_signal_4897 ;
    wire new_AGEMA_signal_4898 ;
    wire new_AGEMA_signal_4899 ;
    wire new_AGEMA_signal_4900 ;
    wire new_AGEMA_signal_4901 ;
    wire new_AGEMA_signal_4902 ;
    wire new_AGEMA_signal_4903 ;
    wire new_AGEMA_signal_4904 ;
    wire new_AGEMA_signal_4905 ;
    wire new_AGEMA_signal_4906 ;
    wire new_AGEMA_signal_4907 ;
    wire new_AGEMA_signal_4908 ;
    wire new_AGEMA_signal_4909 ;
    wire new_AGEMA_signal_4910 ;
    wire new_AGEMA_signal_4911 ;
    wire new_AGEMA_signal_4912 ;
    wire new_AGEMA_signal_4913 ;
    wire new_AGEMA_signal_4914 ;
    wire new_AGEMA_signal_4915 ;
    wire new_AGEMA_signal_4916 ;
    wire new_AGEMA_signal_4917 ;
    wire new_AGEMA_signal_4918 ;
    wire new_AGEMA_signal_4919 ;
    wire new_AGEMA_signal_4920 ;
    wire new_AGEMA_signal_4921 ;
    wire new_AGEMA_signal_4922 ;
    wire new_AGEMA_signal_4923 ;
    wire new_AGEMA_signal_4924 ;
    wire new_AGEMA_signal_4925 ;
    wire new_AGEMA_signal_4926 ;
    wire new_AGEMA_signal_4927 ;
    wire new_AGEMA_signal_4928 ;
    wire new_AGEMA_signal_4929 ;
    wire new_AGEMA_signal_4930 ;
    wire new_AGEMA_signal_4931 ;
    wire new_AGEMA_signal_4932 ;
    wire new_AGEMA_signal_4933 ;
    wire new_AGEMA_signal_4934 ;
    wire new_AGEMA_signal_4935 ;
    wire new_AGEMA_signal_4936 ;
    wire new_AGEMA_signal_4937 ;
    wire new_AGEMA_signal_4938 ;
    wire new_AGEMA_signal_4939 ;
    wire new_AGEMA_signal_4940 ;
    wire new_AGEMA_signal_4941 ;
    wire new_AGEMA_signal_4942 ;
    wire new_AGEMA_signal_4943 ;
    wire new_AGEMA_signal_4944 ;
    wire new_AGEMA_signal_4945 ;
    wire new_AGEMA_signal_4946 ;
    wire new_AGEMA_signal_4947 ;
    wire new_AGEMA_signal_4948 ;
    wire new_AGEMA_signal_4949 ;
    wire new_AGEMA_signal_4950 ;
    wire new_AGEMA_signal_4951 ;
    wire new_AGEMA_signal_4952 ;
    wire new_AGEMA_signal_4953 ;
    wire new_AGEMA_signal_4954 ;
    wire new_AGEMA_signal_4955 ;
    wire new_AGEMA_signal_4956 ;
    wire new_AGEMA_signal_4957 ;
    wire new_AGEMA_signal_4958 ;
    wire new_AGEMA_signal_4959 ;
    wire new_AGEMA_signal_4960 ;
    wire new_AGEMA_signal_4961 ;
    wire new_AGEMA_signal_4962 ;
    wire new_AGEMA_signal_4963 ;
    wire new_AGEMA_signal_4964 ;
    wire new_AGEMA_signal_4965 ;
    wire new_AGEMA_signal_4966 ;
    wire new_AGEMA_signal_4967 ;
    wire new_AGEMA_signal_4968 ;
    wire new_AGEMA_signal_4969 ;
    wire new_AGEMA_signal_4970 ;
    wire new_AGEMA_signal_4971 ;
    wire new_AGEMA_signal_4972 ;
    wire new_AGEMA_signal_4973 ;
    wire new_AGEMA_signal_4974 ;
    wire new_AGEMA_signal_4975 ;
    wire new_AGEMA_signal_4976 ;
    wire new_AGEMA_signal_4977 ;
    wire new_AGEMA_signal_4978 ;
    wire new_AGEMA_signal_4979 ;
    wire new_AGEMA_signal_4980 ;
    wire new_AGEMA_signal_4981 ;
    wire new_AGEMA_signal_4982 ;
    wire new_AGEMA_signal_4983 ;
    wire new_AGEMA_signal_4984 ;
    wire new_AGEMA_signal_4985 ;
    wire new_AGEMA_signal_4986 ;
    wire new_AGEMA_signal_4987 ;
    wire new_AGEMA_signal_4988 ;
    wire new_AGEMA_signal_4989 ;
    wire new_AGEMA_signal_4990 ;
    wire new_AGEMA_signal_4991 ;
    wire new_AGEMA_signal_4992 ;
    wire new_AGEMA_signal_4993 ;
    wire new_AGEMA_signal_4994 ;
    wire new_AGEMA_signal_4995 ;
    wire new_AGEMA_signal_4996 ;
    wire new_AGEMA_signal_4997 ;
    wire new_AGEMA_signal_4998 ;
    wire new_AGEMA_signal_4999 ;
    wire new_AGEMA_signal_5000 ;
    wire new_AGEMA_signal_5001 ;
    wire new_AGEMA_signal_5002 ;
    wire new_AGEMA_signal_5003 ;
    wire new_AGEMA_signal_5004 ;
    wire new_AGEMA_signal_5005 ;
    wire new_AGEMA_signal_5006 ;
    wire new_AGEMA_signal_5007 ;
    wire new_AGEMA_signal_5008 ;
    wire new_AGEMA_signal_5009 ;
    wire new_AGEMA_signal_5010 ;
    wire new_AGEMA_signal_5011 ;
    wire new_AGEMA_signal_5012 ;
    wire new_AGEMA_signal_5013 ;
    wire new_AGEMA_signal_5014 ;
    wire new_AGEMA_signal_5015 ;
    wire new_AGEMA_signal_5016 ;
    wire new_AGEMA_signal_5017 ;
    wire new_AGEMA_signal_5018 ;
    wire new_AGEMA_signal_5019 ;
    wire new_AGEMA_signal_5020 ;
    wire new_AGEMA_signal_5021 ;
    wire new_AGEMA_signal_5022 ;
    wire new_AGEMA_signal_5023 ;
    wire new_AGEMA_signal_5024 ;
    wire new_AGEMA_signal_5025 ;
    wire new_AGEMA_signal_5026 ;
    wire new_AGEMA_signal_5027 ;
    wire new_AGEMA_signal_5028 ;
    wire new_AGEMA_signal_5029 ;
    wire new_AGEMA_signal_5030 ;
    wire new_AGEMA_signal_5031 ;
    wire new_AGEMA_signal_5032 ;
    wire new_AGEMA_signal_5033 ;
    wire new_AGEMA_signal_5034 ;
    wire new_AGEMA_signal_5035 ;
    wire new_AGEMA_signal_5036 ;
    wire new_AGEMA_signal_5037 ;
    wire new_AGEMA_signal_5038 ;
    wire new_AGEMA_signal_5039 ;
    wire new_AGEMA_signal_5040 ;
    wire new_AGEMA_signal_5041 ;
    wire new_AGEMA_signal_5042 ;
    wire new_AGEMA_signal_5043 ;
    wire new_AGEMA_signal_5044 ;
    wire new_AGEMA_signal_5045 ;
    wire new_AGEMA_signal_5046 ;
    wire new_AGEMA_signal_5047 ;
    wire new_AGEMA_signal_5048 ;
    wire new_AGEMA_signal_5049 ;
    wire new_AGEMA_signal_5050 ;
    wire new_AGEMA_signal_5051 ;
    wire new_AGEMA_signal_5052 ;
    wire new_AGEMA_signal_5053 ;
    wire new_AGEMA_signal_5054 ;
    wire new_AGEMA_signal_5055 ;
    wire new_AGEMA_signal_5056 ;
    wire new_AGEMA_signal_5057 ;
    wire new_AGEMA_signal_5058 ;
    wire new_AGEMA_signal_5059 ;
    wire new_AGEMA_signal_5060 ;
    wire new_AGEMA_signal_5061 ;
    wire new_AGEMA_signal_5062 ;
    wire new_AGEMA_signal_5063 ;
    wire new_AGEMA_signal_5064 ;
    wire new_AGEMA_signal_5065 ;
    wire new_AGEMA_signal_5066 ;
    wire new_AGEMA_signal_5067 ;
    wire new_AGEMA_signal_5068 ;
    wire new_AGEMA_signal_5069 ;
    wire new_AGEMA_signal_5070 ;
    wire new_AGEMA_signal_5071 ;
    wire new_AGEMA_signal_5072 ;
    wire new_AGEMA_signal_5073 ;
    wire new_AGEMA_signal_5074 ;
    wire new_AGEMA_signal_5075 ;
    wire new_AGEMA_signal_5076 ;
    wire new_AGEMA_signal_5077 ;
    wire new_AGEMA_signal_5078 ;
    wire new_AGEMA_signal_5079 ;
    wire new_AGEMA_signal_5080 ;
    wire new_AGEMA_signal_5081 ;
    wire new_AGEMA_signal_5082 ;
    wire new_AGEMA_signal_5083 ;
    wire new_AGEMA_signal_5084 ;
    wire new_AGEMA_signal_5085 ;
    wire new_AGEMA_signal_5086 ;
    wire new_AGEMA_signal_5087 ;
    wire new_AGEMA_signal_5088 ;
    wire new_AGEMA_signal_5089 ;
    wire new_AGEMA_signal_5090 ;
    wire new_AGEMA_signal_5091 ;
    wire new_AGEMA_signal_5092 ;
    wire new_AGEMA_signal_5093 ;
    wire new_AGEMA_signal_5094 ;
    wire new_AGEMA_signal_5095 ;
    wire new_AGEMA_signal_5096 ;
    wire new_AGEMA_signal_5097 ;
    wire new_AGEMA_signal_5098 ;
    wire new_AGEMA_signal_5099 ;
    wire new_AGEMA_signal_5100 ;
    wire new_AGEMA_signal_5101 ;
    wire new_AGEMA_signal_5102 ;
    wire new_AGEMA_signal_5103 ;
    wire new_AGEMA_signal_5104 ;
    wire new_AGEMA_signal_5105 ;
    wire new_AGEMA_signal_5106 ;
    wire new_AGEMA_signal_5107 ;
    wire new_AGEMA_signal_5108 ;
    wire new_AGEMA_signal_5109 ;
    wire new_AGEMA_signal_5110 ;
    wire new_AGEMA_signal_5111 ;
    wire new_AGEMA_signal_5112 ;
    wire new_AGEMA_signal_5113 ;
    wire new_AGEMA_signal_5114 ;
    wire new_AGEMA_signal_5115 ;
    wire new_AGEMA_signal_5116 ;
    wire new_AGEMA_signal_5117 ;
    wire new_AGEMA_signal_5118 ;
    wire new_AGEMA_signal_5119 ;
    wire new_AGEMA_signal_5120 ;
    wire new_AGEMA_signal_5121 ;
    wire new_AGEMA_signal_5122 ;
    wire new_AGEMA_signal_5123 ;
    wire new_AGEMA_signal_5124 ;
    wire new_AGEMA_signal_5125 ;
    wire new_AGEMA_signal_5126 ;
    wire new_AGEMA_signal_5127 ;
    wire new_AGEMA_signal_5128 ;
    wire new_AGEMA_signal_5129 ;
    wire new_AGEMA_signal_5130 ;
    wire new_AGEMA_signal_5131 ;
    wire new_AGEMA_signal_5132 ;
    wire new_AGEMA_signal_5133 ;
    wire new_AGEMA_signal_5134 ;
    wire new_AGEMA_signal_5135 ;
    wire new_AGEMA_signal_5136 ;
    wire new_AGEMA_signal_5137 ;
    wire new_AGEMA_signal_5138 ;
    wire new_AGEMA_signal_5139 ;
    wire new_AGEMA_signal_5140 ;
    wire new_AGEMA_signal_5141 ;
    wire new_AGEMA_signal_5142 ;
    wire new_AGEMA_signal_5143 ;
    wire new_AGEMA_signal_5144 ;
    wire new_AGEMA_signal_5145 ;
    wire new_AGEMA_signal_5146 ;
    wire new_AGEMA_signal_5147 ;
    wire new_AGEMA_signal_5148 ;
    wire new_AGEMA_signal_5149 ;
    wire new_AGEMA_signal_5150 ;
    wire new_AGEMA_signal_5151 ;
    wire new_AGEMA_signal_5152 ;
    wire new_AGEMA_signal_5153 ;
    wire new_AGEMA_signal_5154 ;
    wire new_AGEMA_signal_5155 ;
    wire new_AGEMA_signal_5156 ;
    wire new_AGEMA_signal_5157 ;
    wire new_AGEMA_signal_5158 ;
    wire new_AGEMA_signal_5159 ;
    wire new_AGEMA_signal_5160 ;
    wire new_AGEMA_signal_5161 ;
    wire new_AGEMA_signal_5162 ;
    wire new_AGEMA_signal_5163 ;
    wire new_AGEMA_signal_5164 ;
    wire new_AGEMA_signal_5165 ;
    wire new_AGEMA_signal_5166 ;
    wire new_AGEMA_signal_5167 ;
    wire new_AGEMA_signal_5168 ;
    wire new_AGEMA_signal_5169 ;
    wire new_AGEMA_signal_5170 ;
    wire new_AGEMA_signal_5171 ;
    wire new_AGEMA_signal_5172 ;
    wire new_AGEMA_signal_5173 ;
    wire new_AGEMA_signal_5174 ;
    wire new_AGEMA_signal_5175 ;
    wire new_AGEMA_signal_5176 ;
    wire new_AGEMA_signal_5177 ;
    wire new_AGEMA_signal_5178 ;
    wire new_AGEMA_signal_5179 ;
    wire new_AGEMA_signal_5180 ;
    wire new_AGEMA_signal_5181 ;
    wire new_AGEMA_signal_5182 ;
    wire new_AGEMA_signal_5183 ;
    wire new_AGEMA_signal_5184 ;
    wire new_AGEMA_signal_5185 ;
    wire new_AGEMA_signal_5186 ;
    wire new_AGEMA_signal_5187 ;
    wire new_AGEMA_signal_5188 ;
    wire new_AGEMA_signal_5189 ;
    wire new_AGEMA_signal_5190 ;
    wire new_AGEMA_signal_5191 ;
    wire new_AGEMA_signal_5192 ;
    wire new_AGEMA_signal_5193 ;
    wire new_AGEMA_signal_5194 ;
    wire new_AGEMA_signal_5195 ;
    wire new_AGEMA_signal_5196 ;
    wire new_AGEMA_signal_5197 ;
    wire new_AGEMA_signal_5198 ;
    wire new_AGEMA_signal_5199 ;
    wire new_AGEMA_signal_5200 ;
    wire new_AGEMA_signal_5201 ;
    wire new_AGEMA_signal_5202 ;
    wire new_AGEMA_signal_5203 ;
    wire new_AGEMA_signal_5204 ;
    wire new_AGEMA_signal_5205 ;
    wire new_AGEMA_signal_5206 ;
    wire new_AGEMA_signal_5207 ;
    wire new_AGEMA_signal_5208 ;
    wire new_AGEMA_signal_5209 ;
    wire new_AGEMA_signal_5210 ;
    wire new_AGEMA_signal_5211 ;
    wire new_AGEMA_signal_5212 ;
    wire new_AGEMA_signal_5213 ;
    wire new_AGEMA_signal_5214 ;
    wire new_AGEMA_signal_5215 ;
    wire new_AGEMA_signal_5216 ;
    wire new_AGEMA_signal_5217 ;
    wire new_AGEMA_signal_5218 ;
    wire new_AGEMA_signal_5219 ;
    wire new_AGEMA_signal_5220 ;
    wire new_AGEMA_signal_5221 ;
    wire new_AGEMA_signal_5222 ;
    wire new_AGEMA_signal_5223 ;
    wire new_AGEMA_signal_5224 ;
    wire new_AGEMA_signal_5225 ;
    wire new_AGEMA_signal_5226 ;
    wire new_AGEMA_signal_5227 ;
    wire new_AGEMA_signal_5228 ;
    wire new_AGEMA_signal_5229 ;
    wire new_AGEMA_signal_5230 ;
    wire new_AGEMA_signal_5231 ;
    wire new_AGEMA_signal_5232 ;
    wire new_AGEMA_signal_5233 ;
    wire new_AGEMA_signal_5234 ;
    wire new_AGEMA_signal_5235 ;
    wire new_AGEMA_signal_5236 ;
    wire new_AGEMA_signal_5237 ;
    wire new_AGEMA_signal_5238 ;
    wire new_AGEMA_signal_5239 ;
    wire new_AGEMA_signal_5240 ;
    wire new_AGEMA_signal_5241 ;
    wire new_AGEMA_signal_5242 ;
    wire new_AGEMA_signal_5243 ;
    wire new_AGEMA_signal_5244 ;
    wire new_AGEMA_signal_5245 ;
    wire new_AGEMA_signal_5246 ;
    wire new_AGEMA_signal_5247 ;
    wire new_AGEMA_signal_5248 ;
    wire new_AGEMA_signal_5249 ;
    wire new_AGEMA_signal_5250 ;
    wire new_AGEMA_signal_5251 ;
    wire new_AGEMA_signal_5252 ;
    wire new_AGEMA_signal_5253 ;
    wire new_AGEMA_signal_5254 ;
    wire new_AGEMA_signal_5255 ;
    wire new_AGEMA_signal_5256 ;
    wire new_AGEMA_signal_5257 ;
    wire new_AGEMA_signal_5258 ;
    wire new_AGEMA_signal_5259 ;
    wire new_AGEMA_signal_5260 ;
    wire new_AGEMA_signal_5261 ;
    wire new_AGEMA_signal_5262 ;
    wire new_AGEMA_signal_5263 ;
    wire new_AGEMA_signal_5264 ;
    wire new_AGEMA_signal_5265 ;
    wire new_AGEMA_signal_5266 ;
    wire new_AGEMA_signal_5267 ;
    wire new_AGEMA_signal_5268 ;
    wire new_AGEMA_signal_5269 ;
    wire new_AGEMA_signal_5270 ;
    wire new_AGEMA_signal_5271 ;
    wire new_AGEMA_signal_5272 ;
    wire new_AGEMA_signal_5273 ;
    wire new_AGEMA_signal_5274 ;
    wire new_AGEMA_signal_5275 ;
    wire new_AGEMA_signal_5276 ;
    wire new_AGEMA_signal_5277 ;
    wire new_AGEMA_signal_5278 ;
    wire new_AGEMA_signal_5279 ;
    wire new_AGEMA_signal_5280 ;
    wire new_AGEMA_signal_5281 ;
    wire new_AGEMA_signal_5282 ;
    wire new_AGEMA_signal_5283 ;
    wire new_AGEMA_signal_5284 ;
    wire new_AGEMA_signal_5285 ;
    wire new_AGEMA_signal_5286 ;
    wire new_AGEMA_signal_5287 ;
    wire new_AGEMA_signal_5288 ;
    wire new_AGEMA_signal_5289 ;
    wire new_AGEMA_signal_5290 ;
    wire new_AGEMA_signal_5291 ;
    wire new_AGEMA_signal_5292 ;
    wire new_AGEMA_signal_5293 ;
    wire new_AGEMA_signal_5294 ;
    wire new_AGEMA_signal_5295 ;
    wire new_AGEMA_signal_5296 ;
    wire new_AGEMA_signal_5297 ;
    wire new_AGEMA_signal_5298 ;
    wire new_AGEMA_signal_5299 ;
    wire new_AGEMA_signal_5300 ;
    wire new_AGEMA_signal_5301 ;
    wire new_AGEMA_signal_5302 ;
    wire new_AGEMA_signal_5303 ;
    wire new_AGEMA_signal_5304 ;
    wire new_AGEMA_signal_5305 ;
    wire new_AGEMA_signal_5306 ;
    wire new_AGEMA_signal_5307 ;
    wire new_AGEMA_signal_5308 ;
    wire new_AGEMA_signal_5309 ;
    wire new_AGEMA_signal_5310 ;
    wire new_AGEMA_signal_5311 ;
    wire new_AGEMA_signal_5312 ;
    wire new_AGEMA_signal_5313 ;
    wire new_AGEMA_signal_5314 ;
    wire new_AGEMA_signal_5315 ;
    wire new_AGEMA_signal_5316 ;
    wire new_AGEMA_signal_5317 ;
    wire new_AGEMA_signal_5318 ;
    wire new_AGEMA_signal_5319 ;
    wire new_AGEMA_signal_5320 ;
    wire new_AGEMA_signal_5321 ;
    wire new_AGEMA_signal_5322 ;
    wire new_AGEMA_signal_5323 ;
    wire new_AGEMA_signal_5324 ;
    wire new_AGEMA_signal_5325 ;
    wire new_AGEMA_signal_5326 ;
    wire new_AGEMA_signal_5327 ;
    wire new_AGEMA_signal_5328 ;
    wire new_AGEMA_signal_5329 ;
    wire new_AGEMA_signal_5330 ;
    wire new_AGEMA_signal_5331 ;
    wire new_AGEMA_signal_5332 ;
    wire new_AGEMA_signal_5333 ;
    wire new_AGEMA_signal_5334 ;
    wire new_AGEMA_signal_5335 ;
    wire new_AGEMA_signal_5336 ;
    wire new_AGEMA_signal_5337 ;
    wire new_AGEMA_signal_5338 ;
    wire new_AGEMA_signal_5339 ;
    wire new_AGEMA_signal_5340 ;
    wire new_AGEMA_signal_5341 ;
    wire new_AGEMA_signal_5342 ;
    wire new_AGEMA_signal_5343 ;
    wire new_AGEMA_signal_5344 ;
    wire new_AGEMA_signal_5345 ;
    wire new_AGEMA_signal_5346 ;
    wire new_AGEMA_signal_5347 ;
    wire new_AGEMA_signal_5348 ;
    wire new_AGEMA_signal_5349 ;
    wire new_AGEMA_signal_5350 ;
    wire new_AGEMA_signal_5351 ;
    wire new_AGEMA_signal_5352 ;
    wire new_AGEMA_signal_5353 ;
    wire new_AGEMA_signal_5354 ;
    wire new_AGEMA_signal_5355 ;
    wire new_AGEMA_signal_5356 ;
    wire new_AGEMA_signal_5357 ;
    wire new_AGEMA_signal_5358 ;
    wire new_AGEMA_signal_5359 ;
    wire new_AGEMA_signal_5360 ;
    wire new_AGEMA_signal_5361 ;
    wire new_AGEMA_signal_5362 ;
    wire new_AGEMA_signal_5363 ;
    wire new_AGEMA_signal_5364 ;
    wire new_AGEMA_signal_5365 ;
    wire new_AGEMA_signal_5366 ;
    wire new_AGEMA_signal_5367 ;
    wire new_AGEMA_signal_5368 ;
    wire new_AGEMA_signal_5369 ;
    wire new_AGEMA_signal_5370 ;
    wire new_AGEMA_signal_5371 ;
    wire new_AGEMA_signal_5372 ;
    wire new_AGEMA_signal_5373 ;
    wire new_AGEMA_signal_5374 ;
    wire new_AGEMA_signal_5375 ;
    wire new_AGEMA_signal_5376 ;
    wire new_AGEMA_signal_5377 ;
    wire new_AGEMA_signal_5378 ;
    wire new_AGEMA_signal_5379 ;
    wire new_AGEMA_signal_5380 ;
    wire new_AGEMA_signal_5381 ;
    wire new_AGEMA_signal_5382 ;
    wire new_AGEMA_signal_5383 ;
    wire new_AGEMA_signal_5384 ;
    wire new_AGEMA_signal_5385 ;
    wire new_AGEMA_signal_5386 ;
    wire new_AGEMA_signal_5387 ;
    wire new_AGEMA_signal_5391 ;
    wire new_AGEMA_signal_5392 ;
    wire new_AGEMA_signal_5393 ;
    wire new_AGEMA_signal_5394 ;
    wire new_AGEMA_signal_5395 ;
    wire new_AGEMA_signal_5396 ;
    wire new_AGEMA_signal_5397 ;
    wire new_AGEMA_signal_5398 ;
    wire new_AGEMA_signal_5399 ;
    wire new_AGEMA_signal_5400 ;
    wire new_AGEMA_signal_5401 ;
    wire new_AGEMA_signal_5402 ;
    wire new_AGEMA_signal_5403 ;
    wire new_AGEMA_signal_5404 ;
    wire new_AGEMA_signal_5405 ;
    wire new_AGEMA_signal_5406 ;
    wire new_AGEMA_signal_5407 ;
    wire new_AGEMA_signal_5408 ;
    wire new_AGEMA_signal_5412 ;
    wire new_AGEMA_signal_5413 ;
    wire new_AGEMA_signal_5414 ;
    wire new_AGEMA_signal_5415 ;
    wire new_AGEMA_signal_5416 ;
    wire new_AGEMA_signal_5417 ;
    wire new_AGEMA_signal_5418 ;
    wire new_AGEMA_signal_5419 ;
    wire new_AGEMA_signal_5420 ;
    wire new_AGEMA_signal_5421 ;
    wire new_AGEMA_signal_5422 ;
    wire new_AGEMA_signal_5423 ;
    wire new_AGEMA_signal_5424 ;
    wire new_AGEMA_signal_5425 ;
    wire new_AGEMA_signal_5426 ;
    wire new_AGEMA_signal_5427 ;
    wire new_AGEMA_signal_5428 ;
    wire new_AGEMA_signal_5429 ;
    wire new_AGEMA_signal_5430 ;
    wire new_AGEMA_signal_5431 ;
    wire new_AGEMA_signal_5432 ;
    wire new_AGEMA_signal_5433 ;
    wire new_AGEMA_signal_5434 ;
    wire new_AGEMA_signal_5435 ;
    wire new_AGEMA_signal_5436 ;
    wire new_AGEMA_signal_5437 ;
    wire new_AGEMA_signal_5438 ;
    wire new_AGEMA_signal_5439 ;
    wire new_AGEMA_signal_5440 ;
    wire new_AGEMA_signal_5441 ;
    wire new_AGEMA_signal_5442 ;
    wire new_AGEMA_signal_5443 ;
    wire new_AGEMA_signal_5444 ;
    wire new_AGEMA_signal_5445 ;
    wire new_AGEMA_signal_5446 ;
    wire new_AGEMA_signal_5447 ;
    wire new_AGEMA_signal_5448 ;
    wire new_AGEMA_signal_5449 ;
    wire new_AGEMA_signal_5450 ;
    wire new_AGEMA_signal_5451 ;
    wire new_AGEMA_signal_5452 ;
    wire new_AGEMA_signal_5453 ;
    wire new_AGEMA_signal_5454 ;
    wire new_AGEMA_signal_5455 ;
    wire new_AGEMA_signal_5456 ;
    wire new_AGEMA_signal_5457 ;
    wire new_AGEMA_signal_5458 ;
    wire new_AGEMA_signal_5459 ;
    wire new_AGEMA_signal_5460 ;
    wire new_AGEMA_signal_5461 ;
    wire new_AGEMA_signal_5462 ;
    wire new_AGEMA_signal_5463 ;
    wire new_AGEMA_signal_5464 ;
    wire new_AGEMA_signal_5465 ;
    wire new_AGEMA_signal_5466 ;
    wire new_AGEMA_signal_5467 ;
    wire new_AGEMA_signal_5468 ;
    wire new_AGEMA_signal_5469 ;
    wire new_AGEMA_signal_5470 ;
    wire new_AGEMA_signal_5471 ;
    wire new_AGEMA_signal_5472 ;
    wire new_AGEMA_signal_5473 ;
    wire new_AGEMA_signal_5474 ;
    wire new_AGEMA_signal_5475 ;
    wire new_AGEMA_signal_5476 ;
    wire new_AGEMA_signal_5477 ;
    wire new_AGEMA_signal_5478 ;
    wire new_AGEMA_signal_5479 ;
    wire new_AGEMA_signal_5480 ;
    wire new_AGEMA_signal_5481 ;
    wire new_AGEMA_signal_5482 ;
    wire new_AGEMA_signal_5483 ;
    wire new_AGEMA_signal_5484 ;
    wire new_AGEMA_signal_5485 ;
    wire new_AGEMA_signal_5486 ;
    wire new_AGEMA_signal_5487 ;
    wire new_AGEMA_signal_5488 ;
    wire new_AGEMA_signal_5489 ;
    wire new_AGEMA_signal_5490 ;
    wire new_AGEMA_signal_5491 ;
    wire new_AGEMA_signal_5492 ;
    wire new_AGEMA_signal_5493 ;
    wire new_AGEMA_signal_5494 ;
    wire new_AGEMA_signal_5495 ;
    wire new_AGEMA_signal_5499 ;
    wire new_AGEMA_signal_5500 ;
    wire new_AGEMA_signal_5501 ;
    wire new_AGEMA_signal_5502 ;
    wire new_AGEMA_signal_5503 ;
    wire new_AGEMA_signal_5504 ;
    wire new_AGEMA_signal_5505 ;
    wire new_AGEMA_signal_5506 ;
    wire new_AGEMA_signal_5507 ;
    wire new_AGEMA_signal_5508 ;
    wire new_AGEMA_signal_5509 ;
    wire new_AGEMA_signal_5510 ;
    wire new_AGEMA_signal_5511 ;
    wire new_AGEMA_signal_5512 ;
    wire new_AGEMA_signal_5513 ;
    wire new_AGEMA_signal_5514 ;
    wire new_AGEMA_signal_5515 ;
    wire new_AGEMA_signal_5516 ;
    wire new_AGEMA_signal_5517 ;
    wire new_AGEMA_signal_5518 ;
    wire new_AGEMA_signal_5519 ;
    wire new_AGEMA_signal_5520 ;
    wire new_AGEMA_signal_5521 ;
    wire new_AGEMA_signal_5522 ;
    wire new_AGEMA_signal_5523 ;
    wire new_AGEMA_signal_5524 ;
    wire new_AGEMA_signal_5525 ;
    wire new_AGEMA_signal_5526 ;
    wire new_AGEMA_signal_5527 ;
    wire new_AGEMA_signal_5528 ;
    wire new_AGEMA_signal_5529 ;
    wire new_AGEMA_signal_5530 ;
    wire new_AGEMA_signal_5531 ;
    wire new_AGEMA_signal_5532 ;
    wire new_AGEMA_signal_5533 ;
    wire new_AGEMA_signal_5534 ;
    wire new_AGEMA_signal_5538 ;
    wire new_AGEMA_signal_5539 ;
    wire new_AGEMA_signal_5540 ;
    wire new_AGEMA_signal_5541 ;
    wire new_AGEMA_signal_5542 ;
    wire new_AGEMA_signal_5543 ;
    wire new_AGEMA_signal_5544 ;
    wire new_AGEMA_signal_5545 ;
    wire new_AGEMA_signal_5546 ;
    wire new_AGEMA_signal_5547 ;
    wire new_AGEMA_signal_5548 ;
    wire new_AGEMA_signal_5549 ;
    wire new_AGEMA_signal_5550 ;
    wire new_AGEMA_signal_5551 ;
    wire new_AGEMA_signal_5552 ;
    wire new_AGEMA_signal_5553 ;
    wire new_AGEMA_signal_5554 ;
    wire new_AGEMA_signal_5555 ;
    wire new_AGEMA_signal_5556 ;
    wire new_AGEMA_signal_5557 ;
    wire new_AGEMA_signal_5558 ;
    wire new_AGEMA_signal_5559 ;
    wire new_AGEMA_signal_5560 ;
    wire new_AGEMA_signal_5561 ;
    wire new_AGEMA_signal_5562 ;
    wire new_AGEMA_signal_5563 ;
    wire new_AGEMA_signal_5564 ;
    wire new_AGEMA_signal_5565 ;
    wire new_AGEMA_signal_5566 ;
    wire new_AGEMA_signal_5567 ;
    wire new_AGEMA_signal_5568 ;
    wire new_AGEMA_signal_5569 ;
    wire new_AGEMA_signal_5570 ;
    wire new_AGEMA_signal_5574 ;
    wire new_AGEMA_signal_5575 ;
    wire new_AGEMA_signal_5576 ;
    wire new_AGEMA_signal_5577 ;
    wire new_AGEMA_signal_5578 ;
    wire new_AGEMA_signal_5579 ;
    wire new_AGEMA_signal_5580 ;
    wire new_AGEMA_signal_5581 ;
    wire new_AGEMA_signal_5582 ;
    wire new_AGEMA_signal_5583 ;
    wire new_AGEMA_signal_5584 ;
    wire new_AGEMA_signal_5585 ;
    wire new_AGEMA_signal_5586 ;
    wire new_AGEMA_signal_5587 ;
    wire new_AGEMA_signal_5588 ;
    wire new_AGEMA_signal_5589 ;
    wire new_AGEMA_signal_5590 ;
    wire new_AGEMA_signal_5591 ;
    wire new_AGEMA_signal_5592 ;
    wire new_AGEMA_signal_5593 ;
    wire new_AGEMA_signal_5594 ;
    wire new_AGEMA_signal_5595 ;
    wire new_AGEMA_signal_5596 ;
    wire new_AGEMA_signal_5597 ;
    wire new_AGEMA_signal_5598 ;
    wire new_AGEMA_signal_5599 ;
    wire new_AGEMA_signal_5600 ;
    wire new_AGEMA_signal_5601 ;
    wire new_AGEMA_signal_5602 ;
    wire new_AGEMA_signal_5603 ;
    wire new_AGEMA_signal_5604 ;
    wire new_AGEMA_signal_5605 ;
    wire new_AGEMA_signal_5606 ;
    wire new_AGEMA_signal_5607 ;
    wire new_AGEMA_signal_5608 ;
    wire new_AGEMA_signal_5609 ;
    wire new_AGEMA_signal_5610 ;
    wire new_AGEMA_signal_5611 ;
    wire new_AGEMA_signal_5612 ;
    wire new_AGEMA_signal_5613 ;
    wire new_AGEMA_signal_5614 ;
    wire new_AGEMA_signal_5615 ;
    wire new_AGEMA_signal_5616 ;
    wire new_AGEMA_signal_5617 ;
    wire new_AGEMA_signal_5618 ;
    wire new_AGEMA_signal_5619 ;
    wire new_AGEMA_signal_5620 ;
    wire new_AGEMA_signal_5621 ;
    wire new_AGEMA_signal_5622 ;
    wire new_AGEMA_signal_5623 ;
    wire new_AGEMA_signal_5624 ;
    wire new_AGEMA_signal_5625 ;
    wire new_AGEMA_signal_5626 ;
    wire new_AGEMA_signal_5627 ;
    wire new_AGEMA_signal_5628 ;
    wire new_AGEMA_signal_5629 ;
    wire new_AGEMA_signal_5630 ;
    wire new_AGEMA_signal_5631 ;
    wire new_AGEMA_signal_5632 ;
    wire new_AGEMA_signal_5633 ;
    wire new_AGEMA_signal_5634 ;
    wire new_AGEMA_signal_5635 ;
    wire new_AGEMA_signal_5636 ;
    wire new_AGEMA_signal_5637 ;
    wire new_AGEMA_signal_5638 ;
    wire new_AGEMA_signal_5639 ;
    wire new_AGEMA_signal_5640 ;
    wire new_AGEMA_signal_5641 ;
    wire new_AGEMA_signal_5642 ;
    wire new_AGEMA_signal_5643 ;
    wire new_AGEMA_signal_5644 ;
    wire new_AGEMA_signal_5645 ;
    wire new_AGEMA_signal_5646 ;
    wire new_AGEMA_signal_5647 ;
    wire new_AGEMA_signal_5648 ;
    wire new_AGEMA_signal_5649 ;
    wire new_AGEMA_signal_5650 ;
    wire new_AGEMA_signal_5651 ;
    wire new_AGEMA_signal_5652 ;
    wire new_AGEMA_signal_5653 ;
    wire new_AGEMA_signal_5654 ;
    wire new_AGEMA_signal_5655 ;
    wire new_AGEMA_signal_5656 ;
    wire new_AGEMA_signal_5657 ;
    wire new_AGEMA_signal_5658 ;
    wire new_AGEMA_signal_5659 ;
    wire new_AGEMA_signal_5660 ;
    wire new_AGEMA_signal_5661 ;
    wire new_AGEMA_signal_5662 ;
    wire new_AGEMA_signal_5663 ;
    wire new_AGEMA_signal_5664 ;
    wire new_AGEMA_signal_5665 ;
    wire new_AGEMA_signal_5666 ;
    wire new_AGEMA_signal_5667 ;
    wire new_AGEMA_signal_5668 ;
    wire new_AGEMA_signal_5669 ;
    wire new_AGEMA_signal_5670 ;
    wire new_AGEMA_signal_5671 ;
    wire new_AGEMA_signal_5672 ;
    wire new_AGEMA_signal_5676 ;
    wire new_AGEMA_signal_5677 ;
    wire new_AGEMA_signal_5678 ;
    wire new_AGEMA_signal_5679 ;
    wire new_AGEMA_signal_5680 ;
    wire new_AGEMA_signal_5681 ;
    wire new_AGEMA_signal_5682 ;
    wire new_AGEMA_signal_5683 ;
    wire new_AGEMA_signal_5684 ;
    wire new_AGEMA_signal_5685 ;
    wire new_AGEMA_signal_5686 ;
    wire new_AGEMA_signal_5687 ;
    wire new_AGEMA_signal_5688 ;
    wire new_AGEMA_signal_5689 ;
    wire new_AGEMA_signal_5690 ;
    wire new_AGEMA_signal_5691 ;
    wire new_AGEMA_signal_5692 ;
    wire new_AGEMA_signal_5693 ;
    wire new_AGEMA_signal_5694 ;
    wire new_AGEMA_signal_5695 ;
    wire new_AGEMA_signal_5696 ;
    wire new_AGEMA_signal_5697 ;
    wire new_AGEMA_signal_5698 ;
    wire new_AGEMA_signal_5699 ;
    wire new_AGEMA_signal_5700 ;
    wire new_AGEMA_signal_5701 ;
    wire new_AGEMA_signal_5702 ;
    wire new_AGEMA_signal_5703 ;
    wire new_AGEMA_signal_5704 ;
    wire new_AGEMA_signal_5705 ;
    wire new_AGEMA_signal_5709 ;
    wire new_AGEMA_signal_5710 ;
    wire new_AGEMA_signal_5711 ;
    wire new_AGEMA_signal_5712 ;
    wire new_AGEMA_signal_5713 ;
    wire new_AGEMA_signal_5714 ;
    wire new_AGEMA_signal_5715 ;
    wire new_AGEMA_signal_5716 ;
    wire new_AGEMA_signal_5717 ;
    wire new_AGEMA_signal_5718 ;
    wire new_AGEMA_signal_5719 ;
    wire new_AGEMA_signal_5720 ;
    wire new_AGEMA_signal_5721 ;
    wire new_AGEMA_signal_5722 ;
    wire new_AGEMA_signal_5723 ;
    wire new_AGEMA_signal_5724 ;
    wire new_AGEMA_signal_5725 ;
    wire new_AGEMA_signal_5726 ;
    wire new_AGEMA_signal_5727 ;
    wire new_AGEMA_signal_5728 ;
    wire new_AGEMA_signal_5729 ;
    wire new_AGEMA_signal_5730 ;
    wire new_AGEMA_signal_5731 ;
    wire new_AGEMA_signal_5732 ;
    wire new_AGEMA_signal_5733 ;
    wire new_AGEMA_signal_5734 ;
    wire new_AGEMA_signal_5735 ;
    wire new_AGEMA_signal_5739 ;
    wire new_AGEMA_signal_5740 ;
    wire new_AGEMA_signal_5741 ;
    wire new_AGEMA_signal_5742 ;
    wire new_AGEMA_signal_5743 ;
    wire new_AGEMA_signal_5744 ;
    wire new_AGEMA_signal_5745 ;
    wire new_AGEMA_signal_5746 ;
    wire new_AGEMA_signal_5747 ;
    wire new_AGEMA_signal_5748 ;
    wire new_AGEMA_signal_5749 ;
    wire new_AGEMA_signal_5750 ;
    wire new_AGEMA_signal_5751 ;
    wire new_AGEMA_signal_5752 ;
    wire new_AGEMA_signal_5753 ;
    wire new_AGEMA_signal_5754 ;
    wire new_AGEMA_signal_5755 ;
    wire new_AGEMA_signal_5756 ;
    wire new_AGEMA_signal_5757 ;
    wire new_AGEMA_signal_5758 ;
    wire new_AGEMA_signal_5759 ;
    wire new_AGEMA_signal_5760 ;
    wire new_AGEMA_signal_5761 ;
    wire new_AGEMA_signal_5762 ;
    wire new_AGEMA_signal_5763 ;
    wire new_AGEMA_signal_5764 ;
    wire new_AGEMA_signal_5765 ;
    wire new_AGEMA_signal_5766 ;
    wire new_AGEMA_signal_5767 ;
    wire new_AGEMA_signal_5768 ;
    wire new_AGEMA_signal_5769 ;
    wire new_AGEMA_signal_5770 ;
    wire new_AGEMA_signal_5771 ;
    wire new_AGEMA_signal_5772 ;
    wire new_AGEMA_signal_5773 ;
    wire new_AGEMA_signal_5774 ;
    wire new_AGEMA_signal_5775 ;
    wire new_AGEMA_signal_5776 ;
    wire new_AGEMA_signal_5777 ;
    wire new_AGEMA_signal_5778 ;
    wire new_AGEMA_signal_5779 ;
    wire new_AGEMA_signal_5780 ;
    wire new_AGEMA_signal_5781 ;
    wire new_AGEMA_signal_5782 ;
    wire new_AGEMA_signal_5783 ;
    wire new_AGEMA_signal_5784 ;
    wire new_AGEMA_signal_5785 ;
    wire new_AGEMA_signal_5786 ;
    wire new_AGEMA_signal_5787 ;
    wire new_AGEMA_signal_5788 ;
    wire new_AGEMA_signal_5789 ;
    wire new_AGEMA_signal_5790 ;
    wire new_AGEMA_signal_5791 ;
    wire new_AGEMA_signal_5792 ;
    wire new_AGEMA_signal_5793 ;
    wire new_AGEMA_signal_5794 ;
    wire new_AGEMA_signal_5795 ;
    wire new_AGEMA_signal_5796 ;
    wire new_AGEMA_signal_5797 ;
    wire new_AGEMA_signal_5798 ;
    wire new_AGEMA_signal_5799 ;
    wire new_AGEMA_signal_5800 ;
    wire new_AGEMA_signal_5801 ;
    wire new_AGEMA_signal_5802 ;
    wire new_AGEMA_signal_5803 ;
    wire new_AGEMA_signal_5804 ;
    wire new_AGEMA_signal_5805 ;
    wire new_AGEMA_signal_5806 ;
    wire new_AGEMA_signal_5807 ;
    wire new_AGEMA_signal_5808 ;
    wire new_AGEMA_signal_5809 ;
    wire new_AGEMA_signal_5810 ;
    wire new_AGEMA_signal_5811 ;
    wire new_AGEMA_signal_5812 ;
    wire new_AGEMA_signal_5813 ;
    wire new_AGEMA_signal_5814 ;
    wire new_AGEMA_signal_5815 ;
    wire new_AGEMA_signal_5816 ;
    wire new_AGEMA_signal_5817 ;
    wire new_AGEMA_signal_5818 ;
    wire new_AGEMA_signal_5819 ;
    wire new_AGEMA_signal_5820 ;
    wire new_AGEMA_signal_5821 ;
    wire new_AGEMA_signal_5822 ;
    wire new_AGEMA_signal_5823 ;
    wire new_AGEMA_signal_5824 ;
    wire new_AGEMA_signal_5825 ;
    wire new_AGEMA_signal_5826 ;
    wire new_AGEMA_signal_5827 ;
    wire new_AGEMA_signal_5828 ;
    wire new_AGEMA_signal_5829 ;
    wire new_AGEMA_signal_5830 ;
    wire new_AGEMA_signal_5831 ;
    wire new_AGEMA_signal_5832 ;
    wire new_AGEMA_signal_5833 ;
    wire new_AGEMA_signal_5834 ;
    wire new_AGEMA_signal_5835 ;
    wire new_AGEMA_signal_5836 ;
    wire new_AGEMA_signal_5837 ;
    wire new_AGEMA_signal_5838 ;
    wire new_AGEMA_signal_5839 ;
    wire new_AGEMA_signal_5840 ;
    wire new_AGEMA_signal_5841 ;
    wire new_AGEMA_signal_5842 ;
    wire new_AGEMA_signal_5843 ;
    wire new_AGEMA_signal_5844 ;
    wire new_AGEMA_signal_5845 ;
    wire new_AGEMA_signal_5846 ;
    wire new_AGEMA_signal_5847 ;
    wire new_AGEMA_signal_5848 ;
    wire new_AGEMA_signal_5849 ;
    wire new_AGEMA_signal_5850 ;
    wire new_AGEMA_signal_5851 ;
    wire new_AGEMA_signal_5852 ;
    wire new_AGEMA_signal_5853 ;
    wire new_AGEMA_signal_5854 ;
    wire new_AGEMA_signal_5855 ;
    wire new_AGEMA_signal_5856 ;
    wire new_AGEMA_signal_5857 ;
    wire new_AGEMA_signal_5858 ;
    wire new_AGEMA_signal_5859 ;
    wire new_AGEMA_signal_5860 ;
    wire new_AGEMA_signal_5861 ;
    wire new_AGEMA_signal_5862 ;
    wire new_AGEMA_signal_5863 ;
    wire new_AGEMA_signal_5864 ;
    wire new_AGEMA_signal_5865 ;
    wire new_AGEMA_signal_5866 ;
    wire new_AGEMA_signal_5867 ;
    wire new_AGEMA_signal_5868 ;
    wire new_AGEMA_signal_5869 ;
    wire new_AGEMA_signal_5870 ;
    wire new_AGEMA_signal_5871 ;
    wire new_AGEMA_signal_5872 ;
    wire new_AGEMA_signal_5873 ;
    wire new_AGEMA_signal_5874 ;
    wire new_AGEMA_signal_5875 ;
    wire new_AGEMA_signal_5876 ;
    wire new_AGEMA_signal_5877 ;
    wire new_AGEMA_signal_5878 ;
    wire new_AGEMA_signal_5879 ;
    wire new_AGEMA_signal_5880 ;
    wire new_AGEMA_signal_5881 ;
    wire new_AGEMA_signal_5882 ;
    wire new_AGEMA_signal_5883 ;
    wire new_AGEMA_signal_5884 ;
    wire new_AGEMA_signal_5885 ;
    wire new_AGEMA_signal_5886 ;
    wire new_AGEMA_signal_5887 ;
    wire new_AGEMA_signal_5888 ;
    wire new_AGEMA_signal_5889 ;
    wire new_AGEMA_signal_5890 ;
    wire new_AGEMA_signal_5891 ;
    wire new_AGEMA_signal_5892 ;
    wire new_AGEMA_signal_5893 ;
    wire new_AGEMA_signal_5894 ;
    wire new_AGEMA_signal_5895 ;
    wire new_AGEMA_signal_5896 ;
    wire new_AGEMA_signal_5897 ;
    wire new_AGEMA_signal_5898 ;
    wire new_AGEMA_signal_5899 ;
    wire new_AGEMA_signal_5900 ;
    wire new_AGEMA_signal_5901 ;
    wire new_AGEMA_signal_5902 ;
    wire new_AGEMA_signal_5903 ;
    wire new_AGEMA_signal_5904 ;
    wire new_AGEMA_signal_5905 ;
    wire new_AGEMA_signal_5906 ;
    wire new_AGEMA_signal_5907 ;
    wire new_AGEMA_signal_5908 ;
    wire new_AGEMA_signal_5909 ;
    wire new_AGEMA_signal_5910 ;
    wire new_AGEMA_signal_5911 ;
    wire new_AGEMA_signal_5912 ;
    wire new_AGEMA_signal_5913 ;
    wire new_AGEMA_signal_5914 ;
    wire new_AGEMA_signal_5915 ;
    wire new_AGEMA_signal_5916 ;
    wire new_AGEMA_signal_5917 ;
    wire new_AGEMA_signal_5918 ;
    wire new_AGEMA_signal_5919 ;
    wire new_AGEMA_signal_5920 ;
    wire new_AGEMA_signal_5921 ;
    wire new_AGEMA_signal_5922 ;
    wire new_AGEMA_signal_5923 ;
    wire new_AGEMA_signal_5924 ;
    wire new_AGEMA_signal_5925 ;
    wire new_AGEMA_signal_5926 ;
    wire new_AGEMA_signal_5927 ;
    wire new_AGEMA_signal_5928 ;
    wire new_AGEMA_signal_5929 ;
    wire new_AGEMA_signal_5930 ;
    wire new_AGEMA_signal_5931 ;
    wire new_AGEMA_signal_5932 ;
    wire new_AGEMA_signal_5933 ;
    wire new_AGEMA_signal_5934 ;
    wire new_AGEMA_signal_5935 ;
    wire new_AGEMA_signal_5936 ;
    wire new_AGEMA_signal_5937 ;
    wire new_AGEMA_signal_5938 ;
    wire new_AGEMA_signal_5939 ;
    wire new_AGEMA_signal_5940 ;
    wire new_AGEMA_signal_5941 ;
    wire new_AGEMA_signal_5942 ;
    wire new_AGEMA_signal_5943 ;
    wire new_AGEMA_signal_5944 ;
    wire new_AGEMA_signal_5945 ;
    wire new_AGEMA_signal_5946 ;
    wire new_AGEMA_signal_5947 ;
    wire new_AGEMA_signal_5948 ;
    wire new_AGEMA_signal_5949 ;
    wire new_AGEMA_signal_5950 ;
    wire new_AGEMA_signal_5951 ;
    wire new_AGEMA_signal_5952 ;
    wire new_AGEMA_signal_5953 ;
    wire new_AGEMA_signal_5954 ;
    wire new_AGEMA_signal_5955 ;
    wire new_AGEMA_signal_5956 ;
    wire new_AGEMA_signal_5957 ;
    wire new_AGEMA_signal_5958 ;
    wire new_AGEMA_signal_5959 ;
    wire new_AGEMA_signal_5960 ;
    wire new_AGEMA_signal_5961 ;
    wire new_AGEMA_signal_5962 ;
    wire new_AGEMA_signal_5963 ;
    wire new_AGEMA_signal_5964 ;
    wire new_AGEMA_signal_5965 ;
    wire new_AGEMA_signal_5966 ;
    wire new_AGEMA_signal_5967 ;
    wire new_AGEMA_signal_5968 ;
    wire new_AGEMA_signal_5969 ;
    wire new_AGEMA_signal_5970 ;
    wire new_AGEMA_signal_5971 ;
    wire new_AGEMA_signal_5972 ;
    wire new_AGEMA_signal_5973 ;
    wire new_AGEMA_signal_5974 ;
    wire new_AGEMA_signal_5975 ;
    wire new_AGEMA_signal_5976 ;
    wire new_AGEMA_signal_5977 ;
    wire new_AGEMA_signal_5978 ;
    wire new_AGEMA_signal_5979 ;
    wire new_AGEMA_signal_5980 ;
    wire new_AGEMA_signal_5981 ;
    wire new_AGEMA_signal_5982 ;
    wire new_AGEMA_signal_5983 ;
    wire new_AGEMA_signal_5984 ;
    wire new_AGEMA_signal_5985 ;
    wire new_AGEMA_signal_5986 ;
    wire new_AGEMA_signal_5987 ;
    wire new_AGEMA_signal_5988 ;
    wire new_AGEMA_signal_5989 ;
    wire new_AGEMA_signal_5990 ;
    wire new_AGEMA_signal_5991 ;
    wire new_AGEMA_signal_5992 ;
    wire new_AGEMA_signal_5993 ;
    wire new_AGEMA_signal_5994 ;
    wire new_AGEMA_signal_5995 ;
    wire new_AGEMA_signal_5996 ;
    wire new_AGEMA_signal_5997 ;
    wire new_AGEMA_signal_5998 ;
    wire new_AGEMA_signal_5999 ;
    wire new_AGEMA_signal_6000 ;
    wire new_AGEMA_signal_6001 ;
    wire new_AGEMA_signal_6002 ;
    wire new_AGEMA_signal_6003 ;
    wire new_AGEMA_signal_6004 ;
    wire new_AGEMA_signal_6005 ;
    wire new_AGEMA_signal_6006 ;
    wire new_AGEMA_signal_6007 ;
    wire new_AGEMA_signal_6008 ;
    wire new_AGEMA_signal_6009 ;
    wire new_AGEMA_signal_6010 ;
    wire new_AGEMA_signal_6011 ;
    wire new_AGEMA_signal_6012 ;
    wire new_AGEMA_signal_6013 ;
    wire new_AGEMA_signal_6014 ;
    wire new_AGEMA_signal_6015 ;
    wire new_AGEMA_signal_6016 ;
    wire new_AGEMA_signal_6017 ;
    wire new_AGEMA_signal_6018 ;
    wire new_AGEMA_signal_6019 ;
    wire new_AGEMA_signal_6020 ;
    wire new_AGEMA_signal_6021 ;
    wire new_AGEMA_signal_6022 ;
    wire new_AGEMA_signal_6023 ;
    wire new_AGEMA_signal_6024 ;
    wire new_AGEMA_signal_6025 ;
    wire new_AGEMA_signal_6026 ;
    wire new_AGEMA_signal_6027 ;
    wire new_AGEMA_signal_6028 ;
    wire new_AGEMA_signal_6029 ;
    wire new_AGEMA_signal_6030 ;
    wire new_AGEMA_signal_6031 ;
    wire new_AGEMA_signal_6032 ;
    wire new_AGEMA_signal_6033 ;
    wire new_AGEMA_signal_6034 ;
    wire new_AGEMA_signal_6035 ;
    wire new_AGEMA_signal_6036 ;
    wire new_AGEMA_signal_6037 ;
    wire new_AGEMA_signal_6038 ;
    wire new_AGEMA_signal_6039 ;
    wire new_AGEMA_signal_6040 ;
    wire new_AGEMA_signal_6041 ;
    wire new_AGEMA_signal_6042 ;
    wire new_AGEMA_signal_6043 ;
    wire new_AGEMA_signal_6044 ;
    wire new_AGEMA_signal_6045 ;
    wire new_AGEMA_signal_6046 ;
    wire new_AGEMA_signal_6047 ;
    wire new_AGEMA_signal_6048 ;
    wire new_AGEMA_signal_6049 ;
    wire new_AGEMA_signal_6050 ;
    wire new_AGEMA_signal_6051 ;
    wire new_AGEMA_signal_6052 ;
    wire new_AGEMA_signal_6053 ;
    wire new_AGEMA_signal_6054 ;
    wire new_AGEMA_signal_6055 ;
    wire new_AGEMA_signal_6056 ;
    wire new_AGEMA_signal_6057 ;
    wire new_AGEMA_signal_6058 ;
    wire new_AGEMA_signal_6059 ;
    wire new_AGEMA_signal_6060 ;
    wire new_AGEMA_signal_6061 ;
    wire new_AGEMA_signal_6062 ;
    wire new_AGEMA_signal_6063 ;
    wire new_AGEMA_signal_6064 ;
    wire new_AGEMA_signal_6065 ;
    wire new_AGEMA_signal_6066 ;
    wire new_AGEMA_signal_6067 ;
    wire new_AGEMA_signal_6068 ;
    wire new_AGEMA_signal_6069 ;
    wire new_AGEMA_signal_6070 ;
    wire new_AGEMA_signal_6071 ;
    wire new_AGEMA_signal_6072 ;
    wire new_AGEMA_signal_6073 ;
    wire new_AGEMA_signal_6074 ;
    wire new_AGEMA_signal_6075 ;
    wire new_AGEMA_signal_6076 ;
    wire new_AGEMA_signal_6077 ;
    wire new_AGEMA_signal_6078 ;
    wire new_AGEMA_signal_6079 ;
    wire new_AGEMA_signal_6080 ;
    wire new_AGEMA_signal_6081 ;
    wire new_AGEMA_signal_6082 ;
    wire new_AGEMA_signal_6083 ;
    wire new_AGEMA_signal_6084 ;
    wire new_AGEMA_signal_6085 ;
    wire new_AGEMA_signal_6086 ;
    wire new_AGEMA_signal_6087 ;
    wire new_AGEMA_signal_6088 ;
    wire new_AGEMA_signal_6089 ;
    wire new_AGEMA_signal_6090 ;
    wire new_AGEMA_signal_6091 ;
    wire new_AGEMA_signal_6092 ;
    wire new_AGEMA_signal_6093 ;
    wire new_AGEMA_signal_6094 ;
    wire new_AGEMA_signal_6095 ;
    wire new_AGEMA_signal_6096 ;
    wire new_AGEMA_signal_6097 ;
    wire new_AGEMA_signal_6098 ;
    wire new_AGEMA_signal_6099 ;
    wire new_AGEMA_signal_6100 ;
    wire new_AGEMA_signal_6101 ;
    wire new_AGEMA_signal_6102 ;
    wire new_AGEMA_signal_6103 ;
    wire new_AGEMA_signal_6104 ;
    wire new_AGEMA_signal_6105 ;
    wire new_AGEMA_signal_6106 ;
    wire new_AGEMA_signal_6107 ;
    wire new_AGEMA_signal_6108 ;
    wire new_AGEMA_signal_6109 ;
    wire new_AGEMA_signal_6110 ;
    wire new_AGEMA_signal_6111 ;
    wire new_AGEMA_signal_6112 ;
    wire new_AGEMA_signal_6113 ;
    wire new_AGEMA_signal_6114 ;
    wire new_AGEMA_signal_6115 ;
    wire new_AGEMA_signal_6116 ;
    wire new_AGEMA_signal_6117 ;
    wire new_AGEMA_signal_6118 ;
    wire new_AGEMA_signal_6119 ;
    wire new_AGEMA_signal_6120 ;
    wire new_AGEMA_signal_6121 ;
    wire new_AGEMA_signal_6122 ;
    wire new_AGEMA_signal_6123 ;
    wire new_AGEMA_signal_6124 ;
    wire new_AGEMA_signal_6125 ;
    wire new_AGEMA_signal_6126 ;
    wire new_AGEMA_signal_6127 ;
    wire new_AGEMA_signal_6128 ;
    wire new_AGEMA_signal_6129 ;
    wire new_AGEMA_signal_6130 ;
    wire new_AGEMA_signal_6131 ;
    wire new_AGEMA_signal_6132 ;
    wire new_AGEMA_signal_6133 ;
    wire new_AGEMA_signal_6134 ;
    wire new_AGEMA_signal_6135 ;
    wire new_AGEMA_signal_6136 ;
    wire new_AGEMA_signal_6137 ;
    wire new_AGEMA_signal_6138 ;
    wire new_AGEMA_signal_6139 ;
    wire new_AGEMA_signal_6140 ;
    wire new_AGEMA_signal_6141 ;
    wire new_AGEMA_signal_6142 ;
    wire new_AGEMA_signal_6143 ;
    wire new_AGEMA_signal_6144 ;
    wire new_AGEMA_signal_6145 ;
    wire new_AGEMA_signal_6146 ;
    wire new_AGEMA_signal_6147 ;
    wire new_AGEMA_signal_6148 ;
    wire new_AGEMA_signal_6149 ;
    wire new_AGEMA_signal_6150 ;
    wire new_AGEMA_signal_6151 ;
    wire new_AGEMA_signal_6152 ;
    wire new_AGEMA_signal_6153 ;
    wire new_AGEMA_signal_6154 ;
    wire new_AGEMA_signal_6155 ;
    wire new_AGEMA_signal_6156 ;
    wire new_AGEMA_signal_6157 ;
    wire new_AGEMA_signal_6158 ;
    wire new_AGEMA_signal_6159 ;
    wire new_AGEMA_signal_6160 ;
    wire new_AGEMA_signal_6161 ;
    wire new_AGEMA_signal_6162 ;
    wire new_AGEMA_signal_6163 ;
    wire new_AGEMA_signal_6164 ;
    wire new_AGEMA_signal_6165 ;
    wire new_AGEMA_signal_6166 ;
    wire new_AGEMA_signal_6167 ;
    wire new_AGEMA_signal_6168 ;
    wire new_AGEMA_signal_6169 ;
    wire new_AGEMA_signal_6170 ;
    wire new_AGEMA_signal_6171 ;
    wire new_AGEMA_signal_6172 ;
    wire new_AGEMA_signal_6173 ;
    wire new_AGEMA_signal_6174 ;
    wire new_AGEMA_signal_6175 ;
    wire new_AGEMA_signal_6176 ;
    wire new_AGEMA_signal_6177 ;
    wire new_AGEMA_signal_6178 ;
    wire new_AGEMA_signal_6179 ;
    wire new_AGEMA_signal_6180 ;
    wire new_AGEMA_signal_6181 ;
    wire new_AGEMA_signal_6182 ;
    wire new_AGEMA_signal_6183 ;
    wire new_AGEMA_signal_6184 ;
    wire new_AGEMA_signal_6185 ;
    wire new_AGEMA_signal_6186 ;
    wire new_AGEMA_signal_6187 ;
    wire new_AGEMA_signal_6188 ;
    wire new_AGEMA_signal_6189 ;
    wire new_AGEMA_signal_6190 ;
    wire new_AGEMA_signal_6191 ;
    wire new_AGEMA_signal_6192 ;
    wire new_AGEMA_signal_6193 ;
    wire new_AGEMA_signal_6194 ;
    wire new_AGEMA_signal_6195 ;
    wire new_AGEMA_signal_6196 ;
    wire new_AGEMA_signal_6197 ;
    wire new_AGEMA_signal_6198 ;
    wire new_AGEMA_signal_6199 ;
    wire new_AGEMA_signal_6200 ;
    wire new_AGEMA_signal_6201 ;
    wire new_AGEMA_signal_6202 ;
    wire new_AGEMA_signal_6203 ;
    wire new_AGEMA_signal_6204 ;
    wire new_AGEMA_signal_6205 ;
    wire new_AGEMA_signal_6206 ;
    wire new_AGEMA_signal_6207 ;
    wire new_AGEMA_signal_6208 ;
    wire new_AGEMA_signal_6209 ;
    wire new_AGEMA_signal_6210 ;
    wire new_AGEMA_signal_6211 ;
    wire new_AGEMA_signal_6212 ;
    wire new_AGEMA_signal_6213 ;
    wire new_AGEMA_signal_6214 ;
    wire new_AGEMA_signal_6215 ;
    wire new_AGEMA_signal_6216 ;
    wire new_AGEMA_signal_6217 ;
    wire new_AGEMA_signal_6218 ;
    wire new_AGEMA_signal_6219 ;
    wire new_AGEMA_signal_6220 ;
    wire new_AGEMA_signal_6221 ;
    wire new_AGEMA_signal_6222 ;
    wire new_AGEMA_signal_6223 ;
    wire new_AGEMA_signal_6224 ;
    wire new_AGEMA_signal_6225 ;
    wire new_AGEMA_signal_6226 ;
    wire new_AGEMA_signal_6227 ;
    wire new_AGEMA_signal_6228 ;
    wire new_AGEMA_signal_6229 ;
    wire new_AGEMA_signal_6230 ;
    wire new_AGEMA_signal_6231 ;
    wire new_AGEMA_signal_6232 ;
    wire new_AGEMA_signal_6233 ;
    wire new_AGEMA_signal_6234 ;
    wire new_AGEMA_signal_6235 ;
    wire new_AGEMA_signal_6236 ;
    wire new_AGEMA_signal_6237 ;
    wire new_AGEMA_signal_6238 ;
    wire new_AGEMA_signal_6239 ;
    wire new_AGEMA_signal_6240 ;
    wire new_AGEMA_signal_6241 ;
    wire new_AGEMA_signal_6242 ;
    wire new_AGEMA_signal_6243 ;
    wire new_AGEMA_signal_6244 ;
    wire new_AGEMA_signal_6245 ;
    wire new_AGEMA_signal_6246 ;
    wire new_AGEMA_signal_6247 ;
    wire new_AGEMA_signal_6248 ;
    wire new_AGEMA_signal_6249 ;
    wire new_AGEMA_signal_6250 ;
    wire new_AGEMA_signal_6251 ;
    wire new_AGEMA_signal_6252 ;
    wire new_AGEMA_signal_6253 ;
    wire new_AGEMA_signal_6254 ;
    wire new_AGEMA_signal_6255 ;
    wire new_AGEMA_signal_6256 ;
    wire new_AGEMA_signal_6257 ;
    wire new_AGEMA_signal_6258 ;
    wire new_AGEMA_signal_6259 ;
    wire new_AGEMA_signal_6260 ;
    wire new_AGEMA_signal_6261 ;
    wire new_AGEMA_signal_6262 ;
    wire new_AGEMA_signal_6263 ;
    wire new_AGEMA_signal_6264 ;
    wire new_AGEMA_signal_6265 ;
    wire new_AGEMA_signal_6266 ;
    wire new_AGEMA_signal_6267 ;
    wire new_AGEMA_signal_6268 ;
    wire new_AGEMA_signal_6269 ;
    wire new_AGEMA_signal_6270 ;
    wire new_AGEMA_signal_6271 ;
    wire new_AGEMA_signal_6272 ;
    wire new_AGEMA_signal_6273 ;
    wire new_AGEMA_signal_6274 ;
    wire new_AGEMA_signal_6275 ;
    wire new_AGEMA_signal_6276 ;
    wire new_AGEMA_signal_6277 ;
    wire new_AGEMA_signal_6278 ;
    wire new_AGEMA_signal_6279 ;
    wire new_AGEMA_signal_6280 ;
    wire new_AGEMA_signal_6281 ;
    wire new_AGEMA_signal_6282 ;
    wire new_AGEMA_signal_6283 ;
    wire new_AGEMA_signal_6284 ;
    wire new_AGEMA_signal_6285 ;
    wire new_AGEMA_signal_6286 ;
    wire new_AGEMA_signal_6287 ;
    wire new_AGEMA_signal_6288 ;
    wire new_AGEMA_signal_6289 ;
    wire new_AGEMA_signal_6290 ;
    wire new_AGEMA_signal_6291 ;
    wire new_AGEMA_signal_6292 ;
    wire new_AGEMA_signal_6293 ;
    wire new_AGEMA_signal_6294 ;
    wire new_AGEMA_signal_6295 ;
    wire new_AGEMA_signal_6296 ;
    wire new_AGEMA_signal_6297 ;
    wire new_AGEMA_signal_6298 ;
    wire new_AGEMA_signal_6299 ;
    wire new_AGEMA_signal_6300 ;
    wire new_AGEMA_signal_6301 ;
    wire new_AGEMA_signal_6302 ;
    wire new_AGEMA_signal_6303 ;
    wire new_AGEMA_signal_6304 ;
    wire new_AGEMA_signal_6305 ;
    wire new_AGEMA_signal_6306 ;
    wire new_AGEMA_signal_6307 ;
    wire new_AGEMA_signal_6308 ;
    wire new_AGEMA_signal_6309 ;
    wire new_AGEMA_signal_6310 ;
    wire new_AGEMA_signal_6311 ;
    wire new_AGEMA_signal_6312 ;
    wire new_AGEMA_signal_6313 ;
    wire new_AGEMA_signal_6314 ;
    wire new_AGEMA_signal_6315 ;
    wire new_AGEMA_signal_6316 ;
    wire new_AGEMA_signal_6317 ;
    wire new_AGEMA_signal_6318 ;
    wire new_AGEMA_signal_6319 ;
    wire new_AGEMA_signal_6320 ;
    wire new_AGEMA_signal_6321 ;
    wire new_AGEMA_signal_6322 ;
    wire new_AGEMA_signal_6323 ;
    wire new_AGEMA_signal_6324 ;
    wire new_AGEMA_signal_6325 ;
    wire new_AGEMA_signal_6326 ;
    wire new_AGEMA_signal_6327 ;
    wire new_AGEMA_signal_6328 ;
    wire new_AGEMA_signal_6329 ;
    wire new_AGEMA_signal_6330 ;
    wire new_AGEMA_signal_6331 ;
    wire new_AGEMA_signal_6332 ;
    wire new_AGEMA_signal_6333 ;
    wire new_AGEMA_signal_6334 ;
    wire new_AGEMA_signal_6335 ;
    wire new_AGEMA_signal_6336 ;
    wire new_AGEMA_signal_6337 ;
    wire new_AGEMA_signal_6338 ;
    wire new_AGEMA_signal_6339 ;
    wire new_AGEMA_signal_6340 ;
    wire new_AGEMA_signal_6341 ;
    wire new_AGEMA_signal_6342 ;
    wire new_AGEMA_signal_6343 ;
    wire new_AGEMA_signal_6344 ;
    wire new_AGEMA_signal_6345 ;
    wire new_AGEMA_signal_6346 ;
    wire new_AGEMA_signal_6347 ;
    wire new_AGEMA_signal_6348 ;
    wire new_AGEMA_signal_6349 ;
    wire new_AGEMA_signal_6350 ;
    wire new_AGEMA_signal_6351 ;
    wire new_AGEMA_signal_6352 ;
    wire new_AGEMA_signal_6353 ;
    wire new_AGEMA_signal_6354 ;
    wire new_AGEMA_signal_6355 ;
    wire new_AGEMA_signal_6356 ;
    wire new_AGEMA_signal_6357 ;
    wire new_AGEMA_signal_6358 ;
    wire new_AGEMA_signal_6359 ;
    wire new_AGEMA_signal_6360 ;
    wire new_AGEMA_signal_6361 ;
    wire new_AGEMA_signal_6362 ;
    wire new_AGEMA_signal_6363 ;
    wire new_AGEMA_signal_6364 ;
    wire new_AGEMA_signal_6365 ;
    wire new_AGEMA_signal_6366 ;
    wire new_AGEMA_signal_6367 ;
    wire new_AGEMA_signal_6368 ;
    wire new_AGEMA_signal_6369 ;
    wire new_AGEMA_signal_6370 ;
    wire new_AGEMA_signal_6371 ;
    wire new_AGEMA_signal_6372 ;
    wire new_AGEMA_signal_6373 ;
    wire new_AGEMA_signal_6374 ;
    wire new_AGEMA_signal_6375 ;
    wire new_AGEMA_signal_6376 ;
    wire new_AGEMA_signal_6377 ;
    wire new_AGEMA_signal_6378 ;
    wire new_AGEMA_signal_6379 ;
    wire new_AGEMA_signal_6380 ;
    wire new_AGEMA_signal_6381 ;
    wire new_AGEMA_signal_6382 ;
    wire new_AGEMA_signal_6383 ;
    wire new_AGEMA_signal_6384 ;
    wire new_AGEMA_signal_6385 ;
    wire new_AGEMA_signal_6386 ;
    wire new_AGEMA_signal_6387 ;
    wire new_AGEMA_signal_6388 ;
    wire new_AGEMA_signal_6389 ;
    wire new_AGEMA_signal_6390 ;
    wire new_AGEMA_signal_6391 ;
    wire new_AGEMA_signal_6392 ;
    wire new_AGEMA_signal_6393 ;
    wire new_AGEMA_signal_6394 ;
    wire new_AGEMA_signal_6395 ;
    wire new_AGEMA_signal_6396 ;
    wire new_AGEMA_signal_6397 ;
    wire new_AGEMA_signal_6398 ;
    wire new_AGEMA_signal_6399 ;
    wire new_AGEMA_signal_6400 ;
    wire new_AGEMA_signal_6401 ;
    wire new_AGEMA_signal_6402 ;
    wire new_AGEMA_signal_6403 ;
    wire new_AGEMA_signal_6404 ;
    wire new_AGEMA_signal_6405 ;
    wire new_AGEMA_signal_6406 ;
    wire new_AGEMA_signal_6407 ;
    wire new_AGEMA_signal_6408 ;
    wire new_AGEMA_signal_6409 ;
    wire new_AGEMA_signal_6410 ;
    wire new_AGEMA_signal_6411 ;
    wire new_AGEMA_signal_6412 ;
    wire new_AGEMA_signal_6413 ;
    wire new_AGEMA_signal_6414 ;
    wire new_AGEMA_signal_6415 ;
    wire new_AGEMA_signal_6416 ;
    wire new_AGEMA_signal_6417 ;
    wire new_AGEMA_signal_6418 ;
    wire new_AGEMA_signal_6419 ;
    wire new_AGEMA_signal_6420 ;
    wire new_AGEMA_signal_6421 ;
    wire new_AGEMA_signal_6422 ;
    wire new_AGEMA_signal_6423 ;
    wire new_AGEMA_signal_6424 ;
    wire new_AGEMA_signal_6425 ;
    wire new_AGEMA_signal_6426 ;
    wire new_AGEMA_signal_6427 ;
    wire new_AGEMA_signal_6428 ;
    wire new_AGEMA_signal_6429 ;
    wire new_AGEMA_signal_6430 ;
    wire new_AGEMA_signal_6431 ;
    wire new_AGEMA_signal_6432 ;
    wire new_AGEMA_signal_6433 ;
    wire new_AGEMA_signal_6434 ;
    wire new_AGEMA_signal_6435 ;
    wire new_AGEMA_signal_6436 ;
    wire new_AGEMA_signal_6437 ;
    wire new_AGEMA_signal_6438 ;
    wire new_AGEMA_signal_6439 ;

    /* cells in depth 0 */
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) U5 ( .A0_t (Reset_t), .A0_f (Reset_f), .B0_t (Ready_t), .B0_f (Ready_f), .Z0_t (n9), .Z0_f (new_AGEMA_signal_3005) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U400 ( .A0_t (StateOut[199]), .A0_f (new_AGEMA_signal_2448), .A1_t (new_AGEMA_signal_2449), .A1_f (new_AGEMA_signal_2450), .B0_t (THETA_n200), .B0_f (new_AGEMA_signal_3258), .B1_t (new_AGEMA_signal_3259), .B1_f (new_AGEMA_signal_3260), .Z0_t (StateFromRhoPi[165]), .Z0_f (new_AGEMA_signal_3386), .Z1_t (new_AGEMA_signal_3387), .Z1_f (new_AGEMA_signal_3388) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U399 ( .A0_t (StateOut[191]), .A0_f (new_AGEMA_signal_2445), .A1_t (new_AGEMA_signal_2446), .A1_f (new_AGEMA_signal_2447), .B0_t (THETA_n200), .B0_f (new_AGEMA_signal_3258), .B1_t (new_AGEMA_signal_3259), .B1_f (new_AGEMA_signal_3260), .Z0_t (StateFromRhoPi[143]), .Z0_f (new_AGEMA_signal_3389), .Z1_t (new_AGEMA_signal_3390), .Z1_f (new_AGEMA_signal_3391) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U398 ( .A0_t (StateOut[183]), .A0_f (new_AGEMA_signal_3108), .A1_t (new_AGEMA_signal_3109), .A1_f (new_AGEMA_signal_3110), .B0_t (THETA_n200), .B0_f (new_AGEMA_signal_3258), .B1_t (new_AGEMA_signal_3259), .B1_f (new_AGEMA_signal_3260), .Z0_t (StateFromRhoPi[118]), .Z0_f (new_AGEMA_signal_3392), .Z1_t (new_AGEMA_signal_3393), .Z1_f (new_AGEMA_signal_3394) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U397 ( .A0_t (StateOut[175]), .A0_f (new_AGEMA_signal_2436), .A1_t (new_AGEMA_signal_2437), .A1_f (new_AGEMA_signal_2438), .B0_t (THETA_n200), .B0_f (new_AGEMA_signal_3258), .B1_t (new_AGEMA_signal_3259), .B1_f (new_AGEMA_signal_3260), .Z0_t (StateFromRhoPi[51]), .Z0_f (new_AGEMA_signal_3395), .Z1_t (new_AGEMA_signal_3396), .Z1_f (new_AGEMA_signal_3397) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U396 ( .A0_t (StateOut[167]), .A0_f (new_AGEMA_signal_2439), .A1_t (new_AGEMA_signal_2440), .A1_f (new_AGEMA_signal_2441), .B0_t (THETA_n200), .B0_f (new_AGEMA_signal_3258), .B1_t (new_AGEMA_signal_3259), .B1_f (new_AGEMA_signal_3260), .Z0_t (StateFromRhoPi[26]), .Z0_f (new_AGEMA_signal_3398), .Z1_t (new_AGEMA_signal_3399), .Z1_f (new_AGEMA_signal_3400) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U395 ( .A0_t (THETA_n199), .A0_f (new_AGEMA_signal_3015), .A1_t (new_AGEMA_signal_3016), .A1_f (new_AGEMA_signal_3017), .B0_t (THETA_n198), .B0_f (new_AGEMA_signal_3009), .B1_t (new_AGEMA_signal_3010), .B1_f (new_AGEMA_signal_3011), .Z0_t (THETA_n200), .Z0_f (new_AGEMA_signal_3258), .Z1_t (new_AGEMA_signal_3259), .Z1_f (new_AGEMA_signal_3260) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U394 ( .A0_t (StateOut[78]), .A0_f (new_AGEMA_signal_2466), .A1_t (new_AGEMA_signal_2467), .A1_f (new_AGEMA_signal_2468), .B0_t (THETA_n197), .B0_f (new_AGEMA_signal_3261), .B1_t (new_AGEMA_signal_3262), .B1_f (new_AGEMA_signal_3263), .Z0_t (StateFromRhoPi[192]), .Z0_f (new_AGEMA_signal_3401), .Z1_t (new_AGEMA_signal_3402), .Z1_f (new_AGEMA_signal_3403) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U393 ( .A0_t (StateOut[70]), .A0_f (new_AGEMA_signal_2463), .A1_t (new_AGEMA_signal_2464), .A1_f (new_AGEMA_signal_2465), .B0_t (THETA_n197), .B0_f (new_AGEMA_signal_3261), .B1_t (new_AGEMA_signal_3262), .B1_f (new_AGEMA_signal_3263), .Z0_t (StateFromRhoPi[131]), .Z0_f (new_AGEMA_signal_3404), .Z1_t (new_AGEMA_signal_3405), .Z1_f (new_AGEMA_signal_3406) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U392 ( .A0_t (StateOut[62]), .A0_f (new_AGEMA_signal_3114), .A1_t (new_AGEMA_signal_3115), .A1_f (new_AGEMA_signal_3116), .B0_t (THETA_n197), .B0_f (new_AGEMA_signal_3261), .B1_t (new_AGEMA_signal_3262), .B1_f (new_AGEMA_signal_3263), .Z0_t (StateFromRhoPi[104]), .Z0_f (new_AGEMA_signal_3407), .Z1_t (new_AGEMA_signal_3408), .Z1_f (new_AGEMA_signal_3409) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U391 ( .A0_t (StateOut[54]), .A0_f (new_AGEMA_signal_2454), .A1_t (new_AGEMA_signal_2455), .A1_f (new_AGEMA_signal_2456), .B0_t (THETA_n197), .B0_f (new_AGEMA_signal_3261), .B1_t (new_AGEMA_signal_3262), .B1_f (new_AGEMA_signal_3263), .Z0_t (StateFromRhoPi[42]), .Z0_f (new_AGEMA_signal_3410), .Z1_t (new_AGEMA_signal_3411), .Z1_f (new_AGEMA_signal_3412) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U390 ( .A0_t (StateOut[46]), .A0_f (new_AGEMA_signal_2457), .A1_t (new_AGEMA_signal_2458), .A1_f (new_AGEMA_signal_2459), .B0_t (THETA_n197), .B0_f (new_AGEMA_signal_3261), .B1_t (new_AGEMA_signal_3262), .B1_f (new_AGEMA_signal_3263), .Z0_t (StateFromRhoPi[23]), .Z0_f (new_AGEMA_signal_3413), .Z1_t (new_AGEMA_signal_3414), .Z1_f (new_AGEMA_signal_3415) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U389 ( .A0_t (THETA_n196), .A0_f (new_AGEMA_signal_3207), .A1_t (new_AGEMA_signal_3208), .A1_f (new_AGEMA_signal_3209), .B0_t (THETA_n198), .B0_f (new_AGEMA_signal_3009), .B1_t (new_AGEMA_signal_3010), .B1_f (new_AGEMA_signal_3011), .Z0_t (THETA_n197), .Z0_f (new_AGEMA_signal_3261), .Z1_t (new_AGEMA_signal_3262), .Z1_f (new_AGEMA_signal_3263) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U388 ( .A0_t (OutData_s0_t[6]), .A0_f (OutData_s0_f[6]), .A1_t (OutData_s1_t[6]), .A1_f (OutData_s1_f[6]), .B0_t (THETA_n195), .B0_f (new_AGEMA_signal_2868), .B1_t (new_AGEMA_signal_2869), .B1_f (new_AGEMA_signal_2870), .Z0_t (THETA_n198), .Z0_f (new_AGEMA_signal_3009), .Z1_t (new_AGEMA_signal_3010), .Z1_f (new_AGEMA_signal_3011) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U387 ( .A0_t (THETA_n194), .A0_f (new_AGEMA_signal_2145), .A1_t (new_AGEMA_signal_2146), .A1_f (new_AGEMA_signal_2147), .B0_t (THETA_n193), .B0_f (new_AGEMA_signal_2136), .B1_t (new_AGEMA_signal_2137), .B1_f (new_AGEMA_signal_2138), .Z0_t (THETA_n195), .Z0_f (new_AGEMA_signal_2868), .Z1_t (new_AGEMA_signal_2869), .Z1_f (new_AGEMA_signal_2870) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U386 ( .A0_t (StateOut[14]), .A0_f (new_AGEMA_signal_2130), .A1_t (new_AGEMA_signal_2131), .A1_f (new_AGEMA_signal_2132), .B0_t (StateOut[22]), .B0_f (new_AGEMA_signal_2133), .B1_t (new_AGEMA_signal_2134), .B1_f (new_AGEMA_signal_2135), .Z0_t (THETA_n193), .Z0_f (new_AGEMA_signal_2136), .Z1_t (new_AGEMA_signal_2137), .Z1_f (new_AGEMA_signal_2138) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U385 ( .A0_t (StateOut[38]), .A0_f (new_AGEMA_signal_2139), .A1_t (new_AGEMA_signal_2140), .A1_f (new_AGEMA_signal_2141), .B0_t (StateOut[30]), .B0_f (new_AGEMA_signal_2142), .B1_t (new_AGEMA_signal_2143), .B1_f (new_AGEMA_signal_2144), .Z0_t (THETA_n194), .Z0_f (new_AGEMA_signal_2145), .Z1_t (new_AGEMA_signal_2146), .Z1_f (new_AGEMA_signal_2147) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U384 ( .A0_t (StateOut[112]), .A0_f (new_AGEMA_signal_2394), .A1_t (new_AGEMA_signal_2395), .A1_f (new_AGEMA_signal_2396), .B0_t (THETA_n192), .B0_f (new_AGEMA_signal_3264), .B1_t (new_AGEMA_signal_3265), .B1_f (new_AGEMA_signal_3266), .Z0_t (StateFromRhoPi[173]), .Z0_f (new_AGEMA_signal_3416), .Z1_t (new_AGEMA_signal_3417), .Z1_f (new_AGEMA_signal_3418) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U383 ( .A0_t (StateOut[104]), .A0_f (new_AGEMA_signal_2391), .A1_t (new_AGEMA_signal_2392), .A1_f (new_AGEMA_signal_2393), .B0_t (THETA_n192), .B0_f (new_AGEMA_signal_3264), .B1_t (new_AGEMA_signal_3265), .B1_f (new_AGEMA_signal_3266), .Z0_t (StateFromRhoPi[151]), .Z0_f (new_AGEMA_signal_3419), .Z1_t (new_AGEMA_signal_3420), .Z1_f (new_AGEMA_signal_3421) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U382 ( .A0_t (StateOut[96]), .A0_f (new_AGEMA_signal_3090), .A1_t (new_AGEMA_signal_3091), .A1_f (new_AGEMA_signal_3092), .B0_t (THETA_n192), .B0_f (new_AGEMA_signal_3264), .B1_t (new_AGEMA_signal_3265), .B1_f (new_AGEMA_signal_3266), .Z0_t (StateFromRhoPi[83]), .Z0_f (new_AGEMA_signal_3422), .Z1_t (new_AGEMA_signal_3423), .Z1_f (new_AGEMA_signal_3424) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U381 ( .A0_t (StateOut[88]), .A0_f (new_AGEMA_signal_2382), .A1_t (new_AGEMA_signal_2383), .A1_f (new_AGEMA_signal_2384), .B0_t (THETA_n192), .B0_f (new_AGEMA_signal_3264), .B1_t (new_AGEMA_signal_3265), .B1_f (new_AGEMA_signal_3266), .Z0_t (StateFromRhoPi[62]), .Z0_f (new_AGEMA_signal_3425), .Z1_t (new_AGEMA_signal_3426), .Z1_f (new_AGEMA_signal_3427) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U380 ( .A0_t (StateOut[80]), .A0_f (new_AGEMA_signal_2385), .A1_t (new_AGEMA_signal_2386), .A1_f (new_AGEMA_signal_2387), .B0_t (THETA_n192), .B0_f (new_AGEMA_signal_3264), .B1_t (new_AGEMA_signal_3265), .B1_f (new_AGEMA_signal_3266), .Z0_t (StateFromRhoPi[38]), .Z0_f (new_AGEMA_signal_3428), .Z1_t (new_AGEMA_signal_3429), .Z1_f (new_AGEMA_signal_3430) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U379 ( .A0_t (THETA_n191), .A0_f (new_AGEMA_signal_3051), .A1_t (new_AGEMA_signal_3052), .A1_f (new_AGEMA_signal_3053), .B0_t (THETA_n199), .B0_f (new_AGEMA_signal_3015), .B1_t (new_AGEMA_signal_3016), .B1_f (new_AGEMA_signal_3017), .Z0_t (THETA_n192), .Z0_f (new_AGEMA_signal_3264), .Z1_t (new_AGEMA_signal_3265), .Z1_f (new_AGEMA_signal_3266) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U378 ( .A0_t (StateOut[127]), .A0_f (new_AGEMA_signal_3012), .A1_t (new_AGEMA_signal_3013), .A1_f (new_AGEMA_signal_3014), .B0_t (THETA_n190), .B0_f (new_AGEMA_signal_2871), .B1_t (new_AGEMA_signal_2872), .B1_f (new_AGEMA_signal_2873), .Z0_t (THETA_n199), .Z0_f (new_AGEMA_signal_3015), .Z1_t (new_AGEMA_signal_3016), .Z1_f (new_AGEMA_signal_3017) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U377 ( .A0_t (THETA_n189), .A0_f (new_AGEMA_signal_2163), .A1_t (new_AGEMA_signal_2164), .A1_f (new_AGEMA_signal_2165), .B0_t (THETA_n188), .B0_f (new_AGEMA_signal_2154), .B1_t (new_AGEMA_signal_2155), .B1_f (new_AGEMA_signal_2156), .Z0_t (THETA_n190), .Z0_f (new_AGEMA_signal_2871), .Z1_t (new_AGEMA_signal_2872), .Z1_f (new_AGEMA_signal_2873) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U376 ( .A0_t (StateOut[135]), .A0_f (new_AGEMA_signal_2148), .A1_t (new_AGEMA_signal_2149), .A1_f (new_AGEMA_signal_2150), .B0_t (StateOut[143]), .B0_f (new_AGEMA_signal_2151), .B1_t (new_AGEMA_signal_2152), .B1_f (new_AGEMA_signal_2153), .Z0_t (THETA_n188), .Z0_f (new_AGEMA_signal_2154), .Z1_t (new_AGEMA_signal_2155), .Z1_f (new_AGEMA_signal_2156) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U375 ( .A0_t (StateOut[159]), .A0_f (new_AGEMA_signal_2157), .A1_t (new_AGEMA_signal_2158), .A1_f (new_AGEMA_signal_2159), .B0_t (StateOut[151]), .B0_f (new_AGEMA_signal_2160), .B1_t (new_AGEMA_signal_2161), .B1_f (new_AGEMA_signal_2162), .Z0_t (THETA_n189), .Z0_f (new_AGEMA_signal_2163), .Z1_t (new_AGEMA_signal_2164), .Z1_f (new_AGEMA_signal_2165) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U374 ( .A0_t (StateOut[198]), .A0_f (new_AGEMA_signal_2502), .A1_t (new_AGEMA_signal_2503), .A1_f (new_AGEMA_signal_2504), .B0_t (THETA_n187), .B0_f (new_AGEMA_signal_3267), .B1_t (new_AGEMA_signal_3268), .B1_f (new_AGEMA_signal_3269), .Z0_t (StateFromRhoPi[164]), .Z0_f (new_AGEMA_signal_3431), .Z1_t (new_AGEMA_signal_3432), .Z1_f (new_AGEMA_signal_3433) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U373 ( .A0_t (StateOut[190]), .A0_f (new_AGEMA_signal_2499), .A1_t (new_AGEMA_signal_2500), .A1_f (new_AGEMA_signal_2501), .B0_t (THETA_n187), .B0_f (new_AGEMA_signal_3267), .B1_t (new_AGEMA_signal_3268), .B1_f (new_AGEMA_signal_3269), .Z0_t (StateFromRhoPi[142]), .Z0_f (new_AGEMA_signal_3434), .Z1_t (new_AGEMA_signal_3435), .Z1_f (new_AGEMA_signal_3436) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U372 ( .A0_t (StateOut[182]), .A0_f (new_AGEMA_signal_3126), .A1_t (new_AGEMA_signal_3127), .A1_f (new_AGEMA_signal_3128), .B0_t (THETA_n187), .B0_f (new_AGEMA_signal_3267), .B1_t (new_AGEMA_signal_3268), .B1_f (new_AGEMA_signal_3269), .Z0_t (StateFromRhoPi[117]), .Z0_f (new_AGEMA_signal_3437), .Z1_t (new_AGEMA_signal_3438), .Z1_f (new_AGEMA_signal_3439) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U371 ( .A0_t (StateOut[174]), .A0_f (new_AGEMA_signal_2490), .A1_t (new_AGEMA_signal_2491), .A1_f (new_AGEMA_signal_2492), .B0_t (THETA_n187), .B0_f (new_AGEMA_signal_3267), .B1_t (new_AGEMA_signal_3268), .B1_f (new_AGEMA_signal_3269), .Z0_t (StateFromRhoPi[50]), .Z0_f (new_AGEMA_signal_3440), .Z1_t (new_AGEMA_signal_3441), .Z1_f (new_AGEMA_signal_3442) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U370 ( .A0_t (StateOut[166]), .A0_f (new_AGEMA_signal_2493), .A1_t (new_AGEMA_signal_2494), .A1_f (new_AGEMA_signal_2495), .B0_t (THETA_n187), .B0_f (new_AGEMA_signal_3267), .B1_t (new_AGEMA_signal_3268), .B1_f (new_AGEMA_signal_3269), .Z0_t (StateFromRhoPi[25]), .Z0_f (new_AGEMA_signal_3443), .Z1_t (new_AGEMA_signal_3444), .Z1_f (new_AGEMA_signal_3445) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U369 ( .A0_t (THETA_n186), .A0_f (new_AGEMA_signal_3177), .A1_t (new_AGEMA_signal_3178), .A1_f (new_AGEMA_signal_3179), .B0_t (THETA_n185), .B0_f (new_AGEMA_signal_3021), .B1_t (new_AGEMA_signal_3022), .B1_f (new_AGEMA_signal_3023), .Z0_t (THETA_n187), .Z0_f (new_AGEMA_signal_3267), .Z1_t (new_AGEMA_signal_3268), .Z1_f (new_AGEMA_signal_3269) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U368 ( .A0_t (StateOut[119]), .A0_f (new_AGEMA_signal_2484), .A1_t (new_AGEMA_signal_2485), .A1_f (new_AGEMA_signal_2486), .B0_t (THETA_n184), .B0_f (new_AGEMA_signal_3270), .B1_t (new_AGEMA_signal_3271), .B1_f (new_AGEMA_signal_3272), .Z0_t (StateFromRhoPi[172]), .Z0_f (new_AGEMA_signal_3446), .Z1_t (new_AGEMA_signal_3447), .Z1_f (new_AGEMA_signal_3448) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U367 ( .A0_t (StateOut[111]), .A0_f (new_AGEMA_signal_2481), .A1_t (new_AGEMA_signal_2482), .A1_f (new_AGEMA_signal_2483), .B0_t (THETA_n184), .B0_f (new_AGEMA_signal_3270), .B1_t (new_AGEMA_signal_3271), .B1_f (new_AGEMA_signal_3272), .Z0_t (StateFromRhoPi[150]), .Z0_f (new_AGEMA_signal_3449), .Z1_t (new_AGEMA_signal_3450), .Z1_f (new_AGEMA_signal_3451) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U366 ( .A0_t (StateOut[103]), .A0_f (new_AGEMA_signal_3120), .A1_t (new_AGEMA_signal_3121), .A1_f (new_AGEMA_signal_3122), .B0_t (THETA_n184), .B0_f (new_AGEMA_signal_3270), .B1_t (new_AGEMA_signal_3271), .B1_f (new_AGEMA_signal_3272), .Z0_t (StateFromRhoPi[82]), .Z0_f (new_AGEMA_signal_3452), .Z1_t (new_AGEMA_signal_3453), .Z1_f (new_AGEMA_signal_3454) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U365 ( .A0_t (StateOut[95]), .A0_f (new_AGEMA_signal_2472), .A1_t (new_AGEMA_signal_2473), .A1_f (new_AGEMA_signal_2474), .B0_t (THETA_n184), .B0_f (new_AGEMA_signal_3270), .B1_t (new_AGEMA_signal_3271), .B1_f (new_AGEMA_signal_3272), .Z0_t (StateFromRhoPi[61]), .Z0_f (new_AGEMA_signal_3455), .Z1_t (new_AGEMA_signal_3456), .Z1_f (new_AGEMA_signal_3457) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U364 ( .A0_t (StateOut[87]), .A0_f (new_AGEMA_signal_2475), .A1_t (new_AGEMA_signal_2476), .A1_f (new_AGEMA_signal_2477), .B0_t (THETA_n184), .B0_f (new_AGEMA_signal_3270), .B1_t (new_AGEMA_signal_3271), .B1_f (new_AGEMA_signal_3272), .Z0_t (StateFromRhoPi[37]), .Z0_f (new_AGEMA_signal_3458), .Z1_t (new_AGEMA_signal_3459), .Z1_f (new_AGEMA_signal_3460) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U363 ( .A0_t (THETA_n183), .A0_f (new_AGEMA_signal_3075), .A1_t (new_AGEMA_signal_3076), .A1_f (new_AGEMA_signal_3077), .B0_t (THETA_n185), .B0_f (new_AGEMA_signal_3021), .B1_t (new_AGEMA_signal_3022), .B1_f (new_AGEMA_signal_3023), .Z0_t (THETA_n184), .Z0_f (new_AGEMA_signal_3270), .Z1_t (new_AGEMA_signal_3271), .Z1_f (new_AGEMA_signal_3272) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U362 ( .A0_t (StateOut[126]), .A0_f (new_AGEMA_signal_3018), .A1_t (new_AGEMA_signal_3019), .A1_f (new_AGEMA_signal_3020), .B0_t (THETA_n182), .B0_f (new_AGEMA_signal_2874), .B1_t (new_AGEMA_signal_2875), .B1_f (new_AGEMA_signal_2876), .Z0_t (THETA_n185), .Z0_f (new_AGEMA_signal_3021), .Z1_t (new_AGEMA_signal_3022), .Z1_f (new_AGEMA_signal_3023) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U361 ( .A0_t (THETA_n181), .A0_f (new_AGEMA_signal_2181), .A1_t (new_AGEMA_signal_2182), .A1_f (new_AGEMA_signal_2183), .B0_t (THETA_n180), .B0_f (new_AGEMA_signal_2172), .B1_t (new_AGEMA_signal_2173), .B1_f (new_AGEMA_signal_2174), .Z0_t (THETA_n182), .Z0_f (new_AGEMA_signal_2874), .Z1_t (new_AGEMA_signal_2875), .Z1_f (new_AGEMA_signal_2876) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U360 ( .A0_t (StateOut[134]), .A0_f (new_AGEMA_signal_2166), .A1_t (new_AGEMA_signal_2167), .A1_f (new_AGEMA_signal_2168), .B0_t (StateOut[142]), .B0_f (new_AGEMA_signal_2169), .B1_t (new_AGEMA_signal_2170), .B1_f (new_AGEMA_signal_2171), .Z0_t (THETA_n180), .Z0_f (new_AGEMA_signal_2172), .Z1_t (new_AGEMA_signal_2173), .Z1_f (new_AGEMA_signal_2174) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U359 ( .A0_t (StateOut[158]), .A0_f (new_AGEMA_signal_2175), .A1_t (new_AGEMA_signal_2176), .A1_f (new_AGEMA_signal_2177), .B0_t (StateOut[150]), .B0_f (new_AGEMA_signal_2178), .B1_t (new_AGEMA_signal_2179), .B1_f (new_AGEMA_signal_2180), .Z0_t (THETA_n181), .Z0_f (new_AGEMA_signal_2181), .Z1_t (new_AGEMA_signal_2182), .Z1_f (new_AGEMA_signal_2183) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U358 ( .A0_t (StateOut[196]), .A0_f (new_AGEMA_signal_2718), .A1_t (new_AGEMA_signal_2719), .A1_f (new_AGEMA_signal_2720), .B0_t (THETA_n179), .B0_f (new_AGEMA_signal_3273), .B1_t (new_AGEMA_signal_3274), .B1_f (new_AGEMA_signal_3275), .Z0_t (StateFromRhoPi[162]), .Z0_f (new_AGEMA_signal_3461), .Z1_t (new_AGEMA_signal_3462), .Z1_f (new_AGEMA_signal_3463) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U357 ( .A0_t (StateOut[188]), .A0_f (new_AGEMA_signal_2715), .A1_t (new_AGEMA_signal_2716), .A1_f (new_AGEMA_signal_2717), .B0_t (THETA_n179), .B0_f (new_AGEMA_signal_3273), .B1_t (new_AGEMA_signal_3274), .B1_f (new_AGEMA_signal_3275), .Z0_t (StateFromRhoPi[140]), .Z0_f (new_AGEMA_signal_3464), .Z1_t (new_AGEMA_signal_3465), .Z1_f (new_AGEMA_signal_3466) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U356 ( .A0_t (StateOut[180]), .A0_f (new_AGEMA_signal_3198), .A1_t (new_AGEMA_signal_3199), .A1_f (new_AGEMA_signal_3200), .B0_t (THETA_n179), .B0_f (new_AGEMA_signal_3273), .B1_t (new_AGEMA_signal_3274), .B1_f (new_AGEMA_signal_3275), .Z0_t (StateFromRhoPi[115]), .Z0_f (new_AGEMA_signal_3467), .Z1_t (new_AGEMA_signal_3468), .Z1_f (new_AGEMA_signal_3469) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U355 ( .A0_t (StateOut[172]), .A0_f (new_AGEMA_signal_2706), .A1_t (new_AGEMA_signal_2707), .A1_f (new_AGEMA_signal_2708), .B0_t (THETA_n179), .B0_f (new_AGEMA_signal_3273), .B1_t (new_AGEMA_signal_3274), .B1_f (new_AGEMA_signal_3275), .Z0_t (StateFromRhoPi[48]), .Z0_f (new_AGEMA_signal_3470), .Z1_t (new_AGEMA_signal_3471), .Z1_f (new_AGEMA_signal_3472) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U354 ( .A0_t (StateOut[164]), .A0_f (new_AGEMA_signal_2709), .A1_t (new_AGEMA_signal_2710), .A1_f (new_AGEMA_signal_2711), .B0_t (THETA_n179), .B0_f (new_AGEMA_signal_3273), .B1_t (new_AGEMA_signal_3274), .B1_f (new_AGEMA_signal_3275), .Z0_t (StateFromRhoPi[31]), .Z0_f (new_AGEMA_signal_3473), .Z1_t (new_AGEMA_signal_3474), .Z1_f (new_AGEMA_signal_3475) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U353 ( .A0_t (THETA_n178), .A0_f (new_AGEMA_signal_3087), .A1_t (new_AGEMA_signal_3088), .A1_f (new_AGEMA_signal_3089), .B0_t (THETA_n177), .B0_f (new_AGEMA_signal_3027), .B1_t (new_AGEMA_signal_3028), .B1_f (new_AGEMA_signal_3029), .Z0_t (THETA_n179), .Z0_f (new_AGEMA_signal_3273), .Z1_t (new_AGEMA_signal_3274), .Z1_f (new_AGEMA_signal_3275) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U352 ( .A0_t (StateOut[75]), .A0_f (new_AGEMA_signal_2628), .A1_t (new_AGEMA_signal_2629), .A1_f (new_AGEMA_signal_2630), .B0_t (THETA_n176), .B0_f (new_AGEMA_signal_3276), .B1_t (new_AGEMA_signal_3277), .B1_f (new_AGEMA_signal_3278), .Z0_t (StateFromRhoPi[197]), .Z0_f (new_AGEMA_signal_3476), .Z1_t (new_AGEMA_signal_3477), .Z1_f (new_AGEMA_signal_3478) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U351 ( .A0_t (StateOut[67]), .A0_f (new_AGEMA_signal_2625), .A1_t (new_AGEMA_signal_2626), .A1_f (new_AGEMA_signal_2627), .B0_t (THETA_n176), .B0_f (new_AGEMA_signal_3276), .B1_t (new_AGEMA_signal_3277), .B1_f (new_AGEMA_signal_3278), .Z0_t (StateFromRhoPi[128]), .Z0_f (new_AGEMA_signal_3479), .Z1_t (new_AGEMA_signal_3480), .Z1_f (new_AGEMA_signal_3481) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U350 ( .A0_t (StateOut[59]), .A0_f (new_AGEMA_signal_3168), .A1_t (new_AGEMA_signal_3169), .A1_f (new_AGEMA_signal_3170), .B0_t (THETA_n176), .B0_f (new_AGEMA_signal_3276), .B1_t (new_AGEMA_signal_3277), .B1_f (new_AGEMA_signal_3278), .Z0_t (StateFromRhoPi[109]), .Z0_f (new_AGEMA_signal_3482), .Z1_t (new_AGEMA_signal_3483), .Z1_f (new_AGEMA_signal_3484) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U349 ( .A0_t (StateOut[51]), .A0_f (new_AGEMA_signal_2616), .A1_t (new_AGEMA_signal_2617), .A1_f (new_AGEMA_signal_2618), .B0_t (THETA_n176), .B0_f (new_AGEMA_signal_3276), .B1_t (new_AGEMA_signal_3277), .B1_f (new_AGEMA_signal_3278), .Z0_t (StateFromRhoPi[47]), .Z0_f (new_AGEMA_signal_3485), .Z1_t (new_AGEMA_signal_3486), .Z1_f (new_AGEMA_signal_3487) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U348 ( .A0_t (StateOut[43]), .A0_f (new_AGEMA_signal_2619), .A1_t (new_AGEMA_signal_2620), .A1_f (new_AGEMA_signal_2621), .B0_t (THETA_n176), .B0_f (new_AGEMA_signal_3276), .B1_t (new_AGEMA_signal_3277), .B1_f (new_AGEMA_signal_3278), .Z0_t (StateFromRhoPi[20]), .Z0_f (new_AGEMA_signal_3488), .Z1_t (new_AGEMA_signal_3489), .Z1_f (new_AGEMA_signal_3490) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U347 ( .A0_t (THETA_n175), .A0_f (new_AGEMA_signal_3039), .A1_t (new_AGEMA_signal_3040), .A1_f (new_AGEMA_signal_3041), .B0_t (THETA_n177), .B0_f (new_AGEMA_signal_3027), .B1_t (new_AGEMA_signal_3028), .B1_f (new_AGEMA_signal_3029), .Z0_t (THETA_n176), .Z0_f (new_AGEMA_signal_3276), .Z1_t (new_AGEMA_signal_3277), .Z1_f (new_AGEMA_signal_3278) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U346 ( .A0_t (OutData_s0_t[3]), .A0_f (OutData_s0_f[3]), .A1_t (OutData_s1_t[3]), .A1_f (OutData_s1_f[3]), .B0_t (THETA_n174), .B0_f (new_AGEMA_signal_2877), .B1_t (new_AGEMA_signal_2878), .B1_f (new_AGEMA_signal_2879), .Z0_t (THETA_n177), .Z0_f (new_AGEMA_signal_3027), .Z1_t (new_AGEMA_signal_3028), .Z1_f (new_AGEMA_signal_3029) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U345 ( .A0_t (THETA_n173), .A0_f (new_AGEMA_signal_2199), .A1_t (new_AGEMA_signal_2200), .A1_f (new_AGEMA_signal_2201), .B0_t (THETA_n172), .B0_f (new_AGEMA_signal_2190), .B1_t (new_AGEMA_signal_2191), .B1_f (new_AGEMA_signal_2192), .Z0_t (THETA_n174), .Z0_f (new_AGEMA_signal_2877), .Z1_t (new_AGEMA_signal_2878), .Z1_f (new_AGEMA_signal_2879) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U344 ( .A0_t (StateOut[11]), .A0_f (new_AGEMA_signal_2184), .A1_t (new_AGEMA_signal_2185), .A1_f (new_AGEMA_signal_2186), .B0_t (StateOut[19]), .B0_f (new_AGEMA_signal_2187), .B1_t (new_AGEMA_signal_2188), .B1_f (new_AGEMA_signal_2189), .Z0_t (THETA_n172), .Z0_f (new_AGEMA_signal_2190), .Z1_t (new_AGEMA_signal_2191), .Z1_f (new_AGEMA_signal_2192) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U343 ( .A0_t (StateOut[35]), .A0_f (new_AGEMA_signal_2193), .A1_t (new_AGEMA_signal_2194), .A1_f (new_AGEMA_signal_2195), .B0_t (StateOut[27]), .B0_f (new_AGEMA_signal_2196), .B1_t (new_AGEMA_signal_2197), .B1_f (new_AGEMA_signal_2198), .Z0_t (THETA_n173), .Z0_f (new_AGEMA_signal_2199), .Z1_t (new_AGEMA_signal_2200), .Z1_f (new_AGEMA_signal_2201) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U342 ( .A0_t (StateOut[193]), .A0_f (new_AGEMA_signal_2250), .A1_t (new_AGEMA_signal_2251), .A1_f (new_AGEMA_signal_2252), .B0_t (THETA_n171), .B0_f (new_AGEMA_signal_3279), .B1_t (new_AGEMA_signal_3280), .B1_f (new_AGEMA_signal_3281), .Z0_t (StateFromRhoPi[167]), .Z0_f (new_AGEMA_signal_3491), .Z1_t (new_AGEMA_signal_3492), .Z1_f (new_AGEMA_signal_3493) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U341 ( .A0_t (StateOut[185]), .A0_f (new_AGEMA_signal_2247), .A1_t (new_AGEMA_signal_2248), .A1_f (new_AGEMA_signal_2249), .B0_t (THETA_n171), .B0_f (new_AGEMA_signal_3279), .B1_t (new_AGEMA_signal_3280), .B1_f (new_AGEMA_signal_3281), .Z0_t (StateFromRhoPi[137]), .Z0_f (new_AGEMA_signal_3494), .Z1_t (new_AGEMA_signal_3495), .Z1_f (new_AGEMA_signal_3496) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U340 ( .A0_t (StateOut[177]), .A0_f (new_AGEMA_signal_3042), .A1_t (new_AGEMA_signal_3043), .A1_f (new_AGEMA_signal_3044), .B0_t (THETA_n171), .B0_f (new_AGEMA_signal_3279), .B1_t (new_AGEMA_signal_3280), .B1_f (new_AGEMA_signal_3281), .Z0_t (StateFromRhoPi[112]), .Z0_f (new_AGEMA_signal_3497), .Z1_t (new_AGEMA_signal_3498), .Z1_f (new_AGEMA_signal_3499) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U339 ( .A0_t (StateOut[169]), .A0_f (new_AGEMA_signal_2238), .A1_t (new_AGEMA_signal_2239), .A1_f (new_AGEMA_signal_2240), .B0_t (THETA_n171), .B0_f (new_AGEMA_signal_3279), .B1_t (new_AGEMA_signal_3280), .B1_f (new_AGEMA_signal_3281), .Z0_t (StateFromRhoPi[53]), .Z0_f (new_AGEMA_signal_3500), .Z1_t (new_AGEMA_signal_3501), .Z1_f (new_AGEMA_signal_3502) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U338 ( .A0_t (StateOut[161]), .A0_f (new_AGEMA_signal_2241), .A1_t (new_AGEMA_signal_2242), .A1_f (new_AGEMA_signal_2243), .B0_t (THETA_n171), .B0_f (new_AGEMA_signal_3279), .B1_t (new_AGEMA_signal_3280), .B1_f (new_AGEMA_signal_3281), .Z0_t (StateFromRhoPi[28]), .Z0_f (new_AGEMA_signal_3503), .Z1_t (new_AGEMA_signal_3504), .Z1_f (new_AGEMA_signal_3505) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U337 ( .A0_t (THETA_n170), .A0_f (new_AGEMA_signal_3057), .A1_t (new_AGEMA_signal_3058), .A1_f (new_AGEMA_signal_3059), .B0_t (THETA_n169), .B0_f (new_AGEMA_signal_3033), .B1_t (new_AGEMA_signal_3034), .B1_f (new_AGEMA_signal_3035), .Z0_t (THETA_n171), .Z0_f (new_AGEMA_signal_3279), .Z1_t (new_AGEMA_signal_3280), .Z1_f (new_AGEMA_signal_3281) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U336 ( .A0_t (StateOut[72]), .A0_f (new_AGEMA_signal_2265), .A1_t (new_AGEMA_signal_2266), .A1_f (new_AGEMA_signal_2267), .B0_t (THETA_n168), .B0_f (new_AGEMA_signal_3282), .B1_t (new_AGEMA_signal_3283), .B1_f (new_AGEMA_signal_3284), .Z0_t (StateFromRhoPi[194]), .Z0_f (new_AGEMA_signal_3506), .Z1_t (new_AGEMA_signal_3507), .Z1_f (new_AGEMA_signal_3508) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U335 ( .A0_t (StateOut[64]), .A0_f (new_AGEMA_signal_3048), .A1_t (new_AGEMA_signal_3049), .A1_f (new_AGEMA_signal_3050), .B0_t (THETA_n168), .B0_f (new_AGEMA_signal_3282), .B1_t (new_AGEMA_signal_3283), .B1_f (new_AGEMA_signal_3284), .Z0_t (StateFromRhoPi[133]), .Z0_f (new_AGEMA_signal_3509), .Z1_t (new_AGEMA_signal_3510), .Z1_f (new_AGEMA_signal_3511) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U334 ( .A0_t (StateOut[56]), .A0_f (new_AGEMA_signal_2268), .A1_t (new_AGEMA_signal_2269), .A1_f (new_AGEMA_signal_2270), .B0_t (THETA_n168), .B0_f (new_AGEMA_signal_3282), .B1_t (new_AGEMA_signal_3283), .B1_f (new_AGEMA_signal_3284), .Z0_t (StateFromRhoPi[106]), .Z0_f (new_AGEMA_signal_3512), .Z1_t (new_AGEMA_signal_3513), .Z1_f (new_AGEMA_signal_3514) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U333 ( .A0_t (StateOut[48]), .A0_f (new_AGEMA_signal_2256), .A1_t (new_AGEMA_signal_2257), .A1_f (new_AGEMA_signal_2258), .B0_t (THETA_n168), .B0_f (new_AGEMA_signal_3282), .B1_t (new_AGEMA_signal_3283), .B1_f (new_AGEMA_signal_3284), .Z0_t (StateFromRhoPi[44]), .Z0_f (new_AGEMA_signal_3515), .Z1_t (new_AGEMA_signal_3516), .Z1_f (new_AGEMA_signal_3517) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U332 ( .A0_t (StateOut[40]), .A0_f (new_AGEMA_signal_2259), .A1_t (new_AGEMA_signal_2260), .A1_f (new_AGEMA_signal_2261), .B0_t (THETA_n168), .B0_f (new_AGEMA_signal_3282), .B1_t (new_AGEMA_signal_3283), .B1_f (new_AGEMA_signal_3284), .Z0_t (StateFromRhoPi[17]), .Z0_f (new_AGEMA_signal_3518), .Z1_t (new_AGEMA_signal_3519), .Z1_f (new_AGEMA_signal_3520) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U331 ( .A0_t (THETA_n167), .A0_f (new_AGEMA_signal_3123), .A1_t (new_AGEMA_signal_3124), .A1_f (new_AGEMA_signal_3125), .B0_t (THETA_n169), .B0_f (new_AGEMA_signal_3033), .B1_t (new_AGEMA_signal_3034), .B1_f (new_AGEMA_signal_3035), .Z0_t (THETA_n168), .Z0_f (new_AGEMA_signal_3282), .Z1_t (new_AGEMA_signal_3283), .Z1_f (new_AGEMA_signal_3284) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U330 ( .A0_t (OutData_s0_t[0]), .A0_f (OutData_s0_f[0]), .A1_t (OutData_s1_t[0]), .A1_f (OutData_s1_f[0]), .B0_t (THETA_n166), .B0_f (new_AGEMA_signal_2880), .B1_t (new_AGEMA_signal_2881), .B1_f (new_AGEMA_signal_2882), .Z0_t (THETA_n169), .Z0_f (new_AGEMA_signal_3033), .Z1_t (new_AGEMA_signal_3034), .Z1_f (new_AGEMA_signal_3035) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U329 ( .A0_t (THETA_n165), .A0_f (new_AGEMA_signal_2217), .A1_t (new_AGEMA_signal_2218), .A1_f (new_AGEMA_signal_2219), .B0_t (THETA_n164), .B0_f (new_AGEMA_signal_2208), .B1_t (new_AGEMA_signal_2209), .B1_f (new_AGEMA_signal_2210), .Z0_t (THETA_n166), .Z0_f (new_AGEMA_signal_2880), .Z1_t (new_AGEMA_signal_2881), .Z1_f (new_AGEMA_signal_2882) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U328 ( .A0_t (StateOut[8]), .A0_f (new_AGEMA_signal_2202), .A1_t (new_AGEMA_signal_2203), .A1_f (new_AGEMA_signal_2204), .B0_t (StateOut[16]), .B0_f (new_AGEMA_signal_2205), .B1_t (new_AGEMA_signal_2206), .B1_f (new_AGEMA_signal_2207), .Z0_t (THETA_n164), .Z0_f (new_AGEMA_signal_2208), .Z1_t (new_AGEMA_signal_2209), .Z1_f (new_AGEMA_signal_2210) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U327 ( .A0_t (StateOut[32]), .A0_f (new_AGEMA_signal_2211), .A1_t (new_AGEMA_signal_2212), .A1_f (new_AGEMA_signal_2213), .B0_t (StateOut[24]), .B0_f (new_AGEMA_signal_2214), .B1_t (new_AGEMA_signal_2215), .B1_f (new_AGEMA_signal_2216), .Z0_t (THETA_n165), .Z0_f (new_AGEMA_signal_2217), .Z1_t (new_AGEMA_signal_2218), .Z1_f (new_AGEMA_signal_2219) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U326 ( .A0_t (StateOut[154]), .A0_f (new_AGEMA_signal_2754), .A1_t (new_AGEMA_signal_2755), .A1_f (new_AGEMA_signal_2756), .B0_t (THETA_n163), .B0_f (new_AGEMA_signal_3285), .B1_t (new_AGEMA_signal_3286), .B1_f (new_AGEMA_signal_3287), .Z0_t (StateFromRhoPi[186]), .Z0_f (new_AGEMA_signal_3521), .Z1_t (new_AGEMA_signal_3522), .Z1_f (new_AGEMA_signal_3523) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U325 ( .A0_t (StateOut[146]), .A0_f (new_AGEMA_signal_2751), .A1_t (new_AGEMA_signal_2752), .A1_f (new_AGEMA_signal_2753), .B0_t (THETA_n163), .B0_f (new_AGEMA_signal_3285), .B1_t (new_AGEMA_signal_3286), .B1_f (new_AGEMA_signal_3287), .Z0_t (StateFromRhoPi[127]), .Z0_f (new_AGEMA_signal_3524), .Z1_t (new_AGEMA_signal_3525), .Z1_f (new_AGEMA_signal_3526) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U324 ( .A0_t (StateOut[138]), .A0_f (new_AGEMA_signal_3210), .A1_t (new_AGEMA_signal_3211), .A1_f (new_AGEMA_signal_3212), .B0_t (THETA_n163), .B0_f (new_AGEMA_signal_3285), .B1_t (new_AGEMA_signal_3286), .B1_f (new_AGEMA_signal_3287), .Z0_t (StateFromRhoPi[99]), .Z0_f (new_AGEMA_signal_3527), .Z1_t (new_AGEMA_signal_3528), .Z1_f (new_AGEMA_signal_3529) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U323 ( .A0_t (StateOut[130]), .A0_f (new_AGEMA_signal_2742), .A1_t (new_AGEMA_signal_2743), .A1_f (new_AGEMA_signal_2744), .B0_t (THETA_n163), .B0_f (new_AGEMA_signal_3285), .B1_t (new_AGEMA_signal_3286), .B1_f (new_AGEMA_signal_3287), .Z0_t (StateFromRhoPi[73]), .Z0_f (new_AGEMA_signal_3530), .Z1_t (new_AGEMA_signal_3531), .Z1_f (new_AGEMA_signal_3532) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U322 ( .A0_t (StateOut[122]), .A0_f (new_AGEMA_signal_2745), .A1_t (new_AGEMA_signal_2746), .A1_f (new_AGEMA_signal_2747), .B0_t (THETA_n163), .B0_f (new_AGEMA_signal_3285), .B1_t (new_AGEMA_signal_3286), .B1_f (new_AGEMA_signal_3287), .Z0_t (StateFromRhoPi[14]), .Z0_f (new_AGEMA_signal_3533), .Z1_t (new_AGEMA_signal_3534), .Z1_f (new_AGEMA_signal_3535) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U321 ( .A0_t (THETA_n162), .A0_f (new_AGEMA_signal_3045), .A1_t (new_AGEMA_signal_3046), .A1_f (new_AGEMA_signal_3047), .B0_t (THETA_n175), .B0_f (new_AGEMA_signal_3039), .B1_t (new_AGEMA_signal_3040), .B1_f (new_AGEMA_signal_3041), .Z0_t (THETA_n163), .Z0_f (new_AGEMA_signal_3285), .Z1_t (new_AGEMA_signal_3286), .Z1_f (new_AGEMA_signal_3287) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U320 ( .A0_t (StateOut[82]), .A0_f (new_AGEMA_signal_3036), .A1_t (new_AGEMA_signal_3037), .A1_f (new_AGEMA_signal_3038), .B0_t (THETA_n161), .B0_f (new_AGEMA_signal_2883), .B1_t (new_AGEMA_signal_2884), .B1_f (new_AGEMA_signal_2885), .Z0_t (THETA_n175), .Z0_f (new_AGEMA_signal_3039), .Z1_t (new_AGEMA_signal_3040), .Z1_f (new_AGEMA_signal_3041) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U319 ( .A0_t (THETA_n160), .A0_f (new_AGEMA_signal_2235), .A1_t (new_AGEMA_signal_2236), .A1_f (new_AGEMA_signal_2237), .B0_t (THETA_n159), .B0_f (new_AGEMA_signal_2226), .B1_t (new_AGEMA_signal_2227), .B1_f (new_AGEMA_signal_2228), .Z0_t (THETA_n161), .Z0_f (new_AGEMA_signal_2883), .Z1_t (new_AGEMA_signal_2884), .Z1_f (new_AGEMA_signal_2885) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U318 ( .A0_t (StateOut[90]), .A0_f (new_AGEMA_signal_2220), .A1_t (new_AGEMA_signal_2221), .A1_f (new_AGEMA_signal_2222), .B0_t (StateOut[98]), .B0_f (new_AGEMA_signal_2223), .B1_t (new_AGEMA_signal_2224), .B1_f (new_AGEMA_signal_2225), .Z0_t (THETA_n159), .Z0_f (new_AGEMA_signal_2226), .Z1_t (new_AGEMA_signal_2227), .Z1_f (new_AGEMA_signal_2228) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U317 ( .A0_t (StateOut[114]), .A0_f (new_AGEMA_signal_2229), .A1_t (new_AGEMA_signal_2230), .A1_f (new_AGEMA_signal_2231), .B0_t (StateOut[106]), .B0_f (new_AGEMA_signal_2232), .B1_t (new_AGEMA_signal_2233), .B1_f (new_AGEMA_signal_2234), .Z0_t (THETA_n160), .Z0_f (new_AGEMA_signal_2235), .Z1_t (new_AGEMA_signal_2236), .Z1_f (new_AGEMA_signal_2237) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U316 ( .A0_t (StateOut[33]), .A0_f (new_AGEMA_signal_2772), .A1_t (new_AGEMA_signal_2773), .A1_f (new_AGEMA_signal_2774), .B0_t (THETA_n158), .B0_f (new_AGEMA_signal_3288), .B1_t (new_AGEMA_signal_3289), .B1_f (new_AGEMA_signal_3290), .Z0_t (StateFromRhoPi[179]), .Z0_f (new_AGEMA_signal_3536), .Z1_t (new_AGEMA_signal_3537), .Z1_f (new_AGEMA_signal_3538) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U315 ( .A0_t (StateOut[25]), .A0_f (new_AGEMA_signal_2769), .A1_t (new_AGEMA_signal_2770), .A1_f (new_AGEMA_signal_2771), .B0_t (THETA_n158), .B0_f (new_AGEMA_signal_3288), .B1_t (new_AGEMA_signal_3289), .B1_f (new_AGEMA_signal_3290), .Z0_t (StateFromRhoPi[154]), .Z0_f (new_AGEMA_signal_3539), .Z1_t (new_AGEMA_signal_3540), .Z1_f (new_AGEMA_signal_3541) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U314 ( .A0_t (StateOut[17]), .A0_f (new_AGEMA_signal_3216), .A1_t (new_AGEMA_signal_3217), .A1_f (new_AGEMA_signal_3218), .B0_t (THETA_n158), .B0_f (new_AGEMA_signal_3288), .B1_t (new_AGEMA_signal_3289), .B1_f (new_AGEMA_signal_3290), .Z0_t (StateFromRhoPi[92]), .Z0_f (new_AGEMA_signal_3542), .Z1_t (new_AGEMA_signal_3543), .Z1_f (new_AGEMA_signal_3544) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U313 ( .A0_t (StateOut[9]), .A0_f (new_AGEMA_signal_2760), .A1_t (new_AGEMA_signal_2761), .A1_f (new_AGEMA_signal_2762), .B0_t (THETA_n158), .B0_f (new_AGEMA_signal_3288), .B1_t (new_AGEMA_signal_3289), .B1_f (new_AGEMA_signal_3290), .Z0_t (StateFromRhoPi[69]), .Z0_f (new_AGEMA_signal_3545), .Z1_t (new_AGEMA_signal_3546), .Z1_f (new_AGEMA_signal_3547) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U312 ( .A0_t (OutData_s0_t[1]), .A0_f (OutData_s0_f[1]), .A1_t (OutData_s1_t[1]), .A1_f (OutData_s1_f[1]), .B0_t (THETA_n158), .B0_f (new_AGEMA_signal_3288), .B1_t (new_AGEMA_signal_3289), .B1_f (new_AGEMA_signal_3290), .Z0_t (StateFromRhoPi[1]), .Z0_f (new_AGEMA_signal_3548), .Z1_t (new_AGEMA_signal_3549), .Z1_f (new_AGEMA_signal_3550) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U311 ( .A0_t (THETA_n191), .A0_f (new_AGEMA_signal_3051), .A1_t (new_AGEMA_signal_3052), .A1_f (new_AGEMA_signal_3053), .B0_t (THETA_n162), .B0_f (new_AGEMA_signal_3045), .B1_t (new_AGEMA_signal_3046), .B1_f (new_AGEMA_signal_3047), .Z0_t (THETA_n158), .Z0_f (new_AGEMA_signal_3288), .Z1_t (new_AGEMA_signal_3289), .Z1_f (new_AGEMA_signal_3290) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U310 ( .A0_t (StateOut[177]), .A0_f (new_AGEMA_signal_3042), .A1_t (new_AGEMA_signal_3043), .A1_f (new_AGEMA_signal_3044), .B0_t (THETA_n157), .B0_f (new_AGEMA_signal_2886), .B1_t (new_AGEMA_signal_2887), .B1_f (new_AGEMA_signal_2888), .Z0_t (THETA_n162), .Z0_f (new_AGEMA_signal_3045), .Z1_t (new_AGEMA_signal_3046), .Z1_f (new_AGEMA_signal_3047) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U309 ( .A0_t (THETA_n156), .A0_f (new_AGEMA_signal_2253), .A1_t (new_AGEMA_signal_2254), .A1_f (new_AGEMA_signal_2255), .B0_t (THETA_n155), .B0_f (new_AGEMA_signal_2244), .B1_t (new_AGEMA_signal_2245), .B1_f (new_AGEMA_signal_2246), .Z0_t (THETA_n157), .Z0_f (new_AGEMA_signal_2886), .Z1_t (new_AGEMA_signal_2887), .Z1_f (new_AGEMA_signal_2888) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U308 ( .A0_t (StateOut[169]), .A0_f (new_AGEMA_signal_2238), .A1_t (new_AGEMA_signal_2239), .A1_f (new_AGEMA_signal_2240), .B0_t (StateOut[161]), .B0_f (new_AGEMA_signal_2241), .B1_t (new_AGEMA_signal_2242), .B1_f (new_AGEMA_signal_2243), .Z0_t (THETA_n155), .Z0_f (new_AGEMA_signal_2244), .Z1_t (new_AGEMA_signal_2245), .Z1_f (new_AGEMA_signal_2246) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U307 ( .A0_t (StateOut[185]), .A0_f (new_AGEMA_signal_2247), .A1_t (new_AGEMA_signal_2248), .A1_f (new_AGEMA_signal_2249), .B0_t (StateOut[193]), .B0_f (new_AGEMA_signal_2250), .B1_t (new_AGEMA_signal_2251), .B1_f (new_AGEMA_signal_2252), .Z0_t (THETA_n156), .Z0_f (new_AGEMA_signal_2253), .Z1_t (new_AGEMA_signal_2254), .Z1_f (new_AGEMA_signal_2255) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U306 ( .A0_t (StateOut[64]), .A0_f (new_AGEMA_signal_3048), .A1_t (new_AGEMA_signal_3049), .A1_f (new_AGEMA_signal_3050), .B0_t (THETA_n154), .B0_f (new_AGEMA_signal_2889), .B1_t (new_AGEMA_signal_2890), .B1_f (new_AGEMA_signal_2891), .Z0_t (THETA_n191), .Z0_f (new_AGEMA_signal_3051), .Z1_t (new_AGEMA_signal_3052), .Z1_f (new_AGEMA_signal_3053) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U305 ( .A0_t (THETA_n153), .A0_f (new_AGEMA_signal_2271), .A1_t (new_AGEMA_signal_2272), .A1_f (new_AGEMA_signal_2273), .B0_t (THETA_n152), .B0_f (new_AGEMA_signal_2262), .B1_t (new_AGEMA_signal_2263), .B1_f (new_AGEMA_signal_2264), .Z0_t (THETA_n154), .Z0_f (new_AGEMA_signal_2889), .Z1_t (new_AGEMA_signal_2890), .Z1_f (new_AGEMA_signal_2891) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U304 ( .A0_t (StateOut[48]), .A0_f (new_AGEMA_signal_2256), .A1_t (new_AGEMA_signal_2257), .A1_f (new_AGEMA_signal_2258), .B0_t (StateOut[40]), .B0_f (new_AGEMA_signal_2259), .B1_t (new_AGEMA_signal_2260), .B1_f (new_AGEMA_signal_2261), .Z0_t (THETA_n152), .Z0_f (new_AGEMA_signal_2262), .Z1_t (new_AGEMA_signal_2263), .Z1_f (new_AGEMA_signal_2264) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U303 ( .A0_t (StateOut[72]), .A0_f (new_AGEMA_signal_2265), .A1_t (new_AGEMA_signal_2266), .A1_f (new_AGEMA_signal_2267), .B0_t (StateOut[56]), .B0_f (new_AGEMA_signal_2268), .B1_t (new_AGEMA_signal_2269), .B1_f (new_AGEMA_signal_2270), .Z0_t (THETA_n153), .Z0_f (new_AGEMA_signal_2271), .Z1_t (new_AGEMA_signal_2272), .Z1_f (new_AGEMA_signal_2273) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U302 ( .A0_t (StateOut[114]), .A0_f (new_AGEMA_signal_2229), .A1_t (new_AGEMA_signal_2230), .A1_f (new_AGEMA_signal_2231), .B0_t (THETA_n151), .B0_f (new_AGEMA_signal_3291), .B1_t (new_AGEMA_signal_3292), .B1_f (new_AGEMA_signal_3293), .Z0_t (StateFromRhoPi[175]), .Z0_f (new_AGEMA_signal_3551), .Z1_t (new_AGEMA_signal_3552), .Z1_f (new_AGEMA_signal_3553) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U301 ( .A0_t (StateOut[106]), .A0_f (new_AGEMA_signal_2232), .A1_t (new_AGEMA_signal_2233), .A1_f (new_AGEMA_signal_2234), .B0_t (THETA_n151), .B0_f (new_AGEMA_signal_3291), .B1_t (new_AGEMA_signal_3292), .B1_f (new_AGEMA_signal_3293), .Z0_t (StateFromRhoPi[145]), .Z0_f (new_AGEMA_signal_3554), .Z1_t (new_AGEMA_signal_3555), .Z1_f (new_AGEMA_signal_3556) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U300 ( .A0_t (StateOut[98]), .A0_f (new_AGEMA_signal_2223), .A1_t (new_AGEMA_signal_2224), .A1_f (new_AGEMA_signal_2225), .B0_t (THETA_n151), .B0_f (new_AGEMA_signal_3291), .B1_t (new_AGEMA_signal_3292), .B1_f (new_AGEMA_signal_3293), .Z0_t (StateFromRhoPi[85]), .Z0_f (new_AGEMA_signal_3557), .Z1_t (new_AGEMA_signal_3558), .Z1_f (new_AGEMA_signal_3559) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U299 ( .A0_t (StateOut[90]), .A0_f (new_AGEMA_signal_2220), .A1_t (new_AGEMA_signal_2221), .A1_f (new_AGEMA_signal_2222), .B0_t (THETA_n151), .B0_f (new_AGEMA_signal_3291), .B1_t (new_AGEMA_signal_3292), .B1_f (new_AGEMA_signal_3293), .Z0_t (StateFromRhoPi[56]), .Z0_f (new_AGEMA_signal_3560), .Z1_t (new_AGEMA_signal_3561), .Z1_f (new_AGEMA_signal_3562) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U298 ( .A0_t (StateOut[82]), .A0_f (new_AGEMA_signal_3036), .A1_t (new_AGEMA_signal_3037), .A1_f (new_AGEMA_signal_3038), .B0_t (THETA_n151), .B0_f (new_AGEMA_signal_3291), .B1_t (new_AGEMA_signal_3292), .B1_f (new_AGEMA_signal_3293), .Z0_t (StateFromRhoPi[32]), .Z0_f (new_AGEMA_signal_3563), .Z1_t (new_AGEMA_signal_3564), .Z1_f (new_AGEMA_signal_3565) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U297 ( .A0_t (THETA_n150), .A0_f (new_AGEMA_signal_3183), .A1_t (new_AGEMA_signal_3184), .A1_f (new_AGEMA_signal_3185), .B0_t (THETA_n170), .B0_f (new_AGEMA_signal_3057), .B1_t (new_AGEMA_signal_3058), .B1_f (new_AGEMA_signal_3059), .Z0_t (THETA_n151), .Z0_f (new_AGEMA_signal_3291), .Z1_t (new_AGEMA_signal_3292), .Z1_f (new_AGEMA_signal_3293) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U296 ( .A0_t (StateOut[121]), .A0_f (new_AGEMA_signal_3054), .A1_t (new_AGEMA_signal_3055), .A1_f (new_AGEMA_signal_3056), .B0_t (THETA_n149), .B0_f (new_AGEMA_signal_2892), .B1_t (new_AGEMA_signal_2893), .B1_f (new_AGEMA_signal_2894), .Z0_t (THETA_n170), .Z0_f (new_AGEMA_signal_3057), .Z1_t (new_AGEMA_signal_3058), .Z1_f (new_AGEMA_signal_3059) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U295 ( .A0_t (THETA_n148), .A0_f (new_AGEMA_signal_2289), .A1_t (new_AGEMA_signal_2290), .A1_f (new_AGEMA_signal_2291), .B0_t (THETA_n147), .B0_f (new_AGEMA_signal_2280), .B1_t (new_AGEMA_signal_2281), .B1_f (new_AGEMA_signal_2282), .Z0_t (THETA_n149), .Z0_f (new_AGEMA_signal_2892), .Z1_t (new_AGEMA_signal_2893), .Z1_f (new_AGEMA_signal_2894) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U294 ( .A0_t (StateOut[129]), .A0_f (new_AGEMA_signal_2274), .A1_t (new_AGEMA_signal_2275), .A1_f (new_AGEMA_signal_2276), .B0_t (StateOut[137]), .B0_f (new_AGEMA_signal_2277), .B1_t (new_AGEMA_signal_2278), .B1_f (new_AGEMA_signal_2279), .Z0_t (THETA_n147), .Z0_f (new_AGEMA_signal_2280), .Z1_t (new_AGEMA_signal_2281), .Z1_f (new_AGEMA_signal_2282) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U293 ( .A0_t (StateOut[153]), .A0_f (new_AGEMA_signal_2283), .A1_t (new_AGEMA_signal_2284), .A1_f (new_AGEMA_signal_2285), .B0_t (StateOut[145]), .B0_f (new_AGEMA_signal_2286), .B1_t (new_AGEMA_signal_2287), .B1_f (new_AGEMA_signal_2288), .Z0_t (THETA_n148), .Z0_f (new_AGEMA_signal_2289), .Z1_t (new_AGEMA_signal_2290), .Z1_f (new_AGEMA_signal_2291) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U292 ( .A0_t (StateOut[153]), .A0_f (new_AGEMA_signal_2283), .A1_t (new_AGEMA_signal_2284), .A1_f (new_AGEMA_signal_2285), .B0_t (THETA_n146), .B0_f (new_AGEMA_signal_3294), .B1_t (new_AGEMA_signal_3295), .B1_f (new_AGEMA_signal_3296), .Z0_t (StateFromRhoPi[185]), .Z0_f (new_AGEMA_signal_3566), .Z1_t (new_AGEMA_signal_3567), .Z1_f (new_AGEMA_signal_3568) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U291 ( .A0_t (StateOut[145]), .A0_f (new_AGEMA_signal_2286), .A1_t (new_AGEMA_signal_2287), .A1_f (new_AGEMA_signal_2288), .B0_t (THETA_n146), .B0_f (new_AGEMA_signal_3294), .B1_t (new_AGEMA_signal_3295), .B1_f (new_AGEMA_signal_3296), .Z0_t (StateFromRhoPi[126]), .Z0_f (new_AGEMA_signal_3569), .Z1_t (new_AGEMA_signal_3570), .Z1_f (new_AGEMA_signal_3571) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U290 ( .A0_t (StateOut[137]), .A0_f (new_AGEMA_signal_2277), .A1_t (new_AGEMA_signal_2278), .A1_f (new_AGEMA_signal_2279), .B0_t (THETA_n146), .B0_f (new_AGEMA_signal_3294), .B1_t (new_AGEMA_signal_3295), .B1_f (new_AGEMA_signal_3296), .Z0_t (StateFromRhoPi[98]), .Z0_f (new_AGEMA_signal_3572), .Z1_t (new_AGEMA_signal_3573), .Z1_f (new_AGEMA_signal_3574) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U289 ( .A0_t (StateOut[129]), .A0_f (new_AGEMA_signal_2274), .A1_t (new_AGEMA_signal_2275), .A1_f (new_AGEMA_signal_2276), .B0_t (THETA_n146), .B0_f (new_AGEMA_signal_3294), .B1_t (new_AGEMA_signal_3295), .B1_f (new_AGEMA_signal_3296), .Z0_t (StateFromRhoPi[72]), .Z0_f (new_AGEMA_signal_3575), .Z1_t (new_AGEMA_signal_3576), .Z1_f (new_AGEMA_signal_3577) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U288 ( .A0_t (StateOut[121]), .A0_f (new_AGEMA_signal_3054), .A1_t (new_AGEMA_signal_3055), .A1_f (new_AGEMA_signal_3056), .B0_t (THETA_n146), .B0_f (new_AGEMA_signal_3294), .B1_t (new_AGEMA_signal_3295), .B1_f (new_AGEMA_signal_3296), .Z0_t (StateFromRhoPi[13]), .Z0_f (new_AGEMA_signal_3578), .Z1_t (new_AGEMA_signal_3579), .Z1_f (new_AGEMA_signal_3580) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U287 ( .A0_t (THETA_n145), .A0_f (new_AGEMA_signal_3069), .A1_t (new_AGEMA_signal_3070), .A1_f (new_AGEMA_signal_3071), .B0_t (THETA_n144), .B0_f (new_AGEMA_signal_3063), .B1_t (new_AGEMA_signal_3064), .B1_f (new_AGEMA_signal_3065), .Z0_t (THETA_n146), .Z0_f (new_AGEMA_signal_3294), .Z1_t (new_AGEMA_signal_3295), .Z1_f (new_AGEMA_signal_3296) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U286 ( .A0_t (StateOut[74]), .A0_f (new_AGEMA_signal_2661), .A1_t (new_AGEMA_signal_2662), .A1_f (new_AGEMA_signal_2663), .B0_t (THETA_n143), .B0_f (new_AGEMA_signal_3297), .B1_t (new_AGEMA_signal_3298), .B1_f (new_AGEMA_signal_3299), .Z0_t (StateFromRhoPi[196]), .Z0_f (new_AGEMA_signal_3581), .Z1_t (new_AGEMA_signal_3582), .Z1_f (new_AGEMA_signal_3583) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U285 ( .A0_t (StateOut[66]), .A0_f (new_AGEMA_signal_3180), .A1_t (new_AGEMA_signal_3181), .A1_f (new_AGEMA_signal_3182), .B0_t (THETA_n143), .B0_f (new_AGEMA_signal_3297), .B1_t (new_AGEMA_signal_3298), .B1_f (new_AGEMA_signal_3299), .Z0_t (StateFromRhoPi[135]), .Z0_f (new_AGEMA_signal_3584), .Z1_t (new_AGEMA_signal_3585), .Z1_f (new_AGEMA_signal_3586) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U284 ( .A0_t (StateOut[58]), .A0_f (new_AGEMA_signal_2664), .A1_t (new_AGEMA_signal_2665), .A1_f (new_AGEMA_signal_2666), .B0_t (THETA_n143), .B0_f (new_AGEMA_signal_3297), .B1_t (new_AGEMA_signal_3298), .B1_f (new_AGEMA_signal_3299), .Z0_t (StateFromRhoPi[108]), .Z0_f (new_AGEMA_signal_3587), .Z1_t (new_AGEMA_signal_3588), .Z1_f (new_AGEMA_signal_3589) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U283 ( .A0_t (StateOut[50]), .A0_f (new_AGEMA_signal_2652), .A1_t (new_AGEMA_signal_2653), .A1_f (new_AGEMA_signal_2654), .B0_t (THETA_n143), .B0_f (new_AGEMA_signal_3297), .B1_t (new_AGEMA_signal_3298), .B1_f (new_AGEMA_signal_3299), .Z0_t (StateFromRhoPi[46]), .Z0_f (new_AGEMA_signal_3590), .Z1_t (new_AGEMA_signal_3591), .Z1_f (new_AGEMA_signal_3592) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U282 ( .A0_t (StateOut[42]), .A0_f (new_AGEMA_signal_2655), .A1_t (new_AGEMA_signal_2656), .A1_f (new_AGEMA_signal_2657), .B0_t (THETA_n143), .B0_f (new_AGEMA_signal_3297), .B1_t (new_AGEMA_signal_3298), .B1_f (new_AGEMA_signal_3299), .Z0_t (StateFromRhoPi[19]), .Z0_f (new_AGEMA_signal_3593), .Z1_t (new_AGEMA_signal_3594), .Z1_f (new_AGEMA_signal_3595) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U281 ( .A0_t (THETA_n142), .A0_f (new_AGEMA_signal_3141), .A1_t (new_AGEMA_signal_3142), .A1_f (new_AGEMA_signal_3143), .B0_t (THETA_n144), .B0_f (new_AGEMA_signal_3063), .B1_t (new_AGEMA_signal_3064), .B1_f (new_AGEMA_signal_3065), .Z0_t (THETA_n143), .Z0_f (new_AGEMA_signal_3297), .Z1_t (new_AGEMA_signal_3298), .Z1_f (new_AGEMA_signal_3299) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U280 ( .A0_t (StateOut[81]), .A0_f (new_AGEMA_signal_3060), .A1_t (new_AGEMA_signal_3061), .A1_f (new_AGEMA_signal_3062), .B0_t (THETA_n141), .B0_f (new_AGEMA_signal_2895), .B1_t (new_AGEMA_signal_2896), .B1_f (new_AGEMA_signal_2897), .Z0_t (THETA_n144), .Z0_f (new_AGEMA_signal_3063), .Z1_t (new_AGEMA_signal_3064), .Z1_f (new_AGEMA_signal_3065) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U279 ( .A0_t (THETA_n140), .A0_f (new_AGEMA_signal_2307), .A1_t (new_AGEMA_signal_2308), .A1_f (new_AGEMA_signal_2309), .B0_t (THETA_n139), .B0_f (new_AGEMA_signal_2298), .B1_t (new_AGEMA_signal_2299), .B1_f (new_AGEMA_signal_2300), .Z0_t (THETA_n141), .Z0_f (new_AGEMA_signal_2895), .Z1_t (new_AGEMA_signal_2896), .Z1_f (new_AGEMA_signal_2897) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U278 ( .A0_t (StateOut[89]), .A0_f (new_AGEMA_signal_2292), .A1_t (new_AGEMA_signal_2293), .A1_f (new_AGEMA_signal_2294), .B0_t (StateOut[97]), .B0_f (new_AGEMA_signal_2295), .B1_t (new_AGEMA_signal_2296), .B1_f (new_AGEMA_signal_2297), .Z0_t (THETA_n139), .Z0_f (new_AGEMA_signal_2298), .Z1_t (new_AGEMA_signal_2299), .Z1_f (new_AGEMA_signal_2300) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U277 ( .A0_t (StateOut[113]), .A0_f (new_AGEMA_signal_2301), .A1_t (new_AGEMA_signal_2302), .A1_f (new_AGEMA_signal_2303), .B0_t (StateOut[105]), .B0_f (new_AGEMA_signal_2304), .B1_t (new_AGEMA_signal_2305), .B1_f (new_AGEMA_signal_2306), .Z0_t (THETA_n140), .Z0_f (new_AGEMA_signal_2307), .Z1_t (new_AGEMA_signal_2308), .Z1_f (new_AGEMA_signal_2309) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U276 ( .A0_t (StateOut[32]), .A0_f (new_AGEMA_signal_2211), .A1_t (new_AGEMA_signal_2212), .A1_f (new_AGEMA_signal_2213), .B0_t (THETA_n138), .B0_f (new_AGEMA_signal_3300), .B1_t (new_AGEMA_signal_3301), .B1_f (new_AGEMA_signal_3302), .Z0_t (StateFromRhoPi[178]), .Z0_f (new_AGEMA_signal_3596), .Z1_t (new_AGEMA_signal_3597), .Z1_f (new_AGEMA_signal_3598) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U275 ( .A0_t (StateOut[24]), .A0_f (new_AGEMA_signal_2214), .A1_t (new_AGEMA_signal_2215), .A1_f (new_AGEMA_signal_2216), .B0_t (THETA_n138), .B0_f (new_AGEMA_signal_3300), .B1_t (new_AGEMA_signal_3301), .B1_f (new_AGEMA_signal_3302), .Z0_t (StateFromRhoPi[153]), .Z0_f (new_AGEMA_signal_3599), .Z1_t (new_AGEMA_signal_3600), .Z1_f (new_AGEMA_signal_3601) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U274 ( .A0_t (StateOut[16]), .A0_f (new_AGEMA_signal_2205), .A1_t (new_AGEMA_signal_2206), .A1_f (new_AGEMA_signal_2207), .B0_t (THETA_n138), .B0_f (new_AGEMA_signal_3300), .B1_t (new_AGEMA_signal_3301), .B1_f (new_AGEMA_signal_3302), .Z0_t (StateFromRhoPi[91]), .Z0_f (new_AGEMA_signal_3602), .Z1_t (new_AGEMA_signal_3603), .Z1_f (new_AGEMA_signal_3604) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U273 ( .A0_t (StateOut[8]), .A0_f (new_AGEMA_signal_2202), .A1_t (new_AGEMA_signal_2203), .A1_f (new_AGEMA_signal_2204), .B0_t (THETA_n138), .B0_f (new_AGEMA_signal_3300), .B1_t (new_AGEMA_signal_3301), .B1_f (new_AGEMA_signal_3302), .Z0_t (StateFromRhoPi[68]), .Z0_f (new_AGEMA_signal_3605), .Z1_t (new_AGEMA_signal_3606), .Z1_f (new_AGEMA_signal_3607) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U272 ( .A0_t (OutData_s0_t[0]), .A0_f (OutData_s0_f[0]), .A1_t (OutData_s1_t[0]), .A1_f (OutData_s1_f[0]), .B0_t (THETA_n138), .B0_f (new_AGEMA_signal_3300), .B1_t (new_AGEMA_signal_3301), .B1_f (new_AGEMA_signal_3302), .Z0_t (StateFromRhoPi[0]), .Z0_f (new_AGEMA_signal_3608), .Z1_t (new_AGEMA_signal_3609), .Z1_f (new_AGEMA_signal_3610) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U271 ( .A0_t (THETA_n183), .A0_f (new_AGEMA_signal_3075), .A1_t (new_AGEMA_signal_3076), .A1_f (new_AGEMA_signal_3077), .B0_t (THETA_n145), .B0_f (new_AGEMA_signal_3069), .B1_t (new_AGEMA_signal_3070), .B1_f (new_AGEMA_signal_3071), .Z0_t (THETA_n138), .Z0_f (new_AGEMA_signal_3300), .Z1_t (new_AGEMA_signal_3301), .Z1_f (new_AGEMA_signal_3302) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U270 ( .A0_t (StateOut[160]), .A0_f (new_AGEMA_signal_3066), .A1_t (new_AGEMA_signal_3067), .A1_f (new_AGEMA_signal_3068), .B0_t (THETA_n137), .B0_f (new_AGEMA_signal_2898), .B1_t (new_AGEMA_signal_2899), .B1_f (new_AGEMA_signal_2900), .Z0_t (THETA_n145), .Z0_f (new_AGEMA_signal_3069), .Z1_t (new_AGEMA_signal_3070), .Z1_f (new_AGEMA_signal_3071) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U269 ( .A0_t (THETA_n136), .A0_f (new_AGEMA_signal_2325), .A1_t (new_AGEMA_signal_2326), .A1_f (new_AGEMA_signal_2327), .B0_t (THETA_n135), .B0_f (new_AGEMA_signal_2316), .B1_t (new_AGEMA_signal_2317), .B1_f (new_AGEMA_signal_2318), .Z0_t (THETA_n137), .Z0_f (new_AGEMA_signal_2898), .Z1_t (new_AGEMA_signal_2899), .Z1_f (new_AGEMA_signal_2900) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U268 ( .A0_t (StateOut[168]), .A0_f (new_AGEMA_signal_2310), .A1_t (new_AGEMA_signal_2311), .A1_f (new_AGEMA_signal_2312), .B0_t (StateOut[176]), .B0_f (new_AGEMA_signal_2313), .B1_t (new_AGEMA_signal_2314), .B1_f (new_AGEMA_signal_2315), .Z0_t (THETA_n135), .Z0_f (new_AGEMA_signal_2316), .Z1_t (new_AGEMA_signal_2317), .Z1_f (new_AGEMA_signal_2318) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U267 ( .A0_t (StateOut[192]), .A0_f (new_AGEMA_signal_2319), .A1_t (new_AGEMA_signal_2320), .A1_f (new_AGEMA_signal_2321), .B0_t (StateOut[184]), .B0_f (new_AGEMA_signal_2322), .B1_t (new_AGEMA_signal_2323), .B1_f (new_AGEMA_signal_2324), .Z0_t (THETA_n136), .Z0_f (new_AGEMA_signal_2325), .Z1_t (new_AGEMA_signal_2326), .Z1_f (new_AGEMA_signal_2327) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U266 ( .A0_t (StateOut[47]), .A0_f (new_AGEMA_signal_3072), .A1_t (new_AGEMA_signal_3073), .A1_f (new_AGEMA_signal_3074), .B0_t (THETA_n134), .B0_f (new_AGEMA_signal_2901), .B1_t (new_AGEMA_signal_2902), .B1_f (new_AGEMA_signal_2903), .Z0_t (THETA_n183), .Z0_f (new_AGEMA_signal_3075), .Z1_t (new_AGEMA_signal_3076), .Z1_f (new_AGEMA_signal_3077) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U265 ( .A0_t (THETA_n133), .A0_f (new_AGEMA_signal_2343), .A1_t (new_AGEMA_signal_2344), .A1_f (new_AGEMA_signal_2345), .B0_t (THETA_n132), .B0_f (new_AGEMA_signal_2334), .B1_t (new_AGEMA_signal_2335), .B1_f (new_AGEMA_signal_2336), .Z0_t (THETA_n134), .Z0_f (new_AGEMA_signal_2901), .Z1_t (new_AGEMA_signal_2902), .Z1_f (new_AGEMA_signal_2903) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U264 ( .A0_t (StateOut[55]), .A0_f (new_AGEMA_signal_2328), .A1_t (new_AGEMA_signal_2329), .A1_f (new_AGEMA_signal_2330), .B0_t (StateOut[63]), .B0_f (new_AGEMA_signal_2331), .B1_t (new_AGEMA_signal_2332), .B1_f (new_AGEMA_signal_2333), .Z0_t (THETA_n132), .Z0_f (new_AGEMA_signal_2334), .Z1_t (new_AGEMA_signal_2335), .Z1_f (new_AGEMA_signal_2336) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U263 ( .A0_t (StateOut[79]), .A0_f (new_AGEMA_signal_2337), .A1_t (new_AGEMA_signal_2338), .A1_f (new_AGEMA_signal_2339), .B0_t (StateOut[71]), .B0_f (new_AGEMA_signal_2340), .B1_t (new_AGEMA_signal_2341), .B1_f (new_AGEMA_signal_2342), .Z0_t (THETA_n133), .Z0_f (new_AGEMA_signal_2343), .Z1_t (new_AGEMA_signal_2344), .Z1_f (new_AGEMA_signal_2345) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U262 ( .A0_t (StateOut[192]), .A0_f (new_AGEMA_signal_2319), .A1_t (new_AGEMA_signal_2320), .A1_f (new_AGEMA_signal_2321), .B0_t (THETA_n131), .B0_f (new_AGEMA_signal_3303), .B1_t (new_AGEMA_signal_3304), .B1_f (new_AGEMA_signal_3305), .Z0_t (StateFromRhoPi[166]), .Z0_f (new_AGEMA_signal_3611), .Z1_t (new_AGEMA_signal_3612), .Z1_f (new_AGEMA_signal_3613) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U261 ( .A0_t (StateOut[184]), .A0_f (new_AGEMA_signal_2322), .A1_t (new_AGEMA_signal_2323), .A1_f (new_AGEMA_signal_2324), .B0_t (THETA_n131), .B0_f (new_AGEMA_signal_3303), .B1_t (new_AGEMA_signal_3304), .B1_f (new_AGEMA_signal_3305), .Z0_t (StateFromRhoPi[136]), .Z0_f (new_AGEMA_signal_3614), .Z1_t (new_AGEMA_signal_3615), .Z1_f (new_AGEMA_signal_3616) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U260 ( .A0_t (StateOut[176]), .A0_f (new_AGEMA_signal_2313), .A1_t (new_AGEMA_signal_2314), .A1_f (new_AGEMA_signal_2315), .B0_t (THETA_n131), .B0_f (new_AGEMA_signal_3303), .B1_t (new_AGEMA_signal_3304), .B1_f (new_AGEMA_signal_3305), .Z0_t (StateFromRhoPi[119]), .Z0_f (new_AGEMA_signal_3617), .Z1_t (new_AGEMA_signal_3618), .Z1_f (new_AGEMA_signal_3619) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U259 ( .A0_t (StateOut[168]), .A0_f (new_AGEMA_signal_2310), .A1_t (new_AGEMA_signal_2311), .A1_f (new_AGEMA_signal_2312), .B0_t (THETA_n131), .B0_f (new_AGEMA_signal_3303), .B1_t (new_AGEMA_signal_3304), .B1_f (new_AGEMA_signal_3305), .Z0_t (StateFromRhoPi[52]), .Z0_f (new_AGEMA_signal_3620), .Z1_t (new_AGEMA_signal_3621), .Z1_f (new_AGEMA_signal_3622) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U258 ( .A0_t (StateOut[160]), .A0_f (new_AGEMA_signal_3066), .A1_t (new_AGEMA_signal_3067), .A1_f (new_AGEMA_signal_3068), .B0_t (THETA_n131), .B0_f (new_AGEMA_signal_3303), .B1_t (new_AGEMA_signal_3304), .B1_f (new_AGEMA_signal_3305), .Z0_t (StateFromRhoPi[27]), .Z0_f (new_AGEMA_signal_3623), .Z1_t (new_AGEMA_signal_3624), .Z1_f (new_AGEMA_signal_3625) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U257 ( .A0_t (THETA_n130), .A0_f (new_AGEMA_signal_3099), .A1_t (new_AGEMA_signal_3100), .A1_f (new_AGEMA_signal_3101), .B0_t (THETA_n129), .B0_f (new_AGEMA_signal_3081), .B1_t (new_AGEMA_signal_3082), .B1_f (new_AGEMA_signal_3083), .Z0_t (THETA_n131), .Z0_f (new_AGEMA_signal_3303), .Z1_t (new_AGEMA_signal_3304), .Z1_f (new_AGEMA_signal_3305) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U256 ( .A0_t (StateOut[79]), .A0_f (new_AGEMA_signal_2337), .A1_t (new_AGEMA_signal_2338), .A1_f (new_AGEMA_signal_2339), .B0_t (THETA_n128), .B0_f (new_AGEMA_signal_3306), .B1_t (new_AGEMA_signal_3307), .B1_f (new_AGEMA_signal_3308), .Z0_t (StateFromRhoPi[193]), .Z0_f (new_AGEMA_signal_3626), .Z1_t (new_AGEMA_signal_3627), .Z1_f (new_AGEMA_signal_3628) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U255 ( .A0_t (StateOut[71]), .A0_f (new_AGEMA_signal_2340), .A1_t (new_AGEMA_signal_2341), .A1_f (new_AGEMA_signal_2342), .B0_t (THETA_n128), .B0_f (new_AGEMA_signal_3306), .B1_t (new_AGEMA_signal_3307), .B1_f (new_AGEMA_signal_3308), .Z0_t (StateFromRhoPi[132]), .Z0_f (new_AGEMA_signal_3629), .Z1_t (new_AGEMA_signal_3630), .Z1_f (new_AGEMA_signal_3631) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U254 ( .A0_t (StateOut[63]), .A0_f (new_AGEMA_signal_2331), .A1_t (new_AGEMA_signal_2332), .A1_f (new_AGEMA_signal_2333), .B0_t (THETA_n128), .B0_f (new_AGEMA_signal_3306), .B1_t (new_AGEMA_signal_3307), .B1_f (new_AGEMA_signal_3308), .Z0_t (StateFromRhoPi[105]), .Z0_f (new_AGEMA_signal_3632), .Z1_t (new_AGEMA_signal_3633), .Z1_f (new_AGEMA_signal_3634) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U253 ( .A0_t (StateOut[55]), .A0_f (new_AGEMA_signal_2328), .A1_t (new_AGEMA_signal_2329), .A1_f (new_AGEMA_signal_2330), .B0_t (THETA_n128), .B0_f (new_AGEMA_signal_3306), .B1_t (new_AGEMA_signal_3307), .B1_f (new_AGEMA_signal_3308), .Z0_t (StateFromRhoPi[43]), .Z0_f (new_AGEMA_signal_3635), .Z1_t (new_AGEMA_signal_3636), .Z1_f (new_AGEMA_signal_3637) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U252 ( .A0_t (StateOut[47]), .A0_f (new_AGEMA_signal_3072), .A1_t (new_AGEMA_signal_3073), .A1_f (new_AGEMA_signal_3074), .B0_t (THETA_n128), .B0_f (new_AGEMA_signal_3306), .B1_t (new_AGEMA_signal_3307), .B1_f (new_AGEMA_signal_3308), .Z0_t (StateFromRhoPi[16]), .Z0_f (new_AGEMA_signal_3638), .Z1_t (new_AGEMA_signal_3639), .Z1_f (new_AGEMA_signal_3640) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U251 ( .A0_t (THETA_n127), .A0_f (new_AGEMA_signal_3195), .A1_t (new_AGEMA_signal_3196), .A1_f (new_AGEMA_signal_3197), .B0_t (THETA_n129), .B0_f (new_AGEMA_signal_3081), .B1_t (new_AGEMA_signal_3082), .B1_f (new_AGEMA_signal_3083), .Z0_t (THETA_n128), .Z0_f (new_AGEMA_signal_3306), .Z1_t (new_AGEMA_signal_3307), .Z1_f (new_AGEMA_signal_3308) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U250 ( .A0_t (OutData_s0_t[7]), .A0_f (OutData_s0_f[7]), .A1_t (OutData_s1_t[7]), .A1_f (OutData_s1_f[7]), .B0_t (THETA_n126), .B0_f (new_AGEMA_signal_2904), .B1_t (new_AGEMA_signal_2905), .B1_f (new_AGEMA_signal_2906), .Z0_t (THETA_n129), .Z0_f (new_AGEMA_signal_3081), .Z1_t (new_AGEMA_signal_3082), .Z1_f (new_AGEMA_signal_3083) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U249 ( .A0_t (THETA_n125), .A0_f (new_AGEMA_signal_2361), .A1_t (new_AGEMA_signal_2362), .A1_f (new_AGEMA_signal_2363), .B0_t (THETA_n124), .B0_f (new_AGEMA_signal_2352), .B1_t (new_AGEMA_signal_2353), .B1_f (new_AGEMA_signal_2354), .Z0_t (THETA_n126), .Z0_f (new_AGEMA_signal_2904), .Z1_t (new_AGEMA_signal_2905), .Z1_f (new_AGEMA_signal_2906) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U248 ( .A0_t (StateOut[15]), .A0_f (new_AGEMA_signal_2346), .A1_t (new_AGEMA_signal_2347), .A1_f (new_AGEMA_signal_2348), .B0_t (StateOut[23]), .B0_f (new_AGEMA_signal_2349), .B1_t (new_AGEMA_signal_2350), .B1_f (new_AGEMA_signal_2351), .Z0_t (THETA_n124), .Z0_f (new_AGEMA_signal_2352), .Z1_t (new_AGEMA_signal_2353), .Z1_f (new_AGEMA_signal_2354) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U247 ( .A0_t (StateOut[39]), .A0_f (new_AGEMA_signal_2355), .A1_t (new_AGEMA_signal_2356), .A1_f (new_AGEMA_signal_2357), .B0_t (StateOut[31]), .B0_f (new_AGEMA_signal_2358), .B1_t (new_AGEMA_signal_2359), .B1_f (new_AGEMA_signal_2360), .Z0_t (THETA_n125), .Z0_f (new_AGEMA_signal_2361), .Z1_t (new_AGEMA_signal_2362), .Z1_f (new_AGEMA_signal_2363) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U246 ( .A0_t (StateOut[117]), .A0_f (new_AGEMA_signal_2733), .A1_t (new_AGEMA_signal_2734), .A1_f (new_AGEMA_signal_2735), .B0_t (THETA_n123), .B0_f (new_AGEMA_signal_3309), .B1_t (new_AGEMA_signal_3310), .B1_f (new_AGEMA_signal_3311), .Z0_t (StateFromRhoPi[170]), .Z0_f (new_AGEMA_signal_3641), .Z1_t (new_AGEMA_signal_3642), .Z1_f (new_AGEMA_signal_3643) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U245 ( .A0_t (StateOut[109]), .A0_f (new_AGEMA_signal_3204), .A1_t (new_AGEMA_signal_3205), .A1_f (new_AGEMA_signal_3206), .B0_t (THETA_n123), .B0_f (new_AGEMA_signal_3309), .B1_t (new_AGEMA_signal_3310), .B1_f (new_AGEMA_signal_3311), .Z0_t (StateFromRhoPi[148]), .Z0_f (new_AGEMA_signal_3644), .Z1_t (new_AGEMA_signal_3645), .Z1_f (new_AGEMA_signal_3646) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U244 ( .A0_t (StateOut[101]), .A0_f (new_AGEMA_signal_2736), .A1_t (new_AGEMA_signal_2737), .A1_f (new_AGEMA_signal_2738), .B0_t (THETA_n123), .B0_f (new_AGEMA_signal_3309), .B1_t (new_AGEMA_signal_3310), .B1_f (new_AGEMA_signal_3311), .Z0_t (StateFromRhoPi[80]), .Z0_f (new_AGEMA_signal_3647), .Z1_t (new_AGEMA_signal_3648), .Z1_f (new_AGEMA_signal_3649) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U243 ( .A0_t (StateOut[93]), .A0_f (new_AGEMA_signal_2724), .A1_t (new_AGEMA_signal_2725), .A1_f (new_AGEMA_signal_2726), .B0_t (THETA_n123), .B0_f (new_AGEMA_signal_3309), .B1_t (new_AGEMA_signal_3310), .B1_f (new_AGEMA_signal_3311), .Z0_t (StateFromRhoPi[59]), .Z0_f (new_AGEMA_signal_3650), .Z1_t (new_AGEMA_signal_3651), .Z1_f (new_AGEMA_signal_3652) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U242 ( .A0_t (StateOut[85]), .A0_f (new_AGEMA_signal_2727), .A1_t (new_AGEMA_signal_2728), .A1_f (new_AGEMA_signal_2729), .B0_t (THETA_n123), .B0_f (new_AGEMA_signal_3309), .B1_t (new_AGEMA_signal_3310), .B1_f (new_AGEMA_signal_3311), .Z0_t (StateFromRhoPi[35]), .Z0_f (new_AGEMA_signal_3653), .Z1_t (new_AGEMA_signal_3654), .Z1_f (new_AGEMA_signal_3655) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U241 ( .A0_t (THETA_n122), .A0_f (new_AGEMA_signal_3135), .A1_t (new_AGEMA_signal_3136), .A1_f (new_AGEMA_signal_3137), .B0_t (THETA_n178), .B0_f (new_AGEMA_signal_3087), .B1_t (new_AGEMA_signal_3088), .B1_f (new_AGEMA_signal_3089), .Z0_t (THETA_n123), .Z0_f (new_AGEMA_signal_3309), .Z1_t (new_AGEMA_signal_3310), .Z1_f (new_AGEMA_signal_3311) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U240 ( .A0_t (StateOut[124]), .A0_f (new_AGEMA_signal_3084), .A1_t (new_AGEMA_signal_3085), .A1_f (new_AGEMA_signal_3086), .B0_t (THETA_n121), .B0_f (new_AGEMA_signal_2907), .B1_t (new_AGEMA_signal_2908), .B1_f (new_AGEMA_signal_2909), .Z0_t (THETA_n178), .Z0_f (new_AGEMA_signal_3087), .Z1_t (new_AGEMA_signal_3088), .Z1_f (new_AGEMA_signal_3089) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U239 ( .A0_t (THETA_n120), .A0_f (new_AGEMA_signal_2379), .A1_t (new_AGEMA_signal_2380), .A1_f (new_AGEMA_signal_2381), .B0_t (THETA_n119), .B0_f (new_AGEMA_signal_2370), .B1_t (new_AGEMA_signal_2371), .B1_f (new_AGEMA_signal_2372), .Z0_t (THETA_n121), .Z0_f (new_AGEMA_signal_2907), .Z1_t (new_AGEMA_signal_2908), .Z1_f (new_AGEMA_signal_2909) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U238 ( .A0_t (StateOut[132]), .A0_f (new_AGEMA_signal_2364), .A1_t (new_AGEMA_signal_2365), .A1_f (new_AGEMA_signal_2366), .B0_t (StateOut[140]), .B0_f (new_AGEMA_signal_2367), .B1_t (new_AGEMA_signal_2368), .B1_f (new_AGEMA_signal_2369), .Z0_t (THETA_n119), .Z0_f (new_AGEMA_signal_2370), .Z1_t (new_AGEMA_signal_2371), .Z1_f (new_AGEMA_signal_2372) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U237 ( .A0_t (StateOut[156]), .A0_f (new_AGEMA_signal_2373), .A1_t (new_AGEMA_signal_2374), .A1_f (new_AGEMA_signal_2375), .B0_t (StateOut[148]), .B0_f (new_AGEMA_signal_2376), .B1_t (new_AGEMA_signal_2377), .B1_f (new_AGEMA_signal_2378), .Z0_t (THETA_n120), .Z0_f (new_AGEMA_signal_2379), .Z1_t (new_AGEMA_signal_2380), .Z1_f (new_AGEMA_signal_2381) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U236 ( .A0_t (StateOut[152]), .A0_f (new_AGEMA_signal_2409), .A1_t (new_AGEMA_signal_2410), .A1_f (new_AGEMA_signal_2411), .B0_t (THETA_n118), .B0_f (new_AGEMA_signal_3312), .B1_t (new_AGEMA_signal_3313), .B1_f (new_AGEMA_signal_3314), .Z0_t (StateFromRhoPi[184]), .Z0_f (new_AGEMA_signal_3656), .Z1_t (new_AGEMA_signal_3657), .Z1_f (new_AGEMA_signal_3658) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U235 ( .A0_t (StateOut[144]), .A0_f (new_AGEMA_signal_3096), .A1_t (new_AGEMA_signal_3097), .A1_f (new_AGEMA_signal_3098), .B0_t (THETA_n118), .B0_f (new_AGEMA_signal_3312), .B1_t (new_AGEMA_signal_3313), .B1_f (new_AGEMA_signal_3314), .Z0_t (StateFromRhoPi[125]), .Z0_f (new_AGEMA_signal_3659), .Z1_t (new_AGEMA_signal_3660), .Z1_f (new_AGEMA_signal_3661) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U234 ( .A0_t (StateOut[136]), .A0_f (new_AGEMA_signal_2412), .A1_t (new_AGEMA_signal_2413), .A1_f (new_AGEMA_signal_2414), .B0_t (THETA_n118), .B0_f (new_AGEMA_signal_3312), .B1_t (new_AGEMA_signal_3313), .B1_f (new_AGEMA_signal_3314), .Z0_t (StateFromRhoPi[97]), .Z0_f (new_AGEMA_signal_3662), .Z1_t (new_AGEMA_signal_3663), .Z1_f (new_AGEMA_signal_3664) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U233 ( .A0_t (StateOut[128]), .A0_f (new_AGEMA_signal_2400), .A1_t (new_AGEMA_signal_2401), .A1_f (new_AGEMA_signal_2402), .B0_t (THETA_n118), .B0_f (new_AGEMA_signal_3312), .B1_t (new_AGEMA_signal_3313), .B1_f (new_AGEMA_signal_3314), .Z0_t (StateFromRhoPi[79]), .Z0_f (new_AGEMA_signal_3665), .Z1_t (new_AGEMA_signal_3666), .Z1_f (new_AGEMA_signal_3667) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U232 ( .A0_t (StateOut[120]), .A0_f (new_AGEMA_signal_2403), .A1_t (new_AGEMA_signal_2404), .A1_f (new_AGEMA_signal_2405), .B0_t (THETA_n118), .B0_f (new_AGEMA_signal_3312), .B1_t (new_AGEMA_signal_3313), .B1_f (new_AGEMA_signal_3314), .Z0_t (StateFromRhoPi[12]), .Z0_f (new_AGEMA_signal_3668), .Z1_t (new_AGEMA_signal_3669), .Z1_f (new_AGEMA_signal_3670) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U231 ( .A0_t (THETA_n117), .A0_f (new_AGEMA_signal_3111), .A1_t (new_AGEMA_signal_3112), .A1_f (new_AGEMA_signal_3113), .B0_t (THETA_n116), .B0_f (new_AGEMA_signal_3093), .B1_t (new_AGEMA_signal_3094), .B1_f (new_AGEMA_signal_3095), .Z0_t (THETA_n118), .Z0_f (new_AGEMA_signal_3312), .Z1_t (new_AGEMA_signal_3313), .Z1_f (new_AGEMA_signal_3314) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U230 ( .A0_t (StateOut[73]), .A0_f (new_AGEMA_signal_2430), .A1_t (new_AGEMA_signal_2431), .A1_f (new_AGEMA_signal_2432), .B0_t (THETA_n115), .B0_f (new_AGEMA_signal_3315), .B1_t (new_AGEMA_signal_3316), .B1_f (new_AGEMA_signal_3317), .Z0_t (StateFromRhoPi[195]), .Z0_f (new_AGEMA_signal_3671), .Z1_t (new_AGEMA_signal_3672), .Z1_f (new_AGEMA_signal_3673) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U229 ( .A0_t (StateOut[65]), .A0_f (new_AGEMA_signal_2427), .A1_t (new_AGEMA_signal_2428), .A1_f (new_AGEMA_signal_2429), .B0_t (THETA_n115), .B0_f (new_AGEMA_signal_3315), .B1_t (new_AGEMA_signal_3316), .B1_f (new_AGEMA_signal_3317), .Z0_t (StateFromRhoPi[134]), .Z0_f (new_AGEMA_signal_3674), .Z1_t (new_AGEMA_signal_3675), .Z1_f (new_AGEMA_signal_3676) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U228 ( .A0_t (StateOut[57]), .A0_f (new_AGEMA_signal_3102), .A1_t (new_AGEMA_signal_3103), .A1_f (new_AGEMA_signal_3104), .B0_t (THETA_n115), .B0_f (new_AGEMA_signal_3315), .B1_t (new_AGEMA_signal_3316), .B1_f (new_AGEMA_signal_3317), .Z0_t (StateFromRhoPi[107]), .Z0_f (new_AGEMA_signal_3677), .Z1_t (new_AGEMA_signal_3678), .Z1_f (new_AGEMA_signal_3679) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U227 ( .A0_t (StateOut[49]), .A0_f (new_AGEMA_signal_2418), .A1_t (new_AGEMA_signal_2419), .A1_f (new_AGEMA_signal_2420), .B0_t (THETA_n115), .B0_f (new_AGEMA_signal_3315), .B1_t (new_AGEMA_signal_3316), .B1_f (new_AGEMA_signal_3317), .Z0_t (StateFromRhoPi[45]), .Z0_f (new_AGEMA_signal_3680), .Z1_t (new_AGEMA_signal_3681), .Z1_f (new_AGEMA_signal_3682) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U226 ( .A0_t (StateOut[41]), .A0_f (new_AGEMA_signal_2421), .A1_t (new_AGEMA_signal_2422), .A1_f (new_AGEMA_signal_2423), .B0_t (THETA_n115), .B0_f (new_AGEMA_signal_3315), .B1_t (new_AGEMA_signal_3316), .B1_f (new_AGEMA_signal_3317), .Z0_t (StateFromRhoPi[18]), .Z0_f (new_AGEMA_signal_3683), .Z1_t (new_AGEMA_signal_3684), .Z1_f (new_AGEMA_signal_3685) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U225 ( .A0_t (THETA_n114), .A0_f (new_AGEMA_signal_3219), .A1_t (new_AGEMA_signal_3220), .A1_f (new_AGEMA_signal_3221), .B0_t (THETA_n116), .B0_f (new_AGEMA_signal_3093), .B1_t (new_AGEMA_signal_3094), .B1_f (new_AGEMA_signal_3095), .Z0_t (THETA_n115), .Z0_f (new_AGEMA_signal_3315), .Z1_t (new_AGEMA_signal_3316), .Z1_f (new_AGEMA_signal_3317) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U224 ( .A0_t (StateOut[96]), .A0_f (new_AGEMA_signal_3090), .A1_t (new_AGEMA_signal_3091), .A1_f (new_AGEMA_signal_3092), .B0_t (THETA_n113), .B0_f (new_AGEMA_signal_2910), .B1_t (new_AGEMA_signal_2911), .B1_f (new_AGEMA_signal_2912), .Z0_t (THETA_n116), .Z0_f (new_AGEMA_signal_3093), .Z1_t (new_AGEMA_signal_3094), .Z1_f (new_AGEMA_signal_3095) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U223 ( .A0_t (THETA_n112), .A0_f (new_AGEMA_signal_2397), .A1_t (new_AGEMA_signal_2398), .A1_f (new_AGEMA_signal_2399), .B0_t (THETA_n111), .B0_f (new_AGEMA_signal_2388), .B1_t (new_AGEMA_signal_2389), .B1_f (new_AGEMA_signal_2390), .Z0_t (THETA_n113), .Z0_f (new_AGEMA_signal_2910), .Z1_t (new_AGEMA_signal_2911), .Z1_f (new_AGEMA_signal_2912) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U222 ( .A0_t (StateOut[88]), .A0_f (new_AGEMA_signal_2382), .A1_t (new_AGEMA_signal_2383), .A1_f (new_AGEMA_signal_2384), .B0_t (StateOut[80]), .B0_f (new_AGEMA_signal_2385), .B1_t (new_AGEMA_signal_2386), .B1_f (new_AGEMA_signal_2387), .Z0_t (THETA_n111), .Z0_f (new_AGEMA_signal_2388), .Z1_t (new_AGEMA_signal_2389), .Z1_f (new_AGEMA_signal_2390) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U221 ( .A0_t (StateOut[104]), .A0_f (new_AGEMA_signal_2391), .A1_t (new_AGEMA_signal_2392), .A1_f (new_AGEMA_signal_2393), .B0_t (StateOut[112]), .B0_f (new_AGEMA_signal_2394), .B1_t (new_AGEMA_signal_2395), .B1_f (new_AGEMA_signal_2396), .Z0_t (THETA_n112), .Z0_f (new_AGEMA_signal_2397), .Z1_t (new_AGEMA_signal_2398), .Z1_f (new_AGEMA_signal_2399) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U220 ( .A0_t (StateOut[113]), .A0_f (new_AGEMA_signal_2301), .A1_t (new_AGEMA_signal_2302), .A1_f (new_AGEMA_signal_2303), .B0_t (THETA_n110), .B0_f (new_AGEMA_signal_3318), .B1_t (new_AGEMA_signal_3319), .B1_f (new_AGEMA_signal_3320), .Z0_t (StateFromRhoPi[174]), .Z0_f (new_AGEMA_signal_3686), .Z1_t (new_AGEMA_signal_3687), .Z1_f (new_AGEMA_signal_3688) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U219 ( .A0_t (StateOut[105]), .A0_f (new_AGEMA_signal_2304), .A1_t (new_AGEMA_signal_2305), .A1_f (new_AGEMA_signal_2306), .B0_t (THETA_n110), .B0_f (new_AGEMA_signal_3318), .B1_t (new_AGEMA_signal_3319), .B1_f (new_AGEMA_signal_3320), .Z0_t (StateFromRhoPi[144]), .Z0_f (new_AGEMA_signal_3689), .Z1_t (new_AGEMA_signal_3690), .Z1_f (new_AGEMA_signal_3691) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U218 ( .A0_t (StateOut[97]), .A0_f (new_AGEMA_signal_2295), .A1_t (new_AGEMA_signal_2296), .A1_f (new_AGEMA_signal_2297), .B0_t (THETA_n110), .B0_f (new_AGEMA_signal_3318), .B1_t (new_AGEMA_signal_3319), .B1_f (new_AGEMA_signal_3320), .Z0_t (StateFromRhoPi[84]), .Z0_f (new_AGEMA_signal_3692), .Z1_t (new_AGEMA_signal_3693), .Z1_f (new_AGEMA_signal_3694) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U217 ( .A0_t (StateOut[89]), .A0_f (new_AGEMA_signal_2292), .A1_t (new_AGEMA_signal_2293), .A1_f (new_AGEMA_signal_2294), .B0_t (THETA_n110), .B0_f (new_AGEMA_signal_3318), .B1_t (new_AGEMA_signal_3319), .B1_f (new_AGEMA_signal_3320), .Z0_t (StateFromRhoPi[63]), .Z0_f (new_AGEMA_signal_3695), .Z1_t (new_AGEMA_signal_3696), .Z1_f (new_AGEMA_signal_3697) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U216 ( .A0_t (StateOut[81]), .A0_f (new_AGEMA_signal_3060), .A1_t (new_AGEMA_signal_3061), .A1_f (new_AGEMA_signal_3062), .B0_t (THETA_n110), .B0_f (new_AGEMA_signal_3318), .B1_t (new_AGEMA_signal_3319), .B1_f (new_AGEMA_signal_3320), .Z0_t (StateFromRhoPi[39]), .Z0_f (new_AGEMA_signal_3698), .Z1_t (new_AGEMA_signal_3699), .Z1_f (new_AGEMA_signal_3700) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U215 ( .A0_t (THETA_n109), .A0_f (new_AGEMA_signal_3105), .A1_t (new_AGEMA_signal_3106), .A1_f (new_AGEMA_signal_3107), .B0_t (THETA_n130), .B0_f (new_AGEMA_signal_3099), .B1_t (new_AGEMA_signal_3100), .B1_f (new_AGEMA_signal_3101), .Z0_t (THETA_n110), .Z0_f (new_AGEMA_signal_3318), .Z1_t (new_AGEMA_signal_3319), .Z1_f (new_AGEMA_signal_3320) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U214 ( .A0_t (StateOut[144]), .A0_f (new_AGEMA_signal_3096), .A1_t (new_AGEMA_signal_3097), .A1_f (new_AGEMA_signal_3098), .B0_t (THETA_n108), .B0_f (new_AGEMA_signal_2913), .B1_t (new_AGEMA_signal_2914), .B1_f (new_AGEMA_signal_2915), .Z0_t (THETA_n130), .Z0_f (new_AGEMA_signal_3099), .Z1_t (new_AGEMA_signal_3100), .Z1_f (new_AGEMA_signal_3101) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U213 ( .A0_t (THETA_n107), .A0_f (new_AGEMA_signal_2415), .A1_t (new_AGEMA_signal_2416), .A1_f (new_AGEMA_signal_2417), .B0_t (THETA_n106), .B0_f (new_AGEMA_signal_2406), .B1_t (new_AGEMA_signal_2407), .B1_f (new_AGEMA_signal_2408), .Z0_t (THETA_n108), .Z0_f (new_AGEMA_signal_2913), .Z1_t (new_AGEMA_signal_2914), .Z1_f (new_AGEMA_signal_2915) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U212 ( .A0_t (StateOut[128]), .A0_f (new_AGEMA_signal_2400), .A1_t (new_AGEMA_signal_2401), .A1_f (new_AGEMA_signal_2402), .B0_t (StateOut[120]), .B0_f (new_AGEMA_signal_2403), .B1_t (new_AGEMA_signal_2404), .B1_f (new_AGEMA_signal_2405), .Z0_t (THETA_n106), .Z0_f (new_AGEMA_signal_2406), .Z1_t (new_AGEMA_signal_2407), .Z1_f (new_AGEMA_signal_2408) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U211 ( .A0_t (StateOut[152]), .A0_f (new_AGEMA_signal_2409), .A1_t (new_AGEMA_signal_2410), .A1_f (new_AGEMA_signal_2411), .B0_t (StateOut[136]), .B0_f (new_AGEMA_signal_2412), .B1_t (new_AGEMA_signal_2413), .B1_f (new_AGEMA_signal_2414), .Z0_t (THETA_n107), .Z0_f (new_AGEMA_signal_2415), .Z1_t (new_AGEMA_signal_2416), .Z1_f (new_AGEMA_signal_2417) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U210 ( .A0_t (StateOut[34]), .A0_f (new_AGEMA_signal_2535), .A1_t (new_AGEMA_signal_2536), .A1_f (new_AGEMA_signal_2537), .B0_t (THETA_n105), .B0_f (new_AGEMA_signal_3321), .B1_t (new_AGEMA_signal_3322), .B1_f (new_AGEMA_signal_3323), .Z0_t (StateFromRhoPi[180]), .Z0_f (new_AGEMA_signal_3701), .Z1_t (new_AGEMA_signal_3702), .Z1_f (new_AGEMA_signal_3703) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U209 ( .A0_t (StateOut[26]), .A0_f (new_AGEMA_signal_3138), .A1_t (new_AGEMA_signal_3139), .A1_f (new_AGEMA_signal_3140), .B0_t (THETA_n105), .B0_f (new_AGEMA_signal_3321), .B1_t (new_AGEMA_signal_3322), .B1_f (new_AGEMA_signal_3323), .Z0_t (StateFromRhoPi[155]), .Z0_f (new_AGEMA_signal_3704), .Z1_t (new_AGEMA_signal_3705), .Z1_f (new_AGEMA_signal_3706) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U208 ( .A0_t (StateOut[18]), .A0_f (new_AGEMA_signal_2538), .A1_t (new_AGEMA_signal_2539), .A1_f (new_AGEMA_signal_2540), .B0_t (THETA_n105), .B0_f (new_AGEMA_signal_3321), .B1_t (new_AGEMA_signal_3322), .B1_f (new_AGEMA_signal_3323), .Z0_t (StateFromRhoPi[93]), .Z0_f (new_AGEMA_signal_3707), .Z1_t (new_AGEMA_signal_3708), .Z1_f (new_AGEMA_signal_3709) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U207 ( .A0_t (StateOut[10]), .A0_f (new_AGEMA_signal_2526), .A1_t (new_AGEMA_signal_2527), .A1_f (new_AGEMA_signal_2528), .B0_t (THETA_n105), .B0_f (new_AGEMA_signal_3321), .B1_t (new_AGEMA_signal_3322), .B1_f (new_AGEMA_signal_3323), .Z0_t (StateFromRhoPi[70]), .Z0_f (new_AGEMA_signal_3710), .Z1_t (new_AGEMA_signal_3711), .Z1_f (new_AGEMA_signal_3712) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U206 ( .A0_t (OutData_s0_t[2]), .A0_f (OutData_s0_f[2]), .A1_t (OutData_s1_t[2]), .A1_f (OutData_s1_f[2]), .B0_t (THETA_n105), .B0_f (new_AGEMA_signal_3321), .B1_t (new_AGEMA_signal_3322), .B1_f (new_AGEMA_signal_3323), .Z0_t (StateFromRhoPi[2]), .Z0_f (new_AGEMA_signal_3713), .Z1_t (new_AGEMA_signal_3714), .Z1_f (new_AGEMA_signal_3715) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U205 ( .A0_t (THETA_n104), .A0_f (new_AGEMA_signal_3243), .A1_t (new_AGEMA_signal_3244), .A1_f (new_AGEMA_signal_3245), .B0_t (THETA_n109), .B0_f (new_AGEMA_signal_3105), .B1_t (new_AGEMA_signal_3106), .B1_f (new_AGEMA_signal_3107), .Z0_t (THETA_n105), .Z0_f (new_AGEMA_signal_3321), .Z1_t (new_AGEMA_signal_3322), .Z1_f (new_AGEMA_signal_3323) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U204 ( .A0_t (StateOut[57]), .A0_f (new_AGEMA_signal_3102), .A1_t (new_AGEMA_signal_3103), .A1_f (new_AGEMA_signal_3104), .B0_t (THETA_n103), .B0_f (new_AGEMA_signal_2916), .B1_t (new_AGEMA_signal_2917), .B1_f (new_AGEMA_signal_2918), .Z0_t (THETA_n109), .Z0_f (new_AGEMA_signal_3105), .Z1_t (new_AGEMA_signal_3106), .Z1_f (new_AGEMA_signal_3107) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U203 ( .A0_t (THETA_n102), .A0_f (new_AGEMA_signal_2433), .A1_t (new_AGEMA_signal_2434), .A1_f (new_AGEMA_signal_2435), .B0_t (THETA_n101), .B0_f (new_AGEMA_signal_2424), .B1_t (new_AGEMA_signal_2425), .B1_f (new_AGEMA_signal_2426), .Z0_t (THETA_n103), .Z0_f (new_AGEMA_signal_2916), .Z1_t (new_AGEMA_signal_2917), .Z1_f (new_AGEMA_signal_2918) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U202 ( .A0_t (StateOut[49]), .A0_f (new_AGEMA_signal_2418), .A1_t (new_AGEMA_signal_2419), .A1_f (new_AGEMA_signal_2420), .B0_t (StateOut[41]), .B0_f (new_AGEMA_signal_2421), .B1_t (new_AGEMA_signal_2422), .B1_f (new_AGEMA_signal_2423), .Z0_t (THETA_n101), .Z0_f (new_AGEMA_signal_2424), .Z1_t (new_AGEMA_signal_2425), .Z1_f (new_AGEMA_signal_2426) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U201 ( .A0_t (StateOut[65]), .A0_f (new_AGEMA_signal_2427), .A1_t (new_AGEMA_signal_2428), .A1_f (new_AGEMA_signal_2429), .B0_t (StateOut[73]), .B0_f (new_AGEMA_signal_2430), .B1_t (new_AGEMA_signal_2431), .B1_f (new_AGEMA_signal_2432), .Z0_t (THETA_n102), .Z0_f (new_AGEMA_signal_2433), .Z1_t (new_AGEMA_signal_2434), .Z1_f (new_AGEMA_signal_2435) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U200 ( .A0_t (StateOut[39]), .A0_f (new_AGEMA_signal_2355), .A1_t (new_AGEMA_signal_2356), .A1_f (new_AGEMA_signal_2357), .B0_t (THETA_n100), .B0_f (new_AGEMA_signal_3324), .B1_t (new_AGEMA_signal_3325), .B1_f (new_AGEMA_signal_3326), .Z0_t (StateFromRhoPi[177]), .Z0_f (new_AGEMA_signal_3716), .Z1_t (new_AGEMA_signal_3717), .Z1_f (new_AGEMA_signal_3718) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U199 ( .A0_t (StateOut[31]), .A0_f (new_AGEMA_signal_2358), .A1_t (new_AGEMA_signal_2359), .A1_f (new_AGEMA_signal_2360), .B0_t (THETA_n100), .B0_f (new_AGEMA_signal_3324), .B1_t (new_AGEMA_signal_3325), .B1_f (new_AGEMA_signal_3326), .Z0_t (StateFromRhoPi[152]), .Z0_f (new_AGEMA_signal_3719), .Z1_t (new_AGEMA_signal_3720), .Z1_f (new_AGEMA_signal_3721) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U198 ( .A0_t (StateOut[23]), .A0_f (new_AGEMA_signal_2349), .A1_t (new_AGEMA_signal_2350), .A1_f (new_AGEMA_signal_2351), .B0_t (THETA_n100), .B0_f (new_AGEMA_signal_3324), .B1_t (new_AGEMA_signal_3325), .B1_f (new_AGEMA_signal_3326), .Z0_t (StateFromRhoPi[90]), .Z0_f (new_AGEMA_signal_3722), .Z1_t (new_AGEMA_signal_3723), .Z1_f (new_AGEMA_signal_3724) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U197 ( .A0_t (StateOut[15]), .A0_f (new_AGEMA_signal_2346), .A1_t (new_AGEMA_signal_2347), .A1_f (new_AGEMA_signal_2348), .B0_t (THETA_n100), .B0_f (new_AGEMA_signal_3324), .B1_t (new_AGEMA_signal_3325), .B1_f (new_AGEMA_signal_3326), .Z0_t (StateFromRhoPi[67]), .Z0_f (new_AGEMA_signal_3725), .Z1_t (new_AGEMA_signal_3726), .Z1_f (new_AGEMA_signal_3727) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U196 ( .A0_t (OutData_s0_t[7]), .A0_f (OutData_s0_f[7]), .A1_t (OutData_s1_t[7]), .A1_f (OutData_s1_f[7]), .B0_t (THETA_n100), .B0_f (new_AGEMA_signal_3324), .B1_t (new_AGEMA_signal_3325), .B1_f (new_AGEMA_signal_3326), .Z0_t (StateFromRhoPi[7]), .Z0_f (new_AGEMA_signal_3728), .Z1_t (new_AGEMA_signal_3729), .Z1_f (new_AGEMA_signal_3730) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U195 ( .A0_t (THETA_n99), .A0_f (new_AGEMA_signal_3117), .A1_t (new_AGEMA_signal_3118), .A1_f (new_AGEMA_signal_3119), .B0_t (THETA_n117), .B0_f (new_AGEMA_signal_3111), .B1_t (new_AGEMA_signal_3112), .B1_f (new_AGEMA_signal_3113), .Z0_t (THETA_n100), .Z0_f (new_AGEMA_signal_3324), .Z1_t (new_AGEMA_signal_3325), .Z1_f (new_AGEMA_signal_3326) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U194 ( .A0_t (StateOut[183]), .A0_f (new_AGEMA_signal_3108), .A1_t (new_AGEMA_signal_3109), .A1_f (new_AGEMA_signal_3110), .B0_t (THETA_n98), .B0_f (new_AGEMA_signal_2919), .B1_t (new_AGEMA_signal_2920), .B1_f (new_AGEMA_signal_2921), .Z0_t (THETA_n117), .Z0_f (new_AGEMA_signal_3111), .Z1_t (new_AGEMA_signal_3112), .Z1_f (new_AGEMA_signal_3113) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U193 ( .A0_t (THETA_n97), .A0_f (new_AGEMA_signal_2451), .A1_t (new_AGEMA_signal_2452), .A1_f (new_AGEMA_signal_2453), .B0_t (THETA_n96), .B0_f (new_AGEMA_signal_2442), .B1_t (new_AGEMA_signal_2443), .B1_f (new_AGEMA_signal_2444), .Z0_t (THETA_n98), .Z0_f (new_AGEMA_signal_2919), .Z1_t (new_AGEMA_signal_2920), .Z1_f (new_AGEMA_signal_2921) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U192 ( .A0_t (StateOut[175]), .A0_f (new_AGEMA_signal_2436), .A1_t (new_AGEMA_signal_2437), .A1_f (new_AGEMA_signal_2438), .B0_t (StateOut[167]), .B0_f (new_AGEMA_signal_2439), .B1_t (new_AGEMA_signal_2440), .B1_f (new_AGEMA_signal_2441), .Z0_t (THETA_n96), .Z0_f (new_AGEMA_signal_2442), .Z1_t (new_AGEMA_signal_2443), .Z1_f (new_AGEMA_signal_2444) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U191 ( .A0_t (StateOut[191]), .A0_f (new_AGEMA_signal_2445), .A1_t (new_AGEMA_signal_2446), .A1_f (new_AGEMA_signal_2447), .B0_t (StateOut[199]), .B0_f (new_AGEMA_signal_2448), .B1_t (new_AGEMA_signal_2449), .B1_f (new_AGEMA_signal_2450), .Z0_t (THETA_n97), .Z0_f (new_AGEMA_signal_2451), .Z1_t (new_AGEMA_signal_2452), .Z1_f (new_AGEMA_signal_2453) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U190 ( .A0_t (StateOut[118]), .A0_f (new_AGEMA_signal_2697), .A1_t (new_AGEMA_signal_2698), .A1_f (new_AGEMA_signal_2699), .B0_t (THETA_n95), .B0_f (new_AGEMA_signal_3327), .B1_t (new_AGEMA_signal_3328), .B1_f (new_AGEMA_signal_3329), .Z0_t (StateFromRhoPi[171]), .Z0_f (new_AGEMA_signal_3731), .Z1_t (new_AGEMA_signal_3732), .Z1_f (new_AGEMA_signal_3733) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U189 ( .A0_t (StateOut[110]), .A0_f (new_AGEMA_signal_3192), .A1_t (new_AGEMA_signal_3193), .A1_f (new_AGEMA_signal_3194), .B0_t (THETA_n95), .B0_f (new_AGEMA_signal_3327), .B1_t (new_AGEMA_signal_3328), .B1_f (new_AGEMA_signal_3329), .Z0_t (StateFromRhoPi[149]), .Z0_f (new_AGEMA_signal_3734), .Z1_t (new_AGEMA_signal_3735), .Z1_f (new_AGEMA_signal_3736) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U188 ( .A0_t (StateOut[102]), .A0_f (new_AGEMA_signal_2700), .A1_t (new_AGEMA_signal_2701), .A1_f (new_AGEMA_signal_2702), .B0_t (THETA_n95), .B0_f (new_AGEMA_signal_3327), .B1_t (new_AGEMA_signal_3328), .B1_f (new_AGEMA_signal_3329), .Z0_t (StateFromRhoPi[81]), .Z0_f (new_AGEMA_signal_3737), .Z1_t (new_AGEMA_signal_3738), .Z1_f (new_AGEMA_signal_3739) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U187 ( .A0_t (StateOut[94]), .A0_f (new_AGEMA_signal_2688), .A1_t (new_AGEMA_signal_2689), .A1_f (new_AGEMA_signal_2690), .B0_t (THETA_n95), .B0_f (new_AGEMA_signal_3327), .B1_t (new_AGEMA_signal_3328), .B1_f (new_AGEMA_signal_3329), .Z0_t (StateFromRhoPi[60]), .Z0_f (new_AGEMA_signal_3740), .Z1_t (new_AGEMA_signal_3741), .Z1_f (new_AGEMA_signal_3742) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U186 ( .A0_t (StateOut[86]), .A0_f (new_AGEMA_signal_2691), .A1_t (new_AGEMA_signal_2692), .A1_f (new_AGEMA_signal_2693), .B0_t (THETA_n95), .B0_f (new_AGEMA_signal_3327), .B1_t (new_AGEMA_signal_3328), .B1_f (new_AGEMA_signal_3329), .Z0_t (StateFromRhoPi[36]), .Z0_f (new_AGEMA_signal_3743), .Z1_t (new_AGEMA_signal_3744), .Z1_f (new_AGEMA_signal_3745) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U185 ( .A0_t (THETA_n94), .A0_f (new_AGEMA_signal_3147), .A1_t (new_AGEMA_signal_3148), .A1_f (new_AGEMA_signal_3149), .B0_t (THETA_n99), .B0_f (new_AGEMA_signal_3117), .B1_t (new_AGEMA_signal_3118), .B1_f (new_AGEMA_signal_3119), .Z0_t (THETA_n95), .Z0_f (new_AGEMA_signal_3327), .Z1_t (new_AGEMA_signal_3328), .Z1_f (new_AGEMA_signal_3329) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U184 ( .A0_t (StateOut[62]), .A0_f (new_AGEMA_signal_3114), .A1_t (new_AGEMA_signal_3115), .A1_f (new_AGEMA_signal_3116), .B0_t (THETA_n93), .B0_f (new_AGEMA_signal_2922), .B1_t (new_AGEMA_signal_2923), .B1_f (new_AGEMA_signal_2924), .Z0_t (THETA_n99), .Z0_f (new_AGEMA_signal_3117), .Z1_t (new_AGEMA_signal_3118), .Z1_f (new_AGEMA_signal_3119) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U183 ( .A0_t (THETA_n92), .A0_f (new_AGEMA_signal_2469), .A1_t (new_AGEMA_signal_2470), .A1_f (new_AGEMA_signal_2471), .B0_t (THETA_n91), .B0_f (new_AGEMA_signal_2460), .B1_t (new_AGEMA_signal_2461), .B1_f (new_AGEMA_signal_2462), .Z0_t (THETA_n93), .Z0_f (new_AGEMA_signal_2922), .Z1_t (new_AGEMA_signal_2923), .Z1_f (new_AGEMA_signal_2924) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U182 ( .A0_t (StateOut[54]), .A0_f (new_AGEMA_signal_2454), .A1_t (new_AGEMA_signal_2455), .A1_f (new_AGEMA_signal_2456), .B0_t (StateOut[46]), .B0_f (new_AGEMA_signal_2457), .B1_t (new_AGEMA_signal_2458), .B1_f (new_AGEMA_signal_2459), .Z0_t (THETA_n91), .Z0_f (new_AGEMA_signal_2460), .Z1_t (new_AGEMA_signal_2461), .Z1_f (new_AGEMA_signal_2462) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U181 ( .A0_t (StateOut[70]), .A0_f (new_AGEMA_signal_2463), .A1_t (new_AGEMA_signal_2464), .A1_f (new_AGEMA_signal_2465), .B0_t (StateOut[78]), .B0_f (new_AGEMA_signal_2466), .B1_t (new_AGEMA_signal_2467), .B1_f (new_AGEMA_signal_2468), .Z0_t (THETA_n92), .Z0_f (new_AGEMA_signal_2469), .Z1_t (new_AGEMA_signal_2470), .Z1_f (new_AGEMA_signal_2471) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U180 ( .A0_t (StateOut[159]), .A0_f (new_AGEMA_signal_2157), .A1_t (new_AGEMA_signal_2158), .A1_f (new_AGEMA_signal_2159), .B0_t (THETA_n90), .B0_f (new_AGEMA_signal_3330), .B1_t (new_AGEMA_signal_3331), .B1_f (new_AGEMA_signal_3332), .Z0_t (StateFromRhoPi[191]), .Z0_f (new_AGEMA_signal_3746), .Z1_t (new_AGEMA_signal_3747), .Z1_f (new_AGEMA_signal_3748) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U179 ( .A0_t (StateOut[151]), .A0_f (new_AGEMA_signal_2160), .A1_t (new_AGEMA_signal_2161), .A1_f (new_AGEMA_signal_2162), .B0_t (THETA_n90), .B0_f (new_AGEMA_signal_3330), .B1_t (new_AGEMA_signal_3331), .B1_f (new_AGEMA_signal_3332), .Z0_t (StateFromRhoPi[124]), .Z0_f (new_AGEMA_signal_3749), .Z1_t (new_AGEMA_signal_3750), .Z1_f (new_AGEMA_signal_3751) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U178 ( .A0_t (StateOut[143]), .A0_f (new_AGEMA_signal_2151), .A1_t (new_AGEMA_signal_2152), .A1_f (new_AGEMA_signal_2153), .B0_t (THETA_n90), .B0_f (new_AGEMA_signal_3330), .B1_t (new_AGEMA_signal_3331), .B1_f (new_AGEMA_signal_3332), .Z0_t (StateFromRhoPi[96]), .Z0_f (new_AGEMA_signal_3752), .Z1_t (new_AGEMA_signal_3753), .Z1_f (new_AGEMA_signal_3754) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U177 ( .A0_t (StateOut[135]), .A0_f (new_AGEMA_signal_2148), .A1_t (new_AGEMA_signal_2149), .A1_f (new_AGEMA_signal_2150), .B0_t (THETA_n90), .B0_f (new_AGEMA_signal_3330), .B1_t (new_AGEMA_signal_3331), .B1_f (new_AGEMA_signal_3332), .Z0_t (StateFromRhoPi[78]), .Z0_f (new_AGEMA_signal_3755), .Z1_t (new_AGEMA_signal_3756), .Z1_f (new_AGEMA_signal_3757) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U176 ( .A0_t (StateOut[127]), .A0_f (new_AGEMA_signal_3012), .A1_t (new_AGEMA_signal_3013), .A1_f (new_AGEMA_signal_3014), .B0_t (THETA_n90), .B0_f (new_AGEMA_signal_3330), .B1_t (new_AGEMA_signal_3331), .B1_f (new_AGEMA_signal_3332), .Z0_t (StateFromRhoPi[11]), .Z0_f (new_AGEMA_signal_3758), .Z1_t (new_AGEMA_signal_3759), .Z1_f (new_AGEMA_signal_3760) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U175 ( .A0_t (THETA_n89), .A0_f (new_AGEMA_signal_3129), .A1_t (new_AGEMA_signal_3130), .A1_f (new_AGEMA_signal_3131), .B0_t (THETA_n167), .B0_f (new_AGEMA_signal_3123), .B1_t (new_AGEMA_signal_3124), .B1_f (new_AGEMA_signal_3125), .Z0_t (THETA_n90), .Z0_f (new_AGEMA_signal_3330), .Z1_t (new_AGEMA_signal_3331), .Z1_f (new_AGEMA_signal_3332) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U174 ( .A0_t (StateOut[103]), .A0_f (new_AGEMA_signal_3120), .A1_t (new_AGEMA_signal_3121), .A1_f (new_AGEMA_signal_3122), .B0_t (THETA_n88), .B0_f (new_AGEMA_signal_2925), .B1_t (new_AGEMA_signal_2926), .B1_f (new_AGEMA_signal_2927), .Z0_t (THETA_n167), .Z0_f (new_AGEMA_signal_3123), .Z1_t (new_AGEMA_signal_3124), .Z1_f (new_AGEMA_signal_3125) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U173 ( .A0_t (THETA_n87), .A0_f (new_AGEMA_signal_2487), .A1_t (new_AGEMA_signal_2488), .A1_f (new_AGEMA_signal_2489), .B0_t (THETA_n86), .B0_f (new_AGEMA_signal_2478), .B1_t (new_AGEMA_signal_2479), .B1_f (new_AGEMA_signal_2480), .Z0_t (THETA_n88), .Z0_f (new_AGEMA_signal_2925), .Z1_t (new_AGEMA_signal_2926), .Z1_f (new_AGEMA_signal_2927) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U172 ( .A0_t (StateOut[95]), .A0_f (new_AGEMA_signal_2472), .A1_t (new_AGEMA_signal_2473), .A1_f (new_AGEMA_signal_2474), .B0_t (StateOut[87]), .B0_f (new_AGEMA_signal_2475), .B1_t (new_AGEMA_signal_2476), .B1_f (new_AGEMA_signal_2477), .Z0_t (THETA_n86), .Z0_f (new_AGEMA_signal_2478), .Z1_t (new_AGEMA_signal_2479), .Z1_f (new_AGEMA_signal_2480) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U171 ( .A0_t (StateOut[111]), .A0_f (new_AGEMA_signal_2481), .A1_t (new_AGEMA_signal_2482), .A1_f (new_AGEMA_signal_2483), .B0_t (StateOut[119]), .B0_f (new_AGEMA_signal_2484), .B1_t (new_AGEMA_signal_2485), .B1_f (new_AGEMA_signal_2486), .Z0_t (THETA_n87), .Z0_f (new_AGEMA_signal_2487), .Z1_t (new_AGEMA_signal_2488), .Z1_f (new_AGEMA_signal_2489) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U170 ( .A0_t (StateOut[38]), .A0_f (new_AGEMA_signal_2139), .A1_t (new_AGEMA_signal_2140), .A1_f (new_AGEMA_signal_2141), .B0_t (THETA_n85), .B0_f (new_AGEMA_signal_3333), .B1_t (new_AGEMA_signal_3334), .B1_f (new_AGEMA_signal_3335), .Z0_t (StateFromRhoPi[176]), .Z0_f (new_AGEMA_signal_3761), .Z1_t (new_AGEMA_signal_3762), .Z1_f (new_AGEMA_signal_3763) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U169 ( .A0_t (StateOut[30]), .A0_f (new_AGEMA_signal_2142), .A1_t (new_AGEMA_signal_2143), .A1_f (new_AGEMA_signal_2144), .B0_t (THETA_n85), .B0_f (new_AGEMA_signal_3333), .B1_t (new_AGEMA_signal_3334), .B1_f (new_AGEMA_signal_3335), .Z0_t (StateFromRhoPi[159]), .Z0_f (new_AGEMA_signal_3764), .Z1_t (new_AGEMA_signal_3765), .Z1_f (new_AGEMA_signal_3766) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U168 ( .A0_t (StateOut[22]), .A0_f (new_AGEMA_signal_2133), .A1_t (new_AGEMA_signal_2134), .A1_f (new_AGEMA_signal_2135), .B0_t (THETA_n85), .B0_f (new_AGEMA_signal_3333), .B1_t (new_AGEMA_signal_3334), .B1_f (new_AGEMA_signal_3335), .Z0_t (StateFromRhoPi[89]), .Z0_f (new_AGEMA_signal_3767), .Z1_t (new_AGEMA_signal_3768), .Z1_f (new_AGEMA_signal_3769) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U167 ( .A0_t (StateOut[14]), .A0_f (new_AGEMA_signal_2130), .A1_t (new_AGEMA_signal_2131), .A1_f (new_AGEMA_signal_2132), .B0_t (THETA_n85), .B0_f (new_AGEMA_signal_3333), .B1_t (new_AGEMA_signal_3334), .B1_f (new_AGEMA_signal_3335), .Z0_t (StateFromRhoPi[66]), .Z0_f (new_AGEMA_signal_3770), .Z1_t (new_AGEMA_signal_3771), .Z1_f (new_AGEMA_signal_3772) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U166 ( .A0_t (OutData_s0_t[6]), .A0_f (OutData_s0_f[6]), .A1_t (OutData_s1_t[6]), .A1_f (OutData_s1_f[6]), .B0_t (THETA_n85), .B0_f (new_AGEMA_signal_3333), .B1_t (new_AGEMA_signal_3334), .B1_f (new_AGEMA_signal_3335), .Z0_t (StateFromRhoPi[6]), .Z0_f (new_AGEMA_signal_3773), .Z1_t (new_AGEMA_signal_3774), .Z1_f (new_AGEMA_signal_3775) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U165 ( .A0_t (THETA_n122), .A0_f (new_AGEMA_signal_3135), .A1_t (new_AGEMA_signal_3136), .A1_f (new_AGEMA_signal_3137), .B0_t (THETA_n89), .B0_f (new_AGEMA_signal_3129), .B1_t (new_AGEMA_signal_3130), .B1_f (new_AGEMA_signal_3131), .Z0_t (THETA_n85), .Z0_f (new_AGEMA_signal_3333), .Z1_t (new_AGEMA_signal_3334), .Z1_f (new_AGEMA_signal_3335) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U164 ( .A0_t (StateOut[182]), .A0_f (new_AGEMA_signal_3126), .A1_t (new_AGEMA_signal_3127), .A1_f (new_AGEMA_signal_3128), .B0_t (THETA_n84), .B0_f (new_AGEMA_signal_2928), .B1_t (new_AGEMA_signal_2929), .B1_f (new_AGEMA_signal_2930), .Z0_t (THETA_n89), .Z0_f (new_AGEMA_signal_3129), .Z1_t (new_AGEMA_signal_3130), .Z1_f (new_AGEMA_signal_3131) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U163 ( .A0_t (THETA_n83), .A0_f (new_AGEMA_signal_2505), .A1_t (new_AGEMA_signal_2506), .A1_f (new_AGEMA_signal_2507), .B0_t (THETA_n82), .B0_f (new_AGEMA_signal_2496), .B1_t (new_AGEMA_signal_2497), .B1_f (new_AGEMA_signal_2498), .Z0_t (THETA_n84), .Z0_f (new_AGEMA_signal_2928), .Z1_t (new_AGEMA_signal_2929), .Z1_f (new_AGEMA_signal_2930) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U162 ( .A0_t (StateOut[174]), .A0_f (new_AGEMA_signal_2490), .A1_t (new_AGEMA_signal_2491), .A1_f (new_AGEMA_signal_2492), .B0_t (StateOut[166]), .B0_f (new_AGEMA_signal_2493), .B1_t (new_AGEMA_signal_2494), .B1_f (new_AGEMA_signal_2495), .Z0_t (THETA_n82), .Z0_f (new_AGEMA_signal_2496), .Z1_t (new_AGEMA_signal_2497), .Z1_f (new_AGEMA_signal_2498) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U161 ( .A0_t (StateOut[190]), .A0_f (new_AGEMA_signal_2499), .A1_t (new_AGEMA_signal_2500), .A1_f (new_AGEMA_signal_2501), .B0_t (StateOut[198]), .B0_f (new_AGEMA_signal_2502), .B1_t (new_AGEMA_signal_2503), .B1_f (new_AGEMA_signal_2504), .Z0_t (THETA_n83), .Z0_f (new_AGEMA_signal_2505), .Z1_t (new_AGEMA_signal_2506), .Z1_f (new_AGEMA_signal_2507) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U160 ( .A0_t (StateOut[45]), .A0_f (new_AGEMA_signal_3132), .A1_t (new_AGEMA_signal_3133), .A1_f (new_AGEMA_signal_3134), .B0_t (THETA_n81), .B0_f (new_AGEMA_signal_2931), .B1_t (new_AGEMA_signal_2932), .B1_f (new_AGEMA_signal_2933), .Z0_t (THETA_n122), .Z0_f (new_AGEMA_signal_3135), .Z1_t (new_AGEMA_signal_3136), .Z1_f (new_AGEMA_signal_3137) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U159 ( .A0_t (THETA_n80), .A0_f (new_AGEMA_signal_2523), .A1_t (new_AGEMA_signal_2524), .A1_f (new_AGEMA_signal_2525), .B0_t (THETA_n79), .B0_f (new_AGEMA_signal_2514), .B1_t (new_AGEMA_signal_2515), .B1_f (new_AGEMA_signal_2516), .Z0_t (THETA_n81), .Z0_f (new_AGEMA_signal_2931), .Z1_t (new_AGEMA_signal_2932), .Z1_f (new_AGEMA_signal_2933) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U158 ( .A0_t (StateOut[53]), .A0_f (new_AGEMA_signal_2508), .A1_t (new_AGEMA_signal_2509), .A1_f (new_AGEMA_signal_2510), .B0_t (StateOut[61]), .B0_f (new_AGEMA_signal_2511), .B1_t (new_AGEMA_signal_2512), .B1_f (new_AGEMA_signal_2513), .Z0_t (THETA_n79), .Z0_f (new_AGEMA_signal_2514), .Z1_t (new_AGEMA_signal_2515), .Z1_f (new_AGEMA_signal_2516) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U157 ( .A0_t (StateOut[77]), .A0_f (new_AGEMA_signal_2517), .A1_t (new_AGEMA_signal_2518), .A1_f (new_AGEMA_signal_2519), .B0_t (StateOut[69]), .B0_f (new_AGEMA_signal_2520), .B1_t (new_AGEMA_signal_2521), .B1_f (new_AGEMA_signal_2522), .Z0_t (THETA_n80), .Z0_f (new_AGEMA_signal_2523), .Z1_t (new_AGEMA_signal_2524), .Z1_f (new_AGEMA_signal_2525) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U156 ( .A0_t (StateOut[195]), .A0_f (new_AGEMA_signal_2790), .A1_t (new_AGEMA_signal_2791), .A1_f (new_AGEMA_signal_2792), .B0_t (THETA_n78), .B0_f (new_AGEMA_signal_3336), .B1_t (new_AGEMA_signal_3337), .B1_f (new_AGEMA_signal_3338), .Z0_t (StateFromRhoPi[161]), .Z0_f (new_AGEMA_signal_3776), .Z1_t (new_AGEMA_signal_3777), .Z1_f (new_AGEMA_signal_3778) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U155 ( .A0_t (StateOut[187]), .A0_f (new_AGEMA_signal_2787), .A1_t (new_AGEMA_signal_2788), .A1_f (new_AGEMA_signal_2789), .B0_t (THETA_n78), .B0_f (new_AGEMA_signal_3336), .B1_t (new_AGEMA_signal_3337), .B1_f (new_AGEMA_signal_3338), .Z0_t (StateFromRhoPi[139]), .Z0_f (new_AGEMA_signal_3779), .Z1_t (new_AGEMA_signal_3780), .Z1_f (new_AGEMA_signal_3781) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U154 ( .A0_t (StateOut[179]), .A0_f (new_AGEMA_signal_3222), .A1_t (new_AGEMA_signal_3223), .A1_f (new_AGEMA_signal_3224), .B0_t (THETA_n78), .B0_f (new_AGEMA_signal_3336), .B1_t (new_AGEMA_signal_3337), .B1_f (new_AGEMA_signal_3338), .Z0_t (StateFromRhoPi[114]), .Z0_f (new_AGEMA_signal_3782), .Z1_t (new_AGEMA_signal_3783), .Z1_f (new_AGEMA_signal_3784) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U153 ( .A0_t (StateOut[171]), .A0_f (new_AGEMA_signal_2778), .A1_t (new_AGEMA_signal_2779), .A1_f (new_AGEMA_signal_2780), .B0_t (THETA_n78), .B0_f (new_AGEMA_signal_3336), .B1_t (new_AGEMA_signal_3337), .B1_f (new_AGEMA_signal_3338), .Z0_t (StateFromRhoPi[55]), .Z0_f (new_AGEMA_signal_3785), .Z1_t (new_AGEMA_signal_3786), .Z1_f (new_AGEMA_signal_3787) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U152 ( .A0_t (StateOut[163]), .A0_f (new_AGEMA_signal_2781), .A1_t (new_AGEMA_signal_2782), .A1_f (new_AGEMA_signal_2783), .B0_t (THETA_n78), .B0_f (new_AGEMA_signal_3336), .B1_t (new_AGEMA_signal_3337), .B1_f (new_AGEMA_signal_3338), .Z0_t (StateFromRhoPi[30]), .Z0_f (new_AGEMA_signal_3788), .Z1_t (new_AGEMA_signal_3789), .Z1_f (new_AGEMA_signal_3790) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U151 ( .A0_t (THETA_n77), .A0_f (new_AGEMA_signal_3159), .A1_t (new_AGEMA_signal_3160), .A1_f (new_AGEMA_signal_3161), .B0_t (THETA_n142), .B0_f (new_AGEMA_signal_3141), .B1_t (new_AGEMA_signal_3142), .B1_f (new_AGEMA_signal_3143), .Z0_t (THETA_n78), .Z0_f (new_AGEMA_signal_3336), .Z1_t (new_AGEMA_signal_3337), .Z1_f (new_AGEMA_signal_3338) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U150 ( .A0_t (StateOut[26]), .A0_f (new_AGEMA_signal_3138), .A1_t (new_AGEMA_signal_3139), .A1_f (new_AGEMA_signal_3140), .B0_t (THETA_n76), .B0_f (new_AGEMA_signal_2934), .B1_t (new_AGEMA_signal_2935), .B1_f (new_AGEMA_signal_2936), .Z0_t (THETA_n142), .Z0_f (new_AGEMA_signal_3141), .Z1_t (new_AGEMA_signal_3142), .Z1_f (new_AGEMA_signal_3143) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U149 ( .A0_t (THETA_n75), .A0_f (new_AGEMA_signal_2541), .A1_t (new_AGEMA_signal_2542), .A1_f (new_AGEMA_signal_2543), .B0_t (THETA_n74), .B0_f (new_AGEMA_signal_2532), .B1_t (new_AGEMA_signal_2533), .B1_f (new_AGEMA_signal_2534), .Z0_t (THETA_n76), .Z0_f (new_AGEMA_signal_2934), .Z1_t (new_AGEMA_signal_2935), .Z1_f (new_AGEMA_signal_2936) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U148 ( .A0_t (StateOut[10]), .A0_f (new_AGEMA_signal_2526), .A1_t (new_AGEMA_signal_2527), .A1_f (new_AGEMA_signal_2528), .B0_t (OutData_s0_t[2]), .B0_f (OutData_s0_f[2]), .B1_t (OutData_s1_t[2]), .B1_f (OutData_s1_f[2]), .Z0_t (THETA_n74), .Z0_f (new_AGEMA_signal_2532), .Z1_t (new_AGEMA_signal_2533), .Z1_f (new_AGEMA_signal_2534) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U147 ( .A0_t (StateOut[34]), .A0_f (new_AGEMA_signal_2535), .A1_t (new_AGEMA_signal_2536), .A1_f (new_AGEMA_signal_2537), .B0_t (StateOut[18]), .B0_f (new_AGEMA_signal_2538), .B1_t (new_AGEMA_signal_2539), .B1_f (new_AGEMA_signal_2540), .Z0_t (THETA_n75), .Z0_f (new_AGEMA_signal_2541), .Z1_t (new_AGEMA_signal_2542), .Z1_f (new_AGEMA_signal_2543) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U146 ( .A0_t (StateOut[197]), .A0_f (new_AGEMA_signal_2682), .A1_t (new_AGEMA_signal_2683), .A1_f (new_AGEMA_signal_2684), .B0_t (THETA_n73), .B0_f (new_AGEMA_signal_3339), .B1_t (new_AGEMA_signal_3340), .B1_f (new_AGEMA_signal_3341), .Z0_t (StateFromRhoPi[163]), .Z0_f (new_AGEMA_signal_3791), .Z1_t (new_AGEMA_signal_3792), .Z1_f (new_AGEMA_signal_3793) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U145 ( .A0_t (StateOut[189]), .A0_f (new_AGEMA_signal_2679), .A1_t (new_AGEMA_signal_2680), .A1_f (new_AGEMA_signal_2681), .B0_t (THETA_n73), .B0_f (new_AGEMA_signal_3339), .B1_t (new_AGEMA_signal_3340), .B1_f (new_AGEMA_signal_3341), .Z0_t (StateFromRhoPi[141]), .Z0_f (new_AGEMA_signal_3794), .Z1_t (new_AGEMA_signal_3795), .Z1_f (new_AGEMA_signal_3796) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U144 ( .A0_t (StateOut[181]), .A0_f (new_AGEMA_signal_3186), .A1_t (new_AGEMA_signal_3187), .A1_f (new_AGEMA_signal_3188), .B0_t (THETA_n73), .B0_f (new_AGEMA_signal_3339), .B1_t (new_AGEMA_signal_3340), .B1_f (new_AGEMA_signal_3341), .Z0_t (StateFromRhoPi[116]), .Z0_f (new_AGEMA_signal_3797), .Z1_t (new_AGEMA_signal_3798), .Z1_f (new_AGEMA_signal_3799) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U143 ( .A0_t (StateOut[173]), .A0_f (new_AGEMA_signal_2670), .A1_t (new_AGEMA_signal_2671), .A1_f (new_AGEMA_signal_2672), .B0_t (THETA_n73), .B0_f (new_AGEMA_signal_3339), .B1_t (new_AGEMA_signal_3340), .B1_f (new_AGEMA_signal_3341), .Z0_t (StateFromRhoPi[49]), .Z0_f (new_AGEMA_signal_3800), .Z1_t (new_AGEMA_signal_3801), .Z1_f (new_AGEMA_signal_3802) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U142 ( .A0_t (StateOut[165]), .A0_f (new_AGEMA_signal_2673), .A1_t (new_AGEMA_signal_2674), .A1_f (new_AGEMA_signal_2675), .B0_t (THETA_n73), .B0_f (new_AGEMA_signal_3339), .B1_t (new_AGEMA_signal_3340), .B1_f (new_AGEMA_signal_3341), .Z0_t (StateFromRhoPi[24]), .Z0_f (new_AGEMA_signal_3803), .Z1_t (new_AGEMA_signal_3804), .Z1_f (new_AGEMA_signal_3805) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U141 ( .A0_t (THETA_n72), .A0_f (new_AGEMA_signal_3153), .A1_t (new_AGEMA_signal_3154), .A1_f (new_AGEMA_signal_3155), .B0_t (THETA_n94), .B0_f (new_AGEMA_signal_3147), .B1_t (new_AGEMA_signal_3148), .B1_f (new_AGEMA_signal_3149), .Z0_t (THETA_n73), .Z0_f (new_AGEMA_signal_3339), .Z1_t (new_AGEMA_signal_3340), .Z1_f (new_AGEMA_signal_3341) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U140 ( .A0_t (StateOut[125]), .A0_f (new_AGEMA_signal_3144), .A1_t (new_AGEMA_signal_3145), .A1_f (new_AGEMA_signal_3146), .B0_t (THETA_n71), .B0_f (new_AGEMA_signal_2937), .B1_t (new_AGEMA_signal_2938), .B1_f (new_AGEMA_signal_2939), .Z0_t (THETA_n94), .Z0_f (new_AGEMA_signal_3147), .Z1_t (new_AGEMA_signal_3148), .Z1_f (new_AGEMA_signal_3149) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U139 ( .A0_t (THETA_n70), .A0_f (new_AGEMA_signal_2559), .A1_t (new_AGEMA_signal_2560), .A1_f (new_AGEMA_signal_2561), .B0_t (THETA_n69), .B0_f (new_AGEMA_signal_2550), .B1_t (new_AGEMA_signal_2551), .B1_f (new_AGEMA_signal_2552), .Z0_t (THETA_n71), .Z0_f (new_AGEMA_signal_2937), .Z1_t (new_AGEMA_signal_2938), .Z1_f (new_AGEMA_signal_2939) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U138 ( .A0_t (StateOut[133]), .A0_f (new_AGEMA_signal_2544), .A1_t (new_AGEMA_signal_2545), .A1_f (new_AGEMA_signal_2546), .B0_t (StateOut[141]), .B0_f (new_AGEMA_signal_2547), .B1_t (new_AGEMA_signal_2548), .B1_f (new_AGEMA_signal_2549), .Z0_t (THETA_n69), .Z0_f (new_AGEMA_signal_2550), .Z1_t (new_AGEMA_signal_2551), .Z1_f (new_AGEMA_signal_2552) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U137 ( .A0_t (StateOut[157]), .A0_f (new_AGEMA_signal_2553), .A1_t (new_AGEMA_signal_2554), .A1_f (new_AGEMA_signal_2555), .B0_t (StateOut[149]), .B0_f (new_AGEMA_signal_2556), .B1_t (new_AGEMA_signal_2557), .B1_f (new_AGEMA_signal_2558), .Z0_t (THETA_n70), .Z0_f (new_AGEMA_signal_2559), .Z1_t (new_AGEMA_signal_2560), .Z1_f (new_AGEMA_signal_2561) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U136 ( .A0_t (StateOut[76]), .A0_f (new_AGEMA_signal_2610), .A1_t (new_AGEMA_signal_2611), .A1_f (new_AGEMA_signal_2612), .B0_t (THETA_n68), .B0_f (new_AGEMA_signal_3342), .B1_t (new_AGEMA_signal_3343), .B1_f (new_AGEMA_signal_3344), .Z0_t (StateFromRhoPi[198]), .Z0_f (new_AGEMA_signal_3806), .Z1_t (new_AGEMA_signal_3807), .Z1_f (new_AGEMA_signal_3808) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U135 ( .A0_t (StateOut[68]), .A0_f (new_AGEMA_signal_2607), .A1_t (new_AGEMA_signal_2608), .A1_f (new_AGEMA_signal_2609), .B0_t (THETA_n68), .B0_f (new_AGEMA_signal_3342), .B1_t (new_AGEMA_signal_3343), .B1_f (new_AGEMA_signal_3344), .Z0_t (StateFromRhoPi[129]), .Z0_f (new_AGEMA_signal_3809), .Z1_t (new_AGEMA_signal_3810), .Z1_f (new_AGEMA_signal_3811) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U134 ( .A0_t (StateOut[60]), .A0_f (new_AGEMA_signal_3162), .A1_t (new_AGEMA_signal_3163), .A1_f (new_AGEMA_signal_3164), .B0_t (THETA_n68), .B0_f (new_AGEMA_signal_3342), .B1_t (new_AGEMA_signal_3343), .B1_f (new_AGEMA_signal_3344), .Z0_t (StateFromRhoPi[110]), .Z0_f (new_AGEMA_signal_3812), .Z1_t (new_AGEMA_signal_3813), .Z1_f (new_AGEMA_signal_3814) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U133 ( .A0_t (StateOut[52]), .A0_f (new_AGEMA_signal_2598), .A1_t (new_AGEMA_signal_2599), .A1_f (new_AGEMA_signal_2600), .B0_t (THETA_n68), .B0_f (new_AGEMA_signal_3342), .B1_t (new_AGEMA_signal_3343), .B1_f (new_AGEMA_signal_3344), .Z0_t (StateFromRhoPi[40]), .Z0_f (new_AGEMA_signal_3815), .Z1_t (new_AGEMA_signal_3816), .Z1_f (new_AGEMA_signal_3817) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U132 ( .A0_t (StateOut[44]), .A0_f (new_AGEMA_signal_2601), .A1_t (new_AGEMA_signal_2602), .A1_f (new_AGEMA_signal_2603), .B0_t (THETA_n68), .B0_f (new_AGEMA_signal_3342), .B1_t (new_AGEMA_signal_3343), .B1_f (new_AGEMA_signal_3344), .Z0_t (StateFromRhoPi[21]), .Z0_f (new_AGEMA_signal_3818), .Z1_t (new_AGEMA_signal_3819), .Z1_f (new_AGEMA_signal_3820) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U131 ( .A0_t (THETA_n67), .A0_f (new_AGEMA_signal_3237), .A1_t (new_AGEMA_signal_3238), .A1_f (new_AGEMA_signal_3239), .B0_t (THETA_n72), .B0_f (new_AGEMA_signal_3153), .B1_t (new_AGEMA_signal_3154), .B1_f (new_AGEMA_signal_3155), .Z0_t (THETA_n68), .Z0_f (new_AGEMA_signal_3342), .Z1_t (new_AGEMA_signal_3343), .Z1_f (new_AGEMA_signal_3344) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U130 ( .A0_t (OutData_s0_t[4]), .A0_f (OutData_s0_f[4]), .A1_t (OutData_s1_t[4]), .A1_f (OutData_s1_f[4]), .B0_t (THETA_n66), .B0_f (new_AGEMA_signal_2940), .B1_t (new_AGEMA_signal_2941), .B1_f (new_AGEMA_signal_2942), .Z0_t (THETA_n72), .Z0_f (new_AGEMA_signal_3153), .Z1_t (new_AGEMA_signal_3154), .Z1_f (new_AGEMA_signal_3155) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U129 ( .A0_t (THETA_n65), .A0_f (new_AGEMA_signal_2577), .A1_t (new_AGEMA_signal_2578), .A1_f (new_AGEMA_signal_2579), .B0_t (THETA_n64), .B0_f (new_AGEMA_signal_2568), .B1_t (new_AGEMA_signal_2569), .B1_f (new_AGEMA_signal_2570), .Z0_t (THETA_n66), .Z0_f (new_AGEMA_signal_2940), .Z1_t (new_AGEMA_signal_2941), .Z1_f (new_AGEMA_signal_2942) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U128 ( .A0_t (StateOut[12]), .A0_f (new_AGEMA_signal_2562), .A1_t (new_AGEMA_signal_2563), .A1_f (new_AGEMA_signal_2564), .B0_t (StateOut[20]), .B0_f (new_AGEMA_signal_2565), .B1_t (new_AGEMA_signal_2566), .B1_f (new_AGEMA_signal_2567), .Z0_t (THETA_n64), .Z0_f (new_AGEMA_signal_2568), .Z1_t (new_AGEMA_signal_2569), .Z1_f (new_AGEMA_signal_2570) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U127 ( .A0_t (StateOut[36]), .A0_f (new_AGEMA_signal_2571), .A1_t (new_AGEMA_signal_2572), .A1_f (new_AGEMA_signal_2573), .B0_t (StateOut[28]), .B0_f (new_AGEMA_signal_2574), .B1_t (new_AGEMA_signal_2575), .B1_f (new_AGEMA_signal_2576), .Z0_t (THETA_n65), .Z0_f (new_AGEMA_signal_2577), .Z1_t (new_AGEMA_signal_2578), .Z1_f (new_AGEMA_signal_2579) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U126 ( .A0_t (StateOut[116]), .A0_f (new_AGEMA_signal_2808), .A1_t (new_AGEMA_signal_2809), .A1_f (new_AGEMA_signal_2810), .B0_t (THETA_n63), .B0_f (new_AGEMA_signal_3345), .B1_t (new_AGEMA_signal_3346), .B1_f (new_AGEMA_signal_3347), .Z0_t (StateFromRhoPi[169]), .Z0_f (new_AGEMA_signal_3821), .Z1_t (new_AGEMA_signal_3822), .Z1_f (new_AGEMA_signal_3823) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U125 ( .A0_t (StateOut[108]), .A0_f (new_AGEMA_signal_2805), .A1_t (new_AGEMA_signal_2806), .A1_f (new_AGEMA_signal_2807), .B0_t (THETA_n63), .B0_f (new_AGEMA_signal_3345), .B1_t (new_AGEMA_signal_3346), .B1_f (new_AGEMA_signal_3347), .Z0_t (StateFromRhoPi[147]), .Z0_f (new_AGEMA_signal_3824), .Z1_t (new_AGEMA_signal_3825), .Z1_f (new_AGEMA_signal_3826) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U124 ( .A0_t (StateOut[100]), .A0_f (new_AGEMA_signal_3228), .A1_t (new_AGEMA_signal_3229), .A1_f (new_AGEMA_signal_3230), .B0_t (THETA_n63), .B0_f (new_AGEMA_signal_3345), .B1_t (new_AGEMA_signal_3346), .B1_f (new_AGEMA_signal_3347), .Z0_t (StateFromRhoPi[87]), .Z0_f (new_AGEMA_signal_3827), .Z1_t (new_AGEMA_signal_3828), .Z1_f (new_AGEMA_signal_3829) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U123 ( .A0_t (StateOut[92]), .A0_f (new_AGEMA_signal_2796), .A1_t (new_AGEMA_signal_2797), .A1_f (new_AGEMA_signal_2798), .B0_t (THETA_n63), .B0_f (new_AGEMA_signal_3345), .B1_t (new_AGEMA_signal_3346), .B1_f (new_AGEMA_signal_3347), .Z0_t (StateFromRhoPi[58]), .Z0_f (new_AGEMA_signal_3830), .Z1_t (new_AGEMA_signal_3831), .Z1_f (new_AGEMA_signal_3832) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U122 ( .A0_t (StateOut[84]), .A0_f (new_AGEMA_signal_2799), .A1_t (new_AGEMA_signal_2800), .A1_f (new_AGEMA_signal_2801), .B0_t (THETA_n63), .B0_f (new_AGEMA_signal_3345), .B1_t (new_AGEMA_signal_3346), .B1_f (new_AGEMA_signal_3347), .Z0_t (StateFromRhoPi[34]), .Z0_f (new_AGEMA_signal_3833), .Z1_t (new_AGEMA_signal_3834), .Z1_f (new_AGEMA_signal_3835) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U121 ( .A0_t (THETA_n62), .A0_f (new_AGEMA_signal_3165), .A1_t (new_AGEMA_signal_3166), .A1_f (new_AGEMA_signal_3167), .B0_t (THETA_n77), .B0_f (new_AGEMA_signal_3159), .B1_t (new_AGEMA_signal_3160), .B1_f (new_AGEMA_signal_3161), .Z0_t (THETA_n63), .Z0_f (new_AGEMA_signal_3345), .Z1_t (new_AGEMA_signal_3346), .Z1_f (new_AGEMA_signal_3347) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U120 ( .A0_t (StateOut[123]), .A0_f (new_AGEMA_signal_3156), .A1_t (new_AGEMA_signal_3157), .A1_f (new_AGEMA_signal_3158), .B0_t (THETA_n61), .B0_f (new_AGEMA_signal_2943), .B1_t (new_AGEMA_signal_2944), .B1_f (new_AGEMA_signal_2945), .Z0_t (THETA_n77), .Z0_f (new_AGEMA_signal_3159), .Z1_t (new_AGEMA_signal_3160), .Z1_f (new_AGEMA_signal_3161) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U119 ( .A0_t (THETA_n60), .A0_f (new_AGEMA_signal_2595), .A1_t (new_AGEMA_signal_2596), .A1_f (new_AGEMA_signal_2597), .B0_t (THETA_n59), .B0_f (new_AGEMA_signal_2586), .B1_t (new_AGEMA_signal_2587), .B1_f (new_AGEMA_signal_2588), .Z0_t (THETA_n61), .Z0_f (new_AGEMA_signal_2943), .Z1_t (new_AGEMA_signal_2944), .Z1_f (new_AGEMA_signal_2945) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U118 ( .A0_t (StateOut[131]), .A0_f (new_AGEMA_signal_2580), .A1_t (new_AGEMA_signal_2581), .A1_f (new_AGEMA_signal_2582), .B0_t (StateOut[139]), .B0_f (new_AGEMA_signal_2583), .B1_t (new_AGEMA_signal_2584), .B1_f (new_AGEMA_signal_2585), .Z0_t (THETA_n59), .Z0_f (new_AGEMA_signal_2586), .Z1_t (new_AGEMA_signal_2587), .Z1_f (new_AGEMA_signal_2588) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U117 ( .A0_t (StateOut[155]), .A0_f (new_AGEMA_signal_2589), .A1_t (new_AGEMA_signal_2590), .A1_f (new_AGEMA_signal_2591), .B0_t (StateOut[147]), .B0_f (new_AGEMA_signal_2592), .B1_t (new_AGEMA_signal_2593), .B1_f (new_AGEMA_signal_2594), .Z0_t (THETA_n60), .Z0_f (new_AGEMA_signal_2595), .Z1_t (new_AGEMA_signal_2596), .Z1_f (new_AGEMA_signal_2597) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U116 ( .A0_t (StateOut[37]), .A0_f (new_AGEMA_signal_2643), .A1_t (new_AGEMA_signal_2644), .A1_f (new_AGEMA_signal_2645), .B0_t (THETA_n58), .B0_f (new_AGEMA_signal_3348), .B1_t (new_AGEMA_signal_3349), .B1_f (new_AGEMA_signal_3350), .Z0_t (StateFromRhoPi[183]), .Z0_f (new_AGEMA_signal_3836), .Z1_t (new_AGEMA_signal_3837), .Z1_f (new_AGEMA_signal_3838) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U115 ( .A0_t (StateOut[29]), .A0_f (new_AGEMA_signal_3174), .A1_t (new_AGEMA_signal_3175), .A1_f (new_AGEMA_signal_3176), .B0_t (THETA_n58), .B0_f (new_AGEMA_signal_3348), .B1_t (new_AGEMA_signal_3349), .B1_f (new_AGEMA_signal_3350), .Z0_t (StateFromRhoPi[158]), .Z0_f (new_AGEMA_signal_3839), .Z1_t (new_AGEMA_signal_3840), .Z1_f (new_AGEMA_signal_3841) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U114 ( .A0_t (StateOut[21]), .A0_f (new_AGEMA_signal_2646), .A1_t (new_AGEMA_signal_2647), .A1_f (new_AGEMA_signal_2648), .B0_t (THETA_n58), .B0_f (new_AGEMA_signal_3348), .B1_t (new_AGEMA_signal_3349), .B1_f (new_AGEMA_signal_3350), .Z0_t (StateFromRhoPi[88]), .Z0_f (new_AGEMA_signal_3842), .Z1_t (new_AGEMA_signal_3843), .Z1_f (new_AGEMA_signal_3844) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U113 ( .A0_t (StateOut[13]), .A0_f (new_AGEMA_signal_2634), .A1_t (new_AGEMA_signal_2635), .A1_f (new_AGEMA_signal_2636), .B0_t (THETA_n58), .B0_f (new_AGEMA_signal_3348), .B1_t (new_AGEMA_signal_3349), .B1_f (new_AGEMA_signal_3350), .Z0_t (StateFromRhoPi[65]), .Z0_f (new_AGEMA_signal_3845), .Z1_t (new_AGEMA_signal_3846), .Z1_f (new_AGEMA_signal_3847) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U112 ( .A0_t (OutData_s0_t[5]), .A0_f (OutData_s0_f[5]), .A1_t (OutData_s1_t[5]), .A1_f (OutData_s1_f[5]), .B0_t (THETA_n58), .B0_f (new_AGEMA_signal_3348), .B1_t (new_AGEMA_signal_3349), .B1_f (new_AGEMA_signal_3350), .Z0_t (StateFromRhoPi[5]), .Z0_f (new_AGEMA_signal_3848), .Z1_t (new_AGEMA_signal_3849), .Z1_f (new_AGEMA_signal_3850) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U111 ( .A0_t (THETA_n57), .A0_f (new_AGEMA_signal_3189), .A1_t (new_AGEMA_signal_3190), .A1_f (new_AGEMA_signal_3191), .B0_t (THETA_n62), .B0_f (new_AGEMA_signal_3165), .B1_t (new_AGEMA_signal_3166), .B1_f (new_AGEMA_signal_3167), .Z0_t (THETA_n58), .Z0_f (new_AGEMA_signal_3348), .Z1_t (new_AGEMA_signal_3349), .Z1_f (new_AGEMA_signal_3350) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U110 ( .A0_t (StateOut[60]), .A0_f (new_AGEMA_signal_3162), .A1_t (new_AGEMA_signal_3163), .A1_f (new_AGEMA_signal_3164), .B0_t (THETA_n56), .B0_f (new_AGEMA_signal_2946), .B1_t (new_AGEMA_signal_2947), .B1_f (new_AGEMA_signal_2948), .Z0_t (THETA_n62), .Z0_f (new_AGEMA_signal_3165), .Z1_t (new_AGEMA_signal_3166), .Z1_f (new_AGEMA_signal_3167) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U109 ( .A0_t (THETA_n55), .A0_f (new_AGEMA_signal_2613), .A1_t (new_AGEMA_signal_2614), .A1_f (new_AGEMA_signal_2615), .B0_t (THETA_n54), .B0_f (new_AGEMA_signal_2604), .B1_t (new_AGEMA_signal_2605), .B1_f (new_AGEMA_signal_2606), .Z0_t (THETA_n56), .Z0_f (new_AGEMA_signal_2946), .Z1_t (new_AGEMA_signal_2947), .Z1_f (new_AGEMA_signal_2948) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U108 ( .A0_t (StateOut[52]), .A0_f (new_AGEMA_signal_2598), .A1_t (new_AGEMA_signal_2599), .A1_f (new_AGEMA_signal_2600), .B0_t (StateOut[44]), .B0_f (new_AGEMA_signal_2601), .B1_t (new_AGEMA_signal_2602), .B1_f (new_AGEMA_signal_2603), .Z0_t (THETA_n54), .Z0_f (new_AGEMA_signal_2604), .Z1_t (new_AGEMA_signal_2605), .Z1_f (new_AGEMA_signal_2606) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U107 ( .A0_t (StateOut[68]), .A0_f (new_AGEMA_signal_2607), .A1_t (new_AGEMA_signal_2608), .A1_f (new_AGEMA_signal_2609), .B0_t (StateOut[76]), .B0_f (new_AGEMA_signal_2610), .B1_t (new_AGEMA_signal_2611), .B1_f (new_AGEMA_signal_2612), .Z0_t (THETA_n55), .Z0_f (new_AGEMA_signal_2613), .Z1_t (new_AGEMA_signal_2614), .Z1_f (new_AGEMA_signal_2615) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U106 ( .A0_t (StateOut[115]), .A0_f (new_AGEMA_signal_2823), .A1_t (new_AGEMA_signal_2824), .A1_f (new_AGEMA_signal_2825), .B0_t (THETA_n53), .B0_f (new_AGEMA_signal_3351), .B1_t (new_AGEMA_signal_3352), .B1_f (new_AGEMA_signal_3353), .Z0_t (StateFromRhoPi[168]), .Z0_f (new_AGEMA_signal_3851), .Z1_t (new_AGEMA_signal_3852), .Z1_f (new_AGEMA_signal_3853) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U105 ( .A0_t (StateOut[107]), .A0_f (new_AGEMA_signal_3234), .A1_t (new_AGEMA_signal_3235), .A1_f (new_AGEMA_signal_3236), .B0_t (THETA_n53), .B0_f (new_AGEMA_signal_3351), .B1_t (new_AGEMA_signal_3352), .B1_f (new_AGEMA_signal_3353), .Z0_t (StateFromRhoPi[146]), .Z0_f (new_AGEMA_signal_3854), .Z1_t (new_AGEMA_signal_3855), .Z1_f (new_AGEMA_signal_3856) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U104 ( .A0_t (StateOut[99]), .A0_f (new_AGEMA_signal_2826), .A1_t (new_AGEMA_signal_2827), .A1_f (new_AGEMA_signal_2828), .B0_t (THETA_n53), .B0_f (new_AGEMA_signal_3351), .B1_t (new_AGEMA_signal_3352), .B1_f (new_AGEMA_signal_3353), .Z0_t (StateFromRhoPi[86]), .Z0_f (new_AGEMA_signal_3857), .Z1_t (new_AGEMA_signal_3858), .Z1_f (new_AGEMA_signal_3859) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U103 ( .A0_t (StateOut[91]), .A0_f (new_AGEMA_signal_2814), .A1_t (new_AGEMA_signal_2815), .A1_f (new_AGEMA_signal_2816), .B0_t (THETA_n53), .B0_f (new_AGEMA_signal_3351), .B1_t (new_AGEMA_signal_3352), .B1_f (new_AGEMA_signal_3353), .Z0_t (StateFromRhoPi[57]), .Z0_f (new_AGEMA_signal_3860), .Z1_t (new_AGEMA_signal_3861), .Z1_f (new_AGEMA_signal_3862) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U102 ( .A0_t (StateOut[83]), .A0_f (new_AGEMA_signal_2817), .A1_t (new_AGEMA_signal_2818), .A1_f (new_AGEMA_signal_2819), .B0_t (THETA_n53), .B0_f (new_AGEMA_signal_3351), .B1_t (new_AGEMA_signal_3352), .B1_f (new_AGEMA_signal_3353), .Z0_t (StateFromRhoPi[33]), .Z0_f (new_AGEMA_signal_3863), .Z1_t (new_AGEMA_signal_3864), .Z1_f (new_AGEMA_signal_3865) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U101 ( .A0_t (THETA_n52), .A0_f (new_AGEMA_signal_3213), .A1_t (new_AGEMA_signal_3214), .A1_f (new_AGEMA_signal_3215), .B0_t (THETA_n51), .B0_f (new_AGEMA_signal_3171), .B1_t (new_AGEMA_signal_3172), .B1_f (new_AGEMA_signal_3173), .Z0_t (THETA_n53), .Z0_f (new_AGEMA_signal_3351), .Z1_t (new_AGEMA_signal_3352), .Z1_f (new_AGEMA_signal_3353) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U100 ( .A0_t (StateOut[36]), .A0_f (new_AGEMA_signal_2571), .A1_t (new_AGEMA_signal_2572), .A1_f (new_AGEMA_signal_2573), .B0_t (THETA_n50), .B0_f (new_AGEMA_signal_3354), .B1_t (new_AGEMA_signal_3355), .B1_f (new_AGEMA_signal_3356), .Z0_t (StateFromRhoPi[182]), .Z0_f (new_AGEMA_signal_3866), .Z1_t (new_AGEMA_signal_3867), .Z1_f (new_AGEMA_signal_3868) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U99 ( .A0_t (StateOut[28]), .A0_f (new_AGEMA_signal_2574), .A1_t (new_AGEMA_signal_2575), .A1_f (new_AGEMA_signal_2576), .B0_t (THETA_n50), .B0_f (new_AGEMA_signal_3354), .B1_t (new_AGEMA_signal_3355), .B1_f (new_AGEMA_signal_3356), .Z0_t (StateFromRhoPi[157]), .Z0_f (new_AGEMA_signal_3869), .Z1_t (new_AGEMA_signal_3870), .Z1_f (new_AGEMA_signal_3871) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U98 ( .A0_t (StateOut[20]), .A0_f (new_AGEMA_signal_2565), .A1_t (new_AGEMA_signal_2566), .A1_f (new_AGEMA_signal_2567), .B0_t (THETA_n50), .B0_f (new_AGEMA_signal_3354), .B1_t (new_AGEMA_signal_3355), .B1_f (new_AGEMA_signal_3356), .Z0_t (StateFromRhoPi[95]), .Z0_f (new_AGEMA_signal_3872), .Z1_t (new_AGEMA_signal_3873), .Z1_f (new_AGEMA_signal_3874) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U97 ( .A0_t (StateOut[12]), .A0_f (new_AGEMA_signal_2562), .A1_t (new_AGEMA_signal_2563), .A1_f (new_AGEMA_signal_2564), .B0_t (THETA_n50), .B0_f (new_AGEMA_signal_3354), .B1_t (new_AGEMA_signal_3355), .B1_f (new_AGEMA_signal_3356), .Z0_t (StateFromRhoPi[64]), .Z0_f (new_AGEMA_signal_3875), .Z1_t (new_AGEMA_signal_3876), .Z1_f (new_AGEMA_signal_3877) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U96 ( .A0_t (OutData_s0_t[4]), .A0_f (OutData_s0_f[4]), .A1_t (OutData_s1_t[4]), .A1_f (OutData_s1_f[4]), .B0_t (THETA_n50), .B0_f (new_AGEMA_signal_3354), .B1_t (new_AGEMA_signal_3355), .B1_f (new_AGEMA_signal_3356), .Z0_t (StateFromRhoPi[4]), .Z0_f (new_AGEMA_signal_3878), .Z1_t (new_AGEMA_signal_3879), .Z1_f (new_AGEMA_signal_3880) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U95 ( .A0_t (THETA_n49), .A0_f (new_AGEMA_signal_3201), .A1_t (new_AGEMA_signal_3202), .A1_f (new_AGEMA_signal_3203), .B0_t (THETA_n51), .B0_f (new_AGEMA_signal_3171), .B1_t (new_AGEMA_signal_3172), .B1_f (new_AGEMA_signal_3173), .Z0_t (THETA_n50), .Z0_f (new_AGEMA_signal_3354), .Z1_t (new_AGEMA_signal_3355), .Z1_f (new_AGEMA_signal_3356) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U94 ( .A0_t (StateOut[59]), .A0_f (new_AGEMA_signal_3168), .A1_t (new_AGEMA_signal_3169), .A1_f (new_AGEMA_signal_3170), .B0_t (THETA_n48), .B0_f (new_AGEMA_signal_2949), .B1_t (new_AGEMA_signal_2950), .B1_f (new_AGEMA_signal_2951), .Z0_t (THETA_n51), .Z0_f (new_AGEMA_signal_3171), .Z1_t (new_AGEMA_signal_3172), .Z1_f (new_AGEMA_signal_3173) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U93 ( .A0_t (THETA_n47), .A0_f (new_AGEMA_signal_2631), .A1_t (new_AGEMA_signal_2632), .A1_f (new_AGEMA_signal_2633), .B0_t (THETA_n46), .B0_f (new_AGEMA_signal_2622), .B1_t (new_AGEMA_signal_2623), .B1_f (new_AGEMA_signal_2624), .Z0_t (THETA_n48), .Z0_f (new_AGEMA_signal_2949), .Z1_t (new_AGEMA_signal_2950), .Z1_f (new_AGEMA_signal_2951) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U92 ( .A0_t (StateOut[51]), .A0_f (new_AGEMA_signal_2616), .A1_t (new_AGEMA_signal_2617), .A1_f (new_AGEMA_signal_2618), .B0_t (StateOut[43]), .B0_f (new_AGEMA_signal_2619), .B1_t (new_AGEMA_signal_2620), .B1_f (new_AGEMA_signal_2621), .Z0_t (THETA_n46), .Z0_f (new_AGEMA_signal_2622), .Z1_t (new_AGEMA_signal_2623), .Z1_f (new_AGEMA_signal_2624) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U91 ( .A0_t (StateOut[67]), .A0_f (new_AGEMA_signal_2625), .A1_t (new_AGEMA_signal_2626), .A1_f (new_AGEMA_signal_2627), .B0_t (StateOut[75]), .B0_f (new_AGEMA_signal_2628), .B1_t (new_AGEMA_signal_2629), .B1_f (new_AGEMA_signal_2630), .Z0_t (THETA_n47), .Z0_f (new_AGEMA_signal_2631), .Z1_t (new_AGEMA_signal_2632), .Z1_f (new_AGEMA_signal_2633) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U90 ( .A0_t (StateOut[77]), .A0_f (new_AGEMA_signal_2517), .A1_t (new_AGEMA_signal_2518), .A1_f (new_AGEMA_signal_2519), .B0_t (THETA_n45), .B0_f (new_AGEMA_signal_3357), .B1_t (new_AGEMA_signal_3358), .B1_f (new_AGEMA_signal_3359), .Z0_t (StateFromRhoPi[199]), .Z0_f (new_AGEMA_signal_3881), .Z1_t (new_AGEMA_signal_3882), .Z1_f (new_AGEMA_signal_3883) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U89 ( .A0_t (StateOut[69]), .A0_f (new_AGEMA_signal_2520), .A1_t (new_AGEMA_signal_2521), .A1_f (new_AGEMA_signal_2522), .B0_t (THETA_n45), .B0_f (new_AGEMA_signal_3357), .B1_t (new_AGEMA_signal_3358), .B1_f (new_AGEMA_signal_3359), .Z0_t (StateFromRhoPi[130]), .Z0_f (new_AGEMA_signal_3884), .Z1_t (new_AGEMA_signal_3885), .Z1_f (new_AGEMA_signal_3886) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U88 ( .A0_t (StateOut[61]), .A0_f (new_AGEMA_signal_2511), .A1_t (new_AGEMA_signal_2512), .A1_f (new_AGEMA_signal_2513), .B0_t (THETA_n45), .B0_f (new_AGEMA_signal_3357), .B1_t (new_AGEMA_signal_3358), .B1_f (new_AGEMA_signal_3359), .Z0_t (StateFromRhoPi[111]), .Z0_f (new_AGEMA_signal_3887), .Z1_t (new_AGEMA_signal_3888), .Z1_f (new_AGEMA_signal_3889) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U87 ( .A0_t (StateOut[53]), .A0_f (new_AGEMA_signal_2508), .A1_t (new_AGEMA_signal_2509), .A1_f (new_AGEMA_signal_2510), .B0_t (THETA_n45), .B0_f (new_AGEMA_signal_3357), .B1_t (new_AGEMA_signal_3358), .B1_f (new_AGEMA_signal_3359), .Z0_t (StateFromRhoPi[41]), .Z0_f (new_AGEMA_signal_3890), .Z1_t (new_AGEMA_signal_3891), .Z1_f (new_AGEMA_signal_3892) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U86 ( .A0_t (StateOut[45]), .A0_f (new_AGEMA_signal_3132), .A1_t (new_AGEMA_signal_3133), .A1_f (new_AGEMA_signal_3134), .B0_t (THETA_n45), .B0_f (new_AGEMA_signal_3357), .B1_t (new_AGEMA_signal_3358), .B1_f (new_AGEMA_signal_3359), .Z0_t (StateFromRhoPi[22]), .Z0_f (new_AGEMA_signal_3893), .Z1_t (new_AGEMA_signal_3894), .Z1_f (new_AGEMA_signal_3895) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U85 ( .A0_t (THETA_n44), .A0_f (new_AGEMA_signal_3231), .A1_t (new_AGEMA_signal_3232), .A1_f (new_AGEMA_signal_3233), .B0_t (THETA_n186), .B0_f (new_AGEMA_signal_3177), .B1_t (new_AGEMA_signal_3178), .B1_f (new_AGEMA_signal_3179), .Z0_t (THETA_n45), .Z0_f (new_AGEMA_signal_3357), .Z1_t (new_AGEMA_signal_3358), .Z1_f (new_AGEMA_signal_3359) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U84 ( .A0_t (StateOut[29]), .A0_f (new_AGEMA_signal_3174), .A1_t (new_AGEMA_signal_3175), .A1_f (new_AGEMA_signal_3176), .B0_t (THETA_n43), .B0_f (new_AGEMA_signal_2952), .B1_t (new_AGEMA_signal_2953), .B1_f (new_AGEMA_signal_2954), .Z0_t (THETA_n186), .Z0_f (new_AGEMA_signal_3177), .Z1_t (new_AGEMA_signal_3178), .Z1_f (new_AGEMA_signal_3179) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U83 ( .A0_t (THETA_n42), .A0_f (new_AGEMA_signal_2649), .A1_t (new_AGEMA_signal_2650), .A1_f (new_AGEMA_signal_2651), .B0_t (THETA_n41), .B0_f (new_AGEMA_signal_2640), .B1_t (new_AGEMA_signal_2641), .B1_f (new_AGEMA_signal_2642), .Z0_t (THETA_n43), .Z0_f (new_AGEMA_signal_2952), .Z1_t (new_AGEMA_signal_2953), .Z1_f (new_AGEMA_signal_2954) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U82 ( .A0_t (StateOut[13]), .A0_f (new_AGEMA_signal_2634), .A1_t (new_AGEMA_signal_2635), .A1_f (new_AGEMA_signal_2636), .B0_t (OutData_s0_t[5]), .B0_f (OutData_s0_f[5]), .B1_t (OutData_s1_t[5]), .B1_f (OutData_s1_f[5]), .Z0_t (THETA_n41), .Z0_f (new_AGEMA_signal_2640), .Z1_t (new_AGEMA_signal_2641), .Z1_f (new_AGEMA_signal_2642) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U81 ( .A0_t (StateOut[37]), .A0_f (new_AGEMA_signal_2643), .A1_t (new_AGEMA_signal_2644), .A1_f (new_AGEMA_signal_2645), .B0_t (StateOut[21]), .B0_f (new_AGEMA_signal_2646), .B1_t (new_AGEMA_signal_2647), .B1_f (new_AGEMA_signal_2648), .Z0_t (THETA_n42), .Z0_f (new_AGEMA_signal_2649), .Z1_t (new_AGEMA_signal_2650), .Z1_f (new_AGEMA_signal_2651) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U80 ( .A0_t (StateOut[35]), .A0_f (new_AGEMA_signal_2193), .A1_t (new_AGEMA_signal_2194), .A1_f (new_AGEMA_signal_2195), .B0_t (THETA_n40), .B0_f (new_AGEMA_signal_3360), .B1_t (new_AGEMA_signal_3361), .B1_f (new_AGEMA_signal_3362), .Z0_t (StateFromRhoPi[181]), .Z0_f (new_AGEMA_signal_3896), .Z1_t (new_AGEMA_signal_3897), .Z1_f (new_AGEMA_signal_3898) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U79 ( .A0_t (StateOut[27]), .A0_f (new_AGEMA_signal_2196), .A1_t (new_AGEMA_signal_2197), .A1_f (new_AGEMA_signal_2198), .B0_t (THETA_n40), .B0_f (new_AGEMA_signal_3360), .B1_t (new_AGEMA_signal_3361), .B1_f (new_AGEMA_signal_3362), .Z0_t (StateFromRhoPi[156]), .Z0_f (new_AGEMA_signal_3899), .Z1_t (new_AGEMA_signal_3900), .Z1_f (new_AGEMA_signal_3901) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U78 ( .A0_t (StateOut[19]), .A0_f (new_AGEMA_signal_2187), .A1_t (new_AGEMA_signal_2188), .A1_f (new_AGEMA_signal_2189), .B0_t (THETA_n40), .B0_f (new_AGEMA_signal_3360), .B1_t (new_AGEMA_signal_3361), .B1_f (new_AGEMA_signal_3362), .Z0_t (StateFromRhoPi[94]), .Z0_f (new_AGEMA_signal_3902), .Z1_t (new_AGEMA_signal_3903), .Z1_f (new_AGEMA_signal_3904) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U77 ( .A0_t (StateOut[11]), .A0_f (new_AGEMA_signal_2184), .A1_t (new_AGEMA_signal_2185), .A1_f (new_AGEMA_signal_2186), .B0_t (THETA_n40), .B0_f (new_AGEMA_signal_3360), .B1_t (new_AGEMA_signal_3361), .B1_f (new_AGEMA_signal_3362), .Z0_t (StateFromRhoPi[71]), .Z0_f (new_AGEMA_signal_3905), .Z1_t (new_AGEMA_signal_3906), .Z1_f (new_AGEMA_signal_3907) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U76 ( .A0_t (OutData_s0_t[3]), .A0_f (OutData_s0_f[3]), .A1_t (OutData_s1_t[3]), .A1_f (OutData_s1_f[3]), .B0_t (THETA_n40), .B0_f (new_AGEMA_signal_3360), .B1_t (new_AGEMA_signal_3361), .B1_f (new_AGEMA_signal_3362), .Z0_t (StateFromRhoPi[3]), .Z0_f (new_AGEMA_signal_3908), .Z1_t (new_AGEMA_signal_3909), .Z1_f (new_AGEMA_signal_3910) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U75 ( .A0_t (THETA_n39), .A0_f (new_AGEMA_signal_3225), .A1_t (new_AGEMA_signal_3226), .A1_f (new_AGEMA_signal_3227), .B0_t (THETA_n150), .B0_f (new_AGEMA_signal_3183), .B1_t (new_AGEMA_signal_3184), .B1_f (new_AGEMA_signal_3185), .Z0_t (THETA_n40), .Z0_f (new_AGEMA_signal_3360), .Z1_t (new_AGEMA_signal_3361), .Z1_f (new_AGEMA_signal_3362) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U74 ( .A0_t (StateOut[66]), .A0_f (new_AGEMA_signal_3180), .A1_t (new_AGEMA_signal_3181), .A1_f (new_AGEMA_signal_3182), .B0_t (THETA_n38), .B0_f (new_AGEMA_signal_2955), .B1_t (new_AGEMA_signal_2956), .B1_f (new_AGEMA_signal_2957), .Z0_t (THETA_n150), .Z0_f (new_AGEMA_signal_3183), .Z1_t (new_AGEMA_signal_3184), .Z1_f (new_AGEMA_signal_3185) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U73 ( .A0_t (THETA_n37), .A0_f (new_AGEMA_signal_2667), .A1_t (new_AGEMA_signal_2668), .A1_f (new_AGEMA_signal_2669), .B0_t (THETA_n36), .B0_f (new_AGEMA_signal_2658), .B1_t (new_AGEMA_signal_2659), .B1_f (new_AGEMA_signal_2660), .Z0_t (THETA_n38), .Z0_f (new_AGEMA_signal_2955), .Z1_t (new_AGEMA_signal_2956), .Z1_f (new_AGEMA_signal_2957) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U72 ( .A0_t (StateOut[50]), .A0_f (new_AGEMA_signal_2652), .A1_t (new_AGEMA_signal_2653), .A1_f (new_AGEMA_signal_2654), .B0_t (StateOut[42]), .B0_f (new_AGEMA_signal_2655), .B1_t (new_AGEMA_signal_2656), .B1_f (new_AGEMA_signal_2657), .Z0_t (THETA_n36), .Z0_f (new_AGEMA_signal_2658), .Z1_t (new_AGEMA_signal_2659), .Z1_f (new_AGEMA_signal_2660) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U71 ( .A0_t (StateOut[74]), .A0_f (new_AGEMA_signal_2661), .A1_t (new_AGEMA_signal_2662), .A1_f (new_AGEMA_signal_2663), .B0_t (StateOut[58]), .B0_f (new_AGEMA_signal_2664), .B1_t (new_AGEMA_signal_2665), .B1_f (new_AGEMA_signal_2666), .Z0_t (THETA_n37), .Z0_f (new_AGEMA_signal_2667), .Z1_t (new_AGEMA_signal_2668), .Z1_f (new_AGEMA_signal_2669) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U70 ( .A0_t (StateOut[158]), .A0_f (new_AGEMA_signal_2175), .A1_t (new_AGEMA_signal_2176), .A1_f (new_AGEMA_signal_2177), .B0_t (THETA_n35), .B0_f (new_AGEMA_signal_3363), .B1_t (new_AGEMA_signal_3364), .B1_f (new_AGEMA_signal_3365), .Z0_t (StateFromRhoPi[190]), .Z0_f (new_AGEMA_signal_3911), .Z1_t (new_AGEMA_signal_3912), .Z1_f (new_AGEMA_signal_3913) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U69 ( .A0_t (StateOut[150]), .A0_f (new_AGEMA_signal_2178), .A1_t (new_AGEMA_signal_2179), .A1_f (new_AGEMA_signal_2180), .B0_t (THETA_n35), .B0_f (new_AGEMA_signal_3363), .B1_t (new_AGEMA_signal_3364), .B1_f (new_AGEMA_signal_3365), .Z0_t (StateFromRhoPi[123]), .Z0_f (new_AGEMA_signal_3914), .Z1_t (new_AGEMA_signal_3915), .Z1_f (new_AGEMA_signal_3916) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U68 ( .A0_t (StateOut[142]), .A0_f (new_AGEMA_signal_2169), .A1_t (new_AGEMA_signal_2170), .A1_f (new_AGEMA_signal_2171), .B0_t (THETA_n35), .B0_f (new_AGEMA_signal_3363), .B1_t (new_AGEMA_signal_3364), .B1_f (new_AGEMA_signal_3365), .Z0_t (StateFromRhoPi[103]), .Z0_f (new_AGEMA_signal_3917), .Z1_t (new_AGEMA_signal_3918), .Z1_f (new_AGEMA_signal_3919) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U67 ( .A0_t (StateOut[134]), .A0_f (new_AGEMA_signal_2166), .A1_t (new_AGEMA_signal_2167), .A1_f (new_AGEMA_signal_2168), .B0_t (THETA_n35), .B0_f (new_AGEMA_signal_3363), .B1_t (new_AGEMA_signal_3364), .B1_f (new_AGEMA_signal_3365), .Z0_t (StateFromRhoPi[77]), .Z0_f (new_AGEMA_signal_3920), .Z1_t (new_AGEMA_signal_3921), .Z1_f (new_AGEMA_signal_3922) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U66 ( .A0_t (StateOut[126]), .A0_f (new_AGEMA_signal_3018), .A1_t (new_AGEMA_signal_3019), .A1_f (new_AGEMA_signal_3020), .B0_t (THETA_n35), .B0_f (new_AGEMA_signal_3363), .B1_t (new_AGEMA_signal_3364), .B1_f (new_AGEMA_signal_3365), .Z0_t (StateFromRhoPi[10]), .Z0_f (new_AGEMA_signal_3923), .Z1_t (new_AGEMA_signal_3924), .Z1_f (new_AGEMA_signal_3925) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U65 ( .A0_t (THETA_n127), .A0_f (new_AGEMA_signal_3195), .A1_t (new_AGEMA_signal_3196), .A1_f (new_AGEMA_signal_3197), .B0_t (THETA_n57), .B0_f (new_AGEMA_signal_3189), .B1_t (new_AGEMA_signal_3190), .B1_f (new_AGEMA_signal_3191), .Z0_t (THETA_n35), .Z0_f (new_AGEMA_signal_3363), .Z1_t (new_AGEMA_signal_3364), .Z1_f (new_AGEMA_signal_3365) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U64 ( .A0_t (StateOut[181]), .A0_f (new_AGEMA_signal_3186), .A1_t (new_AGEMA_signal_3187), .A1_f (new_AGEMA_signal_3188), .B0_t (THETA_n34), .B0_f (new_AGEMA_signal_2958), .B1_t (new_AGEMA_signal_2959), .B1_f (new_AGEMA_signal_2960), .Z0_t (THETA_n57), .Z0_f (new_AGEMA_signal_3189), .Z1_t (new_AGEMA_signal_3190), .Z1_f (new_AGEMA_signal_3191) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U63 ( .A0_t (THETA_n33), .A0_f (new_AGEMA_signal_2685), .A1_t (new_AGEMA_signal_2686), .A1_f (new_AGEMA_signal_2687), .B0_t (THETA_n32), .B0_f (new_AGEMA_signal_2676), .B1_t (new_AGEMA_signal_2677), .B1_f (new_AGEMA_signal_2678), .Z0_t (THETA_n34), .Z0_f (new_AGEMA_signal_2958), .Z1_t (new_AGEMA_signal_2959), .Z1_f (new_AGEMA_signal_2960) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U62 ( .A0_t (StateOut[173]), .A0_f (new_AGEMA_signal_2670), .A1_t (new_AGEMA_signal_2671), .A1_f (new_AGEMA_signal_2672), .B0_t (StateOut[165]), .B0_f (new_AGEMA_signal_2673), .B1_t (new_AGEMA_signal_2674), .B1_f (new_AGEMA_signal_2675), .Z0_t (THETA_n32), .Z0_f (new_AGEMA_signal_2676), .Z1_t (new_AGEMA_signal_2677), .Z1_f (new_AGEMA_signal_2678) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U61 ( .A0_t (StateOut[189]), .A0_f (new_AGEMA_signal_2679), .A1_t (new_AGEMA_signal_2680), .A1_f (new_AGEMA_signal_2681), .B0_t (StateOut[197]), .B0_f (new_AGEMA_signal_2682), .B1_t (new_AGEMA_signal_2683), .B1_f (new_AGEMA_signal_2684), .Z0_t (THETA_n33), .Z0_f (new_AGEMA_signal_2685), .Z1_t (new_AGEMA_signal_2686), .Z1_f (new_AGEMA_signal_2687) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U60 ( .A0_t (StateOut[110]), .A0_f (new_AGEMA_signal_3192), .A1_t (new_AGEMA_signal_3193), .A1_f (new_AGEMA_signal_3194), .B0_t (THETA_n31), .B0_f (new_AGEMA_signal_2961), .B1_t (new_AGEMA_signal_2962), .B1_f (new_AGEMA_signal_2963), .Z0_t (THETA_n127), .Z0_f (new_AGEMA_signal_3195), .Z1_t (new_AGEMA_signal_3196), .Z1_f (new_AGEMA_signal_3197) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U59 ( .A0_t (THETA_n30), .A0_f (new_AGEMA_signal_2703), .A1_t (new_AGEMA_signal_2704), .A1_f (new_AGEMA_signal_2705), .B0_t (THETA_n29), .B0_f (new_AGEMA_signal_2694), .B1_t (new_AGEMA_signal_2695), .B1_f (new_AGEMA_signal_2696), .Z0_t (THETA_n31), .Z0_f (new_AGEMA_signal_2961), .Z1_t (new_AGEMA_signal_2962), .Z1_f (new_AGEMA_signal_2963) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U58 ( .A0_t (StateOut[94]), .A0_f (new_AGEMA_signal_2688), .A1_t (new_AGEMA_signal_2689), .A1_f (new_AGEMA_signal_2690), .B0_t (StateOut[86]), .B0_f (new_AGEMA_signal_2691), .B1_t (new_AGEMA_signal_2692), .B1_f (new_AGEMA_signal_2693), .Z0_t (THETA_n29), .Z0_f (new_AGEMA_signal_2694), .Z1_t (new_AGEMA_signal_2695), .Z1_f (new_AGEMA_signal_2696) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U57 ( .A0_t (StateOut[118]), .A0_f (new_AGEMA_signal_2697), .A1_t (new_AGEMA_signal_2698), .A1_f (new_AGEMA_signal_2699), .B0_t (StateOut[102]), .B0_f (new_AGEMA_signal_2700), .B1_t (new_AGEMA_signal_2701), .B1_f (new_AGEMA_signal_2702), .Z0_t (THETA_n30), .Z0_f (new_AGEMA_signal_2703), .Z1_t (new_AGEMA_signal_2704), .Z1_f (new_AGEMA_signal_2705) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U56 ( .A0_t (StateOut[157]), .A0_f (new_AGEMA_signal_2553), .A1_t (new_AGEMA_signal_2554), .A1_f (new_AGEMA_signal_2555), .B0_t (THETA_n28), .B0_f (new_AGEMA_signal_3366), .B1_t (new_AGEMA_signal_3367), .B1_f (new_AGEMA_signal_3368), .Z0_t (StateFromRhoPi[189]), .Z0_f (new_AGEMA_signal_3926), .Z1_t (new_AGEMA_signal_3927), .Z1_f (new_AGEMA_signal_3928) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U55 ( .A0_t (StateOut[149]), .A0_f (new_AGEMA_signal_2556), .A1_t (new_AGEMA_signal_2557), .A1_f (new_AGEMA_signal_2558), .B0_t (THETA_n28), .B0_f (new_AGEMA_signal_3366), .B1_t (new_AGEMA_signal_3367), .B1_f (new_AGEMA_signal_3368), .Z0_t (StateFromRhoPi[122]), .Z0_f (new_AGEMA_signal_3929), .Z1_t (new_AGEMA_signal_3930), .Z1_f (new_AGEMA_signal_3931) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U54 ( .A0_t (StateOut[141]), .A0_f (new_AGEMA_signal_2547), .A1_t (new_AGEMA_signal_2548), .A1_f (new_AGEMA_signal_2549), .B0_t (THETA_n28), .B0_f (new_AGEMA_signal_3366), .B1_t (new_AGEMA_signal_3367), .B1_f (new_AGEMA_signal_3368), .Z0_t (StateFromRhoPi[102]), .Z0_f (new_AGEMA_signal_3932), .Z1_t (new_AGEMA_signal_3933), .Z1_f (new_AGEMA_signal_3934) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U53 ( .A0_t (StateOut[133]), .A0_f (new_AGEMA_signal_2544), .A1_t (new_AGEMA_signal_2545), .A1_f (new_AGEMA_signal_2546), .B0_t (THETA_n28), .B0_f (new_AGEMA_signal_3366), .B1_t (new_AGEMA_signal_3367), .B1_f (new_AGEMA_signal_3368), .Z0_t (StateFromRhoPi[76]), .Z0_f (new_AGEMA_signal_3935), .Z1_t (new_AGEMA_signal_3936), .Z1_f (new_AGEMA_signal_3937) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U52 ( .A0_t (StateOut[125]), .A0_f (new_AGEMA_signal_3144), .A1_t (new_AGEMA_signal_3145), .A1_f (new_AGEMA_signal_3146), .B0_t (THETA_n28), .B0_f (new_AGEMA_signal_3366), .B1_t (new_AGEMA_signal_3367), .B1_f (new_AGEMA_signal_3368), .Z0_t (StateFromRhoPi[9]), .Z0_f (new_AGEMA_signal_3938), .Z1_t (new_AGEMA_signal_3939), .Z1_f (new_AGEMA_signal_3940) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U51 ( .A0_t (THETA_n196), .A0_f (new_AGEMA_signal_3207), .A1_t (new_AGEMA_signal_3208), .A1_f (new_AGEMA_signal_3209), .B0_t (THETA_n49), .B0_f (new_AGEMA_signal_3201), .B1_t (new_AGEMA_signal_3202), .B1_f (new_AGEMA_signal_3203), .Z0_t (THETA_n28), .Z0_f (new_AGEMA_signal_3366), .Z1_t (new_AGEMA_signal_3367), .Z1_f (new_AGEMA_signal_3368) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U50 ( .A0_t (StateOut[180]), .A0_f (new_AGEMA_signal_3198), .A1_t (new_AGEMA_signal_3199), .A1_f (new_AGEMA_signal_3200), .B0_t (THETA_n27), .B0_f (new_AGEMA_signal_2964), .B1_t (new_AGEMA_signal_2965), .B1_f (new_AGEMA_signal_2966), .Z0_t (THETA_n49), .Z0_f (new_AGEMA_signal_3201), .Z1_t (new_AGEMA_signal_3202), .Z1_f (new_AGEMA_signal_3203) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U49 ( .A0_t (THETA_n26), .A0_f (new_AGEMA_signal_2721), .A1_t (new_AGEMA_signal_2722), .A1_f (new_AGEMA_signal_2723), .B0_t (THETA_n25), .B0_f (new_AGEMA_signal_2712), .B1_t (new_AGEMA_signal_2713), .B1_f (new_AGEMA_signal_2714), .Z0_t (THETA_n27), .Z0_f (new_AGEMA_signal_2964), .Z1_t (new_AGEMA_signal_2965), .Z1_f (new_AGEMA_signal_2966) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U48 ( .A0_t (StateOut[172]), .A0_f (new_AGEMA_signal_2706), .A1_t (new_AGEMA_signal_2707), .A1_f (new_AGEMA_signal_2708), .B0_t (StateOut[164]), .B0_f (new_AGEMA_signal_2709), .B1_t (new_AGEMA_signal_2710), .B1_f (new_AGEMA_signal_2711), .Z0_t (THETA_n25), .Z0_f (new_AGEMA_signal_2712), .Z1_t (new_AGEMA_signal_2713), .Z1_f (new_AGEMA_signal_2714) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U47 ( .A0_t (StateOut[188]), .A0_f (new_AGEMA_signal_2715), .A1_t (new_AGEMA_signal_2716), .A1_f (new_AGEMA_signal_2717), .B0_t (StateOut[196]), .B0_f (new_AGEMA_signal_2718), .B1_t (new_AGEMA_signal_2719), .B1_f (new_AGEMA_signal_2720), .Z0_t (THETA_n26), .Z0_f (new_AGEMA_signal_2721), .Z1_t (new_AGEMA_signal_2722), .Z1_f (new_AGEMA_signal_2723) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U46 ( .A0_t (StateOut[109]), .A0_f (new_AGEMA_signal_3204), .A1_t (new_AGEMA_signal_3205), .A1_f (new_AGEMA_signal_3206), .B0_t (THETA_n24), .B0_f (new_AGEMA_signal_2967), .B1_t (new_AGEMA_signal_2968), .B1_f (new_AGEMA_signal_2969), .Z0_t (THETA_n196), .Z0_f (new_AGEMA_signal_3207), .Z1_t (new_AGEMA_signal_3208), .Z1_f (new_AGEMA_signal_3209) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U45 ( .A0_t (THETA_n23), .A0_f (new_AGEMA_signal_2739), .A1_t (new_AGEMA_signal_2740), .A1_f (new_AGEMA_signal_2741), .B0_t (THETA_n22), .B0_f (new_AGEMA_signal_2730), .B1_t (new_AGEMA_signal_2731), .B1_f (new_AGEMA_signal_2732), .Z0_t (THETA_n24), .Z0_f (new_AGEMA_signal_2967), .Z1_t (new_AGEMA_signal_2968), .Z1_f (new_AGEMA_signal_2969) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U44 ( .A0_t (StateOut[93]), .A0_f (new_AGEMA_signal_2724), .A1_t (new_AGEMA_signal_2725), .A1_f (new_AGEMA_signal_2726), .B0_t (StateOut[85]), .B0_f (new_AGEMA_signal_2727), .B1_t (new_AGEMA_signal_2728), .B1_f (new_AGEMA_signal_2729), .Z0_t (THETA_n22), .Z0_f (new_AGEMA_signal_2730), .Z1_t (new_AGEMA_signal_2731), .Z1_f (new_AGEMA_signal_2732) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U43 ( .A0_t (StateOut[117]), .A0_f (new_AGEMA_signal_2733), .A1_t (new_AGEMA_signal_2734), .A1_f (new_AGEMA_signal_2735), .B0_t (StateOut[101]), .B0_f (new_AGEMA_signal_2736), .B1_t (new_AGEMA_signal_2737), .B1_f (new_AGEMA_signal_2738), .Z0_t (THETA_n23), .Z0_f (new_AGEMA_signal_2739), .Z1_t (new_AGEMA_signal_2740), .Z1_f (new_AGEMA_signal_2741) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U42 ( .A0_t (StateOut[194]), .A0_f (new_AGEMA_signal_2841), .A1_t (new_AGEMA_signal_2842), .A1_f (new_AGEMA_signal_2843), .B0_t (THETA_n21), .B0_f (new_AGEMA_signal_3369), .B1_t (new_AGEMA_signal_3370), .B1_f (new_AGEMA_signal_3371), .Z0_t (StateFromRhoPi[160]), .Z0_f (new_AGEMA_signal_3941), .Z1_t (new_AGEMA_signal_3942), .Z1_f (new_AGEMA_signal_3943) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U41 ( .A0_t (StateOut[186]), .A0_f (new_AGEMA_signal_3240), .A1_t (new_AGEMA_signal_3241), .A1_f (new_AGEMA_signal_3242), .B0_t (THETA_n21), .B0_f (new_AGEMA_signal_3369), .B1_t (new_AGEMA_signal_3370), .B1_f (new_AGEMA_signal_3371), .Z0_t (StateFromRhoPi[138]), .Z0_f (new_AGEMA_signal_3944), .Z1_t (new_AGEMA_signal_3945), .Z1_f (new_AGEMA_signal_3946) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U40 ( .A0_t (StateOut[178]), .A0_f (new_AGEMA_signal_2844), .A1_t (new_AGEMA_signal_2845), .A1_f (new_AGEMA_signal_2846), .B0_t (THETA_n21), .B0_f (new_AGEMA_signal_3369), .B1_t (new_AGEMA_signal_3370), .B1_f (new_AGEMA_signal_3371), .Z0_t (StateFromRhoPi[113]), .Z0_f (new_AGEMA_signal_3947), .Z1_t (new_AGEMA_signal_3948), .Z1_f (new_AGEMA_signal_3949) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U39 ( .A0_t (StateOut[170]), .A0_f (new_AGEMA_signal_2832), .A1_t (new_AGEMA_signal_2833), .A1_f (new_AGEMA_signal_2834), .B0_t (THETA_n21), .B0_f (new_AGEMA_signal_3369), .B1_t (new_AGEMA_signal_3370), .B1_f (new_AGEMA_signal_3371), .Z0_t (StateFromRhoPi[54]), .Z0_f (new_AGEMA_signal_3950), .Z1_t (new_AGEMA_signal_3951), .Z1_f (new_AGEMA_signal_3952) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U38 ( .A0_t (StateOut[162]), .A0_f (new_AGEMA_signal_2835), .A1_t (new_AGEMA_signal_2836), .A1_f (new_AGEMA_signal_2837), .B0_t (THETA_n21), .B0_f (new_AGEMA_signal_3369), .B1_t (new_AGEMA_signal_3370), .B1_f (new_AGEMA_signal_3371), .Z0_t (StateFromRhoPi[29]), .Z0_f (new_AGEMA_signal_3953), .Z1_t (new_AGEMA_signal_3954), .Z1_f (new_AGEMA_signal_3955) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U37 ( .A0_t (THETA_n114), .A0_f (new_AGEMA_signal_3219), .A1_t (new_AGEMA_signal_3220), .A1_f (new_AGEMA_signal_3221), .B0_t (THETA_n52), .B0_f (new_AGEMA_signal_3213), .B1_t (new_AGEMA_signal_3214), .B1_f (new_AGEMA_signal_3215), .Z0_t (THETA_n21), .Z0_f (new_AGEMA_signal_3369), .Z1_t (new_AGEMA_signal_3370), .Z1_f (new_AGEMA_signal_3371) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U36 ( .A0_t (StateOut[138]), .A0_f (new_AGEMA_signal_3210), .A1_t (new_AGEMA_signal_3211), .A1_f (new_AGEMA_signal_3212), .B0_t (THETA_n20), .B0_f (new_AGEMA_signal_2970), .B1_t (new_AGEMA_signal_2971), .B1_f (new_AGEMA_signal_2972), .Z0_t (THETA_n52), .Z0_f (new_AGEMA_signal_3213), .Z1_t (new_AGEMA_signal_3214), .Z1_f (new_AGEMA_signal_3215) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U35 ( .A0_t (THETA_n19), .A0_f (new_AGEMA_signal_2757), .A1_t (new_AGEMA_signal_2758), .A1_f (new_AGEMA_signal_2759), .B0_t (THETA_n18), .B0_f (new_AGEMA_signal_2748), .B1_t (new_AGEMA_signal_2749), .B1_f (new_AGEMA_signal_2750), .Z0_t (THETA_n20), .Z0_f (new_AGEMA_signal_2970), .Z1_t (new_AGEMA_signal_2971), .Z1_f (new_AGEMA_signal_2972) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U34 ( .A0_t (StateOut[130]), .A0_f (new_AGEMA_signal_2742), .A1_t (new_AGEMA_signal_2743), .A1_f (new_AGEMA_signal_2744), .B0_t (StateOut[122]), .B0_f (new_AGEMA_signal_2745), .B1_t (new_AGEMA_signal_2746), .B1_f (new_AGEMA_signal_2747), .Z0_t (THETA_n18), .Z0_f (new_AGEMA_signal_2748), .Z1_t (new_AGEMA_signal_2749), .Z1_f (new_AGEMA_signal_2750) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U33 ( .A0_t (StateOut[146]), .A0_f (new_AGEMA_signal_2751), .A1_t (new_AGEMA_signal_2752), .A1_f (new_AGEMA_signal_2753), .B0_t (StateOut[154]), .B0_f (new_AGEMA_signal_2754), .B1_t (new_AGEMA_signal_2755), .B1_f (new_AGEMA_signal_2756), .Z0_t (THETA_n19), .Z0_f (new_AGEMA_signal_2757), .Z1_t (new_AGEMA_signal_2758), .Z1_f (new_AGEMA_signal_2759) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U32 ( .A0_t (StateOut[17]), .A0_f (new_AGEMA_signal_3216), .A1_t (new_AGEMA_signal_3217), .A1_f (new_AGEMA_signal_3218), .B0_t (THETA_n17), .B0_f (new_AGEMA_signal_2973), .B1_t (new_AGEMA_signal_2974), .B1_f (new_AGEMA_signal_2975), .Z0_t (THETA_n114), .Z0_f (new_AGEMA_signal_3219), .Z1_t (new_AGEMA_signal_3220), .Z1_f (new_AGEMA_signal_3221) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U31 ( .A0_t (THETA_n16), .A0_f (new_AGEMA_signal_2775), .A1_t (new_AGEMA_signal_2776), .A1_f (new_AGEMA_signal_2777), .B0_t (THETA_n15), .B0_f (new_AGEMA_signal_2766), .B1_t (new_AGEMA_signal_2767), .B1_f (new_AGEMA_signal_2768), .Z0_t (THETA_n17), .Z0_f (new_AGEMA_signal_2973), .Z1_t (new_AGEMA_signal_2974), .Z1_f (new_AGEMA_signal_2975) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U30 ( .A0_t (StateOut[9]), .A0_f (new_AGEMA_signal_2760), .A1_t (new_AGEMA_signal_2761), .A1_f (new_AGEMA_signal_2762), .B0_t (OutData_s0_t[1]), .B0_f (OutData_s0_f[1]), .B1_t (OutData_s1_t[1]), .B1_f (OutData_s1_f[1]), .Z0_t (THETA_n15), .Z0_f (new_AGEMA_signal_2766), .Z1_t (new_AGEMA_signal_2767), .Z1_f (new_AGEMA_signal_2768) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U29 ( .A0_t (StateOut[25]), .A0_f (new_AGEMA_signal_2769), .A1_t (new_AGEMA_signal_2770), .A1_f (new_AGEMA_signal_2771), .B0_t (StateOut[33]), .B0_f (new_AGEMA_signal_2772), .B1_t (new_AGEMA_signal_2773), .B1_f (new_AGEMA_signal_2774), .Z0_t (THETA_n16), .Z0_f (new_AGEMA_signal_2775), .Z1_t (new_AGEMA_signal_2776), .Z1_f (new_AGEMA_signal_2777) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U28 ( .A0_t (StateOut[156]), .A0_f (new_AGEMA_signal_2373), .A1_t (new_AGEMA_signal_2374), .A1_f (new_AGEMA_signal_2375), .B0_t (THETA_n14), .B0_f (new_AGEMA_signal_3372), .B1_t (new_AGEMA_signal_3373), .B1_f (new_AGEMA_signal_3374), .Z0_t (StateFromRhoPi[188]), .Z0_f (new_AGEMA_signal_3956), .Z1_t (new_AGEMA_signal_3957), .Z1_f (new_AGEMA_signal_3958) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U27 ( .A0_t (StateOut[148]), .A0_f (new_AGEMA_signal_2376), .A1_t (new_AGEMA_signal_2377), .A1_f (new_AGEMA_signal_2378), .B0_t (THETA_n14), .B0_f (new_AGEMA_signal_3372), .B1_t (new_AGEMA_signal_3373), .B1_f (new_AGEMA_signal_3374), .Z0_t (StateFromRhoPi[121]), .Z0_f (new_AGEMA_signal_3959), .Z1_t (new_AGEMA_signal_3960), .Z1_f (new_AGEMA_signal_3961) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U26 ( .A0_t (StateOut[140]), .A0_f (new_AGEMA_signal_2367), .A1_t (new_AGEMA_signal_2368), .A1_f (new_AGEMA_signal_2369), .B0_t (THETA_n14), .B0_f (new_AGEMA_signal_3372), .B1_t (new_AGEMA_signal_3373), .B1_f (new_AGEMA_signal_3374), .Z0_t (StateFromRhoPi[101]), .Z0_f (new_AGEMA_signal_3962), .Z1_t (new_AGEMA_signal_3963), .Z1_f (new_AGEMA_signal_3964) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U25 ( .A0_t (StateOut[132]), .A0_f (new_AGEMA_signal_2364), .A1_t (new_AGEMA_signal_2365), .A1_f (new_AGEMA_signal_2366), .B0_t (THETA_n14), .B0_f (new_AGEMA_signal_3372), .B1_t (new_AGEMA_signal_3373), .B1_f (new_AGEMA_signal_3374), .Z0_t (StateFromRhoPi[75]), .Z0_f (new_AGEMA_signal_3965), .Z1_t (new_AGEMA_signal_3966), .Z1_f (new_AGEMA_signal_3967) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U24 ( .A0_t (StateOut[124]), .A0_f (new_AGEMA_signal_3084), .A1_t (new_AGEMA_signal_3085), .A1_f (new_AGEMA_signal_3086), .B0_t (THETA_n14), .B0_f (new_AGEMA_signal_3372), .B1_t (new_AGEMA_signal_3373), .B1_f (new_AGEMA_signal_3374), .Z0_t (StateFromRhoPi[8]), .Z0_f (new_AGEMA_signal_3968), .Z1_t (new_AGEMA_signal_3969), .Z1_f (new_AGEMA_signal_3970) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U23 ( .A0_t (THETA_n44), .A0_f (new_AGEMA_signal_3231), .A1_t (new_AGEMA_signal_3232), .A1_f (new_AGEMA_signal_3233), .B0_t (THETA_n39), .B0_f (new_AGEMA_signal_3225), .B1_t (new_AGEMA_signal_3226), .B1_f (new_AGEMA_signal_3227), .Z0_t (THETA_n14), .Z0_f (new_AGEMA_signal_3372), .Z1_t (new_AGEMA_signal_3373), .Z1_f (new_AGEMA_signal_3374) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U22 ( .A0_t (StateOut[179]), .A0_f (new_AGEMA_signal_3222), .A1_t (new_AGEMA_signal_3223), .A1_f (new_AGEMA_signal_3224), .B0_t (THETA_n13), .B0_f (new_AGEMA_signal_2976), .B1_t (new_AGEMA_signal_2977), .B1_f (new_AGEMA_signal_2978), .Z0_t (THETA_n39), .Z0_f (new_AGEMA_signal_3225), .Z1_t (new_AGEMA_signal_3226), .Z1_f (new_AGEMA_signal_3227) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U21 ( .A0_t (THETA_n12), .A0_f (new_AGEMA_signal_2793), .A1_t (new_AGEMA_signal_2794), .A1_f (new_AGEMA_signal_2795), .B0_t (THETA_n11), .B0_f (new_AGEMA_signal_2784), .B1_t (new_AGEMA_signal_2785), .B1_f (new_AGEMA_signal_2786), .Z0_t (THETA_n13), .Z0_f (new_AGEMA_signal_2976), .Z1_t (new_AGEMA_signal_2977), .Z1_f (new_AGEMA_signal_2978) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U20 ( .A0_t (StateOut[171]), .A0_f (new_AGEMA_signal_2778), .A1_t (new_AGEMA_signal_2779), .A1_f (new_AGEMA_signal_2780), .B0_t (StateOut[163]), .B0_f (new_AGEMA_signal_2781), .B1_t (new_AGEMA_signal_2782), .B1_f (new_AGEMA_signal_2783), .Z0_t (THETA_n11), .Z0_f (new_AGEMA_signal_2784), .Z1_t (new_AGEMA_signal_2785), .Z1_f (new_AGEMA_signal_2786) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U19 ( .A0_t (StateOut[187]), .A0_f (new_AGEMA_signal_2787), .A1_t (new_AGEMA_signal_2788), .A1_f (new_AGEMA_signal_2789), .B0_t (StateOut[195]), .B0_f (new_AGEMA_signal_2790), .B1_t (new_AGEMA_signal_2791), .B1_f (new_AGEMA_signal_2792), .Z0_t (THETA_n12), .Z0_f (new_AGEMA_signal_2793), .Z1_t (new_AGEMA_signal_2794), .Z1_f (new_AGEMA_signal_2795) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U18 ( .A0_t (StateOut[100]), .A0_f (new_AGEMA_signal_3228), .A1_t (new_AGEMA_signal_3229), .A1_f (new_AGEMA_signal_3230), .B0_t (THETA_n10), .B0_f (new_AGEMA_signal_2979), .B1_t (new_AGEMA_signal_2980), .B1_f (new_AGEMA_signal_2981), .Z0_t (THETA_n44), .Z0_f (new_AGEMA_signal_3231), .Z1_t (new_AGEMA_signal_3232), .Z1_f (new_AGEMA_signal_3233) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U17 ( .A0_t (THETA_n9), .A0_f (new_AGEMA_signal_2811), .A1_t (new_AGEMA_signal_2812), .A1_f (new_AGEMA_signal_2813), .B0_t (THETA_n8), .B0_f (new_AGEMA_signal_2802), .B1_t (new_AGEMA_signal_2803), .B1_f (new_AGEMA_signal_2804), .Z0_t (THETA_n10), .Z0_f (new_AGEMA_signal_2979), .Z1_t (new_AGEMA_signal_2980), .Z1_f (new_AGEMA_signal_2981) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U16 ( .A0_t (StateOut[92]), .A0_f (new_AGEMA_signal_2796), .A1_t (new_AGEMA_signal_2797), .A1_f (new_AGEMA_signal_2798), .B0_t (StateOut[84]), .B0_f (new_AGEMA_signal_2799), .B1_t (new_AGEMA_signal_2800), .B1_f (new_AGEMA_signal_2801), .Z0_t (THETA_n8), .Z0_f (new_AGEMA_signal_2802), .Z1_t (new_AGEMA_signal_2803), .Z1_f (new_AGEMA_signal_2804) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U15 ( .A0_t (StateOut[108]), .A0_f (new_AGEMA_signal_2805), .A1_t (new_AGEMA_signal_2806), .A1_f (new_AGEMA_signal_2807), .B0_t (StateOut[116]), .B0_f (new_AGEMA_signal_2808), .B1_t (new_AGEMA_signal_2809), .B1_f (new_AGEMA_signal_2810), .Z0_t (THETA_n9), .Z0_f (new_AGEMA_signal_2811), .Z1_t (new_AGEMA_signal_2812), .Z1_f (new_AGEMA_signal_2813) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U14 ( .A0_t (StateOut[155]), .A0_f (new_AGEMA_signal_2589), .A1_t (new_AGEMA_signal_2590), .A1_f (new_AGEMA_signal_2591), .B0_t (THETA_n7), .B0_f (new_AGEMA_signal_3375), .B1_t (new_AGEMA_signal_3376), .B1_f (new_AGEMA_signal_3377), .Z0_t (StateFromRhoPi[187]), .Z0_f (new_AGEMA_signal_3971), .Z1_t (new_AGEMA_signal_3972), .Z1_f (new_AGEMA_signal_3973) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U13 ( .A0_t (StateOut[147]), .A0_f (new_AGEMA_signal_2592), .A1_t (new_AGEMA_signal_2593), .A1_f (new_AGEMA_signal_2594), .B0_t (THETA_n7), .B0_f (new_AGEMA_signal_3375), .B1_t (new_AGEMA_signal_3376), .B1_f (new_AGEMA_signal_3377), .Z0_t (StateFromRhoPi[120]), .Z0_f (new_AGEMA_signal_3974), .Z1_t (new_AGEMA_signal_3975), .Z1_f (new_AGEMA_signal_3976) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U12 ( .A0_t (StateOut[139]), .A0_f (new_AGEMA_signal_2583), .A1_t (new_AGEMA_signal_2584), .A1_f (new_AGEMA_signal_2585), .B0_t (THETA_n7), .B0_f (new_AGEMA_signal_3375), .B1_t (new_AGEMA_signal_3376), .B1_f (new_AGEMA_signal_3377), .Z0_t (StateFromRhoPi[100]), .Z0_f (new_AGEMA_signal_3977), .Z1_t (new_AGEMA_signal_3978), .Z1_f (new_AGEMA_signal_3979) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U11 ( .A0_t (StateOut[131]), .A0_f (new_AGEMA_signal_2580), .A1_t (new_AGEMA_signal_2581), .A1_f (new_AGEMA_signal_2582), .B0_t (THETA_n7), .B0_f (new_AGEMA_signal_3375), .B1_t (new_AGEMA_signal_3376), .B1_f (new_AGEMA_signal_3377), .Z0_t (StateFromRhoPi[74]), .Z0_f (new_AGEMA_signal_3980), .Z1_t (new_AGEMA_signal_3981), .Z1_f (new_AGEMA_signal_3982) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U10 ( .A0_t (StateOut[123]), .A0_f (new_AGEMA_signal_3156), .A1_t (new_AGEMA_signal_3157), .A1_f (new_AGEMA_signal_3158), .B0_t (THETA_n7), .B0_f (new_AGEMA_signal_3375), .B1_t (new_AGEMA_signal_3376), .B1_f (new_AGEMA_signal_3377), .Z0_t (StateFromRhoPi[15]), .Z0_f (new_AGEMA_signal_3983), .Z1_t (new_AGEMA_signal_3984), .Z1_f (new_AGEMA_signal_3985) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U9 ( .A0_t (THETA_n104), .A0_f (new_AGEMA_signal_3243), .A1_t (new_AGEMA_signal_3244), .A1_f (new_AGEMA_signal_3245), .B0_t (THETA_n67), .B0_f (new_AGEMA_signal_3237), .B1_t (new_AGEMA_signal_3238), .B1_f (new_AGEMA_signal_3239), .Z0_t (THETA_n7), .Z0_f (new_AGEMA_signal_3375), .Z1_t (new_AGEMA_signal_3376), .Z1_f (new_AGEMA_signal_3377) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U8 ( .A0_t (StateOut[107]), .A0_f (new_AGEMA_signal_3234), .A1_t (new_AGEMA_signal_3235), .A1_f (new_AGEMA_signal_3236), .B0_t (THETA_n6), .B0_f (new_AGEMA_signal_2982), .B1_t (new_AGEMA_signal_2983), .B1_f (new_AGEMA_signal_2984), .Z0_t (THETA_n67), .Z0_f (new_AGEMA_signal_3237), .Z1_t (new_AGEMA_signal_3238), .Z1_f (new_AGEMA_signal_3239) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U7 ( .A0_t (THETA_n5), .A0_f (new_AGEMA_signal_2829), .A1_t (new_AGEMA_signal_2830), .A1_f (new_AGEMA_signal_2831), .B0_t (THETA_n4), .B0_f (new_AGEMA_signal_2820), .B1_t (new_AGEMA_signal_2821), .B1_f (new_AGEMA_signal_2822), .Z0_t (THETA_n6), .Z0_f (new_AGEMA_signal_2982), .Z1_t (new_AGEMA_signal_2983), .Z1_f (new_AGEMA_signal_2984) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U6 ( .A0_t (StateOut[91]), .A0_f (new_AGEMA_signal_2814), .A1_t (new_AGEMA_signal_2815), .A1_f (new_AGEMA_signal_2816), .B0_t (StateOut[83]), .B0_f (new_AGEMA_signal_2817), .B1_t (new_AGEMA_signal_2818), .B1_f (new_AGEMA_signal_2819), .Z0_t (THETA_n4), .Z0_f (new_AGEMA_signal_2820), .Z1_t (new_AGEMA_signal_2821), .Z1_f (new_AGEMA_signal_2822) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U5 ( .A0_t (StateOut[115]), .A0_f (new_AGEMA_signal_2823), .A1_t (new_AGEMA_signal_2824), .A1_f (new_AGEMA_signal_2825), .B0_t (StateOut[99]), .B0_f (new_AGEMA_signal_2826), .B1_t (new_AGEMA_signal_2827), .B1_f (new_AGEMA_signal_2828), .Z0_t (THETA_n5), .Z0_f (new_AGEMA_signal_2829), .Z1_t (new_AGEMA_signal_2830), .Z1_f (new_AGEMA_signal_2831) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U4 ( .A0_t (StateOut[186]), .A0_f (new_AGEMA_signal_3240), .A1_t (new_AGEMA_signal_3241), .A1_f (new_AGEMA_signal_3242), .B0_t (THETA_n3), .B0_f (new_AGEMA_signal_2985), .B1_t (new_AGEMA_signal_2986), .B1_f (new_AGEMA_signal_2987), .Z0_t (THETA_n104), .Z0_f (new_AGEMA_signal_3243), .Z1_t (new_AGEMA_signal_3244), .Z1_f (new_AGEMA_signal_3245) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U3 ( .A0_t (THETA_n2), .A0_f (new_AGEMA_signal_2847), .A1_t (new_AGEMA_signal_2848), .A1_f (new_AGEMA_signal_2849), .B0_t (THETA_n1), .B0_f (new_AGEMA_signal_2838), .B1_t (new_AGEMA_signal_2839), .B1_f (new_AGEMA_signal_2840), .Z0_t (THETA_n3), .Z0_f (new_AGEMA_signal_2985), .Z1_t (new_AGEMA_signal_2986), .Z1_f (new_AGEMA_signal_2987) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U2 ( .A0_t (StateOut[170]), .A0_f (new_AGEMA_signal_2832), .A1_t (new_AGEMA_signal_2833), .A1_f (new_AGEMA_signal_2834), .B0_t (StateOut[162]), .B0_f (new_AGEMA_signal_2835), .B1_t (new_AGEMA_signal_2836), .B1_f (new_AGEMA_signal_2837), .Z0_t (THETA_n1), .Z0_f (new_AGEMA_signal_2838), .Z1_t (new_AGEMA_signal_2839), .Z1_f (new_AGEMA_signal_2840) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U1 ( .A0_t (StateOut[194]), .A0_f (new_AGEMA_signal_2841), .A1_t (new_AGEMA_signal_2842), .A1_f (new_AGEMA_signal_2843), .B0_t (StateOut[178]), .B0_f (new_AGEMA_signal_2844), .B1_t (new_AGEMA_signal_2845), .B1_f (new_AGEMA_signal_2846), .Z0_t (THETA_n2), .Z0_f (new_AGEMA_signal_2847), .Z1_t (new_AGEMA_signal_2848), .Z1_f (new_AGEMA_signal_2849) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_U4 ( .A0_t (CHI_ChiOut[0]), .A0_f (new_AGEMA_signal_4599), .A1_t (new_AGEMA_signal_4600), .A1_f (new_AGEMA_signal_4601), .B0_t (1'b0), .B0_f (1'b1), .B1_t (IotaRC[0]), .B1_f (new_AGEMA_signal_3990), .Z0_t (StateFromChi[0]), .Z0_f (new_AGEMA_signal_5201), .Z1_t (new_AGEMA_signal_5202), .Z1_f (new_AGEMA_signal_5203) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_U3 ( .A0_t (CHI_ChiOut[1]), .A0_f (new_AGEMA_signal_4674), .A1_t (new_AGEMA_signal_4675), .A1_f (new_AGEMA_signal_4676), .B0_t (1'b0), .B0_f (1'b1), .B1_t (IotaRC[1]), .B1_f (new_AGEMA_signal_6421), .Z0_t (StateFromChi[1]), .Z0_f (new_AGEMA_signal_6431), .Z1_t (new_AGEMA_signal_6432), .Z1_f (new_AGEMA_signal_6433) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_U2 ( .A0_t (CHI_ChiOut_7), .A0_f (new_AGEMA_signal_5124), .A1_t (new_AGEMA_signal_5125), .A1_f (new_AGEMA_signal_5126), .B0_t (1'b0), .B0_f (1'b1), .B1_t (IotaRC_7), .B1_f (new_AGEMA_signal_5199), .Z0_t (StateFromChi[7]), .Z0_f (new_AGEMA_signal_5204), .Z1_t (new_AGEMA_signal_5205), .Z1_f (new_AGEMA_signal_5206) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_U1 ( .A0_t (CHI_ChiOut_3), .A0_f (new_AGEMA_signal_4824), .A1_t (new_AGEMA_signal_4825), .A1_f (new_AGEMA_signal_4826), .B0_t (1'b0), .B0_f (1'b1), .B1_t (IotaRC_3), .B1_f (new_AGEMA_signal_4596), .Z0_t (StateFromChi[3]), .Z0_f (new_AGEMA_signal_5207), .Z1_t (new_AGEMA_signal_5208), .Z1_f (new_AGEMA_signal_5209) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[40]), .A0_f (new_AGEMA_signal_3815), .A1_t (new_AGEMA_signal_3816), .A1_f (new_AGEMA_signal_3817), .B0_t (StateFromRhoPi[80]), .B0_f (new_AGEMA_signal_3647), .B1_t (new_AGEMA_signal_3648), .B1_f (new_AGEMA_signal_3649), .Z0_t (CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_and_xor_inst_a_nxy), .Z0_f (new_AGEMA_signal_3993), .Z1_t (new_AGEMA_signal_3994), .Z1_f (new_AGEMA_signal_3995) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_and_xor_inst_a_nxy), .A0_f (new_AGEMA_signal_3993), .A1_t (new_AGEMA_signal_3994), .A1_f (new_AGEMA_signal_3995), .B0_t (StateFromRhoPi[0]), .B0_f (new_AGEMA_signal_3608), .B1_t (new_AGEMA_signal_3609), .B1_f (new_AGEMA_signal_3610), .Z0_t (CHI_ChiOut[0]), .Z0_f (new_AGEMA_signal_4599), .Z1_t (new_AGEMA_signal_4600), .Z1_f (new_AGEMA_signal_4601) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[80]), .A0_f (new_AGEMA_signal_3647), .A1_t (new_AGEMA_signal_3648), .A1_f (new_AGEMA_signal_3649), .B0_t (StateFromRhoPi[120]), .B0_f (new_AGEMA_signal_3974), .B1_t (new_AGEMA_signal_3975), .B1_f (new_AGEMA_signal_3976), .Z0_t (CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_and_xor_inst_b_nxy), .Z0_f (new_AGEMA_signal_3996), .Z1_t (new_AGEMA_signal_3997), .Z1_f (new_AGEMA_signal_3998) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_and_xor_inst_b_nxy), .A0_f (new_AGEMA_signal_3996), .A1_t (new_AGEMA_signal_3997), .A1_f (new_AGEMA_signal_3998), .B0_t (StateFromRhoPi[40]), .B0_f (new_AGEMA_signal_3815), .B1_t (new_AGEMA_signal_3816), .B1_f (new_AGEMA_signal_3817), .Z0_t (StateFromChi[40]), .Z0_f (new_AGEMA_signal_4602), .Z1_t (new_AGEMA_signal_4603), .Z1_f (new_AGEMA_signal_4604) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[120]), .A0_f (new_AGEMA_signal_3974), .A1_t (new_AGEMA_signal_3975), .A1_f (new_AGEMA_signal_3976), .B0_t (StateFromRhoPi[160]), .B0_f (new_AGEMA_signal_3941), .B1_t (new_AGEMA_signal_3942), .B1_f (new_AGEMA_signal_3943), .Z0_t (CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_and_xor_inst_c_nxy), .Z0_f (new_AGEMA_signal_3999), .Z1_t (new_AGEMA_signal_4000), .Z1_f (new_AGEMA_signal_4001) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_and_xor_inst_c_nxy), .A0_f (new_AGEMA_signal_3999), .A1_t (new_AGEMA_signal_4000), .A1_f (new_AGEMA_signal_4001), .B0_t (StateFromRhoPi[80]), .B0_f (new_AGEMA_signal_3647), .B1_t (new_AGEMA_signal_3648), .B1_f (new_AGEMA_signal_3649), .Z0_t (StateFromChi[80]), .Z0_f (new_AGEMA_signal_4605), .Z1_t (new_AGEMA_signal_4606), .Z1_f (new_AGEMA_signal_4607) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[160]), .A0_f (new_AGEMA_signal_3941), .A1_t (new_AGEMA_signal_3942), .A1_f (new_AGEMA_signal_3943), .B0_t (StateFromRhoPi[0]), .B0_f (new_AGEMA_signal_3608), .B1_t (new_AGEMA_signal_3609), .B1_f (new_AGEMA_signal_3610), .Z0_t (CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_and_xor_inst_d_nxy), .Z0_f (new_AGEMA_signal_4002), .Z1_t (new_AGEMA_signal_4003), .Z1_f (new_AGEMA_signal_4004) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_and_xor_inst_d_nxy), .A0_f (new_AGEMA_signal_4002), .A1_t (new_AGEMA_signal_4003), .A1_f (new_AGEMA_signal_4004), .B0_t (StateFromRhoPi[120]), .B0_f (new_AGEMA_signal_3974), .B1_t (new_AGEMA_signal_3975), .B1_f (new_AGEMA_signal_3976), .Z0_t (StateFromChi[120]), .Z0_f (new_AGEMA_signal_4608), .Z1_t (new_AGEMA_signal_4609), .Z1_f (new_AGEMA_signal_4610) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[0]), .A0_f (new_AGEMA_signal_3608), .A1_t (new_AGEMA_signal_3609), .A1_f (new_AGEMA_signal_3610), .B0_t (StateFromRhoPi[40]), .B0_f (new_AGEMA_signal_3815), .B1_t (new_AGEMA_signal_3816), .B1_f (new_AGEMA_signal_3817), .Z0_t (CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_and_xor_inst_e_nxy), .Z0_f (new_AGEMA_signal_4005), .Z1_t (new_AGEMA_signal_4006), .Z1_f (new_AGEMA_signal_4007) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_and_xor_inst_e_nxy), .A0_f (new_AGEMA_signal_4005), .A1_t (new_AGEMA_signal_4006), .A1_f (new_AGEMA_signal_4007), .B0_t (StateFromRhoPi[160]), .B0_f (new_AGEMA_signal_3941), .B1_t (new_AGEMA_signal_3942), .B1_f (new_AGEMA_signal_3943), .Z0_t (StateFromChi[160]), .Z0_f (new_AGEMA_signal_4611), .Z1_t (new_AGEMA_signal_4612), .Z1_f (new_AGEMA_signal_4613) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[48]), .A0_f (new_AGEMA_signal_3470), .A1_t (new_AGEMA_signal_3471), .A1_f (new_AGEMA_signal_3472), .B0_t (StateFromRhoPi[88]), .B0_f (new_AGEMA_signal_3842), .B1_t (new_AGEMA_signal_3843), .B1_f (new_AGEMA_signal_3844), .Z0_t (CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_and_xor_inst_a_nxy), .Z0_f (new_AGEMA_signal_4008), .Z1_t (new_AGEMA_signal_4009), .Z1_f (new_AGEMA_signal_4010) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_and_xor_inst_a_nxy), .A0_f (new_AGEMA_signal_4008), .A1_t (new_AGEMA_signal_4009), .A1_f (new_AGEMA_signal_4010), .B0_t (StateFromRhoPi[8]), .B0_f (new_AGEMA_signal_3968), .B1_t (new_AGEMA_signal_3969), .B1_f (new_AGEMA_signal_3970), .Z0_t (StateFromChi[8]), .Z0_f (new_AGEMA_signal_4614), .Z1_t (new_AGEMA_signal_4615), .Z1_f (new_AGEMA_signal_4616) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[88]), .A0_f (new_AGEMA_signal_3842), .A1_t (new_AGEMA_signal_3843), .A1_f (new_AGEMA_signal_3844), .B0_t (StateFromRhoPi[128]), .B0_f (new_AGEMA_signal_3479), .B1_t (new_AGEMA_signal_3480), .B1_f (new_AGEMA_signal_3481), .Z0_t (CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_and_xor_inst_b_nxy), .Z0_f (new_AGEMA_signal_4011), .Z1_t (new_AGEMA_signal_4012), .Z1_f (new_AGEMA_signal_4013) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_and_xor_inst_b_nxy), .A0_f (new_AGEMA_signal_4011), .A1_t (new_AGEMA_signal_4012), .A1_f (new_AGEMA_signal_4013), .B0_t (StateFromRhoPi[48]), .B0_f (new_AGEMA_signal_3470), .B1_t (new_AGEMA_signal_3471), .B1_f (new_AGEMA_signal_3472), .Z0_t (StateFromChi[48]), .Z0_f (new_AGEMA_signal_4617), .Z1_t (new_AGEMA_signal_4618), .Z1_f (new_AGEMA_signal_4619) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[128]), .A0_f (new_AGEMA_signal_3479), .A1_t (new_AGEMA_signal_3480), .A1_f (new_AGEMA_signal_3481), .B0_t (StateFromRhoPi[168]), .B0_f (new_AGEMA_signal_3851), .B1_t (new_AGEMA_signal_3852), .B1_f (new_AGEMA_signal_3853), .Z0_t (CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_and_xor_inst_c_nxy), .Z0_f (new_AGEMA_signal_4014), .Z1_t (new_AGEMA_signal_4015), .Z1_f (new_AGEMA_signal_4016) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_and_xor_inst_c_nxy), .A0_f (new_AGEMA_signal_4014), .A1_t (new_AGEMA_signal_4015), .A1_f (new_AGEMA_signal_4016), .B0_t (StateFromRhoPi[88]), .B0_f (new_AGEMA_signal_3842), .B1_t (new_AGEMA_signal_3843), .B1_f (new_AGEMA_signal_3844), .Z0_t (StateFromChi[88]), .Z0_f (new_AGEMA_signal_4620), .Z1_t (new_AGEMA_signal_4621), .Z1_f (new_AGEMA_signal_4622) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[168]), .A0_f (new_AGEMA_signal_3851), .A1_t (new_AGEMA_signal_3852), .A1_f (new_AGEMA_signal_3853), .B0_t (StateFromRhoPi[8]), .B0_f (new_AGEMA_signal_3968), .B1_t (new_AGEMA_signal_3969), .B1_f (new_AGEMA_signal_3970), .Z0_t (CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_and_xor_inst_d_nxy), .Z0_f (new_AGEMA_signal_4017), .Z1_t (new_AGEMA_signal_4018), .Z1_f (new_AGEMA_signal_4019) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_and_xor_inst_d_nxy), .A0_f (new_AGEMA_signal_4017), .A1_t (new_AGEMA_signal_4018), .A1_f (new_AGEMA_signal_4019), .B0_t (StateFromRhoPi[128]), .B0_f (new_AGEMA_signal_3479), .B1_t (new_AGEMA_signal_3480), .B1_f (new_AGEMA_signal_3481), .Z0_t (StateFromChi[128]), .Z0_f (new_AGEMA_signal_4623), .Z1_t (new_AGEMA_signal_4624), .Z1_f (new_AGEMA_signal_4625) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[8]), .A0_f (new_AGEMA_signal_3968), .A1_t (new_AGEMA_signal_3969), .A1_f (new_AGEMA_signal_3970), .B0_t (StateFromRhoPi[48]), .B0_f (new_AGEMA_signal_3470), .B1_t (new_AGEMA_signal_3471), .B1_f (new_AGEMA_signal_3472), .Z0_t (CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_and_xor_inst_e_nxy), .Z0_f (new_AGEMA_signal_4020), .Z1_t (new_AGEMA_signal_4021), .Z1_f (new_AGEMA_signal_4022) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_and_xor_inst_e_nxy), .A0_f (new_AGEMA_signal_4020), .A1_t (new_AGEMA_signal_4021), .A1_f (new_AGEMA_signal_4022), .B0_t (StateFromRhoPi[168]), .B0_f (new_AGEMA_signal_3851), .B1_t (new_AGEMA_signal_3852), .B1_f (new_AGEMA_signal_3853), .Z0_t (StateFromChi[168]), .Z0_f (new_AGEMA_signal_4626), .Z1_t (new_AGEMA_signal_4627), .Z1_f (new_AGEMA_signal_4628) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[56]), .A0_f (new_AGEMA_signal_3560), .A1_t (new_AGEMA_signal_3561), .A1_f (new_AGEMA_signal_3562), .B0_t (StateFromRhoPi[96]), .B0_f (new_AGEMA_signal_3752), .B1_t (new_AGEMA_signal_3753), .B1_f (new_AGEMA_signal_3754), .Z0_t (CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_and_xor_inst_a_nxy), .Z0_f (new_AGEMA_signal_4023), .Z1_t (new_AGEMA_signal_4024), .Z1_f (new_AGEMA_signal_4025) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_and_xor_inst_a_nxy), .A0_f (new_AGEMA_signal_4023), .A1_t (new_AGEMA_signal_4024), .A1_f (new_AGEMA_signal_4025), .B0_t (StateFromRhoPi[16]), .B0_f (new_AGEMA_signal_3638), .B1_t (new_AGEMA_signal_3639), .B1_f (new_AGEMA_signal_3640), .Z0_t (StateFromChi[16]), .Z0_f (new_AGEMA_signal_4629), .Z1_t (new_AGEMA_signal_4630), .Z1_f (new_AGEMA_signal_4631) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[96]), .A0_f (new_AGEMA_signal_3752), .A1_t (new_AGEMA_signal_3753), .A1_f (new_AGEMA_signal_3754), .B0_t (StateFromRhoPi[136]), .B0_f (new_AGEMA_signal_3614), .B1_t (new_AGEMA_signal_3615), .B1_f (new_AGEMA_signal_3616), .Z0_t (CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_and_xor_inst_b_nxy), .Z0_f (new_AGEMA_signal_4026), .Z1_t (new_AGEMA_signal_4027), .Z1_f (new_AGEMA_signal_4028) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_and_xor_inst_b_nxy), .A0_f (new_AGEMA_signal_4026), .A1_t (new_AGEMA_signal_4027), .A1_f (new_AGEMA_signal_4028), .B0_t (StateFromRhoPi[56]), .B0_f (new_AGEMA_signal_3560), .B1_t (new_AGEMA_signal_3561), .B1_f (new_AGEMA_signal_3562), .Z0_t (StateFromChi[56]), .Z0_f (new_AGEMA_signal_4632), .Z1_t (new_AGEMA_signal_4633), .Z1_f (new_AGEMA_signal_4634) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[136]), .A0_f (new_AGEMA_signal_3614), .A1_t (new_AGEMA_signal_3615), .A1_f (new_AGEMA_signal_3616), .B0_t (StateFromRhoPi[176]), .B0_f (new_AGEMA_signal_3761), .B1_t (new_AGEMA_signal_3762), .B1_f (new_AGEMA_signal_3763), .Z0_t (CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_and_xor_inst_c_nxy), .Z0_f (new_AGEMA_signal_4029), .Z1_t (new_AGEMA_signal_4030), .Z1_f (new_AGEMA_signal_4031) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_and_xor_inst_c_nxy), .A0_f (new_AGEMA_signal_4029), .A1_t (new_AGEMA_signal_4030), .A1_f (new_AGEMA_signal_4031), .B0_t (StateFromRhoPi[96]), .B0_f (new_AGEMA_signal_3752), .B1_t (new_AGEMA_signal_3753), .B1_f (new_AGEMA_signal_3754), .Z0_t (StateFromChi[96]), .Z0_f (new_AGEMA_signal_4635), .Z1_t (new_AGEMA_signal_4636), .Z1_f (new_AGEMA_signal_4637) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[176]), .A0_f (new_AGEMA_signal_3761), .A1_t (new_AGEMA_signal_3762), .A1_f (new_AGEMA_signal_3763), .B0_t (StateFromRhoPi[16]), .B0_f (new_AGEMA_signal_3638), .B1_t (new_AGEMA_signal_3639), .B1_f (new_AGEMA_signal_3640), .Z0_t (CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_and_xor_inst_d_nxy), .Z0_f (new_AGEMA_signal_4032), .Z1_t (new_AGEMA_signal_4033), .Z1_f (new_AGEMA_signal_4034) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_and_xor_inst_d_nxy), .A0_f (new_AGEMA_signal_4032), .A1_t (new_AGEMA_signal_4033), .A1_f (new_AGEMA_signal_4034), .B0_t (StateFromRhoPi[136]), .B0_f (new_AGEMA_signal_3614), .B1_t (new_AGEMA_signal_3615), .B1_f (new_AGEMA_signal_3616), .Z0_t (StateFromChi[136]), .Z0_f (new_AGEMA_signal_4638), .Z1_t (new_AGEMA_signal_4639), .Z1_f (new_AGEMA_signal_4640) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[16]), .A0_f (new_AGEMA_signal_3638), .A1_t (new_AGEMA_signal_3639), .A1_f (new_AGEMA_signal_3640), .B0_t (StateFromRhoPi[56]), .B0_f (new_AGEMA_signal_3560), .B1_t (new_AGEMA_signal_3561), .B1_f (new_AGEMA_signal_3562), .Z0_t (CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_and_xor_inst_e_nxy), .Z0_f (new_AGEMA_signal_4035), .Z1_t (new_AGEMA_signal_4036), .Z1_f (new_AGEMA_signal_4037) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_and_xor_inst_e_nxy), .A0_f (new_AGEMA_signal_4035), .A1_t (new_AGEMA_signal_4036), .A1_f (new_AGEMA_signal_4037), .B0_t (StateFromRhoPi[176]), .B0_f (new_AGEMA_signal_3761), .B1_t (new_AGEMA_signal_3762), .B1_f (new_AGEMA_signal_3763), .Z0_t (StateFromChi[176]), .Z0_f (new_AGEMA_signal_4641), .Z1_t (new_AGEMA_signal_4642), .Z1_f (new_AGEMA_signal_4643) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[64]), .A0_f (new_AGEMA_signal_3875), .A1_t (new_AGEMA_signal_3876), .A1_f (new_AGEMA_signal_3877), .B0_t (StateFromRhoPi[104]), .B0_f (new_AGEMA_signal_3407), .B1_t (new_AGEMA_signal_3408), .B1_f (new_AGEMA_signal_3409), .Z0_t (CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_and_xor_inst_a_nxy), .Z0_f (new_AGEMA_signal_4038), .Z1_t (new_AGEMA_signal_4039), .Z1_f (new_AGEMA_signal_4040) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_and_xor_inst_a_nxy), .A0_f (new_AGEMA_signal_4038), .A1_t (new_AGEMA_signal_4039), .A1_f (new_AGEMA_signal_4040), .B0_t (StateFromRhoPi[24]), .B0_f (new_AGEMA_signal_3803), .B1_t (new_AGEMA_signal_3804), .B1_f (new_AGEMA_signal_3805), .Z0_t (StateFromChi[24]), .Z0_f (new_AGEMA_signal_4644), .Z1_t (new_AGEMA_signal_4645), .Z1_f (new_AGEMA_signal_4646) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[104]), .A0_f (new_AGEMA_signal_3407), .A1_t (new_AGEMA_signal_3408), .A1_f (new_AGEMA_signal_3409), .B0_t (StateFromRhoPi[144]), .B0_f (new_AGEMA_signal_3689), .B1_t (new_AGEMA_signal_3690), .B1_f (new_AGEMA_signal_3691), .Z0_t (CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_and_xor_inst_b_nxy), .Z0_f (new_AGEMA_signal_4041), .Z1_t (new_AGEMA_signal_4042), .Z1_f (new_AGEMA_signal_4043) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_and_xor_inst_b_nxy), .A0_f (new_AGEMA_signal_4041), .A1_t (new_AGEMA_signal_4042), .A1_f (new_AGEMA_signal_4043), .B0_t (StateFromRhoPi[64]), .B0_f (new_AGEMA_signal_3875), .B1_t (new_AGEMA_signal_3876), .B1_f (new_AGEMA_signal_3877), .Z0_t (StateFromChi[64]), .Z0_f (new_AGEMA_signal_4647), .Z1_t (new_AGEMA_signal_4648), .Z1_f (new_AGEMA_signal_4649) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[144]), .A0_f (new_AGEMA_signal_3689), .A1_t (new_AGEMA_signal_3690), .A1_f (new_AGEMA_signal_3691), .B0_t (StateFromRhoPi[184]), .B0_f (new_AGEMA_signal_3656), .B1_t (new_AGEMA_signal_3657), .B1_f (new_AGEMA_signal_3658), .Z0_t (CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_and_xor_inst_c_nxy), .Z0_f (new_AGEMA_signal_4044), .Z1_t (new_AGEMA_signal_4045), .Z1_f (new_AGEMA_signal_4046) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_and_xor_inst_c_nxy), .A0_f (new_AGEMA_signal_4044), .A1_t (new_AGEMA_signal_4045), .A1_f (new_AGEMA_signal_4046), .B0_t (StateFromRhoPi[104]), .B0_f (new_AGEMA_signal_3407), .B1_t (new_AGEMA_signal_3408), .B1_f (new_AGEMA_signal_3409), .Z0_t (StateFromChi[104]), .Z0_f (new_AGEMA_signal_4650), .Z1_t (new_AGEMA_signal_4651), .Z1_f (new_AGEMA_signal_4652) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[184]), .A0_f (new_AGEMA_signal_3656), .A1_t (new_AGEMA_signal_3657), .A1_f (new_AGEMA_signal_3658), .B0_t (StateFromRhoPi[24]), .B0_f (new_AGEMA_signal_3803), .B1_t (new_AGEMA_signal_3804), .B1_f (new_AGEMA_signal_3805), .Z0_t (CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_and_xor_inst_d_nxy), .Z0_f (new_AGEMA_signal_4047), .Z1_t (new_AGEMA_signal_4048), .Z1_f (new_AGEMA_signal_4049) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_and_xor_inst_d_nxy), .A0_f (new_AGEMA_signal_4047), .A1_t (new_AGEMA_signal_4048), .A1_f (new_AGEMA_signal_4049), .B0_t (StateFromRhoPi[144]), .B0_f (new_AGEMA_signal_3689), .B1_t (new_AGEMA_signal_3690), .B1_f (new_AGEMA_signal_3691), .Z0_t (StateFromChi[144]), .Z0_f (new_AGEMA_signal_4653), .Z1_t (new_AGEMA_signal_4654), .Z1_f (new_AGEMA_signal_4655) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[24]), .A0_f (new_AGEMA_signal_3803), .A1_t (new_AGEMA_signal_3804), .A1_f (new_AGEMA_signal_3805), .B0_t (StateFromRhoPi[64]), .B0_f (new_AGEMA_signal_3875), .B1_t (new_AGEMA_signal_3876), .B1_f (new_AGEMA_signal_3877), .Z0_t (CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_and_xor_inst_e_nxy), .Z0_f (new_AGEMA_signal_4050), .Z1_t (new_AGEMA_signal_4051), .Z1_f (new_AGEMA_signal_4052) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_and_xor_inst_e_nxy), .A0_f (new_AGEMA_signal_4050), .A1_t (new_AGEMA_signal_4051), .A1_f (new_AGEMA_signal_4052), .B0_t (StateFromRhoPi[184]), .B0_f (new_AGEMA_signal_3656), .B1_t (new_AGEMA_signal_3657), .B1_f (new_AGEMA_signal_3658), .Z0_t (StateFromChi[184]), .Z0_f (new_AGEMA_signal_4656), .Z1_t (new_AGEMA_signal_4657), .Z1_f (new_AGEMA_signal_4658) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[72]), .A0_f (new_AGEMA_signal_3575), .A1_t (new_AGEMA_signal_3576), .A1_f (new_AGEMA_signal_3577), .B0_t (StateFromRhoPi[112]), .B0_f (new_AGEMA_signal_3497), .B1_t (new_AGEMA_signal_3498), .B1_f (new_AGEMA_signal_3499), .Z0_t (CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_and_xor_inst_a_nxy), .Z0_f (new_AGEMA_signal_4053), .Z1_t (new_AGEMA_signal_4054), .Z1_f (new_AGEMA_signal_4055) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_and_xor_inst_a_nxy), .A0_f (new_AGEMA_signal_4053), .A1_t (new_AGEMA_signal_4054), .A1_f (new_AGEMA_signal_4055), .B0_t (StateFromRhoPi[32]), .B0_f (new_AGEMA_signal_3563), .B1_t (new_AGEMA_signal_3564), .B1_f (new_AGEMA_signal_3565), .Z0_t (StateFromChi[32]), .Z0_f (new_AGEMA_signal_4659), .Z1_t (new_AGEMA_signal_4660), .Z1_f (new_AGEMA_signal_4661) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[112]), .A0_f (new_AGEMA_signal_3497), .A1_t (new_AGEMA_signal_3498), .A1_f (new_AGEMA_signal_3499), .B0_t (StateFromRhoPi[152]), .B0_f (new_AGEMA_signal_3719), .B1_t (new_AGEMA_signal_3720), .B1_f (new_AGEMA_signal_3721), .Z0_t (CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_and_xor_inst_b_nxy), .Z0_f (new_AGEMA_signal_4056), .Z1_t (new_AGEMA_signal_4057), .Z1_f (new_AGEMA_signal_4058) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_and_xor_inst_b_nxy), .A0_f (new_AGEMA_signal_4056), .A1_t (new_AGEMA_signal_4057), .A1_f (new_AGEMA_signal_4058), .B0_t (StateFromRhoPi[72]), .B0_f (new_AGEMA_signal_3575), .B1_t (new_AGEMA_signal_3576), .B1_f (new_AGEMA_signal_3577), .Z0_t (StateFromChi[72]), .Z0_f (new_AGEMA_signal_4662), .Z1_t (new_AGEMA_signal_4663), .Z1_f (new_AGEMA_signal_4664) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[152]), .A0_f (new_AGEMA_signal_3719), .A1_t (new_AGEMA_signal_3720), .A1_f (new_AGEMA_signal_3721), .B0_t (StateFromRhoPi[192]), .B0_f (new_AGEMA_signal_3401), .B1_t (new_AGEMA_signal_3402), .B1_f (new_AGEMA_signal_3403), .Z0_t (CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_and_xor_inst_c_nxy), .Z0_f (new_AGEMA_signal_4059), .Z1_t (new_AGEMA_signal_4060), .Z1_f (new_AGEMA_signal_4061) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_and_xor_inst_c_nxy), .A0_f (new_AGEMA_signal_4059), .A1_t (new_AGEMA_signal_4060), .A1_f (new_AGEMA_signal_4061), .B0_t (StateFromRhoPi[112]), .B0_f (new_AGEMA_signal_3497), .B1_t (new_AGEMA_signal_3498), .B1_f (new_AGEMA_signal_3499), .Z0_t (StateFromChi[112]), .Z0_f (new_AGEMA_signal_4665), .Z1_t (new_AGEMA_signal_4666), .Z1_f (new_AGEMA_signal_4667) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[192]), .A0_f (new_AGEMA_signal_3401), .A1_t (new_AGEMA_signal_3402), .A1_f (new_AGEMA_signal_3403), .B0_t (StateFromRhoPi[32]), .B0_f (new_AGEMA_signal_3563), .B1_t (new_AGEMA_signal_3564), .B1_f (new_AGEMA_signal_3565), .Z0_t (CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_and_xor_inst_d_nxy), .Z0_f (new_AGEMA_signal_4062), .Z1_t (new_AGEMA_signal_4063), .Z1_f (new_AGEMA_signal_4064) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_and_xor_inst_d_nxy), .A0_f (new_AGEMA_signal_4062), .A1_t (new_AGEMA_signal_4063), .A1_f (new_AGEMA_signal_4064), .B0_t (StateFromRhoPi[152]), .B0_f (new_AGEMA_signal_3719), .B1_t (new_AGEMA_signal_3720), .B1_f (new_AGEMA_signal_3721), .Z0_t (StateFromChi[152]), .Z0_f (new_AGEMA_signal_4668), .Z1_t (new_AGEMA_signal_4669), .Z1_f (new_AGEMA_signal_4670) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[32]), .A0_f (new_AGEMA_signal_3563), .A1_t (new_AGEMA_signal_3564), .A1_f (new_AGEMA_signal_3565), .B0_t (StateFromRhoPi[72]), .B0_f (new_AGEMA_signal_3575), .B1_t (new_AGEMA_signal_3576), .B1_f (new_AGEMA_signal_3577), .Z0_t (CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_and_xor_inst_e_nxy), .Z0_f (new_AGEMA_signal_4065), .Z1_t (new_AGEMA_signal_4066), .Z1_f (new_AGEMA_signal_4067) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_and_xor_inst_e_nxy), .A0_f (new_AGEMA_signal_4065), .A1_t (new_AGEMA_signal_4066), .A1_f (new_AGEMA_signal_4067), .B0_t (StateFromRhoPi[192]), .B0_f (new_AGEMA_signal_3401), .B1_t (new_AGEMA_signal_3402), .B1_f (new_AGEMA_signal_3403), .Z0_t (StateFromChi[192]), .Z0_f (new_AGEMA_signal_4671), .Z1_t (new_AGEMA_signal_4672), .Z1_f (new_AGEMA_signal_4673) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_0__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[41]), .A0_f (new_AGEMA_signal_3890), .A1_t (new_AGEMA_signal_3891), .A1_f (new_AGEMA_signal_3892), .B0_t (StateFromRhoPi[81]), .B0_f (new_AGEMA_signal_3737), .B1_t (new_AGEMA_signal_3738), .B1_f (new_AGEMA_signal_3739), .Z0_t (CHI_GEN_SLICES_1__GEN_ROWS_0__sbox_and_xor_inst_a_nxy), .Z0_f (new_AGEMA_signal_4068), .Z1_t (new_AGEMA_signal_4069), .Z1_f (new_AGEMA_signal_4070) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_0__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_1__GEN_ROWS_0__sbox_and_xor_inst_a_nxy), .A0_f (new_AGEMA_signal_4068), .A1_t (new_AGEMA_signal_4069), .A1_f (new_AGEMA_signal_4070), .B0_t (StateFromRhoPi[1]), .B0_f (new_AGEMA_signal_3548), .B1_t (new_AGEMA_signal_3549), .B1_f (new_AGEMA_signal_3550), .Z0_t (CHI_ChiOut[1]), .Z0_f (new_AGEMA_signal_4674), .Z1_t (new_AGEMA_signal_4675), .Z1_f (new_AGEMA_signal_4676) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_0__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[81]), .A0_f (new_AGEMA_signal_3737), .A1_t (new_AGEMA_signal_3738), .A1_f (new_AGEMA_signal_3739), .B0_t (StateFromRhoPi[121]), .B0_f (new_AGEMA_signal_3959), .B1_t (new_AGEMA_signal_3960), .B1_f (new_AGEMA_signal_3961), .Z0_t (CHI_GEN_SLICES_1__GEN_ROWS_0__sbox_and_xor_inst_b_nxy), .Z0_f (new_AGEMA_signal_4071), .Z1_t (new_AGEMA_signal_4072), .Z1_f (new_AGEMA_signal_4073) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_0__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_1__GEN_ROWS_0__sbox_and_xor_inst_b_nxy), .A0_f (new_AGEMA_signal_4071), .A1_t (new_AGEMA_signal_4072), .A1_f (new_AGEMA_signal_4073), .B0_t (StateFromRhoPi[41]), .B0_f (new_AGEMA_signal_3890), .B1_t (new_AGEMA_signal_3891), .B1_f (new_AGEMA_signal_3892), .Z0_t (StateFromChi[41]), .Z0_f (new_AGEMA_signal_4677), .Z1_t (new_AGEMA_signal_4678), .Z1_f (new_AGEMA_signal_4679) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_0__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[121]), .A0_f (new_AGEMA_signal_3959), .A1_t (new_AGEMA_signal_3960), .A1_f (new_AGEMA_signal_3961), .B0_t (StateFromRhoPi[161]), .B0_f (new_AGEMA_signal_3776), .B1_t (new_AGEMA_signal_3777), .B1_f (new_AGEMA_signal_3778), .Z0_t (CHI_GEN_SLICES_1__GEN_ROWS_0__sbox_and_xor_inst_c_nxy), .Z0_f (new_AGEMA_signal_4074), .Z1_t (new_AGEMA_signal_4075), .Z1_f (new_AGEMA_signal_4076) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_0__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_1__GEN_ROWS_0__sbox_and_xor_inst_c_nxy), .A0_f (new_AGEMA_signal_4074), .A1_t (new_AGEMA_signal_4075), .A1_f (new_AGEMA_signal_4076), .B0_t (StateFromRhoPi[81]), .B0_f (new_AGEMA_signal_3737), .B1_t (new_AGEMA_signal_3738), .B1_f (new_AGEMA_signal_3739), .Z0_t (StateFromChi[81]), .Z0_f (new_AGEMA_signal_4680), .Z1_t (new_AGEMA_signal_4681), .Z1_f (new_AGEMA_signal_4682) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_0__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[161]), .A0_f (new_AGEMA_signal_3776), .A1_t (new_AGEMA_signal_3777), .A1_f (new_AGEMA_signal_3778), .B0_t (StateFromRhoPi[1]), .B0_f (new_AGEMA_signal_3548), .B1_t (new_AGEMA_signal_3549), .B1_f (new_AGEMA_signal_3550), .Z0_t (CHI_GEN_SLICES_1__GEN_ROWS_0__sbox_and_xor_inst_d_nxy), .Z0_f (new_AGEMA_signal_4077), .Z1_t (new_AGEMA_signal_4078), .Z1_f (new_AGEMA_signal_4079) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_0__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_1__GEN_ROWS_0__sbox_and_xor_inst_d_nxy), .A0_f (new_AGEMA_signal_4077), .A1_t (new_AGEMA_signal_4078), .A1_f (new_AGEMA_signal_4079), .B0_t (StateFromRhoPi[121]), .B0_f (new_AGEMA_signal_3959), .B1_t (new_AGEMA_signal_3960), .B1_f (new_AGEMA_signal_3961), .Z0_t (StateFromChi[121]), .Z0_f (new_AGEMA_signal_4683), .Z1_t (new_AGEMA_signal_4684), .Z1_f (new_AGEMA_signal_4685) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_0__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[1]), .A0_f (new_AGEMA_signal_3548), .A1_t (new_AGEMA_signal_3549), .A1_f (new_AGEMA_signal_3550), .B0_t (StateFromRhoPi[41]), .B0_f (new_AGEMA_signal_3890), .B1_t (new_AGEMA_signal_3891), .B1_f (new_AGEMA_signal_3892), .Z0_t (CHI_GEN_SLICES_1__GEN_ROWS_0__sbox_and_xor_inst_e_nxy), .Z0_f (new_AGEMA_signal_4080), .Z1_t (new_AGEMA_signal_4081), .Z1_f (new_AGEMA_signal_4082) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_0__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_1__GEN_ROWS_0__sbox_and_xor_inst_e_nxy), .A0_f (new_AGEMA_signal_4080), .A1_t (new_AGEMA_signal_4081), .A1_f (new_AGEMA_signal_4082), .B0_t (StateFromRhoPi[161]), .B0_f (new_AGEMA_signal_3776), .B1_t (new_AGEMA_signal_3777), .B1_f (new_AGEMA_signal_3778), .Z0_t (StateFromChi[161]), .Z0_f (new_AGEMA_signal_4686), .Z1_t (new_AGEMA_signal_4687), .Z1_f (new_AGEMA_signal_4688) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_1__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[49]), .A0_f (new_AGEMA_signal_3800), .A1_t (new_AGEMA_signal_3801), .A1_f (new_AGEMA_signal_3802), .B0_t (StateFromRhoPi[89]), .B0_f (new_AGEMA_signal_3767), .B1_t (new_AGEMA_signal_3768), .B1_f (new_AGEMA_signal_3769), .Z0_t (CHI_GEN_SLICES_1__GEN_ROWS_1__sbox_and_xor_inst_a_nxy), .Z0_f (new_AGEMA_signal_4083), .Z1_t (new_AGEMA_signal_4084), .Z1_f (new_AGEMA_signal_4085) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_1__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_1__GEN_ROWS_1__sbox_and_xor_inst_a_nxy), .A0_f (new_AGEMA_signal_4083), .A1_t (new_AGEMA_signal_4084), .A1_f (new_AGEMA_signal_4085), .B0_t (StateFromRhoPi[9]), .B0_f (new_AGEMA_signal_3938), .B1_t (new_AGEMA_signal_3939), .B1_f (new_AGEMA_signal_3940), .Z0_t (StateFromChi[9]), .Z0_f (new_AGEMA_signal_4689), .Z1_t (new_AGEMA_signal_4690), .Z1_f (new_AGEMA_signal_4691) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_1__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[89]), .A0_f (new_AGEMA_signal_3767), .A1_t (new_AGEMA_signal_3768), .A1_f (new_AGEMA_signal_3769), .B0_t (StateFromRhoPi[129]), .B0_f (new_AGEMA_signal_3809), .B1_t (new_AGEMA_signal_3810), .B1_f (new_AGEMA_signal_3811), .Z0_t (CHI_GEN_SLICES_1__GEN_ROWS_1__sbox_and_xor_inst_b_nxy), .Z0_f (new_AGEMA_signal_4086), .Z1_t (new_AGEMA_signal_4087), .Z1_f (new_AGEMA_signal_4088) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_1__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_1__GEN_ROWS_1__sbox_and_xor_inst_b_nxy), .A0_f (new_AGEMA_signal_4086), .A1_t (new_AGEMA_signal_4087), .A1_f (new_AGEMA_signal_4088), .B0_t (StateFromRhoPi[49]), .B0_f (new_AGEMA_signal_3800), .B1_t (new_AGEMA_signal_3801), .B1_f (new_AGEMA_signal_3802), .Z0_t (StateFromChi[49]), .Z0_f (new_AGEMA_signal_4692), .Z1_t (new_AGEMA_signal_4693), .Z1_f (new_AGEMA_signal_4694) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_1__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[129]), .A0_f (new_AGEMA_signal_3809), .A1_t (new_AGEMA_signal_3810), .A1_f (new_AGEMA_signal_3811), .B0_t (StateFromRhoPi[169]), .B0_f (new_AGEMA_signal_3821), .B1_t (new_AGEMA_signal_3822), .B1_f (new_AGEMA_signal_3823), .Z0_t (CHI_GEN_SLICES_1__GEN_ROWS_1__sbox_and_xor_inst_c_nxy), .Z0_f (new_AGEMA_signal_4089), .Z1_t (new_AGEMA_signal_4090), .Z1_f (new_AGEMA_signal_4091) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_1__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_1__GEN_ROWS_1__sbox_and_xor_inst_c_nxy), .A0_f (new_AGEMA_signal_4089), .A1_t (new_AGEMA_signal_4090), .A1_f (new_AGEMA_signal_4091), .B0_t (StateFromRhoPi[89]), .B0_f (new_AGEMA_signal_3767), .B1_t (new_AGEMA_signal_3768), .B1_f (new_AGEMA_signal_3769), .Z0_t (StateFromChi[89]), .Z0_f (new_AGEMA_signal_4695), .Z1_t (new_AGEMA_signal_4696), .Z1_f (new_AGEMA_signal_4697) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_1__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[169]), .A0_f (new_AGEMA_signal_3821), .A1_t (new_AGEMA_signal_3822), .A1_f (new_AGEMA_signal_3823), .B0_t (StateFromRhoPi[9]), .B0_f (new_AGEMA_signal_3938), .B1_t (new_AGEMA_signal_3939), .B1_f (new_AGEMA_signal_3940), .Z0_t (CHI_GEN_SLICES_1__GEN_ROWS_1__sbox_and_xor_inst_d_nxy), .Z0_f (new_AGEMA_signal_4092), .Z1_t (new_AGEMA_signal_4093), .Z1_f (new_AGEMA_signal_4094) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_1__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_1__GEN_ROWS_1__sbox_and_xor_inst_d_nxy), .A0_f (new_AGEMA_signal_4092), .A1_t (new_AGEMA_signal_4093), .A1_f (new_AGEMA_signal_4094), .B0_t (StateFromRhoPi[129]), .B0_f (new_AGEMA_signal_3809), .B1_t (new_AGEMA_signal_3810), .B1_f (new_AGEMA_signal_3811), .Z0_t (StateFromChi[129]), .Z0_f (new_AGEMA_signal_4698), .Z1_t (new_AGEMA_signal_4699), .Z1_f (new_AGEMA_signal_4700) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_1__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[9]), .A0_f (new_AGEMA_signal_3938), .A1_t (new_AGEMA_signal_3939), .A1_f (new_AGEMA_signal_3940), .B0_t (StateFromRhoPi[49]), .B0_f (new_AGEMA_signal_3800), .B1_t (new_AGEMA_signal_3801), .B1_f (new_AGEMA_signal_3802), .Z0_t (CHI_GEN_SLICES_1__GEN_ROWS_1__sbox_and_xor_inst_e_nxy), .Z0_f (new_AGEMA_signal_4095), .Z1_t (new_AGEMA_signal_4096), .Z1_f (new_AGEMA_signal_4097) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_1__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_1__GEN_ROWS_1__sbox_and_xor_inst_e_nxy), .A0_f (new_AGEMA_signal_4095), .A1_t (new_AGEMA_signal_4096), .A1_f (new_AGEMA_signal_4097), .B0_t (StateFromRhoPi[169]), .B0_f (new_AGEMA_signal_3821), .B1_t (new_AGEMA_signal_3822), .B1_f (new_AGEMA_signal_3823), .Z0_t (StateFromChi[169]), .Z0_f (new_AGEMA_signal_4701), .Z1_t (new_AGEMA_signal_4702), .Z1_f (new_AGEMA_signal_4703) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_2__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[57]), .A0_f (new_AGEMA_signal_3860), .A1_t (new_AGEMA_signal_3861), .A1_f (new_AGEMA_signal_3862), .B0_t (StateFromRhoPi[97]), .B0_f (new_AGEMA_signal_3662), .B1_t (new_AGEMA_signal_3663), .B1_f (new_AGEMA_signal_3664), .Z0_t (CHI_GEN_SLICES_1__GEN_ROWS_2__sbox_and_xor_inst_a_nxy), .Z0_f (new_AGEMA_signal_4098), .Z1_t (new_AGEMA_signal_4099), .Z1_f (new_AGEMA_signal_4100) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_2__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_1__GEN_ROWS_2__sbox_and_xor_inst_a_nxy), .A0_f (new_AGEMA_signal_4098), .A1_t (new_AGEMA_signal_4099), .A1_f (new_AGEMA_signal_4100), .B0_t (StateFromRhoPi[17]), .B0_f (new_AGEMA_signal_3518), .B1_t (new_AGEMA_signal_3519), .B1_f (new_AGEMA_signal_3520), .Z0_t (StateFromChi[17]), .Z0_f (new_AGEMA_signal_4704), .Z1_t (new_AGEMA_signal_4705), .Z1_f (new_AGEMA_signal_4706) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_2__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[97]), .A0_f (new_AGEMA_signal_3662), .A1_t (new_AGEMA_signal_3663), .A1_f (new_AGEMA_signal_3664), .B0_t (StateFromRhoPi[137]), .B0_f (new_AGEMA_signal_3494), .B1_t (new_AGEMA_signal_3495), .B1_f (new_AGEMA_signal_3496), .Z0_t (CHI_GEN_SLICES_1__GEN_ROWS_2__sbox_and_xor_inst_b_nxy), .Z0_f (new_AGEMA_signal_4101), .Z1_t (new_AGEMA_signal_4102), .Z1_f (new_AGEMA_signal_4103) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_2__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_1__GEN_ROWS_2__sbox_and_xor_inst_b_nxy), .A0_f (new_AGEMA_signal_4101), .A1_t (new_AGEMA_signal_4102), .A1_f (new_AGEMA_signal_4103), .B0_t (StateFromRhoPi[57]), .B0_f (new_AGEMA_signal_3860), .B1_t (new_AGEMA_signal_3861), .B1_f (new_AGEMA_signal_3862), .Z0_t (StateFromChi[57]), .Z0_f (new_AGEMA_signal_4707), .Z1_t (new_AGEMA_signal_4708), .Z1_f (new_AGEMA_signal_4709) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_2__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[137]), .A0_f (new_AGEMA_signal_3494), .A1_t (new_AGEMA_signal_3495), .A1_f (new_AGEMA_signal_3496), .B0_t (StateFromRhoPi[177]), .B0_f (new_AGEMA_signal_3716), .B1_t (new_AGEMA_signal_3717), .B1_f (new_AGEMA_signal_3718), .Z0_t (CHI_GEN_SLICES_1__GEN_ROWS_2__sbox_and_xor_inst_c_nxy), .Z0_f (new_AGEMA_signal_4104), .Z1_t (new_AGEMA_signal_4105), .Z1_f (new_AGEMA_signal_4106) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_2__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_1__GEN_ROWS_2__sbox_and_xor_inst_c_nxy), .A0_f (new_AGEMA_signal_4104), .A1_t (new_AGEMA_signal_4105), .A1_f (new_AGEMA_signal_4106), .B0_t (StateFromRhoPi[97]), .B0_f (new_AGEMA_signal_3662), .B1_t (new_AGEMA_signal_3663), .B1_f (new_AGEMA_signal_3664), .Z0_t (StateFromChi[97]), .Z0_f (new_AGEMA_signal_4710), .Z1_t (new_AGEMA_signal_4711), .Z1_f (new_AGEMA_signal_4712) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_2__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[177]), .A0_f (new_AGEMA_signal_3716), .A1_t (new_AGEMA_signal_3717), .A1_f (new_AGEMA_signal_3718), .B0_t (StateFromRhoPi[17]), .B0_f (new_AGEMA_signal_3518), .B1_t (new_AGEMA_signal_3519), .B1_f (new_AGEMA_signal_3520), .Z0_t (CHI_GEN_SLICES_1__GEN_ROWS_2__sbox_and_xor_inst_d_nxy), .Z0_f (new_AGEMA_signal_4107), .Z1_t (new_AGEMA_signal_4108), .Z1_f (new_AGEMA_signal_4109) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_2__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_1__GEN_ROWS_2__sbox_and_xor_inst_d_nxy), .A0_f (new_AGEMA_signal_4107), .A1_t (new_AGEMA_signal_4108), .A1_f (new_AGEMA_signal_4109), .B0_t (StateFromRhoPi[137]), .B0_f (new_AGEMA_signal_3494), .B1_t (new_AGEMA_signal_3495), .B1_f (new_AGEMA_signal_3496), .Z0_t (StateFromChi[137]), .Z0_f (new_AGEMA_signal_4713), .Z1_t (new_AGEMA_signal_4714), .Z1_f (new_AGEMA_signal_4715) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_2__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[17]), .A0_f (new_AGEMA_signal_3518), .A1_t (new_AGEMA_signal_3519), .A1_f (new_AGEMA_signal_3520), .B0_t (StateFromRhoPi[57]), .B0_f (new_AGEMA_signal_3860), .B1_t (new_AGEMA_signal_3861), .B1_f (new_AGEMA_signal_3862), .Z0_t (CHI_GEN_SLICES_1__GEN_ROWS_2__sbox_and_xor_inst_e_nxy), .Z0_f (new_AGEMA_signal_4110), .Z1_t (new_AGEMA_signal_4111), .Z1_f (new_AGEMA_signal_4112) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_2__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_1__GEN_ROWS_2__sbox_and_xor_inst_e_nxy), .A0_f (new_AGEMA_signal_4110), .A1_t (new_AGEMA_signal_4111), .A1_f (new_AGEMA_signal_4112), .B0_t (StateFromRhoPi[177]), .B0_f (new_AGEMA_signal_3716), .B1_t (new_AGEMA_signal_3717), .B1_f (new_AGEMA_signal_3718), .Z0_t (StateFromChi[177]), .Z0_f (new_AGEMA_signal_4716), .Z1_t (new_AGEMA_signal_4717), .Z1_f (new_AGEMA_signal_4718) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_3__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[65]), .A0_f (new_AGEMA_signal_3845), .A1_t (new_AGEMA_signal_3846), .A1_f (new_AGEMA_signal_3847), .B0_t (StateFromRhoPi[105]), .B0_f (new_AGEMA_signal_3632), .B1_t (new_AGEMA_signal_3633), .B1_f (new_AGEMA_signal_3634), .Z0_t (CHI_GEN_SLICES_1__GEN_ROWS_3__sbox_and_xor_inst_a_nxy), .Z0_f (new_AGEMA_signal_4113), .Z1_t (new_AGEMA_signal_4114), .Z1_f (new_AGEMA_signal_4115) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_3__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_1__GEN_ROWS_3__sbox_and_xor_inst_a_nxy), .A0_f (new_AGEMA_signal_4113), .A1_t (new_AGEMA_signal_4114), .A1_f (new_AGEMA_signal_4115), .B0_t (StateFromRhoPi[25]), .B0_f (new_AGEMA_signal_3443), .B1_t (new_AGEMA_signal_3444), .B1_f (new_AGEMA_signal_3445), .Z0_t (StateFromChi[25]), .Z0_f (new_AGEMA_signal_4719), .Z1_t (new_AGEMA_signal_4720), .Z1_f (new_AGEMA_signal_4721) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_3__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[105]), .A0_f (new_AGEMA_signal_3632), .A1_t (new_AGEMA_signal_3633), .A1_f (new_AGEMA_signal_3634), .B0_t (StateFromRhoPi[145]), .B0_f (new_AGEMA_signal_3554), .B1_t (new_AGEMA_signal_3555), .B1_f (new_AGEMA_signal_3556), .Z0_t (CHI_GEN_SLICES_1__GEN_ROWS_3__sbox_and_xor_inst_b_nxy), .Z0_f (new_AGEMA_signal_4116), .Z1_t (new_AGEMA_signal_4117), .Z1_f (new_AGEMA_signal_4118) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_3__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_1__GEN_ROWS_3__sbox_and_xor_inst_b_nxy), .A0_f (new_AGEMA_signal_4116), .A1_t (new_AGEMA_signal_4117), .A1_f (new_AGEMA_signal_4118), .B0_t (StateFromRhoPi[65]), .B0_f (new_AGEMA_signal_3845), .B1_t (new_AGEMA_signal_3846), .B1_f (new_AGEMA_signal_3847), .Z0_t (StateFromChi[65]), .Z0_f (new_AGEMA_signal_4722), .Z1_t (new_AGEMA_signal_4723), .Z1_f (new_AGEMA_signal_4724) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_3__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[145]), .A0_f (new_AGEMA_signal_3554), .A1_t (new_AGEMA_signal_3555), .A1_f (new_AGEMA_signal_3556), .B0_t (StateFromRhoPi[185]), .B0_f (new_AGEMA_signal_3566), .B1_t (new_AGEMA_signal_3567), .B1_f (new_AGEMA_signal_3568), .Z0_t (CHI_GEN_SLICES_1__GEN_ROWS_3__sbox_and_xor_inst_c_nxy), .Z0_f (new_AGEMA_signal_4119), .Z1_t (new_AGEMA_signal_4120), .Z1_f (new_AGEMA_signal_4121) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_3__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_1__GEN_ROWS_3__sbox_and_xor_inst_c_nxy), .A0_f (new_AGEMA_signal_4119), .A1_t (new_AGEMA_signal_4120), .A1_f (new_AGEMA_signal_4121), .B0_t (StateFromRhoPi[105]), .B0_f (new_AGEMA_signal_3632), .B1_t (new_AGEMA_signal_3633), .B1_f (new_AGEMA_signal_3634), .Z0_t (StateFromChi[105]), .Z0_f (new_AGEMA_signal_4725), .Z1_t (new_AGEMA_signal_4726), .Z1_f (new_AGEMA_signal_4727) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_3__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[185]), .A0_f (new_AGEMA_signal_3566), .A1_t (new_AGEMA_signal_3567), .A1_f (new_AGEMA_signal_3568), .B0_t (StateFromRhoPi[25]), .B0_f (new_AGEMA_signal_3443), .B1_t (new_AGEMA_signal_3444), .B1_f (new_AGEMA_signal_3445), .Z0_t (CHI_GEN_SLICES_1__GEN_ROWS_3__sbox_and_xor_inst_d_nxy), .Z0_f (new_AGEMA_signal_4122), .Z1_t (new_AGEMA_signal_4123), .Z1_f (new_AGEMA_signal_4124) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_3__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_1__GEN_ROWS_3__sbox_and_xor_inst_d_nxy), .A0_f (new_AGEMA_signal_4122), .A1_t (new_AGEMA_signal_4123), .A1_f (new_AGEMA_signal_4124), .B0_t (StateFromRhoPi[145]), .B0_f (new_AGEMA_signal_3554), .B1_t (new_AGEMA_signal_3555), .B1_f (new_AGEMA_signal_3556), .Z0_t (StateFromChi[145]), .Z0_f (new_AGEMA_signal_4728), .Z1_t (new_AGEMA_signal_4729), .Z1_f (new_AGEMA_signal_4730) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_3__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[25]), .A0_f (new_AGEMA_signal_3443), .A1_t (new_AGEMA_signal_3444), .A1_f (new_AGEMA_signal_3445), .B0_t (StateFromRhoPi[65]), .B0_f (new_AGEMA_signal_3845), .B1_t (new_AGEMA_signal_3846), .B1_f (new_AGEMA_signal_3847), .Z0_t (CHI_GEN_SLICES_1__GEN_ROWS_3__sbox_and_xor_inst_e_nxy), .Z0_f (new_AGEMA_signal_4125), .Z1_t (new_AGEMA_signal_4126), .Z1_f (new_AGEMA_signal_4127) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_3__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_1__GEN_ROWS_3__sbox_and_xor_inst_e_nxy), .A0_f (new_AGEMA_signal_4125), .A1_t (new_AGEMA_signal_4126), .A1_f (new_AGEMA_signal_4127), .B0_t (StateFromRhoPi[185]), .B0_f (new_AGEMA_signal_3566), .B1_t (new_AGEMA_signal_3567), .B1_f (new_AGEMA_signal_3568), .Z0_t (StateFromChi[185]), .Z0_f (new_AGEMA_signal_4731), .Z1_t (new_AGEMA_signal_4732), .Z1_f (new_AGEMA_signal_4733) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_4__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[73]), .A0_f (new_AGEMA_signal_3530), .A1_t (new_AGEMA_signal_3531), .A1_f (new_AGEMA_signal_3532), .B0_t (StateFromRhoPi[113]), .B0_f (new_AGEMA_signal_3947), .B1_t (new_AGEMA_signal_3948), .B1_f (new_AGEMA_signal_3949), .Z0_t (CHI_GEN_SLICES_1__GEN_ROWS_4__sbox_and_xor_inst_a_nxy), .Z0_f (new_AGEMA_signal_4128), .Z1_t (new_AGEMA_signal_4129), .Z1_f (new_AGEMA_signal_4130) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_4__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_1__GEN_ROWS_4__sbox_and_xor_inst_a_nxy), .A0_f (new_AGEMA_signal_4128), .A1_t (new_AGEMA_signal_4129), .A1_f (new_AGEMA_signal_4130), .B0_t (StateFromRhoPi[33]), .B0_f (new_AGEMA_signal_3863), .B1_t (new_AGEMA_signal_3864), .B1_f (new_AGEMA_signal_3865), .Z0_t (StateFromChi[33]), .Z0_f (new_AGEMA_signal_4734), .Z1_t (new_AGEMA_signal_4735), .Z1_f (new_AGEMA_signal_4736) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_4__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[113]), .A0_f (new_AGEMA_signal_3947), .A1_t (new_AGEMA_signal_3948), .A1_f (new_AGEMA_signal_3949), .B0_t (StateFromRhoPi[153]), .B0_f (new_AGEMA_signal_3599), .B1_t (new_AGEMA_signal_3600), .B1_f (new_AGEMA_signal_3601), .Z0_t (CHI_GEN_SLICES_1__GEN_ROWS_4__sbox_and_xor_inst_b_nxy), .Z0_f (new_AGEMA_signal_4131), .Z1_t (new_AGEMA_signal_4132), .Z1_f (new_AGEMA_signal_4133) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_4__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_1__GEN_ROWS_4__sbox_and_xor_inst_b_nxy), .A0_f (new_AGEMA_signal_4131), .A1_t (new_AGEMA_signal_4132), .A1_f (new_AGEMA_signal_4133), .B0_t (StateFromRhoPi[73]), .B0_f (new_AGEMA_signal_3530), .B1_t (new_AGEMA_signal_3531), .B1_f (new_AGEMA_signal_3532), .Z0_t (StateFromChi[73]), .Z0_f (new_AGEMA_signal_4737), .Z1_t (new_AGEMA_signal_4738), .Z1_f (new_AGEMA_signal_4739) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_4__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[153]), .A0_f (new_AGEMA_signal_3599), .A1_t (new_AGEMA_signal_3600), .A1_f (new_AGEMA_signal_3601), .B0_t (StateFromRhoPi[193]), .B0_f (new_AGEMA_signal_3626), .B1_t (new_AGEMA_signal_3627), .B1_f (new_AGEMA_signal_3628), .Z0_t (CHI_GEN_SLICES_1__GEN_ROWS_4__sbox_and_xor_inst_c_nxy), .Z0_f (new_AGEMA_signal_4134), .Z1_t (new_AGEMA_signal_4135), .Z1_f (new_AGEMA_signal_4136) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_4__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_1__GEN_ROWS_4__sbox_and_xor_inst_c_nxy), .A0_f (new_AGEMA_signal_4134), .A1_t (new_AGEMA_signal_4135), .A1_f (new_AGEMA_signal_4136), .B0_t (StateFromRhoPi[113]), .B0_f (new_AGEMA_signal_3947), .B1_t (new_AGEMA_signal_3948), .B1_f (new_AGEMA_signal_3949), .Z0_t (StateFromChi[113]), .Z0_f (new_AGEMA_signal_4740), .Z1_t (new_AGEMA_signal_4741), .Z1_f (new_AGEMA_signal_4742) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_4__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[193]), .A0_f (new_AGEMA_signal_3626), .A1_t (new_AGEMA_signal_3627), .A1_f (new_AGEMA_signal_3628), .B0_t (StateFromRhoPi[33]), .B0_f (new_AGEMA_signal_3863), .B1_t (new_AGEMA_signal_3864), .B1_f (new_AGEMA_signal_3865), .Z0_t (CHI_GEN_SLICES_1__GEN_ROWS_4__sbox_and_xor_inst_d_nxy), .Z0_f (new_AGEMA_signal_4137), .Z1_t (new_AGEMA_signal_4138), .Z1_f (new_AGEMA_signal_4139) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_4__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_1__GEN_ROWS_4__sbox_and_xor_inst_d_nxy), .A0_f (new_AGEMA_signal_4137), .A1_t (new_AGEMA_signal_4138), .A1_f (new_AGEMA_signal_4139), .B0_t (StateFromRhoPi[153]), .B0_f (new_AGEMA_signal_3599), .B1_t (new_AGEMA_signal_3600), .B1_f (new_AGEMA_signal_3601), .Z0_t (StateFromChi[153]), .Z0_f (new_AGEMA_signal_4743), .Z1_t (new_AGEMA_signal_4744), .Z1_f (new_AGEMA_signal_4745) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_4__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[33]), .A0_f (new_AGEMA_signal_3863), .A1_t (new_AGEMA_signal_3864), .A1_f (new_AGEMA_signal_3865), .B0_t (StateFromRhoPi[73]), .B0_f (new_AGEMA_signal_3530), .B1_t (new_AGEMA_signal_3531), .B1_f (new_AGEMA_signal_3532), .Z0_t (CHI_GEN_SLICES_1__GEN_ROWS_4__sbox_and_xor_inst_e_nxy), .Z0_f (new_AGEMA_signal_4140), .Z1_t (new_AGEMA_signal_4141), .Z1_f (new_AGEMA_signal_4142) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_4__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_1__GEN_ROWS_4__sbox_and_xor_inst_e_nxy), .A0_f (new_AGEMA_signal_4140), .A1_t (new_AGEMA_signal_4141), .A1_f (new_AGEMA_signal_4142), .B0_t (StateFromRhoPi[193]), .B0_f (new_AGEMA_signal_3626), .B1_t (new_AGEMA_signal_3627), .B1_f (new_AGEMA_signal_3628), .Z0_t (StateFromChi[193]), .Z0_f (new_AGEMA_signal_4746), .Z1_t (new_AGEMA_signal_4747), .Z1_f (new_AGEMA_signal_4748) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_0__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[42]), .A0_f (new_AGEMA_signal_3410), .A1_t (new_AGEMA_signal_3411), .A1_f (new_AGEMA_signal_3412), .B0_t (StateFromRhoPi[82]), .B0_f (new_AGEMA_signal_3452), .B1_t (new_AGEMA_signal_3453), .B1_f (new_AGEMA_signal_3454), .Z0_t (CHI_GEN_SLICES_2__GEN_ROWS_0__sbox_and_xor_inst_a_nxy), .Z0_f (new_AGEMA_signal_4143), .Z1_t (new_AGEMA_signal_4144), .Z1_f (new_AGEMA_signal_4145) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_0__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_2__GEN_ROWS_0__sbox_and_xor_inst_a_nxy), .A0_f (new_AGEMA_signal_4143), .A1_t (new_AGEMA_signal_4144), .A1_f (new_AGEMA_signal_4145), .B0_t (StateFromRhoPi[2]), .B0_f (new_AGEMA_signal_3713), .B1_t (new_AGEMA_signal_3714), .B1_f (new_AGEMA_signal_3715), .Z0_t (StateFromChi[2]), .Z0_f (new_AGEMA_signal_4749), .Z1_t (new_AGEMA_signal_4750), .Z1_f (new_AGEMA_signal_4751) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_0__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[82]), .A0_f (new_AGEMA_signal_3452), .A1_t (new_AGEMA_signal_3453), .A1_f (new_AGEMA_signal_3454), .B0_t (StateFromRhoPi[122]), .B0_f (new_AGEMA_signal_3929), .B1_t (new_AGEMA_signal_3930), .B1_f (new_AGEMA_signal_3931), .Z0_t (CHI_GEN_SLICES_2__GEN_ROWS_0__sbox_and_xor_inst_b_nxy), .Z0_f (new_AGEMA_signal_4146), .Z1_t (new_AGEMA_signal_4147), .Z1_f (new_AGEMA_signal_4148) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_0__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_2__GEN_ROWS_0__sbox_and_xor_inst_b_nxy), .A0_f (new_AGEMA_signal_4146), .A1_t (new_AGEMA_signal_4147), .A1_f (new_AGEMA_signal_4148), .B0_t (StateFromRhoPi[42]), .B0_f (new_AGEMA_signal_3410), .B1_t (new_AGEMA_signal_3411), .B1_f (new_AGEMA_signal_3412), .Z0_t (StateFromChi[42]), .Z0_f (new_AGEMA_signal_4752), .Z1_t (new_AGEMA_signal_4753), .Z1_f (new_AGEMA_signal_4754) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_0__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[122]), .A0_f (new_AGEMA_signal_3929), .A1_t (new_AGEMA_signal_3930), .A1_f (new_AGEMA_signal_3931), .B0_t (StateFromRhoPi[162]), .B0_f (new_AGEMA_signal_3461), .B1_t (new_AGEMA_signal_3462), .B1_f (new_AGEMA_signal_3463), .Z0_t (CHI_GEN_SLICES_2__GEN_ROWS_0__sbox_and_xor_inst_c_nxy), .Z0_f (new_AGEMA_signal_4149), .Z1_t (new_AGEMA_signal_4150), .Z1_f (new_AGEMA_signal_4151) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_0__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_2__GEN_ROWS_0__sbox_and_xor_inst_c_nxy), .A0_f (new_AGEMA_signal_4149), .A1_t (new_AGEMA_signal_4150), .A1_f (new_AGEMA_signal_4151), .B0_t (StateFromRhoPi[82]), .B0_f (new_AGEMA_signal_3452), .B1_t (new_AGEMA_signal_3453), .B1_f (new_AGEMA_signal_3454), .Z0_t (StateFromChi[82]), .Z0_f (new_AGEMA_signal_4755), .Z1_t (new_AGEMA_signal_4756), .Z1_f (new_AGEMA_signal_4757) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_0__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[162]), .A0_f (new_AGEMA_signal_3461), .A1_t (new_AGEMA_signal_3462), .A1_f (new_AGEMA_signal_3463), .B0_t (StateFromRhoPi[2]), .B0_f (new_AGEMA_signal_3713), .B1_t (new_AGEMA_signal_3714), .B1_f (new_AGEMA_signal_3715), .Z0_t (CHI_GEN_SLICES_2__GEN_ROWS_0__sbox_and_xor_inst_d_nxy), .Z0_f (new_AGEMA_signal_4152), .Z1_t (new_AGEMA_signal_4153), .Z1_f (new_AGEMA_signal_4154) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_0__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_2__GEN_ROWS_0__sbox_and_xor_inst_d_nxy), .A0_f (new_AGEMA_signal_4152), .A1_t (new_AGEMA_signal_4153), .A1_f (new_AGEMA_signal_4154), .B0_t (StateFromRhoPi[122]), .B0_f (new_AGEMA_signal_3929), .B1_t (new_AGEMA_signal_3930), .B1_f (new_AGEMA_signal_3931), .Z0_t (StateFromChi[122]), .Z0_f (new_AGEMA_signal_4758), .Z1_t (new_AGEMA_signal_4759), .Z1_f (new_AGEMA_signal_4760) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_0__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[2]), .A0_f (new_AGEMA_signal_3713), .A1_t (new_AGEMA_signal_3714), .A1_f (new_AGEMA_signal_3715), .B0_t (StateFromRhoPi[42]), .B0_f (new_AGEMA_signal_3410), .B1_t (new_AGEMA_signal_3411), .B1_f (new_AGEMA_signal_3412), .Z0_t (CHI_GEN_SLICES_2__GEN_ROWS_0__sbox_and_xor_inst_e_nxy), .Z0_f (new_AGEMA_signal_4155), .Z1_t (new_AGEMA_signal_4156), .Z1_f (new_AGEMA_signal_4157) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_0__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_2__GEN_ROWS_0__sbox_and_xor_inst_e_nxy), .A0_f (new_AGEMA_signal_4155), .A1_t (new_AGEMA_signal_4156), .A1_f (new_AGEMA_signal_4157), .B0_t (StateFromRhoPi[162]), .B0_f (new_AGEMA_signal_3461), .B1_t (new_AGEMA_signal_3462), .B1_f (new_AGEMA_signal_3463), .Z0_t (StateFromChi[162]), .Z0_f (new_AGEMA_signal_4761), .Z1_t (new_AGEMA_signal_4762), .Z1_f (new_AGEMA_signal_4763) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_1__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[50]), .A0_f (new_AGEMA_signal_3440), .A1_t (new_AGEMA_signal_3441), .A1_f (new_AGEMA_signal_3442), .B0_t (StateFromRhoPi[90]), .B0_f (new_AGEMA_signal_3722), .B1_t (new_AGEMA_signal_3723), .B1_f (new_AGEMA_signal_3724), .Z0_t (CHI_GEN_SLICES_2__GEN_ROWS_1__sbox_and_xor_inst_a_nxy), .Z0_f (new_AGEMA_signal_4158), .Z1_t (new_AGEMA_signal_4159), .Z1_f (new_AGEMA_signal_4160) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_1__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_2__GEN_ROWS_1__sbox_and_xor_inst_a_nxy), .A0_f (new_AGEMA_signal_4158), .A1_t (new_AGEMA_signal_4159), .A1_f (new_AGEMA_signal_4160), .B0_t (StateFromRhoPi[10]), .B0_f (new_AGEMA_signal_3923), .B1_t (new_AGEMA_signal_3924), .B1_f (new_AGEMA_signal_3925), .Z0_t (StateFromChi[10]), .Z0_f (new_AGEMA_signal_4764), .Z1_t (new_AGEMA_signal_4765), .Z1_f (new_AGEMA_signal_4766) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_1__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[90]), .A0_f (new_AGEMA_signal_3722), .A1_t (new_AGEMA_signal_3723), .A1_f (new_AGEMA_signal_3724), .B0_t (StateFromRhoPi[130]), .B0_f (new_AGEMA_signal_3884), .B1_t (new_AGEMA_signal_3885), .B1_f (new_AGEMA_signal_3886), .Z0_t (CHI_GEN_SLICES_2__GEN_ROWS_1__sbox_and_xor_inst_b_nxy), .Z0_f (new_AGEMA_signal_4161), .Z1_t (new_AGEMA_signal_4162), .Z1_f (new_AGEMA_signal_4163) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_1__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_2__GEN_ROWS_1__sbox_and_xor_inst_b_nxy), .A0_f (new_AGEMA_signal_4161), .A1_t (new_AGEMA_signal_4162), .A1_f (new_AGEMA_signal_4163), .B0_t (StateFromRhoPi[50]), .B0_f (new_AGEMA_signal_3440), .B1_t (new_AGEMA_signal_3441), .B1_f (new_AGEMA_signal_3442), .Z0_t (StateFromChi[50]), .Z0_f (new_AGEMA_signal_4767), .Z1_t (new_AGEMA_signal_4768), .Z1_f (new_AGEMA_signal_4769) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_1__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[130]), .A0_f (new_AGEMA_signal_3884), .A1_t (new_AGEMA_signal_3885), .A1_f (new_AGEMA_signal_3886), .B0_t (StateFromRhoPi[170]), .B0_f (new_AGEMA_signal_3641), .B1_t (new_AGEMA_signal_3642), .B1_f (new_AGEMA_signal_3643), .Z0_t (CHI_GEN_SLICES_2__GEN_ROWS_1__sbox_and_xor_inst_c_nxy), .Z0_f (new_AGEMA_signal_4164), .Z1_t (new_AGEMA_signal_4165), .Z1_f (new_AGEMA_signal_4166) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_1__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_2__GEN_ROWS_1__sbox_and_xor_inst_c_nxy), .A0_f (new_AGEMA_signal_4164), .A1_t (new_AGEMA_signal_4165), .A1_f (new_AGEMA_signal_4166), .B0_t (StateFromRhoPi[90]), .B0_f (new_AGEMA_signal_3722), .B1_t (new_AGEMA_signal_3723), .B1_f (new_AGEMA_signal_3724), .Z0_t (StateFromChi[90]), .Z0_f (new_AGEMA_signal_4770), .Z1_t (new_AGEMA_signal_4771), .Z1_f (new_AGEMA_signal_4772) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_1__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[170]), .A0_f (new_AGEMA_signal_3641), .A1_t (new_AGEMA_signal_3642), .A1_f (new_AGEMA_signal_3643), .B0_t (StateFromRhoPi[10]), .B0_f (new_AGEMA_signal_3923), .B1_t (new_AGEMA_signal_3924), .B1_f (new_AGEMA_signal_3925), .Z0_t (CHI_GEN_SLICES_2__GEN_ROWS_1__sbox_and_xor_inst_d_nxy), .Z0_f (new_AGEMA_signal_4167), .Z1_t (new_AGEMA_signal_4168), .Z1_f (new_AGEMA_signal_4169) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_1__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_2__GEN_ROWS_1__sbox_and_xor_inst_d_nxy), .A0_f (new_AGEMA_signal_4167), .A1_t (new_AGEMA_signal_4168), .A1_f (new_AGEMA_signal_4169), .B0_t (StateFromRhoPi[130]), .B0_f (new_AGEMA_signal_3884), .B1_t (new_AGEMA_signal_3885), .B1_f (new_AGEMA_signal_3886), .Z0_t (StateFromChi[130]), .Z0_f (new_AGEMA_signal_4773), .Z1_t (new_AGEMA_signal_4774), .Z1_f (new_AGEMA_signal_4775) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_1__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[10]), .A0_f (new_AGEMA_signal_3923), .A1_t (new_AGEMA_signal_3924), .A1_f (new_AGEMA_signal_3925), .B0_t (StateFromRhoPi[50]), .B0_f (new_AGEMA_signal_3440), .B1_t (new_AGEMA_signal_3441), .B1_f (new_AGEMA_signal_3442), .Z0_t (CHI_GEN_SLICES_2__GEN_ROWS_1__sbox_and_xor_inst_e_nxy), .Z0_f (new_AGEMA_signal_4170), .Z1_t (new_AGEMA_signal_4171), .Z1_f (new_AGEMA_signal_4172) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_1__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_2__GEN_ROWS_1__sbox_and_xor_inst_e_nxy), .A0_f (new_AGEMA_signal_4170), .A1_t (new_AGEMA_signal_4171), .A1_f (new_AGEMA_signal_4172), .B0_t (StateFromRhoPi[170]), .B0_f (new_AGEMA_signal_3641), .B1_t (new_AGEMA_signal_3642), .B1_f (new_AGEMA_signal_3643), .Z0_t (StateFromChi[170]), .Z0_f (new_AGEMA_signal_4776), .Z1_t (new_AGEMA_signal_4777), .Z1_f (new_AGEMA_signal_4778) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_2__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[58]), .A0_f (new_AGEMA_signal_3830), .A1_t (new_AGEMA_signal_3831), .A1_f (new_AGEMA_signal_3832), .B0_t (StateFromRhoPi[98]), .B0_f (new_AGEMA_signal_3572), .B1_t (new_AGEMA_signal_3573), .B1_f (new_AGEMA_signal_3574), .Z0_t (CHI_GEN_SLICES_2__GEN_ROWS_2__sbox_and_xor_inst_a_nxy), .Z0_f (new_AGEMA_signal_4173), .Z1_t (new_AGEMA_signal_4174), .Z1_f (new_AGEMA_signal_4175) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_2__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_2__GEN_ROWS_2__sbox_and_xor_inst_a_nxy), .A0_f (new_AGEMA_signal_4173), .A1_t (new_AGEMA_signal_4174), .A1_f (new_AGEMA_signal_4175), .B0_t (StateFromRhoPi[18]), .B0_f (new_AGEMA_signal_3683), .B1_t (new_AGEMA_signal_3684), .B1_f (new_AGEMA_signal_3685), .Z0_t (StateFromChi[18]), .Z0_f (new_AGEMA_signal_4779), .Z1_t (new_AGEMA_signal_4780), .Z1_f (new_AGEMA_signal_4781) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_2__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[98]), .A0_f (new_AGEMA_signal_3572), .A1_t (new_AGEMA_signal_3573), .A1_f (new_AGEMA_signal_3574), .B0_t (StateFromRhoPi[138]), .B0_f (new_AGEMA_signal_3944), .B1_t (new_AGEMA_signal_3945), .B1_f (new_AGEMA_signal_3946), .Z0_t (CHI_GEN_SLICES_2__GEN_ROWS_2__sbox_and_xor_inst_b_nxy), .Z0_f (new_AGEMA_signal_4176), .Z1_t (new_AGEMA_signal_4177), .Z1_f (new_AGEMA_signal_4178) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_2__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_2__GEN_ROWS_2__sbox_and_xor_inst_b_nxy), .A0_f (new_AGEMA_signal_4176), .A1_t (new_AGEMA_signal_4177), .A1_f (new_AGEMA_signal_4178), .B0_t (StateFromRhoPi[58]), .B0_f (new_AGEMA_signal_3830), .B1_t (new_AGEMA_signal_3831), .B1_f (new_AGEMA_signal_3832), .Z0_t (StateFromChi[58]), .Z0_f (new_AGEMA_signal_4782), .Z1_t (new_AGEMA_signal_4783), .Z1_f (new_AGEMA_signal_4784) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_2__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[138]), .A0_f (new_AGEMA_signal_3944), .A1_t (new_AGEMA_signal_3945), .A1_f (new_AGEMA_signal_3946), .B0_t (StateFromRhoPi[178]), .B0_f (new_AGEMA_signal_3596), .B1_t (new_AGEMA_signal_3597), .B1_f (new_AGEMA_signal_3598), .Z0_t (CHI_GEN_SLICES_2__GEN_ROWS_2__sbox_and_xor_inst_c_nxy), .Z0_f (new_AGEMA_signal_4179), .Z1_t (new_AGEMA_signal_4180), .Z1_f (new_AGEMA_signal_4181) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_2__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_2__GEN_ROWS_2__sbox_and_xor_inst_c_nxy), .A0_f (new_AGEMA_signal_4179), .A1_t (new_AGEMA_signal_4180), .A1_f (new_AGEMA_signal_4181), .B0_t (StateFromRhoPi[98]), .B0_f (new_AGEMA_signal_3572), .B1_t (new_AGEMA_signal_3573), .B1_f (new_AGEMA_signal_3574), .Z0_t (StateFromChi[98]), .Z0_f (new_AGEMA_signal_4785), .Z1_t (new_AGEMA_signal_4786), .Z1_f (new_AGEMA_signal_4787) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_2__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[178]), .A0_f (new_AGEMA_signal_3596), .A1_t (new_AGEMA_signal_3597), .A1_f (new_AGEMA_signal_3598), .B0_t (StateFromRhoPi[18]), .B0_f (new_AGEMA_signal_3683), .B1_t (new_AGEMA_signal_3684), .B1_f (new_AGEMA_signal_3685), .Z0_t (CHI_GEN_SLICES_2__GEN_ROWS_2__sbox_and_xor_inst_d_nxy), .Z0_f (new_AGEMA_signal_4182), .Z1_t (new_AGEMA_signal_4183), .Z1_f (new_AGEMA_signal_4184) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_2__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_2__GEN_ROWS_2__sbox_and_xor_inst_d_nxy), .A0_f (new_AGEMA_signal_4182), .A1_t (new_AGEMA_signal_4183), .A1_f (new_AGEMA_signal_4184), .B0_t (StateFromRhoPi[138]), .B0_f (new_AGEMA_signal_3944), .B1_t (new_AGEMA_signal_3945), .B1_f (new_AGEMA_signal_3946), .Z0_t (StateFromChi[138]), .Z0_f (new_AGEMA_signal_4788), .Z1_t (new_AGEMA_signal_4789), .Z1_f (new_AGEMA_signal_4790) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_2__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[18]), .A0_f (new_AGEMA_signal_3683), .A1_t (new_AGEMA_signal_3684), .A1_f (new_AGEMA_signal_3685), .B0_t (StateFromRhoPi[58]), .B0_f (new_AGEMA_signal_3830), .B1_t (new_AGEMA_signal_3831), .B1_f (new_AGEMA_signal_3832), .Z0_t (CHI_GEN_SLICES_2__GEN_ROWS_2__sbox_and_xor_inst_e_nxy), .Z0_f (new_AGEMA_signal_4185), .Z1_t (new_AGEMA_signal_4186), .Z1_f (new_AGEMA_signal_4187) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_2__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_2__GEN_ROWS_2__sbox_and_xor_inst_e_nxy), .A0_f (new_AGEMA_signal_4185), .A1_t (new_AGEMA_signal_4186), .A1_f (new_AGEMA_signal_4187), .B0_t (StateFromRhoPi[178]), .B0_f (new_AGEMA_signal_3596), .B1_t (new_AGEMA_signal_3597), .B1_f (new_AGEMA_signal_3598), .Z0_t (StateFromChi[178]), .Z0_f (new_AGEMA_signal_4791), .Z1_t (new_AGEMA_signal_4792), .Z1_f (new_AGEMA_signal_4793) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_3__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[66]), .A0_f (new_AGEMA_signal_3770), .A1_t (new_AGEMA_signal_3771), .A1_f (new_AGEMA_signal_3772), .B0_t (StateFromRhoPi[106]), .B0_f (new_AGEMA_signal_3512), .B1_t (new_AGEMA_signal_3513), .B1_f (new_AGEMA_signal_3514), .Z0_t (CHI_GEN_SLICES_2__GEN_ROWS_3__sbox_and_xor_inst_a_nxy), .Z0_f (new_AGEMA_signal_4188), .Z1_t (new_AGEMA_signal_4189), .Z1_f (new_AGEMA_signal_4190) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_3__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_2__GEN_ROWS_3__sbox_and_xor_inst_a_nxy), .A0_f (new_AGEMA_signal_4188), .A1_t (new_AGEMA_signal_4189), .A1_f (new_AGEMA_signal_4190), .B0_t (StateFromRhoPi[26]), .B0_f (new_AGEMA_signal_3398), .B1_t (new_AGEMA_signal_3399), .B1_f (new_AGEMA_signal_3400), .Z0_t (StateFromChi[26]), .Z0_f (new_AGEMA_signal_4794), .Z1_t (new_AGEMA_signal_4795), .Z1_f (new_AGEMA_signal_4796) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_3__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[106]), .A0_f (new_AGEMA_signal_3512), .A1_t (new_AGEMA_signal_3513), .A1_f (new_AGEMA_signal_3514), .B0_t (StateFromRhoPi[146]), .B0_f (new_AGEMA_signal_3854), .B1_t (new_AGEMA_signal_3855), .B1_f (new_AGEMA_signal_3856), .Z0_t (CHI_GEN_SLICES_2__GEN_ROWS_3__sbox_and_xor_inst_b_nxy), .Z0_f (new_AGEMA_signal_4191), .Z1_t (new_AGEMA_signal_4192), .Z1_f (new_AGEMA_signal_4193) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_3__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_2__GEN_ROWS_3__sbox_and_xor_inst_b_nxy), .A0_f (new_AGEMA_signal_4191), .A1_t (new_AGEMA_signal_4192), .A1_f (new_AGEMA_signal_4193), .B0_t (StateFromRhoPi[66]), .B0_f (new_AGEMA_signal_3770), .B1_t (new_AGEMA_signal_3771), .B1_f (new_AGEMA_signal_3772), .Z0_t (StateFromChi[66]), .Z0_f (new_AGEMA_signal_4797), .Z1_t (new_AGEMA_signal_4798), .Z1_f (new_AGEMA_signal_4799) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_3__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[146]), .A0_f (new_AGEMA_signal_3854), .A1_t (new_AGEMA_signal_3855), .A1_f (new_AGEMA_signal_3856), .B0_t (StateFromRhoPi[186]), .B0_f (new_AGEMA_signal_3521), .B1_t (new_AGEMA_signal_3522), .B1_f (new_AGEMA_signal_3523), .Z0_t (CHI_GEN_SLICES_2__GEN_ROWS_3__sbox_and_xor_inst_c_nxy), .Z0_f (new_AGEMA_signal_4194), .Z1_t (new_AGEMA_signal_4195), .Z1_f (new_AGEMA_signal_4196) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_3__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_2__GEN_ROWS_3__sbox_and_xor_inst_c_nxy), .A0_f (new_AGEMA_signal_4194), .A1_t (new_AGEMA_signal_4195), .A1_f (new_AGEMA_signal_4196), .B0_t (StateFromRhoPi[106]), .B0_f (new_AGEMA_signal_3512), .B1_t (new_AGEMA_signal_3513), .B1_f (new_AGEMA_signal_3514), .Z0_t (StateFromChi[106]), .Z0_f (new_AGEMA_signal_4800), .Z1_t (new_AGEMA_signal_4801), .Z1_f (new_AGEMA_signal_4802) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_3__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[186]), .A0_f (new_AGEMA_signal_3521), .A1_t (new_AGEMA_signal_3522), .A1_f (new_AGEMA_signal_3523), .B0_t (StateFromRhoPi[26]), .B0_f (new_AGEMA_signal_3398), .B1_t (new_AGEMA_signal_3399), .B1_f (new_AGEMA_signal_3400), .Z0_t (CHI_GEN_SLICES_2__GEN_ROWS_3__sbox_and_xor_inst_d_nxy), .Z0_f (new_AGEMA_signal_4197), .Z1_t (new_AGEMA_signal_4198), .Z1_f (new_AGEMA_signal_4199) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_3__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_2__GEN_ROWS_3__sbox_and_xor_inst_d_nxy), .A0_f (new_AGEMA_signal_4197), .A1_t (new_AGEMA_signal_4198), .A1_f (new_AGEMA_signal_4199), .B0_t (StateFromRhoPi[146]), .B0_f (new_AGEMA_signal_3854), .B1_t (new_AGEMA_signal_3855), .B1_f (new_AGEMA_signal_3856), .Z0_t (StateFromChi[146]), .Z0_f (new_AGEMA_signal_4803), .Z1_t (new_AGEMA_signal_4804), .Z1_f (new_AGEMA_signal_4805) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_3__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[26]), .A0_f (new_AGEMA_signal_3398), .A1_t (new_AGEMA_signal_3399), .A1_f (new_AGEMA_signal_3400), .B0_t (StateFromRhoPi[66]), .B0_f (new_AGEMA_signal_3770), .B1_t (new_AGEMA_signal_3771), .B1_f (new_AGEMA_signal_3772), .Z0_t (CHI_GEN_SLICES_2__GEN_ROWS_3__sbox_and_xor_inst_e_nxy), .Z0_f (new_AGEMA_signal_4200), .Z1_t (new_AGEMA_signal_4201), .Z1_f (new_AGEMA_signal_4202) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_3__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_2__GEN_ROWS_3__sbox_and_xor_inst_e_nxy), .A0_f (new_AGEMA_signal_4200), .A1_t (new_AGEMA_signal_4201), .A1_f (new_AGEMA_signal_4202), .B0_t (StateFromRhoPi[186]), .B0_f (new_AGEMA_signal_3521), .B1_t (new_AGEMA_signal_3522), .B1_f (new_AGEMA_signal_3523), .Z0_t (StateFromChi[186]), .Z0_f (new_AGEMA_signal_4806), .Z1_t (new_AGEMA_signal_4807), .Z1_f (new_AGEMA_signal_4808) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_4__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[74]), .A0_f (new_AGEMA_signal_3980), .A1_t (new_AGEMA_signal_3981), .A1_f (new_AGEMA_signal_3982), .B0_t (StateFromRhoPi[114]), .B0_f (new_AGEMA_signal_3782), .B1_t (new_AGEMA_signal_3783), .B1_f (new_AGEMA_signal_3784), .Z0_t (CHI_GEN_SLICES_2__GEN_ROWS_4__sbox_and_xor_inst_a_nxy), .Z0_f (new_AGEMA_signal_4203), .Z1_t (new_AGEMA_signal_4204), .Z1_f (new_AGEMA_signal_4205) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_4__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_2__GEN_ROWS_4__sbox_and_xor_inst_a_nxy), .A0_f (new_AGEMA_signal_4203), .A1_t (new_AGEMA_signal_4204), .A1_f (new_AGEMA_signal_4205), .B0_t (StateFromRhoPi[34]), .B0_f (new_AGEMA_signal_3833), .B1_t (new_AGEMA_signal_3834), .B1_f (new_AGEMA_signal_3835), .Z0_t (StateFromChi[34]), .Z0_f (new_AGEMA_signal_4809), .Z1_t (new_AGEMA_signal_4810), .Z1_f (new_AGEMA_signal_4811) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_4__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[114]), .A0_f (new_AGEMA_signal_3782), .A1_t (new_AGEMA_signal_3783), .A1_f (new_AGEMA_signal_3784), .B0_t (StateFromRhoPi[154]), .B0_f (new_AGEMA_signal_3539), .B1_t (new_AGEMA_signal_3540), .B1_f (new_AGEMA_signal_3541), .Z0_t (CHI_GEN_SLICES_2__GEN_ROWS_4__sbox_and_xor_inst_b_nxy), .Z0_f (new_AGEMA_signal_4206), .Z1_t (new_AGEMA_signal_4207), .Z1_f (new_AGEMA_signal_4208) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_4__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_2__GEN_ROWS_4__sbox_and_xor_inst_b_nxy), .A0_f (new_AGEMA_signal_4206), .A1_t (new_AGEMA_signal_4207), .A1_f (new_AGEMA_signal_4208), .B0_t (StateFromRhoPi[74]), .B0_f (new_AGEMA_signal_3980), .B1_t (new_AGEMA_signal_3981), .B1_f (new_AGEMA_signal_3982), .Z0_t (StateFromChi[74]), .Z0_f (new_AGEMA_signal_4812), .Z1_t (new_AGEMA_signal_4813), .Z1_f (new_AGEMA_signal_4814) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_4__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[154]), .A0_f (new_AGEMA_signal_3539), .A1_t (new_AGEMA_signal_3540), .A1_f (new_AGEMA_signal_3541), .B0_t (StateFromRhoPi[194]), .B0_f (new_AGEMA_signal_3506), .B1_t (new_AGEMA_signal_3507), .B1_f (new_AGEMA_signal_3508), .Z0_t (CHI_GEN_SLICES_2__GEN_ROWS_4__sbox_and_xor_inst_c_nxy), .Z0_f (new_AGEMA_signal_4209), .Z1_t (new_AGEMA_signal_4210), .Z1_f (new_AGEMA_signal_4211) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_4__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_2__GEN_ROWS_4__sbox_and_xor_inst_c_nxy), .A0_f (new_AGEMA_signal_4209), .A1_t (new_AGEMA_signal_4210), .A1_f (new_AGEMA_signal_4211), .B0_t (StateFromRhoPi[114]), .B0_f (new_AGEMA_signal_3782), .B1_t (new_AGEMA_signal_3783), .B1_f (new_AGEMA_signal_3784), .Z0_t (StateFromChi[114]), .Z0_f (new_AGEMA_signal_4815), .Z1_t (new_AGEMA_signal_4816), .Z1_f (new_AGEMA_signal_4817) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_4__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[194]), .A0_f (new_AGEMA_signal_3506), .A1_t (new_AGEMA_signal_3507), .A1_f (new_AGEMA_signal_3508), .B0_t (StateFromRhoPi[34]), .B0_f (new_AGEMA_signal_3833), .B1_t (new_AGEMA_signal_3834), .B1_f (new_AGEMA_signal_3835), .Z0_t (CHI_GEN_SLICES_2__GEN_ROWS_4__sbox_and_xor_inst_d_nxy), .Z0_f (new_AGEMA_signal_4212), .Z1_t (new_AGEMA_signal_4213), .Z1_f (new_AGEMA_signal_4214) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_4__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_2__GEN_ROWS_4__sbox_and_xor_inst_d_nxy), .A0_f (new_AGEMA_signal_4212), .A1_t (new_AGEMA_signal_4213), .A1_f (new_AGEMA_signal_4214), .B0_t (StateFromRhoPi[154]), .B0_f (new_AGEMA_signal_3539), .B1_t (new_AGEMA_signal_3540), .B1_f (new_AGEMA_signal_3541), .Z0_t (StateFromChi[154]), .Z0_f (new_AGEMA_signal_4818), .Z1_t (new_AGEMA_signal_4819), .Z1_f (new_AGEMA_signal_4820) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_4__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[34]), .A0_f (new_AGEMA_signal_3833), .A1_t (new_AGEMA_signal_3834), .A1_f (new_AGEMA_signal_3835), .B0_t (StateFromRhoPi[74]), .B0_f (new_AGEMA_signal_3980), .B1_t (new_AGEMA_signal_3981), .B1_f (new_AGEMA_signal_3982), .Z0_t (CHI_GEN_SLICES_2__GEN_ROWS_4__sbox_and_xor_inst_e_nxy), .Z0_f (new_AGEMA_signal_4215), .Z1_t (new_AGEMA_signal_4216), .Z1_f (new_AGEMA_signal_4217) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_4__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_2__GEN_ROWS_4__sbox_and_xor_inst_e_nxy), .A0_f (new_AGEMA_signal_4215), .A1_t (new_AGEMA_signal_4216), .A1_f (new_AGEMA_signal_4217), .B0_t (StateFromRhoPi[194]), .B0_f (new_AGEMA_signal_3506), .B1_t (new_AGEMA_signal_3507), .B1_f (new_AGEMA_signal_3508), .Z0_t (StateFromChi[194]), .Z0_f (new_AGEMA_signal_4821), .Z1_t (new_AGEMA_signal_4822), .Z1_f (new_AGEMA_signal_4823) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_0__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[43]), .A0_f (new_AGEMA_signal_3635), .A1_t (new_AGEMA_signal_3636), .A1_f (new_AGEMA_signal_3637), .B0_t (StateFromRhoPi[83]), .B0_f (new_AGEMA_signal_3422), .B1_t (new_AGEMA_signal_3423), .B1_f (new_AGEMA_signal_3424), .Z0_t (CHI_GEN_SLICES_3__GEN_ROWS_0__sbox_and_xor_inst_a_nxy), .Z0_f (new_AGEMA_signal_4218), .Z1_t (new_AGEMA_signal_4219), .Z1_f (new_AGEMA_signal_4220) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_0__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_3__GEN_ROWS_0__sbox_and_xor_inst_a_nxy), .A0_f (new_AGEMA_signal_4218), .A1_t (new_AGEMA_signal_4219), .A1_f (new_AGEMA_signal_4220), .B0_t (StateFromRhoPi[3]), .B0_f (new_AGEMA_signal_3908), .B1_t (new_AGEMA_signal_3909), .B1_f (new_AGEMA_signal_3910), .Z0_t (CHI_ChiOut_3), .Z0_f (new_AGEMA_signal_4824), .Z1_t (new_AGEMA_signal_4825), .Z1_f (new_AGEMA_signal_4826) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_0__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[83]), .A0_f (new_AGEMA_signal_3422), .A1_t (new_AGEMA_signal_3423), .A1_f (new_AGEMA_signal_3424), .B0_t (StateFromRhoPi[123]), .B0_f (new_AGEMA_signal_3914), .B1_t (new_AGEMA_signal_3915), .B1_f (new_AGEMA_signal_3916), .Z0_t (CHI_GEN_SLICES_3__GEN_ROWS_0__sbox_and_xor_inst_b_nxy), .Z0_f (new_AGEMA_signal_4221), .Z1_t (new_AGEMA_signal_4222), .Z1_f (new_AGEMA_signal_4223) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_0__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_3__GEN_ROWS_0__sbox_and_xor_inst_b_nxy), .A0_f (new_AGEMA_signal_4221), .A1_t (new_AGEMA_signal_4222), .A1_f (new_AGEMA_signal_4223), .B0_t (StateFromRhoPi[43]), .B0_f (new_AGEMA_signal_3635), .B1_t (new_AGEMA_signal_3636), .B1_f (new_AGEMA_signal_3637), .Z0_t (StateFromChi[43]), .Z0_f (new_AGEMA_signal_4827), .Z1_t (new_AGEMA_signal_4828), .Z1_f (new_AGEMA_signal_4829) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_0__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[123]), .A0_f (new_AGEMA_signal_3914), .A1_t (new_AGEMA_signal_3915), .A1_f (new_AGEMA_signal_3916), .B0_t (StateFromRhoPi[163]), .B0_f (new_AGEMA_signal_3791), .B1_t (new_AGEMA_signal_3792), .B1_f (new_AGEMA_signal_3793), .Z0_t (CHI_GEN_SLICES_3__GEN_ROWS_0__sbox_and_xor_inst_c_nxy), .Z0_f (new_AGEMA_signal_4224), .Z1_t (new_AGEMA_signal_4225), .Z1_f (new_AGEMA_signal_4226) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_0__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_3__GEN_ROWS_0__sbox_and_xor_inst_c_nxy), .A0_f (new_AGEMA_signal_4224), .A1_t (new_AGEMA_signal_4225), .A1_f (new_AGEMA_signal_4226), .B0_t (StateFromRhoPi[83]), .B0_f (new_AGEMA_signal_3422), .B1_t (new_AGEMA_signal_3423), .B1_f (new_AGEMA_signal_3424), .Z0_t (StateFromChi[83]), .Z0_f (new_AGEMA_signal_4830), .Z1_t (new_AGEMA_signal_4831), .Z1_f (new_AGEMA_signal_4832) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_0__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[163]), .A0_f (new_AGEMA_signal_3791), .A1_t (new_AGEMA_signal_3792), .A1_f (new_AGEMA_signal_3793), .B0_t (StateFromRhoPi[3]), .B0_f (new_AGEMA_signal_3908), .B1_t (new_AGEMA_signal_3909), .B1_f (new_AGEMA_signal_3910), .Z0_t (CHI_GEN_SLICES_3__GEN_ROWS_0__sbox_and_xor_inst_d_nxy), .Z0_f (new_AGEMA_signal_4227), .Z1_t (new_AGEMA_signal_4228), .Z1_f (new_AGEMA_signal_4229) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_0__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_3__GEN_ROWS_0__sbox_and_xor_inst_d_nxy), .A0_f (new_AGEMA_signal_4227), .A1_t (new_AGEMA_signal_4228), .A1_f (new_AGEMA_signal_4229), .B0_t (StateFromRhoPi[123]), .B0_f (new_AGEMA_signal_3914), .B1_t (new_AGEMA_signal_3915), .B1_f (new_AGEMA_signal_3916), .Z0_t (StateFromChi[123]), .Z0_f (new_AGEMA_signal_4833), .Z1_t (new_AGEMA_signal_4834), .Z1_f (new_AGEMA_signal_4835) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_0__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[3]), .A0_f (new_AGEMA_signal_3908), .A1_t (new_AGEMA_signal_3909), .A1_f (new_AGEMA_signal_3910), .B0_t (StateFromRhoPi[43]), .B0_f (new_AGEMA_signal_3635), .B1_t (new_AGEMA_signal_3636), .B1_f (new_AGEMA_signal_3637), .Z0_t (CHI_GEN_SLICES_3__GEN_ROWS_0__sbox_and_xor_inst_e_nxy), .Z0_f (new_AGEMA_signal_4230), .Z1_t (new_AGEMA_signal_4231), .Z1_f (new_AGEMA_signal_4232) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_0__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_3__GEN_ROWS_0__sbox_and_xor_inst_e_nxy), .A0_f (new_AGEMA_signal_4230), .A1_t (new_AGEMA_signal_4231), .A1_f (new_AGEMA_signal_4232), .B0_t (StateFromRhoPi[163]), .B0_f (new_AGEMA_signal_3791), .B1_t (new_AGEMA_signal_3792), .B1_f (new_AGEMA_signal_3793), .Z0_t (StateFromChi[163]), .Z0_f (new_AGEMA_signal_4836), .Z1_t (new_AGEMA_signal_4837), .Z1_f (new_AGEMA_signal_4838) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_1__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[51]), .A0_f (new_AGEMA_signal_3395), .A1_t (new_AGEMA_signal_3396), .A1_f (new_AGEMA_signal_3397), .B0_t (StateFromRhoPi[91]), .B0_f (new_AGEMA_signal_3602), .B1_t (new_AGEMA_signal_3603), .B1_f (new_AGEMA_signal_3604), .Z0_t (CHI_GEN_SLICES_3__GEN_ROWS_1__sbox_and_xor_inst_a_nxy), .Z0_f (new_AGEMA_signal_4233), .Z1_t (new_AGEMA_signal_4234), .Z1_f (new_AGEMA_signal_4235) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_1__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_3__GEN_ROWS_1__sbox_and_xor_inst_a_nxy), .A0_f (new_AGEMA_signal_4233), .A1_t (new_AGEMA_signal_4234), .A1_f (new_AGEMA_signal_4235), .B0_t (StateFromRhoPi[11]), .B0_f (new_AGEMA_signal_3758), .B1_t (new_AGEMA_signal_3759), .B1_f (new_AGEMA_signal_3760), .Z0_t (StateFromChi[11]), .Z0_f (new_AGEMA_signal_4839), .Z1_t (new_AGEMA_signal_4840), .Z1_f (new_AGEMA_signal_4841) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_1__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[91]), .A0_f (new_AGEMA_signal_3602), .A1_t (new_AGEMA_signal_3603), .A1_f (new_AGEMA_signal_3604), .B0_t (StateFromRhoPi[131]), .B0_f (new_AGEMA_signal_3404), .B1_t (new_AGEMA_signal_3405), .B1_f (new_AGEMA_signal_3406), .Z0_t (CHI_GEN_SLICES_3__GEN_ROWS_1__sbox_and_xor_inst_b_nxy), .Z0_f (new_AGEMA_signal_4236), .Z1_t (new_AGEMA_signal_4237), .Z1_f (new_AGEMA_signal_4238) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_1__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_3__GEN_ROWS_1__sbox_and_xor_inst_b_nxy), .A0_f (new_AGEMA_signal_4236), .A1_t (new_AGEMA_signal_4237), .A1_f (new_AGEMA_signal_4238), .B0_t (StateFromRhoPi[51]), .B0_f (new_AGEMA_signal_3395), .B1_t (new_AGEMA_signal_3396), .B1_f (new_AGEMA_signal_3397), .Z0_t (StateFromChi[51]), .Z0_f (new_AGEMA_signal_4842), .Z1_t (new_AGEMA_signal_4843), .Z1_f (new_AGEMA_signal_4844) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_1__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[131]), .A0_f (new_AGEMA_signal_3404), .A1_t (new_AGEMA_signal_3405), .A1_f (new_AGEMA_signal_3406), .B0_t (StateFromRhoPi[171]), .B0_f (new_AGEMA_signal_3731), .B1_t (new_AGEMA_signal_3732), .B1_f (new_AGEMA_signal_3733), .Z0_t (CHI_GEN_SLICES_3__GEN_ROWS_1__sbox_and_xor_inst_c_nxy), .Z0_f (new_AGEMA_signal_4239), .Z1_t (new_AGEMA_signal_4240), .Z1_f (new_AGEMA_signal_4241) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_1__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_3__GEN_ROWS_1__sbox_and_xor_inst_c_nxy), .A0_f (new_AGEMA_signal_4239), .A1_t (new_AGEMA_signal_4240), .A1_f (new_AGEMA_signal_4241), .B0_t (StateFromRhoPi[91]), .B0_f (new_AGEMA_signal_3602), .B1_t (new_AGEMA_signal_3603), .B1_f (new_AGEMA_signal_3604), .Z0_t (StateFromChi[91]), .Z0_f (new_AGEMA_signal_4845), .Z1_t (new_AGEMA_signal_4846), .Z1_f (new_AGEMA_signal_4847) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_1__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[171]), .A0_f (new_AGEMA_signal_3731), .A1_t (new_AGEMA_signal_3732), .A1_f (new_AGEMA_signal_3733), .B0_t (StateFromRhoPi[11]), .B0_f (new_AGEMA_signal_3758), .B1_t (new_AGEMA_signal_3759), .B1_f (new_AGEMA_signal_3760), .Z0_t (CHI_GEN_SLICES_3__GEN_ROWS_1__sbox_and_xor_inst_d_nxy), .Z0_f (new_AGEMA_signal_4242), .Z1_t (new_AGEMA_signal_4243), .Z1_f (new_AGEMA_signal_4244) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_1__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_3__GEN_ROWS_1__sbox_and_xor_inst_d_nxy), .A0_f (new_AGEMA_signal_4242), .A1_t (new_AGEMA_signal_4243), .A1_f (new_AGEMA_signal_4244), .B0_t (StateFromRhoPi[131]), .B0_f (new_AGEMA_signal_3404), .B1_t (new_AGEMA_signal_3405), .B1_f (new_AGEMA_signal_3406), .Z0_t (StateFromChi[131]), .Z0_f (new_AGEMA_signal_4848), .Z1_t (new_AGEMA_signal_4849), .Z1_f (new_AGEMA_signal_4850) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_1__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[11]), .A0_f (new_AGEMA_signal_3758), .A1_t (new_AGEMA_signal_3759), .A1_f (new_AGEMA_signal_3760), .B0_t (StateFromRhoPi[51]), .B0_f (new_AGEMA_signal_3395), .B1_t (new_AGEMA_signal_3396), .B1_f (new_AGEMA_signal_3397), .Z0_t (CHI_GEN_SLICES_3__GEN_ROWS_1__sbox_and_xor_inst_e_nxy), .Z0_f (new_AGEMA_signal_4245), .Z1_t (new_AGEMA_signal_4246), .Z1_f (new_AGEMA_signal_4247) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_1__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_3__GEN_ROWS_1__sbox_and_xor_inst_e_nxy), .A0_f (new_AGEMA_signal_4245), .A1_t (new_AGEMA_signal_4246), .A1_f (new_AGEMA_signal_4247), .B0_t (StateFromRhoPi[171]), .B0_f (new_AGEMA_signal_3731), .B1_t (new_AGEMA_signal_3732), .B1_f (new_AGEMA_signal_3733), .Z0_t (StateFromChi[171]), .Z0_f (new_AGEMA_signal_4851), .Z1_t (new_AGEMA_signal_4852), .Z1_f (new_AGEMA_signal_4853) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_2__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[59]), .A0_f (new_AGEMA_signal_3650), .A1_t (new_AGEMA_signal_3651), .A1_f (new_AGEMA_signal_3652), .B0_t (StateFromRhoPi[99]), .B0_f (new_AGEMA_signal_3527), .B1_t (new_AGEMA_signal_3528), .B1_f (new_AGEMA_signal_3529), .Z0_t (CHI_GEN_SLICES_3__GEN_ROWS_2__sbox_and_xor_inst_a_nxy), .Z0_f (new_AGEMA_signal_4248), .Z1_t (new_AGEMA_signal_4249), .Z1_f (new_AGEMA_signal_4250) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_2__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_3__GEN_ROWS_2__sbox_and_xor_inst_a_nxy), .A0_f (new_AGEMA_signal_4248), .A1_t (new_AGEMA_signal_4249), .A1_f (new_AGEMA_signal_4250), .B0_t (StateFromRhoPi[19]), .B0_f (new_AGEMA_signal_3593), .B1_t (new_AGEMA_signal_3594), .B1_f (new_AGEMA_signal_3595), .Z0_t (StateFromChi[19]), .Z0_f (new_AGEMA_signal_4854), .Z1_t (new_AGEMA_signal_4855), .Z1_f (new_AGEMA_signal_4856) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_2__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[99]), .A0_f (new_AGEMA_signal_3527), .A1_t (new_AGEMA_signal_3528), .A1_f (new_AGEMA_signal_3529), .B0_t (StateFromRhoPi[139]), .B0_f (new_AGEMA_signal_3779), .B1_t (new_AGEMA_signal_3780), .B1_f (new_AGEMA_signal_3781), .Z0_t (CHI_GEN_SLICES_3__GEN_ROWS_2__sbox_and_xor_inst_b_nxy), .Z0_f (new_AGEMA_signal_4251), .Z1_t (new_AGEMA_signal_4252), .Z1_f (new_AGEMA_signal_4253) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_2__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_3__GEN_ROWS_2__sbox_and_xor_inst_b_nxy), .A0_f (new_AGEMA_signal_4251), .A1_t (new_AGEMA_signal_4252), .A1_f (new_AGEMA_signal_4253), .B0_t (StateFromRhoPi[59]), .B0_f (new_AGEMA_signal_3650), .B1_t (new_AGEMA_signal_3651), .B1_f (new_AGEMA_signal_3652), .Z0_t (StateFromChi[59]), .Z0_f (new_AGEMA_signal_4857), .Z1_t (new_AGEMA_signal_4858), .Z1_f (new_AGEMA_signal_4859) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_2__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[139]), .A0_f (new_AGEMA_signal_3779), .A1_t (new_AGEMA_signal_3780), .A1_f (new_AGEMA_signal_3781), .B0_t (StateFromRhoPi[179]), .B0_f (new_AGEMA_signal_3536), .B1_t (new_AGEMA_signal_3537), .B1_f (new_AGEMA_signal_3538), .Z0_t (CHI_GEN_SLICES_3__GEN_ROWS_2__sbox_and_xor_inst_c_nxy), .Z0_f (new_AGEMA_signal_4254), .Z1_t (new_AGEMA_signal_4255), .Z1_f (new_AGEMA_signal_4256) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_2__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_3__GEN_ROWS_2__sbox_and_xor_inst_c_nxy), .A0_f (new_AGEMA_signal_4254), .A1_t (new_AGEMA_signal_4255), .A1_f (new_AGEMA_signal_4256), .B0_t (StateFromRhoPi[99]), .B0_f (new_AGEMA_signal_3527), .B1_t (new_AGEMA_signal_3528), .B1_f (new_AGEMA_signal_3529), .Z0_t (StateFromChi[99]), .Z0_f (new_AGEMA_signal_4860), .Z1_t (new_AGEMA_signal_4861), .Z1_f (new_AGEMA_signal_4862) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_2__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[179]), .A0_f (new_AGEMA_signal_3536), .A1_t (new_AGEMA_signal_3537), .A1_f (new_AGEMA_signal_3538), .B0_t (StateFromRhoPi[19]), .B0_f (new_AGEMA_signal_3593), .B1_t (new_AGEMA_signal_3594), .B1_f (new_AGEMA_signal_3595), .Z0_t (CHI_GEN_SLICES_3__GEN_ROWS_2__sbox_and_xor_inst_d_nxy), .Z0_f (new_AGEMA_signal_4257), .Z1_t (new_AGEMA_signal_4258), .Z1_f (new_AGEMA_signal_4259) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_2__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_3__GEN_ROWS_2__sbox_and_xor_inst_d_nxy), .A0_f (new_AGEMA_signal_4257), .A1_t (new_AGEMA_signal_4258), .A1_f (new_AGEMA_signal_4259), .B0_t (StateFromRhoPi[139]), .B0_f (new_AGEMA_signal_3779), .B1_t (new_AGEMA_signal_3780), .B1_f (new_AGEMA_signal_3781), .Z0_t (StateFromChi[139]), .Z0_f (new_AGEMA_signal_4863), .Z1_t (new_AGEMA_signal_4864), .Z1_f (new_AGEMA_signal_4865) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_2__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[19]), .A0_f (new_AGEMA_signal_3593), .A1_t (new_AGEMA_signal_3594), .A1_f (new_AGEMA_signal_3595), .B0_t (StateFromRhoPi[59]), .B0_f (new_AGEMA_signal_3650), .B1_t (new_AGEMA_signal_3651), .B1_f (new_AGEMA_signal_3652), .Z0_t (CHI_GEN_SLICES_3__GEN_ROWS_2__sbox_and_xor_inst_e_nxy), .Z0_f (new_AGEMA_signal_4260), .Z1_t (new_AGEMA_signal_4261), .Z1_f (new_AGEMA_signal_4262) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_2__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_3__GEN_ROWS_2__sbox_and_xor_inst_e_nxy), .A0_f (new_AGEMA_signal_4260), .A1_t (new_AGEMA_signal_4261), .A1_f (new_AGEMA_signal_4262), .B0_t (StateFromRhoPi[179]), .B0_f (new_AGEMA_signal_3536), .B1_t (new_AGEMA_signal_3537), .B1_f (new_AGEMA_signal_3538), .Z0_t (StateFromChi[179]), .Z0_f (new_AGEMA_signal_4866), .Z1_t (new_AGEMA_signal_4867), .Z1_f (new_AGEMA_signal_4868) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_3__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[67]), .A0_f (new_AGEMA_signal_3725), .A1_t (new_AGEMA_signal_3726), .A1_f (new_AGEMA_signal_3727), .B0_t (StateFromRhoPi[107]), .B0_f (new_AGEMA_signal_3677), .B1_t (new_AGEMA_signal_3678), .B1_f (new_AGEMA_signal_3679), .Z0_t (CHI_GEN_SLICES_3__GEN_ROWS_3__sbox_and_xor_inst_a_nxy), .Z0_f (new_AGEMA_signal_4263), .Z1_t (new_AGEMA_signal_4264), .Z1_f (new_AGEMA_signal_4265) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_3__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_3__GEN_ROWS_3__sbox_and_xor_inst_a_nxy), .A0_f (new_AGEMA_signal_4263), .A1_t (new_AGEMA_signal_4264), .A1_f (new_AGEMA_signal_4265), .B0_t (StateFromRhoPi[27]), .B0_f (new_AGEMA_signal_3623), .B1_t (new_AGEMA_signal_3624), .B1_f (new_AGEMA_signal_3625), .Z0_t (StateFromChi[27]), .Z0_f (new_AGEMA_signal_4869), .Z1_t (new_AGEMA_signal_4870), .Z1_f (new_AGEMA_signal_4871) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_3__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[107]), .A0_f (new_AGEMA_signal_3677), .A1_t (new_AGEMA_signal_3678), .A1_f (new_AGEMA_signal_3679), .B0_t (StateFromRhoPi[147]), .B0_f (new_AGEMA_signal_3824), .B1_t (new_AGEMA_signal_3825), .B1_f (new_AGEMA_signal_3826), .Z0_t (CHI_GEN_SLICES_3__GEN_ROWS_3__sbox_and_xor_inst_b_nxy), .Z0_f (new_AGEMA_signal_4266), .Z1_t (new_AGEMA_signal_4267), .Z1_f (new_AGEMA_signal_4268) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_3__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_3__GEN_ROWS_3__sbox_and_xor_inst_b_nxy), .A0_f (new_AGEMA_signal_4266), .A1_t (new_AGEMA_signal_4267), .A1_f (new_AGEMA_signal_4268), .B0_t (StateFromRhoPi[67]), .B0_f (new_AGEMA_signal_3725), .B1_t (new_AGEMA_signal_3726), .B1_f (new_AGEMA_signal_3727), .Z0_t (StateFromChi[67]), .Z0_f (new_AGEMA_signal_4872), .Z1_t (new_AGEMA_signal_4873), .Z1_f (new_AGEMA_signal_4874) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_3__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[147]), .A0_f (new_AGEMA_signal_3824), .A1_t (new_AGEMA_signal_3825), .A1_f (new_AGEMA_signal_3826), .B0_t (StateFromRhoPi[187]), .B0_f (new_AGEMA_signal_3971), .B1_t (new_AGEMA_signal_3972), .B1_f (new_AGEMA_signal_3973), .Z0_t (CHI_GEN_SLICES_3__GEN_ROWS_3__sbox_and_xor_inst_c_nxy), .Z0_f (new_AGEMA_signal_4269), .Z1_t (new_AGEMA_signal_4270), .Z1_f (new_AGEMA_signal_4271) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_3__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_3__GEN_ROWS_3__sbox_and_xor_inst_c_nxy), .A0_f (new_AGEMA_signal_4269), .A1_t (new_AGEMA_signal_4270), .A1_f (new_AGEMA_signal_4271), .B0_t (StateFromRhoPi[107]), .B0_f (new_AGEMA_signal_3677), .B1_t (new_AGEMA_signal_3678), .B1_f (new_AGEMA_signal_3679), .Z0_t (StateFromChi[107]), .Z0_f (new_AGEMA_signal_4875), .Z1_t (new_AGEMA_signal_4876), .Z1_f (new_AGEMA_signal_4877) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_3__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[187]), .A0_f (new_AGEMA_signal_3971), .A1_t (new_AGEMA_signal_3972), .A1_f (new_AGEMA_signal_3973), .B0_t (StateFromRhoPi[27]), .B0_f (new_AGEMA_signal_3623), .B1_t (new_AGEMA_signal_3624), .B1_f (new_AGEMA_signal_3625), .Z0_t (CHI_GEN_SLICES_3__GEN_ROWS_3__sbox_and_xor_inst_d_nxy), .Z0_f (new_AGEMA_signal_4272), .Z1_t (new_AGEMA_signal_4273), .Z1_f (new_AGEMA_signal_4274) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_3__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_3__GEN_ROWS_3__sbox_and_xor_inst_d_nxy), .A0_f (new_AGEMA_signal_4272), .A1_t (new_AGEMA_signal_4273), .A1_f (new_AGEMA_signal_4274), .B0_t (StateFromRhoPi[147]), .B0_f (new_AGEMA_signal_3824), .B1_t (new_AGEMA_signal_3825), .B1_f (new_AGEMA_signal_3826), .Z0_t (StateFromChi[147]), .Z0_f (new_AGEMA_signal_4878), .Z1_t (new_AGEMA_signal_4879), .Z1_f (new_AGEMA_signal_4880) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_3__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[27]), .A0_f (new_AGEMA_signal_3623), .A1_t (new_AGEMA_signal_3624), .A1_f (new_AGEMA_signal_3625), .B0_t (StateFromRhoPi[67]), .B0_f (new_AGEMA_signal_3725), .B1_t (new_AGEMA_signal_3726), .B1_f (new_AGEMA_signal_3727), .Z0_t (CHI_GEN_SLICES_3__GEN_ROWS_3__sbox_and_xor_inst_e_nxy), .Z0_f (new_AGEMA_signal_4275), .Z1_t (new_AGEMA_signal_4276), .Z1_f (new_AGEMA_signal_4277) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_3__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_3__GEN_ROWS_3__sbox_and_xor_inst_e_nxy), .A0_f (new_AGEMA_signal_4275), .A1_t (new_AGEMA_signal_4276), .A1_f (new_AGEMA_signal_4277), .B0_t (StateFromRhoPi[187]), .B0_f (new_AGEMA_signal_3971), .B1_t (new_AGEMA_signal_3972), .B1_f (new_AGEMA_signal_3973), .Z0_t (StateFromChi[187]), .Z0_f (new_AGEMA_signal_4881), .Z1_t (new_AGEMA_signal_4882), .Z1_f (new_AGEMA_signal_4883) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_4__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[75]), .A0_f (new_AGEMA_signal_3965), .A1_t (new_AGEMA_signal_3966), .A1_f (new_AGEMA_signal_3967), .B0_t (StateFromRhoPi[115]), .B0_f (new_AGEMA_signal_3467), .B1_t (new_AGEMA_signal_3468), .B1_f (new_AGEMA_signal_3469), .Z0_t (CHI_GEN_SLICES_3__GEN_ROWS_4__sbox_and_xor_inst_a_nxy), .Z0_f (new_AGEMA_signal_4278), .Z1_t (new_AGEMA_signal_4279), .Z1_f (new_AGEMA_signal_4280) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_4__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_3__GEN_ROWS_4__sbox_and_xor_inst_a_nxy), .A0_f (new_AGEMA_signal_4278), .A1_t (new_AGEMA_signal_4279), .A1_f (new_AGEMA_signal_4280), .B0_t (StateFromRhoPi[35]), .B0_f (new_AGEMA_signal_3653), .B1_t (new_AGEMA_signal_3654), .B1_f (new_AGEMA_signal_3655), .Z0_t (StateFromChi[35]), .Z0_f (new_AGEMA_signal_4884), .Z1_t (new_AGEMA_signal_4885), .Z1_f (new_AGEMA_signal_4886) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_4__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[115]), .A0_f (new_AGEMA_signal_3467), .A1_t (new_AGEMA_signal_3468), .A1_f (new_AGEMA_signal_3469), .B0_t (StateFromRhoPi[155]), .B0_f (new_AGEMA_signal_3704), .B1_t (new_AGEMA_signal_3705), .B1_f (new_AGEMA_signal_3706), .Z0_t (CHI_GEN_SLICES_3__GEN_ROWS_4__sbox_and_xor_inst_b_nxy), .Z0_f (new_AGEMA_signal_4281), .Z1_t (new_AGEMA_signal_4282), .Z1_f (new_AGEMA_signal_4283) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_4__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_3__GEN_ROWS_4__sbox_and_xor_inst_b_nxy), .A0_f (new_AGEMA_signal_4281), .A1_t (new_AGEMA_signal_4282), .A1_f (new_AGEMA_signal_4283), .B0_t (StateFromRhoPi[75]), .B0_f (new_AGEMA_signal_3965), .B1_t (new_AGEMA_signal_3966), .B1_f (new_AGEMA_signal_3967), .Z0_t (StateFromChi[75]), .Z0_f (new_AGEMA_signal_4887), .Z1_t (new_AGEMA_signal_4888), .Z1_f (new_AGEMA_signal_4889) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_4__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[155]), .A0_f (new_AGEMA_signal_3704), .A1_t (new_AGEMA_signal_3705), .A1_f (new_AGEMA_signal_3706), .B0_t (StateFromRhoPi[195]), .B0_f (new_AGEMA_signal_3671), .B1_t (new_AGEMA_signal_3672), .B1_f (new_AGEMA_signal_3673), .Z0_t (CHI_GEN_SLICES_3__GEN_ROWS_4__sbox_and_xor_inst_c_nxy), .Z0_f (new_AGEMA_signal_4284), .Z1_t (new_AGEMA_signal_4285), .Z1_f (new_AGEMA_signal_4286) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_4__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_3__GEN_ROWS_4__sbox_and_xor_inst_c_nxy), .A0_f (new_AGEMA_signal_4284), .A1_t (new_AGEMA_signal_4285), .A1_f (new_AGEMA_signal_4286), .B0_t (StateFromRhoPi[115]), .B0_f (new_AGEMA_signal_3467), .B1_t (new_AGEMA_signal_3468), .B1_f (new_AGEMA_signal_3469), .Z0_t (StateFromChi[115]), .Z0_f (new_AGEMA_signal_4890), .Z1_t (new_AGEMA_signal_4891), .Z1_f (new_AGEMA_signal_4892) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_4__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[195]), .A0_f (new_AGEMA_signal_3671), .A1_t (new_AGEMA_signal_3672), .A1_f (new_AGEMA_signal_3673), .B0_t (StateFromRhoPi[35]), .B0_f (new_AGEMA_signal_3653), .B1_t (new_AGEMA_signal_3654), .B1_f (new_AGEMA_signal_3655), .Z0_t (CHI_GEN_SLICES_3__GEN_ROWS_4__sbox_and_xor_inst_d_nxy), .Z0_f (new_AGEMA_signal_4287), .Z1_t (new_AGEMA_signal_4288), .Z1_f (new_AGEMA_signal_4289) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_4__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_3__GEN_ROWS_4__sbox_and_xor_inst_d_nxy), .A0_f (new_AGEMA_signal_4287), .A1_t (new_AGEMA_signal_4288), .A1_f (new_AGEMA_signal_4289), .B0_t (StateFromRhoPi[155]), .B0_f (new_AGEMA_signal_3704), .B1_t (new_AGEMA_signal_3705), .B1_f (new_AGEMA_signal_3706), .Z0_t (StateFromChi[155]), .Z0_f (new_AGEMA_signal_4893), .Z1_t (new_AGEMA_signal_4894), .Z1_f (new_AGEMA_signal_4895) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_4__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[35]), .A0_f (new_AGEMA_signal_3653), .A1_t (new_AGEMA_signal_3654), .A1_f (new_AGEMA_signal_3655), .B0_t (StateFromRhoPi[75]), .B0_f (new_AGEMA_signal_3965), .B1_t (new_AGEMA_signal_3966), .B1_f (new_AGEMA_signal_3967), .Z0_t (CHI_GEN_SLICES_3__GEN_ROWS_4__sbox_and_xor_inst_e_nxy), .Z0_f (new_AGEMA_signal_4290), .Z1_t (new_AGEMA_signal_4291), .Z1_f (new_AGEMA_signal_4292) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_4__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_3__GEN_ROWS_4__sbox_and_xor_inst_e_nxy), .A0_f (new_AGEMA_signal_4290), .A1_t (new_AGEMA_signal_4291), .A1_f (new_AGEMA_signal_4292), .B0_t (StateFromRhoPi[195]), .B0_f (new_AGEMA_signal_3671), .B1_t (new_AGEMA_signal_3672), .B1_f (new_AGEMA_signal_3673), .Z0_t (StateFromChi[195]), .Z0_f (new_AGEMA_signal_4896), .Z1_t (new_AGEMA_signal_4897), .Z1_f (new_AGEMA_signal_4898) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_0__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[44]), .A0_f (new_AGEMA_signal_3515), .A1_t (new_AGEMA_signal_3516), .A1_f (new_AGEMA_signal_3517), .B0_t (StateFromRhoPi[84]), .B0_f (new_AGEMA_signal_3692), .B1_t (new_AGEMA_signal_3693), .B1_f (new_AGEMA_signal_3694), .Z0_t (CHI_GEN_SLICES_4__GEN_ROWS_0__sbox_and_xor_inst_a_nxy), .Z0_f (new_AGEMA_signal_4293), .Z1_t (new_AGEMA_signal_4294), .Z1_f (new_AGEMA_signal_4295) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_0__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_4__GEN_ROWS_0__sbox_and_xor_inst_a_nxy), .A0_f (new_AGEMA_signal_4293), .A1_t (new_AGEMA_signal_4294), .A1_f (new_AGEMA_signal_4295), .B0_t (StateFromRhoPi[4]), .B0_f (new_AGEMA_signal_3878), .B1_t (new_AGEMA_signal_3879), .B1_f (new_AGEMA_signal_3880), .Z0_t (StateFromChi[4]), .Z0_f (new_AGEMA_signal_4899), .Z1_t (new_AGEMA_signal_4900), .Z1_f (new_AGEMA_signal_4901) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_0__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[84]), .A0_f (new_AGEMA_signal_3692), .A1_t (new_AGEMA_signal_3693), .A1_f (new_AGEMA_signal_3694), .B0_t (StateFromRhoPi[124]), .B0_f (new_AGEMA_signal_3749), .B1_t (new_AGEMA_signal_3750), .B1_f (new_AGEMA_signal_3751), .Z0_t (CHI_GEN_SLICES_4__GEN_ROWS_0__sbox_and_xor_inst_b_nxy), .Z0_f (new_AGEMA_signal_4296), .Z1_t (new_AGEMA_signal_4297), .Z1_f (new_AGEMA_signal_4298) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_0__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_4__GEN_ROWS_0__sbox_and_xor_inst_b_nxy), .A0_f (new_AGEMA_signal_4296), .A1_t (new_AGEMA_signal_4297), .A1_f (new_AGEMA_signal_4298), .B0_t (StateFromRhoPi[44]), .B0_f (new_AGEMA_signal_3515), .B1_t (new_AGEMA_signal_3516), .B1_f (new_AGEMA_signal_3517), .Z0_t (StateFromChi[44]), .Z0_f (new_AGEMA_signal_4902), .Z1_t (new_AGEMA_signal_4903), .Z1_f (new_AGEMA_signal_4904) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_0__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[124]), .A0_f (new_AGEMA_signal_3749), .A1_t (new_AGEMA_signal_3750), .A1_f (new_AGEMA_signal_3751), .B0_t (StateFromRhoPi[164]), .B0_f (new_AGEMA_signal_3431), .B1_t (new_AGEMA_signal_3432), .B1_f (new_AGEMA_signal_3433), .Z0_t (CHI_GEN_SLICES_4__GEN_ROWS_0__sbox_and_xor_inst_c_nxy), .Z0_f (new_AGEMA_signal_4299), .Z1_t (new_AGEMA_signal_4300), .Z1_f (new_AGEMA_signal_4301) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_0__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_4__GEN_ROWS_0__sbox_and_xor_inst_c_nxy), .A0_f (new_AGEMA_signal_4299), .A1_t (new_AGEMA_signal_4300), .A1_f (new_AGEMA_signal_4301), .B0_t (StateFromRhoPi[84]), .B0_f (new_AGEMA_signal_3692), .B1_t (new_AGEMA_signal_3693), .B1_f (new_AGEMA_signal_3694), .Z0_t (StateFromChi[84]), .Z0_f (new_AGEMA_signal_4905), .Z1_t (new_AGEMA_signal_4906), .Z1_f (new_AGEMA_signal_4907) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_0__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[164]), .A0_f (new_AGEMA_signal_3431), .A1_t (new_AGEMA_signal_3432), .A1_f (new_AGEMA_signal_3433), .B0_t (StateFromRhoPi[4]), .B0_f (new_AGEMA_signal_3878), .B1_t (new_AGEMA_signal_3879), .B1_f (new_AGEMA_signal_3880), .Z0_t (CHI_GEN_SLICES_4__GEN_ROWS_0__sbox_and_xor_inst_d_nxy), .Z0_f (new_AGEMA_signal_4302), .Z1_t (new_AGEMA_signal_4303), .Z1_f (new_AGEMA_signal_4304) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_0__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_4__GEN_ROWS_0__sbox_and_xor_inst_d_nxy), .A0_f (new_AGEMA_signal_4302), .A1_t (new_AGEMA_signal_4303), .A1_f (new_AGEMA_signal_4304), .B0_t (StateFromRhoPi[124]), .B0_f (new_AGEMA_signal_3749), .B1_t (new_AGEMA_signal_3750), .B1_f (new_AGEMA_signal_3751), .Z0_t (StateFromChi[124]), .Z0_f (new_AGEMA_signal_4908), .Z1_t (new_AGEMA_signal_4909), .Z1_f (new_AGEMA_signal_4910) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_0__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[4]), .A0_f (new_AGEMA_signal_3878), .A1_t (new_AGEMA_signal_3879), .A1_f (new_AGEMA_signal_3880), .B0_t (StateFromRhoPi[44]), .B0_f (new_AGEMA_signal_3515), .B1_t (new_AGEMA_signal_3516), .B1_f (new_AGEMA_signal_3517), .Z0_t (CHI_GEN_SLICES_4__GEN_ROWS_0__sbox_and_xor_inst_e_nxy), .Z0_f (new_AGEMA_signal_4305), .Z1_t (new_AGEMA_signal_4306), .Z1_f (new_AGEMA_signal_4307) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_0__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_4__GEN_ROWS_0__sbox_and_xor_inst_e_nxy), .A0_f (new_AGEMA_signal_4305), .A1_t (new_AGEMA_signal_4306), .A1_f (new_AGEMA_signal_4307), .B0_t (StateFromRhoPi[164]), .B0_f (new_AGEMA_signal_3431), .B1_t (new_AGEMA_signal_3432), .B1_f (new_AGEMA_signal_3433), .Z0_t (StateFromChi[164]), .Z0_f (new_AGEMA_signal_4911), .Z1_t (new_AGEMA_signal_4912), .Z1_f (new_AGEMA_signal_4913) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_1__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[52]), .A0_f (new_AGEMA_signal_3620), .A1_t (new_AGEMA_signal_3621), .A1_f (new_AGEMA_signal_3622), .B0_t (StateFromRhoPi[92]), .B0_f (new_AGEMA_signal_3542), .B1_t (new_AGEMA_signal_3543), .B1_f (new_AGEMA_signal_3544), .Z0_t (CHI_GEN_SLICES_4__GEN_ROWS_1__sbox_and_xor_inst_a_nxy), .Z0_f (new_AGEMA_signal_4308), .Z1_t (new_AGEMA_signal_4309), .Z1_f (new_AGEMA_signal_4310) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_1__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_4__GEN_ROWS_1__sbox_and_xor_inst_a_nxy), .A0_f (new_AGEMA_signal_4308), .A1_t (new_AGEMA_signal_4309), .A1_f (new_AGEMA_signal_4310), .B0_t (StateFromRhoPi[12]), .B0_f (new_AGEMA_signal_3668), .B1_t (new_AGEMA_signal_3669), .B1_f (new_AGEMA_signal_3670), .Z0_t (StateFromChi[12]), .Z0_f (new_AGEMA_signal_4914), .Z1_t (new_AGEMA_signal_4915), .Z1_f (new_AGEMA_signal_4916) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_1__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[92]), .A0_f (new_AGEMA_signal_3542), .A1_t (new_AGEMA_signal_3543), .A1_f (new_AGEMA_signal_3544), .B0_t (StateFromRhoPi[132]), .B0_f (new_AGEMA_signal_3629), .B1_t (new_AGEMA_signal_3630), .B1_f (new_AGEMA_signal_3631), .Z0_t (CHI_GEN_SLICES_4__GEN_ROWS_1__sbox_and_xor_inst_b_nxy), .Z0_f (new_AGEMA_signal_4311), .Z1_t (new_AGEMA_signal_4312), .Z1_f (new_AGEMA_signal_4313) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_1__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_4__GEN_ROWS_1__sbox_and_xor_inst_b_nxy), .A0_f (new_AGEMA_signal_4311), .A1_t (new_AGEMA_signal_4312), .A1_f (new_AGEMA_signal_4313), .B0_t (StateFromRhoPi[52]), .B0_f (new_AGEMA_signal_3620), .B1_t (new_AGEMA_signal_3621), .B1_f (new_AGEMA_signal_3622), .Z0_t (StateFromChi[52]), .Z0_f (new_AGEMA_signal_4917), .Z1_t (new_AGEMA_signal_4918), .Z1_f (new_AGEMA_signal_4919) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_1__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[132]), .A0_f (new_AGEMA_signal_3629), .A1_t (new_AGEMA_signal_3630), .A1_f (new_AGEMA_signal_3631), .B0_t (StateFromRhoPi[172]), .B0_f (new_AGEMA_signal_3446), .B1_t (new_AGEMA_signal_3447), .B1_f (new_AGEMA_signal_3448), .Z0_t (CHI_GEN_SLICES_4__GEN_ROWS_1__sbox_and_xor_inst_c_nxy), .Z0_f (new_AGEMA_signal_4314), .Z1_t (new_AGEMA_signal_4315), .Z1_f (new_AGEMA_signal_4316) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_1__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_4__GEN_ROWS_1__sbox_and_xor_inst_c_nxy), .A0_f (new_AGEMA_signal_4314), .A1_t (new_AGEMA_signal_4315), .A1_f (new_AGEMA_signal_4316), .B0_t (StateFromRhoPi[92]), .B0_f (new_AGEMA_signal_3542), .B1_t (new_AGEMA_signal_3543), .B1_f (new_AGEMA_signal_3544), .Z0_t (StateFromChi[92]), .Z0_f (new_AGEMA_signal_4920), .Z1_t (new_AGEMA_signal_4921), .Z1_f (new_AGEMA_signal_4922) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_1__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[172]), .A0_f (new_AGEMA_signal_3446), .A1_t (new_AGEMA_signal_3447), .A1_f (new_AGEMA_signal_3448), .B0_t (StateFromRhoPi[12]), .B0_f (new_AGEMA_signal_3668), .B1_t (new_AGEMA_signal_3669), .B1_f (new_AGEMA_signal_3670), .Z0_t (CHI_GEN_SLICES_4__GEN_ROWS_1__sbox_and_xor_inst_d_nxy), .Z0_f (new_AGEMA_signal_4317), .Z1_t (new_AGEMA_signal_4318), .Z1_f (new_AGEMA_signal_4319) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_1__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_4__GEN_ROWS_1__sbox_and_xor_inst_d_nxy), .A0_f (new_AGEMA_signal_4317), .A1_t (new_AGEMA_signal_4318), .A1_f (new_AGEMA_signal_4319), .B0_t (StateFromRhoPi[132]), .B0_f (new_AGEMA_signal_3629), .B1_t (new_AGEMA_signal_3630), .B1_f (new_AGEMA_signal_3631), .Z0_t (StateFromChi[132]), .Z0_f (new_AGEMA_signal_4923), .Z1_t (new_AGEMA_signal_4924), .Z1_f (new_AGEMA_signal_4925) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_1__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[12]), .A0_f (new_AGEMA_signal_3668), .A1_t (new_AGEMA_signal_3669), .A1_f (new_AGEMA_signal_3670), .B0_t (StateFromRhoPi[52]), .B0_f (new_AGEMA_signal_3620), .B1_t (new_AGEMA_signal_3621), .B1_f (new_AGEMA_signal_3622), .Z0_t (CHI_GEN_SLICES_4__GEN_ROWS_1__sbox_and_xor_inst_e_nxy), .Z0_f (new_AGEMA_signal_4320), .Z1_t (new_AGEMA_signal_4321), .Z1_f (new_AGEMA_signal_4322) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_1__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_4__GEN_ROWS_1__sbox_and_xor_inst_e_nxy), .A0_f (new_AGEMA_signal_4320), .A1_t (new_AGEMA_signal_4321), .A1_f (new_AGEMA_signal_4322), .B0_t (StateFromRhoPi[172]), .B0_f (new_AGEMA_signal_3446), .B1_t (new_AGEMA_signal_3447), .B1_f (new_AGEMA_signal_3448), .Z0_t (StateFromChi[172]), .Z0_f (new_AGEMA_signal_4926), .Z1_t (new_AGEMA_signal_4927), .Z1_f (new_AGEMA_signal_4928) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_2__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[60]), .A0_f (new_AGEMA_signal_3740), .A1_t (new_AGEMA_signal_3741), .A1_f (new_AGEMA_signal_3742), .B0_t (StateFromRhoPi[100]), .B0_f (new_AGEMA_signal_3977), .B1_t (new_AGEMA_signal_3978), .B1_f (new_AGEMA_signal_3979), .Z0_t (CHI_GEN_SLICES_4__GEN_ROWS_2__sbox_and_xor_inst_a_nxy), .Z0_f (new_AGEMA_signal_4323), .Z1_t (new_AGEMA_signal_4324), .Z1_f (new_AGEMA_signal_4325) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_2__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_4__GEN_ROWS_2__sbox_and_xor_inst_a_nxy), .A0_f (new_AGEMA_signal_4323), .A1_t (new_AGEMA_signal_4324), .A1_f (new_AGEMA_signal_4325), .B0_t (StateFromRhoPi[20]), .B0_f (new_AGEMA_signal_3488), .B1_t (new_AGEMA_signal_3489), .B1_f (new_AGEMA_signal_3490), .Z0_t (StateFromChi[20]), .Z0_f (new_AGEMA_signal_4929), .Z1_t (new_AGEMA_signal_4930), .Z1_f (new_AGEMA_signal_4931) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_2__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[100]), .A0_f (new_AGEMA_signal_3977), .A1_t (new_AGEMA_signal_3978), .A1_f (new_AGEMA_signal_3979), .B0_t (StateFromRhoPi[140]), .B0_f (new_AGEMA_signal_3464), .B1_t (new_AGEMA_signal_3465), .B1_f (new_AGEMA_signal_3466), .Z0_t (CHI_GEN_SLICES_4__GEN_ROWS_2__sbox_and_xor_inst_b_nxy), .Z0_f (new_AGEMA_signal_4326), .Z1_t (new_AGEMA_signal_4327), .Z1_f (new_AGEMA_signal_4328) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_2__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_4__GEN_ROWS_2__sbox_and_xor_inst_b_nxy), .A0_f (new_AGEMA_signal_4326), .A1_t (new_AGEMA_signal_4327), .A1_f (new_AGEMA_signal_4328), .B0_t (StateFromRhoPi[60]), .B0_f (new_AGEMA_signal_3740), .B1_t (new_AGEMA_signal_3741), .B1_f (new_AGEMA_signal_3742), .Z0_t (StateFromChi[60]), .Z0_f (new_AGEMA_signal_4932), .Z1_t (new_AGEMA_signal_4933), .Z1_f (new_AGEMA_signal_4934) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_2__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[140]), .A0_f (new_AGEMA_signal_3464), .A1_t (new_AGEMA_signal_3465), .A1_f (new_AGEMA_signal_3466), .B0_t (StateFromRhoPi[180]), .B0_f (new_AGEMA_signal_3701), .B1_t (new_AGEMA_signal_3702), .B1_f (new_AGEMA_signal_3703), .Z0_t (CHI_GEN_SLICES_4__GEN_ROWS_2__sbox_and_xor_inst_c_nxy), .Z0_f (new_AGEMA_signal_4329), .Z1_t (new_AGEMA_signal_4330), .Z1_f (new_AGEMA_signal_4331) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_2__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_4__GEN_ROWS_2__sbox_and_xor_inst_c_nxy), .A0_f (new_AGEMA_signal_4329), .A1_t (new_AGEMA_signal_4330), .A1_f (new_AGEMA_signal_4331), .B0_t (StateFromRhoPi[100]), .B0_f (new_AGEMA_signal_3977), .B1_t (new_AGEMA_signal_3978), .B1_f (new_AGEMA_signal_3979), .Z0_t (StateFromChi[100]), .Z0_f (new_AGEMA_signal_4935), .Z1_t (new_AGEMA_signal_4936), .Z1_f (new_AGEMA_signal_4937) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_2__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[180]), .A0_f (new_AGEMA_signal_3701), .A1_t (new_AGEMA_signal_3702), .A1_f (new_AGEMA_signal_3703), .B0_t (StateFromRhoPi[20]), .B0_f (new_AGEMA_signal_3488), .B1_t (new_AGEMA_signal_3489), .B1_f (new_AGEMA_signal_3490), .Z0_t (CHI_GEN_SLICES_4__GEN_ROWS_2__sbox_and_xor_inst_d_nxy), .Z0_f (new_AGEMA_signal_4332), .Z1_t (new_AGEMA_signal_4333), .Z1_f (new_AGEMA_signal_4334) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_2__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_4__GEN_ROWS_2__sbox_and_xor_inst_d_nxy), .A0_f (new_AGEMA_signal_4332), .A1_t (new_AGEMA_signal_4333), .A1_f (new_AGEMA_signal_4334), .B0_t (StateFromRhoPi[140]), .B0_f (new_AGEMA_signal_3464), .B1_t (new_AGEMA_signal_3465), .B1_f (new_AGEMA_signal_3466), .Z0_t (StateFromChi[140]), .Z0_f (new_AGEMA_signal_4938), .Z1_t (new_AGEMA_signal_4939), .Z1_f (new_AGEMA_signal_4940) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_2__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[20]), .A0_f (new_AGEMA_signal_3488), .A1_t (new_AGEMA_signal_3489), .A1_f (new_AGEMA_signal_3490), .B0_t (StateFromRhoPi[60]), .B0_f (new_AGEMA_signal_3740), .B1_t (new_AGEMA_signal_3741), .B1_f (new_AGEMA_signal_3742), .Z0_t (CHI_GEN_SLICES_4__GEN_ROWS_2__sbox_and_xor_inst_e_nxy), .Z0_f (new_AGEMA_signal_4335), .Z1_t (new_AGEMA_signal_4336), .Z1_f (new_AGEMA_signal_4337) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_2__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_4__GEN_ROWS_2__sbox_and_xor_inst_e_nxy), .A0_f (new_AGEMA_signal_4335), .A1_t (new_AGEMA_signal_4336), .A1_f (new_AGEMA_signal_4337), .B0_t (StateFromRhoPi[180]), .B0_f (new_AGEMA_signal_3701), .B1_t (new_AGEMA_signal_3702), .B1_f (new_AGEMA_signal_3703), .Z0_t (StateFromChi[180]), .Z0_f (new_AGEMA_signal_4941), .Z1_t (new_AGEMA_signal_4942), .Z1_f (new_AGEMA_signal_4943) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_3__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[68]), .A0_f (new_AGEMA_signal_3605), .A1_t (new_AGEMA_signal_3606), .A1_f (new_AGEMA_signal_3607), .B0_t (StateFromRhoPi[108]), .B0_f (new_AGEMA_signal_3587), .B1_t (new_AGEMA_signal_3588), .B1_f (new_AGEMA_signal_3589), .Z0_t (CHI_GEN_SLICES_4__GEN_ROWS_3__sbox_and_xor_inst_a_nxy), .Z0_f (new_AGEMA_signal_4338), .Z1_t (new_AGEMA_signal_4339), .Z1_f (new_AGEMA_signal_4340) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_3__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_4__GEN_ROWS_3__sbox_and_xor_inst_a_nxy), .A0_f (new_AGEMA_signal_4338), .A1_t (new_AGEMA_signal_4339), .A1_f (new_AGEMA_signal_4340), .B0_t (StateFromRhoPi[28]), .B0_f (new_AGEMA_signal_3503), .B1_t (new_AGEMA_signal_3504), .B1_f (new_AGEMA_signal_3505), .Z0_t (StateFromChi[28]), .Z0_f (new_AGEMA_signal_4944), .Z1_t (new_AGEMA_signal_4945), .Z1_f (new_AGEMA_signal_4946) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_3__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[108]), .A0_f (new_AGEMA_signal_3587), .A1_t (new_AGEMA_signal_3588), .A1_f (new_AGEMA_signal_3589), .B0_t (StateFromRhoPi[148]), .B0_f (new_AGEMA_signal_3644), .B1_t (new_AGEMA_signal_3645), .B1_f (new_AGEMA_signal_3646), .Z0_t (CHI_GEN_SLICES_4__GEN_ROWS_3__sbox_and_xor_inst_b_nxy), .Z0_f (new_AGEMA_signal_4341), .Z1_t (new_AGEMA_signal_4342), .Z1_f (new_AGEMA_signal_4343) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_3__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_4__GEN_ROWS_3__sbox_and_xor_inst_b_nxy), .A0_f (new_AGEMA_signal_4341), .A1_t (new_AGEMA_signal_4342), .A1_f (new_AGEMA_signal_4343), .B0_t (StateFromRhoPi[68]), .B0_f (new_AGEMA_signal_3605), .B1_t (new_AGEMA_signal_3606), .B1_f (new_AGEMA_signal_3607), .Z0_t (StateFromChi[68]), .Z0_f (new_AGEMA_signal_4947), .Z1_t (new_AGEMA_signal_4948), .Z1_f (new_AGEMA_signal_4949) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_3__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[148]), .A0_f (new_AGEMA_signal_3644), .A1_t (new_AGEMA_signal_3645), .A1_f (new_AGEMA_signal_3646), .B0_t (StateFromRhoPi[188]), .B0_f (new_AGEMA_signal_3956), .B1_t (new_AGEMA_signal_3957), .B1_f (new_AGEMA_signal_3958), .Z0_t (CHI_GEN_SLICES_4__GEN_ROWS_3__sbox_and_xor_inst_c_nxy), .Z0_f (new_AGEMA_signal_4344), .Z1_t (new_AGEMA_signal_4345), .Z1_f (new_AGEMA_signal_4346) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_3__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_4__GEN_ROWS_3__sbox_and_xor_inst_c_nxy), .A0_f (new_AGEMA_signal_4344), .A1_t (new_AGEMA_signal_4345), .A1_f (new_AGEMA_signal_4346), .B0_t (StateFromRhoPi[108]), .B0_f (new_AGEMA_signal_3587), .B1_t (new_AGEMA_signal_3588), .B1_f (new_AGEMA_signal_3589), .Z0_t (StateFromChi[108]), .Z0_f (new_AGEMA_signal_4950), .Z1_t (new_AGEMA_signal_4951), .Z1_f (new_AGEMA_signal_4952) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_3__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[188]), .A0_f (new_AGEMA_signal_3956), .A1_t (new_AGEMA_signal_3957), .A1_f (new_AGEMA_signal_3958), .B0_t (StateFromRhoPi[28]), .B0_f (new_AGEMA_signal_3503), .B1_t (new_AGEMA_signal_3504), .B1_f (new_AGEMA_signal_3505), .Z0_t (CHI_GEN_SLICES_4__GEN_ROWS_3__sbox_and_xor_inst_d_nxy), .Z0_f (new_AGEMA_signal_4347), .Z1_t (new_AGEMA_signal_4348), .Z1_f (new_AGEMA_signal_4349) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_3__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_4__GEN_ROWS_3__sbox_and_xor_inst_d_nxy), .A0_f (new_AGEMA_signal_4347), .A1_t (new_AGEMA_signal_4348), .A1_f (new_AGEMA_signal_4349), .B0_t (StateFromRhoPi[148]), .B0_f (new_AGEMA_signal_3644), .B1_t (new_AGEMA_signal_3645), .B1_f (new_AGEMA_signal_3646), .Z0_t (StateFromChi[148]), .Z0_f (new_AGEMA_signal_4953), .Z1_t (new_AGEMA_signal_4954), .Z1_f (new_AGEMA_signal_4955) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_3__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[28]), .A0_f (new_AGEMA_signal_3503), .A1_t (new_AGEMA_signal_3504), .A1_f (new_AGEMA_signal_3505), .B0_t (StateFromRhoPi[68]), .B0_f (new_AGEMA_signal_3605), .B1_t (new_AGEMA_signal_3606), .B1_f (new_AGEMA_signal_3607), .Z0_t (CHI_GEN_SLICES_4__GEN_ROWS_3__sbox_and_xor_inst_e_nxy), .Z0_f (new_AGEMA_signal_4350), .Z1_t (new_AGEMA_signal_4351), .Z1_f (new_AGEMA_signal_4352) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_3__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_4__GEN_ROWS_3__sbox_and_xor_inst_e_nxy), .A0_f (new_AGEMA_signal_4350), .A1_t (new_AGEMA_signal_4351), .A1_f (new_AGEMA_signal_4352), .B0_t (StateFromRhoPi[188]), .B0_f (new_AGEMA_signal_3956), .B1_t (new_AGEMA_signal_3957), .B1_f (new_AGEMA_signal_3958), .Z0_t (StateFromChi[188]), .Z0_f (new_AGEMA_signal_4956), .Z1_t (new_AGEMA_signal_4957), .Z1_f (new_AGEMA_signal_4958) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_4__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[76]), .A0_f (new_AGEMA_signal_3935), .A1_t (new_AGEMA_signal_3936), .A1_f (new_AGEMA_signal_3937), .B0_t (StateFromRhoPi[116]), .B0_f (new_AGEMA_signal_3797), .B1_t (new_AGEMA_signal_3798), .B1_f (new_AGEMA_signal_3799), .Z0_t (CHI_GEN_SLICES_4__GEN_ROWS_4__sbox_and_xor_inst_a_nxy), .Z0_f (new_AGEMA_signal_4353), .Z1_t (new_AGEMA_signal_4354), .Z1_f (new_AGEMA_signal_4355) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_4__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_4__GEN_ROWS_4__sbox_and_xor_inst_a_nxy), .A0_f (new_AGEMA_signal_4353), .A1_t (new_AGEMA_signal_4354), .A1_f (new_AGEMA_signal_4355), .B0_t (StateFromRhoPi[36]), .B0_f (new_AGEMA_signal_3743), .B1_t (new_AGEMA_signal_3744), .B1_f (new_AGEMA_signal_3745), .Z0_t (StateFromChi[36]), .Z0_f (new_AGEMA_signal_4959), .Z1_t (new_AGEMA_signal_4960), .Z1_f (new_AGEMA_signal_4961) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_4__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[116]), .A0_f (new_AGEMA_signal_3797), .A1_t (new_AGEMA_signal_3798), .A1_f (new_AGEMA_signal_3799), .B0_t (StateFromRhoPi[156]), .B0_f (new_AGEMA_signal_3899), .B1_t (new_AGEMA_signal_3900), .B1_f (new_AGEMA_signal_3901), .Z0_t (CHI_GEN_SLICES_4__GEN_ROWS_4__sbox_and_xor_inst_b_nxy), .Z0_f (new_AGEMA_signal_4356), .Z1_t (new_AGEMA_signal_4357), .Z1_f (new_AGEMA_signal_4358) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_4__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_4__GEN_ROWS_4__sbox_and_xor_inst_b_nxy), .A0_f (new_AGEMA_signal_4356), .A1_t (new_AGEMA_signal_4357), .A1_f (new_AGEMA_signal_4358), .B0_t (StateFromRhoPi[76]), .B0_f (new_AGEMA_signal_3935), .B1_t (new_AGEMA_signal_3936), .B1_f (new_AGEMA_signal_3937), .Z0_t (StateFromChi[76]), .Z0_f (new_AGEMA_signal_4962), .Z1_t (new_AGEMA_signal_4963), .Z1_f (new_AGEMA_signal_4964) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_4__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[156]), .A0_f (new_AGEMA_signal_3899), .A1_t (new_AGEMA_signal_3900), .A1_f (new_AGEMA_signal_3901), .B0_t (StateFromRhoPi[196]), .B0_f (new_AGEMA_signal_3581), .B1_t (new_AGEMA_signal_3582), .B1_f (new_AGEMA_signal_3583), .Z0_t (CHI_GEN_SLICES_4__GEN_ROWS_4__sbox_and_xor_inst_c_nxy), .Z0_f (new_AGEMA_signal_4359), .Z1_t (new_AGEMA_signal_4360), .Z1_f (new_AGEMA_signal_4361) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_4__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_4__GEN_ROWS_4__sbox_and_xor_inst_c_nxy), .A0_f (new_AGEMA_signal_4359), .A1_t (new_AGEMA_signal_4360), .A1_f (new_AGEMA_signal_4361), .B0_t (StateFromRhoPi[116]), .B0_f (new_AGEMA_signal_3797), .B1_t (new_AGEMA_signal_3798), .B1_f (new_AGEMA_signal_3799), .Z0_t (StateFromChi[116]), .Z0_f (new_AGEMA_signal_4965), .Z1_t (new_AGEMA_signal_4966), .Z1_f (new_AGEMA_signal_4967) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_4__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[196]), .A0_f (new_AGEMA_signal_3581), .A1_t (new_AGEMA_signal_3582), .A1_f (new_AGEMA_signal_3583), .B0_t (StateFromRhoPi[36]), .B0_f (new_AGEMA_signal_3743), .B1_t (new_AGEMA_signal_3744), .B1_f (new_AGEMA_signal_3745), .Z0_t (CHI_GEN_SLICES_4__GEN_ROWS_4__sbox_and_xor_inst_d_nxy), .Z0_f (new_AGEMA_signal_4362), .Z1_t (new_AGEMA_signal_4363), .Z1_f (new_AGEMA_signal_4364) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_4__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_4__GEN_ROWS_4__sbox_and_xor_inst_d_nxy), .A0_f (new_AGEMA_signal_4362), .A1_t (new_AGEMA_signal_4363), .A1_f (new_AGEMA_signal_4364), .B0_t (StateFromRhoPi[156]), .B0_f (new_AGEMA_signal_3899), .B1_t (new_AGEMA_signal_3900), .B1_f (new_AGEMA_signal_3901), .Z0_t (StateFromChi[156]), .Z0_f (new_AGEMA_signal_4968), .Z1_t (new_AGEMA_signal_4969), .Z1_f (new_AGEMA_signal_4970) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_4__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[36]), .A0_f (new_AGEMA_signal_3743), .A1_t (new_AGEMA_signal_3744), .A1_f (new_AGEMA_signal_3745), .B0_t (StateFromRhoPi[76]), .B0_f (new_AGEMA_signal_3935), .B1_t (new_AGEMA_signal_3936), .B1_f (new_AGEMA_signal_3937), .Z0_t (CHI_GEN_SLICES_4__GEN_ROWS_4__sbox_and_xor_inst_e_nxy), .Z0_f (new_AGEMA_signal_4365), .Z1_t (new_AGEMA_signal_4366), .Z1_f (new_AGEMA_signal_4367) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_4__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_4__GEN_ROWS_4__sbox_and_xor_inst_e_nxy), .A0_f (new_AGEMA_signal_4365), .A1_t (new_AGEMA_signal_4366), .A1_f (new_AGEMA_signal_4367), .B0_t (StateFromRhoPi[196]), .B0_f (new_AGEMA_signal_3581), .B1_t (new_AGEMA_signal_3582), .B1_f (new_AGEMA_signal_3583), .Z0_t (StateFromChi[196]), .Z0_f (new_AGEMA_signal_4971), .Z1_t (new_AGEMA_signal_4972), .Z1_f (new_AGEMA_signal_4973) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_0__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[45]), .A0_f (new_AGEMA_signal_3680), .A1_t (new_AGEMA_signal_3681), .A1_f (new_AGEMA_signal_3682), .B0_t (StateFromRhoPi[85]), .B0_f (new_AGEMA_signal_3557), .B1_t (new_AGEMA_signal_3558), .B1_f (new_AGEMA_signal_3559), .Z0_t (CHI_GEN_SLICES_5__GEN_ROWS_0__sbox_and_xor_inst_a_nxy), .Z0_f (new_AGEMA_signal_4368), .Z1_t (new_AGEMA_signal_4369), .Z1_f (new_AGEMA_signal_4370) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_0__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_5__GEN_ROWS_0__sbox_and_xor_inst_a_nxy), .A0_f (new_AGEMA_signal_4368), .A1_t (new_AGEMA_signal_4369), .A1_f (new_AGEMA_signal_4370), .B0_t (StateFromRhoPi[5]), .B0_f (new_AGEMA_signal_3848), .B1_t (new_AGEMA_signal_3849), .B1_f (new_AGEMA_signal_3850), .Z0_t (StateFromChi[5]), .Z0_f (new_AGEMA_signal_4974), .Z1_t (new_AGEMA_signal_4975), .Z1_f (new_AGEMA_signal_4976) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_0__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[85]), .A0_f (new_AGEMA_signal_3557), .A1_t (new_AGEMA_signal_3558), .A1_f (new_AGEMA_signal_3559), .B0_t (StateFromRhoPi[125]), .B0_f (new_AGEMA_signal_3659), .B1_t (new_AGEMA_signal_3660), .B1_f (new_AGEMA_signal_3661), .Z0_t (CHI_GEN_SLICES_5__GEN_ROWS_0__sbox_and_xor_inst_b_nxy), .Z0_f (new_AGEMA_signal_4371), .Z1_t (new_AGEMA_signal_4372), .Z1_f (new_AGEMA_signal_4373) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_0__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_5__GEN_ROWS_0__sbox_and_xor_inst_b_nxy), .A0_f (new_AGEMA_signal_4371), .A1_t (new_AGEMA_signal_4372), .A1_f (new_AGEMA_signal_4373), .B0_t (StateFromRhoPi[45]), .B0_f (new_AGEMA_signal_3680), .B1_t (new_AGEMA_signal_3681), .B1_f (new_AGEMA_signal_3682), .Z0_t (StateFromChi[45]), .Z0_f (new_AGEMA_signal_4977), .Z1_t (new_AGEMA_signal_4978), .Z1_f (new_AGEMA_signal_4979) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_0__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[125]), .A0_f (new_AGEMA_signal_3659), .A1_t (new_AGEMA_signal_3660), .A1_f (new_AGEMA_signal_3661), .B0_t (StateFromRhoPi[165]), .B0_f (new_AGEMA_signal_3386), .B1_t (new_AGEMA_signal_3387), .B1_f (new_AGEMA_signal_3388), .Z0_t (CHI_GEN_SLICES_5__GEN_ROWS_0__sbox_and_xor_inst_c_nxy), .Z0_f (new_AGEMA_signal_4374), .Z1_t (new_AGEMA_signal_4375), .Z1_f (new_AGEMA_signal_4376) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_0__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_5__GEN_ROWS_0__sbox_and_xor_inst_c_nxy), .A0_f (new_AGEMA_signal_4374), .A1_t (new_AGEMA_signal_4375), .A1_f (new_AGEMA_signal_4376), .B0_t (StateFromRhoPi[85]), .B0_f (new_AGEMA_signal_3557), .B1_t (new_AGEMA_signal_3558), .B1_f (new_AGEMA_signal_3559), .Z0_t (StateFromChi[85]), .Z0_f (new_AGEMA_signal_4980), .Z1_t (new_AGEMA_signal_4981), .Z1_f (new_AGEMA_signal_4982) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_0__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[165]), .A0_f (new_AGEMA_signal_3386), .A1_t (new_AGEMA_signal_3387), .A1_f (new_AGEMA_signal_3388), .B0_t (StateFromRhoPi[5]), .B0_f (new_AGEMA_signal_3848), .B1_t (new_AGEMA_signal_3849), .B1_f (new_AGEMA_signal_3850), .Z0_t (CHI_GEN_SLICES_5__GEN_ROWS_0__sbox_and_xor_inst_d_nxy), .Z0_f (new_AGEMA_signal_4377), .Z1_t (new_AGEMA_signal_4378), .Z1_f (new_AGEMA_signal_4379) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_0__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_5__GEN_ROWS_0__sbox_and_xor_inst_d_nxy), .A0_f (new_AGEMA_signal_4377), .A1_t (new_AGEMA_signal_4378), .A1_f (new_AGEMA_signal_4379), .B0_t (StateFromRhoPi[125]), .B0_f (new_AGEMA_signal_3659), .B1_t (new_AGEMA_signal_3660), .B1_f (new_AGEMA_signal_3661), .Z0_t (StateFromChi[125]), .Z0_f (new_AGEMA_signal_4983), .Z1_t (new_AGEMA_signal_4984), .Z1_f (new_AGEMA_signal_4985) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_0__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[5]), .A0_f (new_AGEMA_signal_3848), .A1_t (new_AGEMA_signal_3849), .A1_f (new_AGEMA_signal_3850), .B0_t (StateFromRhoPi[45]), .B0_f (new_AGEMA_signal_3680), .B1_t (new_AGEMA_signal_3681), .B1_f (new_AGEMA_signal_3682), .Z0_t (CHI_GEN_SLICES_5__GEN_ROWS_0__sbox_and_xor_inst_e_nxy), .Z0_f (new_AGEMA_signal_4380), .Z1_t (new_AGEMA_signal_4381), .Z1_f (new_AGEMA_signal_4382) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_0__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_5__GEN_ROWS_0__sbox_and_xor_inst_e_nxy), .A0_f (new_AGEMA_signal_4380), .A1_t (new_AGEMA_signal_4381), .A1_f (new_AGEMA_signal_4382), .B0_t (StateFromRhoPi[165]), .B0_f (new_AGEMA_signal_3386), .B1_t (new_AGEMA_signal_3387), .B1_f (new_AGEMA_signal_3388), .Z0_t (StateFromChi[165]), .Z0_f (new_AGEMA_signal_4986), .Z1_t (new_AGEMA_signal_4987), .Z1_f (new_AGEMA_signal_4988) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_1__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[53]), .A0_f (new_AGEMA_signal_3500), .A1_t (new_AGEMA_signal_3501), .A1_f (new_AGEMA_signal_3502), .B0_t (StateFromRhoPi[93]), .B0_f (new_AGEMA_signal_3707), .B1_t (new_AGEMA_signal_3708), .B1_f (new_AGEMA_signal_3709), .Z0_t (CHI_GEN_SLICES_5__GEN_ROWS_1__sbox_and_xor_inst_a_nxy), .Z0_f (new_AGEMA_signal_4383), .Z1_t (new_AGEMA_signal_4384), .Z1_f (new_AGEMA_signal_4385) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_1__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_5__GEN_ROWS_1__sbox_and_xor_inst_a_nxy), .A0_f (new_AGEMA_signal_4383), .A1_t (new_AGEMA_signal_4384), .A1_f (new_AGEMA_signal_4385), .B0_t (StateFromRhoPi[13]), .B0_f (new_AGEMA_signal_3578), .B1_t (new_AGEMA_signal_3579), .B1_f (new_AGEMA_signal_3580), .Z0_t (StateFromChi[13]), .Z0_f (new_AGEMA_signal_4989), .Z1_t (new_AGEMA_signal_4990), .Z1_f (new_AGEMA_signal_4991) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_1__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[93]), .A0_f (new_AGEMA_signal_3707), .A1_t (new_AGEMA_signal_3708), .A1_f (new_AGEMA_signal_3709), .B0_t (StateFromRhoPi[133]), .B0_f (new_AGEMA_signal_3509), .B1_t (new_AGEMA_signal_3510), .B1_f (new_AGEMA_signal_3511), .Z0_t (CHI_GEN_SLICES_5__GEN_ROWS_1__sbox_and_xor_inst_b_nxy), .Z0_f (new_AGEMA_signal_4386), .Z1_t (new_AGEMA_signal_4387), .Z1_f (new_AGEMA_signal_4388) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_1__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_5__GEN_ROWS_1__sbox_and_xor_inst_b_nxy), .A0_f (new_AGEMA_signal_4386), .A1_t (new_AGEMA_signal_4387), .A1_f (new_AGEMA_signal_4388), .B0_t (StateFromRhoPi[53]), .B0_f (new_AGEMA_signal_3500), .B1_t (new_AGEMA_signal_3501), .B1_f (new_AGEMA_signal_3502), .Z0_t (StateFromChi[53]), .Z0_f (new_AGEMA_signal_4992), .Z1_t (new_AGEMA_signal_4993), .Z1_f (new_AGEMA_signal_4994) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_1__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[133]), .A0_f (new_AGEMA_signal_3509), .A1_t (new_AGEMA_signal_3510), .A1_f (new_AGEMA_signal_3511), .B0_t (StateFromRhoPi[173]), .B0_f (new_AGEMA_signal_3416), .B1_t (new_AGEMA_signal_3417), .B1_f (new_AGEMA_signal_3418), .Z0_t (CHI_GEN_SLICES_5__GEN_ROWS_1__sbox_and_xor_inst_c_nxy), .Z0_f (new_AGEMA_signal_4389), .Z1_t (new_AGEMA_signal_4390), .Z1_f (new_AGEMA_signal_4391) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_1__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_5__GEN_ROWS_1__sbox_and_xor_inst_c_nxy), .A0_f (new_AGEMA_signal_4389), .A1_t (new_AGEMA_signal_4390), .A1_f (new_AGEMA_signal_4391), .B0_t (StateFromRhoPi[93]), .B0_f (new_AGEMA_signal_3707), .B1_t (new_AGEMA_signal_3708), .B1_f (new_AGEMA_signal_3709), .Z0_t (StateFromChi[93]), .Z0_f (new_AGEMA_signal_4995), .Z1_t (new_AGEMA_signal_4996), .Z1_f (new_AGEMA_signal_4997) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_1__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[173]), .A0_f (new_AGEMA_signal_3416), .A1_t (new_AGEMA_signal_3417), .A1_f (new_AGEMA_signal_3418), .B0_t (StateFromRhoPi[13]), .B0_f (new_AGEMA_signal_3578), .B1_t (new_AGEMA_signal_3579), .B1_f (new_AGEMA_signal_3580), .Z0_t (CHI_GEN_SLICES_5__GEN_ROWS_1__sbox_and_xor_inst_d_nxy), .Z0_f (new_AGEMA_signal_4392), .Z1_t (new_AGEMA_signal_4393), .Z1_f (new_AGEMA_signal_4394) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_1__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_5__GEN_ROWS_1__sbox_and_xor_inst_d_nxy), .A0_f (new_AGEMA_signal_4392), .A1_t (new_AGEMA_signal_4393), .A1_f (new_AGEMA_signal_4394), .B0_t (StateFromRhoPi[133]), .B0_f (new_AGEMA_signal_3509), .B1_t (new_AGEMA_signal_3510), .B1_f (new_AGEMA_signal_3511), .Z0_t (StateFromChi[133]), .Z0_f (new_AGEMA_signal_4998), .Z1_t (new_AGEMA_signal_4999), .Z1_f (new_AGEMA_signal_5000) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_1__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[13]), .A0_f (new_AGEMA_signal_3578), .A1_t (new_AGEMA_signal_3579), .A1_f (new_AGEMA_signal_3580), .B0_t (StateFromRhoPi[53]), .B0_f (new_AGEMA_signal_3500), .B1_t (new_AGEMA_signal_3501), .B1_f (new_AGEMA_signal_3502), .Z0_t (CHI_GEN_SLICES_5__GEN_ROWS_1__sbox_and_xor_inst_e_nxy), .Z0_f (new_AGEMA_signal_4395), .Z1_t (new_AGEMA_signal_4396), .Z1_f (new_AGEMA_signal_4397) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_1__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_5__GEN_ROWS_1__sbox_and_xor_inst_e_nxy), .A0_f (new_AGEMA_signal_4395), .A1_t (new_AGEMA_signal_4396), .A1_f (new_AGEMA_signal_4397), .B0_t (StateFromRhoPi[173]), .B0_f (new_AGEMA_signal_3416), .B1_t (new_AGEMA_signal_3417), .B1_f (new_AGEMA_signal_3418), .Z0_t (StateFromChi[173]), .Z0_f (new_AGEMA_signal_5001), .Z1_t (new_AGEMA_signal_5002), .Z1_f (new_AGEMA_signal_5003) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_2__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[61]), .A0_f (new_AGEMA_signal_3455), .A1_t (new_AGEMA_signal_3456), .A1_f (new_AGEMA_signal_3457), .B0_t (StateFromRhoPi[101]), .B0_f (new_AGEMA_signal_3962), .B1_t (new_AGEMA_signal_3963), .B1_f (new_AGEMA_signal_3964), .Z0_t (CHI_GEN_SLICES_5__GEN_ROWS_2__sbox_and_xor_inst_a_nxy), .Z0_f (new_AGEMA_signal_4398), .Z1_t (new_AGEMA_signal_4399), .Z1_f (new_AGEMA_signal_4400) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_2__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_5__GEN_ROWS_2__sbox_and_xor_inst_a_nxy), .A0_f (new_AGEMA_signal_4398), .A1_t (new_AGEMA_signal_4399), .A1_f (new_AGEMA_signal_4400), .B0_t (StateFromRhoPi[21]), .B0_f (new_AGEMA_signal_3818), .B1_t (new_AGEMA_signal_3819), .B1_f (new_AGEMA_signal_3820), .Z0_t (StateFromChi[21]), .Z0_f (new_AGEMA_signal_5004), .Z1_t (new_AGEMA_signal_5005), .Z1_f (new_AGEMA_signal_5006) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_2__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[101]), .A0_f (new_AGEMA_signal_3962), .A1_t (new_AGEMA_signal_3963), .A1_f (new_AGEMA_signal_3964), .B0_t (StateFromRhoPi[141]), .B0_f (new_AGEMA_signal_3794), .B1_t (new_AGEMA_signal_3795), .B1_f (new_AGEMA_signal_3796), .Z0_t (CHI_GEN_SLICES_5__GEN_ROWS_2__sbox_and_xor_inst_b_nxy), .Z0_f (new_AGEMA_signal_4401), .Z1_t (new_AGEMA_signal_4402), .Z1_f (new_AGEMA_signal_4403) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_2__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_5__GEN_ROWS_2__sbox_and_xor_inst_b_nxy), .A0_f (new_AGEMA_signal_4401), .A1_t (new_AGEMA_signal_4402), .A1_f (new_AGEMA_signal_4403), .B0_t (StateFromRhoPi[61]), .B0_f (new_AGEMA_signal_3455), .B1_t (new_AGEMA_signal_3456), .B1_f (new_AGEMA_signal_3457), .Z0_t (StateFromChi[61]), .Z0_f (new_AGEMA_signal_5007), .Z1_t (new_AGEMA_signal_5008), .Z1_f (new_AGEMA_signal_5009) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_2__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[141]), .A0_f (new_AGEMA_signal_3794), .A1_t (new_AGEMA_signal_3795), .A1_f (new_AGEMA_signal_3796), .B0_t (StateFromRhoPi[181]), .B0_f (new_AGEMA_signal_3896), .B1_t (new_AGEMA_signal_3897), .B1_f (new_AGEMA_signal_3898), .Z0_t (CHI_GEN_SLICES_5__GEN_ROWS_2__sbox_and_xor_inst_c_nxy), .Z0_f (new_AGEMA_signal_4404), .Z1_t (new_AGEMA_signal_4405), .Z1_f (new_AGEMA_signal_4406) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_2__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_5__GEN_ROWS_2__sbox_and_xor_inst_c_nxy), .A0_f (new_AGEMA_signal_4404), .A1_t (new_AGEMA_signal_4405), .A1_f (new_AGEMA_signal_4406), .B0_t (StateFromRhoPi[101]), .B0_f (new_AGEMA_signal_3962), .B1_t (new_AGEMA_signal_3963), .B1_f (new_AGEMA_signal_3964), .Z0_t (StateFromChi[101]), .Z0_f (new_AGEMA_signal_5010), .Z1_t (new_AGEMA_signal_5011), .Z1_f (new_AGEMA_signal_5012) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_2__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[181]), .A0_f (new_AGEMA_signal_3896), .A1_t (new_AGEMA_signal_3897), .A1_f (new_AGEMA_signal_3898), .B0_t (StateFromRhoPi[21]), .B0_f (new_AGEMA_signal_3818), .B1_t (new_AGEMA_signal_3819), .B1_f (new_AGEMA_signal_3820), .Z0_t (CHI_GEN_SLICES_5__GEN_ROWS_2__sbox_and_xor_inst_d_nxy), .Z0_f (new_AGEMA_signal_4407), .Z1_t (new_AGEMA_signal_4408), .Z1_f (new_AGEMA_signal_4409) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_2__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_5__GEN_ROWS_2__sbox_and_xor_inst_d_nxy), .A0_f (new_AGEMA_signal_4407), .A1_t (new_AGEMA_signal_4408), .A1_f (new_AGEMA_signal_4409), .B0_t (StateFromRhoPi[141]), .B0_f (new_AGEMA_signal_3794), .B1_t (new_AGEMA_signal_3795), .B1_f (new_AGEMA_signal_3796), .Z0_t (StateFromChi[141]), .Z0_f (new_AGEMA_signal_5013), .Z1_t (new_AGEMA_signal_5014), .Z1_f (new_AGEMA_signal_5015) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_2__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[21]), .A0_f (new_AGEMA_signal_3818), .A1_t (new_AGEMA_signal_3819), .A1_f (new_AGEMA_signal_3820), .B0_t (StateFromRhoPi[61]), .B0_f (new_AGEMA_signal_3455), .B1_t (new_AGEMA_signal_3456), .B1_f (new_AGEMA_signal_3457), .Z0_t (CHI_GEN_SLICES_5__GEN_ROWS_2__sbox_and_xor_inst_e_nxy), .Z0_f (new_AGEMA_signal_4410), .Z1_t (new_AGEMA_signal_4411), .Z1_f (new_AGEMA_signal_4412) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_2__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_5__GEN_ROWS_2__sbox_and_xor_inst_e_nxy), .A0_f (new_AGEMA_signal_4410), .A1_t (new_AGEMA_signal_4411), .A1_f (new_AGEMA_signal_4412), .B0_t (StateFromRhoPi[181]), .B0_f (new_AGEMA_signal_3896), .B1_t (new_AGEMA_signal_3897), .B1_f (new_AGEMA_signal_3898), .Z0_t (StateFromChi[181]), .Z0_f (new_AGEMA_signal_5016), .Z1_t (new_AGEMA_signal_5017), .Z1_f (new_AGEMA_signal_5018) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_3__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[69]), .A0_f (new_AGEMA_signal_3545), .A1_t (new_AGEMA_signal_3546), .A1_f (new_AGEMA_signal_3547), .B0_t (StateFromRhoPi[109]), .B0_f (new_AGEMA_signal_3482), .B1_t (new_AGEMA_signal_3483), .B1_f (new_AGEMA_signal_3484), .Z0_t (CHI_GEN_SLICES_5__GEN_ROWS_3__sbox_and_xor_inst_a_nxy), .Z0_f (new_AGEMA_signal_4413), .Z1_t (new_AGEMA_signal_4414), .Z1_f (new_AGEMA_signal_4415) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_3__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_5__GEN_ROWS_3__sbox_and_xor_inst_a_nxy), .A0_f (new_AGEMA_signal_4413), .A1_t (new_AGEMA_signal_4414), .A1_f (new_AGEMA_signal_4415), .B0_t (StateFromRhoPi[29]), .B0_f (new_AGEMA_signal_3953), .B1_t (new_AGEMA_signal_3954), .B1_f (new_AGEMA_signal_3955), .Z0_t (StateFromChi[29]), .Z0_f (new_AGEMA_signal_5019), .Z1_t (new_AGEMA_signal_5020), .Z1_f (new_AGEMA_signal_5021) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_3__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[109]), .A0_f (new_AGEMA_signal_3482), .A1_t (new_AGEMA_signal_3483), .A1_f (new_AGEMA_signal_3484), .B0_t (StateFromRhoPi[149]), .B0_f (new_AGEMA_signal_3734), .B1_t (new_AGEMA_signal_3735), .B1_f (new_AGEMA_signal_3736), .Z0_t (CHI_GEN_SLICES_5__GEN_ROWS_3__sbox_and_xor_inst_b_nxy), .Z0_f (new_AGEMA_signal_4416), .Z1_t (new_AGEMA_signal_4417), .Z1_f (new_AGEMA_signal_4418) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_3__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_5__GEN_ROWS_3__sbox_and_xor_inst_b_nxy), .A0_f (new_AGEMA_signal_4416), .A1_t (new_AGEMA_signal_4417), .A1_f (new_AGEMA_signal_4418), .B0_t (StateFromRhoPi[69]), .B0_f (new_AGEMA_signal_3545), .B1_t (new_AGEMA_signal_3546), .B1_f (new_AGEMA_signal_3547), .Z0_t (StateFromChi[69]), .Z0_f (new_AGEMA_signal_5022), .Z1_t (new_AGEMA_signal_5023), .Z1_f (new_AGEMA_signal_5024) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_3__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[149]), .A0_f (new_AGEMA_signal_3734), .A1_t (new_AGEMA_signal_3735), .A1_f (new_AGEMA_signal_3736), .B0_t (StateFromRhoPi[189]), .B0_f (new_AGEMA_signal_3926), .B1_t (new_AGEMA_signal_3927), .B1_f (new_AGEMA_signal_3928), .Z0_t (CHI_GEN_SLICES_5__GEN_ROWS_3__sbox_and_xor_inst_c_nxy), .Z0_f (new_AGEMA_signal_4419), .Z1_t (new_AGEMA_signal_4420), .Z1_f (new_AGEMA_signal_4421) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_3__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_5__GEN_ROWS_3__sbox_and_xor_inst_c_nxy), .A0_f (new_AGEMA_signal_4419), .A1_t (new_AGEMA_signal_4420), .A1_f (new_AGEMA_signal_4421), .B0_t (StateFromRhoPi[109]), .B0_f (new_AGEMA_signal_3482), .B1_t (new_AGEMA_signal_3483), .B1_f (new_AGEMA_signal_3484), .Z0_t (StateFromChi[109]), .Z0_f (new_AGEMA_signal_5025), .Z1_t (new_AGEMA_signal_5026), .Z1_f (new_AGEMA_signal_5027) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_3__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[189]), .A0_f (new_AGEMA_signal_3926), .A1_t (new_AGEMA_signal_3927), .A1_f (new_AGEMA_signal_3928), .B0_t (StateFromRhoPi[29]), .B0_f (new_AGEMA_signal_3953), .B1_t (new_AGEMA_signal_3954), .B1_f (new_AGEMA_signal_3955), .Z0_t (CHI_GEN_SLICES_5__GEN_ROWS_3__sbox_and_xor_inst_d_nxy), .Z0_f (new_AGEMA_signal_4422), .Z1_t (new_AGEMA_signal_4423), .Z1_f (new_AGEMA_signal_4424) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_3__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_5__GEN_ROWS_3__sbox_and_xor_inst_d_nxy), .A0_f (new_AGEMA_signal_4422), .A1_t (new_AGEMA_signal_4423), .A1_f (new_AGEMA_signal_4424), .B0_t (StateFromRhoPi[149]), .B0_f (new_AGEMA_signal_3734), .B1_t (new_AGEMA_signal_3735), .B1_f (new_AGEMA_signal_3736), .Z0_t (StateFromChi[149]), .Z0_f (new_AGEMA_signal_5028), .Z1_t (new_AGEMA_signal_5029), .Z1_f (new_AGEMA_signal_5030) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_3__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[29]), .A0_f (new_AGEMA_signal_3953), .A1_t (new_AGEMA_signal_3954), .A1_f (new_AGEMA_signal_3955), .B0_t (StateFromRhoPi[69]), .B0_f (new_AGEMA_signal_3545), .B1_t (new_AGEMA_signal_3546), .B1_f (new_AGEMA_signal_3547), .Z0_t (CHI_GEN_SLICES_5__GEN_ROWS_3__sbox_and_xor_inst_e_nxy), .Z0_f (new_AGEMA_signal_4425), .Z1_t (new_AGEMA_signal_4426), .Z1_f (new_AGEMA_signal_4427) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_3__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_5__GEN_ROWS_3__sbox_and_xor_inst_e_nxy), .A0_f (new_AGEMA_signal_4425), .A1_t (new_AGEMA_signal_4426), .A1_f (new_AGEMA_signal_4427), .B0_t (StateFromRhoPi[189]), .B0_f (new_AGEMA_signal_3926), .B1_t (new_AGEMA_signal_3927), .B1_f (new_AGEMA_signal_3928), .Z0_t (StateFromChi[189]), .Z0_f (new_AGEMA_signal_5031), .Z1_t (new_AGEMA_signal_5032), .Z1_f (new_AGEMA_signal_5033) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_4__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[77]), .A0_f (new_AGEMA_signal_3920), .A1_t (new_AGEMA_signal_3921), .A1_f (new_AGEMA_signal_3922), .B0_t (StateFromRhoPi[117]), .B0_f (new_AGEMA_signal_3437), .B1_t (new_AGEMA_signal_3438), .B1_f (new_AGEMA_signal_3439), .Z0_t (CHI_GEN_SLICES_5__GEN_ROWS_4__sbox_and_xor_inst_a_nxy), .Z0_f (new_AGEMA_signal_4428), .Z1_t (new_AGEMA_signal_4429), .Z1_f (new_AGEMA_signal_4430) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_4__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_5__GEN_ROWS_4__sbox_and_xor_inst_a_nxy), .A0_f (new_AGEMA_signal_4428), .A1_t (new_AGEMA_signal_4429), .A1_f (new_AGEMA_signal_4430), .B0_t (StateFromRhoPi[37]), .B0_f (new_AGEMA_signal_3458), .B1_t (new_AGEMA_signal_3459), .B1_f (new_AGEMA_signal_3460), .Z0_t (StateFromChi[37]), .Z0_f (new_AGEMA_signal_5034), .Z1_t (new_AGEMA_signal_5035), .Z1_f (new_AGEMA_signal_5036) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_4__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[117]), .A0_f (new_AGEMA_signal_3437), .A1_t (new_AGEMA_signal_3438), .A1_f (new_AGEMA_signal_3439), .B0_t (StateFromRhoPi[157]), .B0_f (new_AGEMA_signal_3869), .B1_t (new_AGEMA_signal_3870), .B1_f (new_AGEMA_signal_3871), .Z0_t (CHI_GEN_SLICES_5__GEN_ROWS_4__sbox_and_xor_inst_b_nxy), .Z0_f (new_AGEMA_signal_4431), .Z1_t (new_AGEMA_signal_4432), .Z1_f (new_AGEMA_signal_4433) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_4__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_5__GEN_ROWS_4__sbox_and_xor_inst_b_nxy), .A0_f (new_AGEMA_signal_4431), .A1_t (new_AGEMA_signal_4432), .A1_f (new_AGEMA_signal_4433), .B0_t (StateFromRhoPi[77]), .B0_f (new_AGEMA_signal_3920), .B1_t (new_AGEMA_signal_3921), .B1_f (new_AGEMA_signal_3922), .Z0_t (StateFromChi[77]), .Z0_f (new_AGEMA_signal_5037), .Z1_t (new_AGEMA_signal_5038), .Z1_f (new_AGEMA_signal_5039) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_4__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[157]), .A0_f (new_AGEMA_signal_3869), .A1_t (new_AGEMA_signal_3870), .A1_f (new_AGEMA_signal_3871), .B0_t (StateFromRhoPi[197]), .B0_f (new_AGEMA_signal_3476), .B1_t (new_AGEMA_signal_3477), .B1_f (new_AGEMA_signal_3478), .Z0_t (CHI_GEN_SLICES_5__GEN_ROWS_4__sbox_and_xor_inst_c_nxy), .Z0_f (new_AGEMA_signal_4434), .Z1_t (new_AGEMA_signal_4435), .Z1_f (new_AGEMA_signal_4436) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_4__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_5__GEN_ROWS_4__sbox_and_xor_inst_c_nxy), .A0_f (new_AGEMA_signal_4434), .A1_t (new_AGEMA_signal_4435), .A1_f (new_AGEMA_signal_4436), .B0_t (StateFromRhoPi[117]), .B0_f (new_AGEMA_signal_3437), .B1_t (new_AGEMA_signal_3438), .B1_f (new_AGEMA_signal_3439), .Z0_t (StateFromChi[117]), .Z0_f (new_AGEMA_signal_5040), .Z1_t (new_AGEMA_signal_5041), .Z1_f (new_AGEMA_signal_5042) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_4__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[197]), .A0_f (new_AGEMA_signal_3476), .A1_t (new_AGEMA_signal_3477), .A1_f (new_AGEMA_signal_3478), .B0_t (StateFromRhoPi[37]), .B0_f (new_AGEMA_signal_3458), .B1_t (new_AGEMA_signal_3459), .B1_f (new_AGEMA_signal_3460), .Z0_t (CHI_GEN_SLICES_5__GEN_ROWS_4__sbox_and_xor_inst_d_nxy), .Z0_f (new_AGEMA_signal_4437), .Z1_t (new_AGEMA_signal_4438), .Z1_f (new_AGEMA_signal_4439) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_4__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_5__GEN_ROWS_4__sbox_and_xor_inst_d_nxy), .A0_f (new_AGEMA_signal_4437), .A1_t (new_AGEMA_signal_4438), .A1_f (new_AGEMA_signal_4439), .B0_t (StateFromRhoPi[157]), .B0_f (new_AGEMA_signal_3869), .B1_t (new_AGEMA_signal_3870), .B1_f (new_AGEMA_signal_3871), .Z0_t (StateFromChi[157]), .Z0_f (new_AGEMA_signal_5043), .Z1_t (new_AGEMA_signal_5044), .Z1_f (new_AGEMA_signal_5045) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_4__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[37]), .A0_f (new_AGEMA_signal_3458), .A1_t (new_AGEMA_signal_3459), .A1_f (new_AGEMA_signal_3460), .B0_t (StateFromRhoPi[77]), .B0_f (new_AGEMA_signal_3920), .B1_t (new_AGEMA_signal_3921), .B1_f (new_AGEMA_signal_3922), .Z0_t (CHI_GEN_SLICES_5__GEN_ROWS_4__sbox_and_xor_inst_e_nxy), .Z0_f (new_AGEMA_signal_4440), .Z1_t (new_AGEMA_signal_4441), .Z1_f (new_AGEMA_signal_4442) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_4__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_5__GEN_ROWS_4__sbox_and_xor_inst_e_nxy), .A0_f (new_AGEMA_signal_4440), .A1_t (new_AGEMA_signal_4441), .A1_f (new_AGEMA_signal_4442), .B0_t (StateFromRhoPi[197]), .B0_f (new_AGEMA_signal_3476), .B1_t (new_AGEMA_signal_3477), .B1_f (new_AGEMA_signal_3478), .Z0_t (StateFromChi[197]), .Z0_f (new_AGEMA_signal_5046), .Z1_t (new_AGEMA_signal_5047), .Z1_f (new_AGEMA_signal_5048) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_0__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[46]), .A0_f (new_AGEMA_signal_3590), .A1_t (new_AGEMA_signal_3591), .A1_f (new_AGEMA_signal_3592), .B0_t (StateFromRhoPi[86]), .B0_f (new_AGEMA_signal_3857), .B1_t (new_AGEMA_signal_3858), .B1_f (new_AGEMA_signal_3859), .Z0_t (CHI_GEN_SLICES_6__GEN_ROWS_0__sbox_and_xor_inst_a_nxy), .Z0_f (new_AGEMA_signal_4443), .Z1_t (new_AGEMA_signal_4444), .Z1_f (new_AGEMA_signal_4445) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_0__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_6__GEN_ROWS_0__sbox_and_xor_inst_a_nxy), .A0_f (new_AGEMA_signal_4443), .A1_t (new_AGEMA_signal_4444), .A1_f (new_AGEMA_signal_4445), .B0_t (StateFromRhoPi[6]), .B0_f (new_AGEMA_signal_3773), .B1_t (new_AGEMA_signal_3774), .B1_f (new_AGEMA_signal_3775), .Z0_t (StateFromChi[6]), .Z0_f (new_AGEMA_signal_5049), .Z1_t (new_AGEMA_signal_5050), .Z1_f (new_AGEMA_signal_5051) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_0__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[86]), .A0_f (new_AGEMA_signal_3857), .A1_t (new_AGEMA_signal_3858), .A1_f (new_AGEMA_signal_3859), .B0_t (StateFromRhoPi[126]), .B0_f (new_AGEMA_signal_3569), .B1_t (new_AGEMA_signal_3570), .B1_f (new_AGEMA_signal_3571), .Z0_t (CHI_GEN_SLICES_6__GEN_ROWS_0__sbox_and_xor_inst_b_nxy), .Z0_f (new_AGEMA_signal_4446), .Z1_t (new_AGEMA_signal_4447), .Z1_f (new_AGEMA_signal_4448) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_0__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_6__GEN_ROWS_0__sbox_and_xor_inst_b_nxy), .A0_f (new_AGEMA_signal_4446), .A1_t (new_AGEMA_signal_4447), .A1_f (new_AGEMA_signal_4448), .B0_t (StateFromRhoPi[46]), .B0_f (new_AGEMA_signal_3590), .B1_t (new_AGEMA_signal_3591), .B1_f (new_AGEMA_signal_3592), .Z0_t (StateFromChi[46]), .Z0_f (new_AGEMA_signal_5052), .Z1_t (new_AGEMA_signal_5053), .Z1_f (new_AGEMA_signal_5054) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_0__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[126]), .A0_f (new_AGEMA_signal_3569), .A1_t (new_AGEMA_signal_3570), .A1_f (new_AGEMA_signal_3571), .B0_t (StateFromRhoPi[166]), .B0_f (new_AGEMA_signal_3611), .B1_t (new_AGEMA_signal_3612), .B1_f (new_AGEMA_signal_3613), .Z0_t (CHI_GEN_SLICES_6__GEN_ROWS_0__sbox_and_xor_inst_c_nxy), .Z0_f (new_AGEMA_signal_4449), .Z1_t (new_AGEMA_signal_4450), .Z1_f (new_AGEMA_signal_4451) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_0__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_6__GEN_ROWS_0__sbox_and_xor_inst_c_nxy), .A0_f (new_AGEMA_signal_4449), .A1_t (new_AGEMA_signal_4450), .A1_f (new_AGEMA_signal_4451), .B0_t (StateFromRhoPi[86]), .B0_f (new_AGEMA_signal_3857), .B1_t (new_AGEMA_signal_3858), .B1_f (new_AGEMA_signal_3859), .Z0_t (StateFromChi[86]), .Z0_f (new_AGEMA_signal_5055), .Z1_t (new_AGEMA_signal_5056), .Z1_f (new_AGEMA_signal_5057) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_0__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[166]), .A0_f (new_AGEMA_signal_3611), .A1_t (new_AGEMA_signal_3612), .A1_f (new_AGEMA_signal_3613), .B0_t (StateFromRhoPi[6]), .B0_f (new_AGEMA_signal_3773), .B1_t (new_AGEMA_signal_3774), .B1_f (new_AGEMA_signal_3775), .Z0_t (CHI_GEN_SLICES_6__GEN_ROWS_0__sbox_and_xor_inst_d_nxy), .Z0_f (new_AGEMA_signal_4452), .Z1_t (new_AGEMA_signal_4453), .Z1_f (new_AGEMA_signal_4454) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_0__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_6__GEN_ROWS_0__sbox_and_xor_inst_d_nxy), .A0_f (new_AGEMA_signal_4452), .A1_t (new_AGEMA_signal_4453), .A1_f (new_AGEMA_signal_4454), .B0_t (StateFromRhoPi[126]), .B0_f (new_AGEMA_signal_3569), .B1_t (new_AGEMA_signal_3570), .B1_f (new_AGEMA_signal_3571), .Z0_t (StateFromChi[126]), .Z0_f (new_AGEMA_signal_5058), .Z1_t (new_AGEMA_signal_5059), .Z1_f (new_AGEMA_signal_5060) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_0__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[6]), .A0_f (new_AGEMA_signal_3773), .A1_t (new_AGEMA_signal_3774), .A1_f (new_AGEMA_signal_3775), .B0_t (StateFromRhoPi[46]), .B0_f (new_AGEMA_signal_3590), .B1_t (new_AGEMA_signal_3591), .B1_f (new_AGEMA_signal_3592), .Z0_t (CHI_GEN_SLICES_6__GEN_ROWS_0__sbox_and_xor_inst_e_nxy), .Z0_f (new_AGEMA_signal_4455), .Z1_t (new_AGEMA_signal_4456), .Z1_f (new_AGEMA_signal_4457) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_0__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_6__GEN_ROWS_0__sbox_and_xor_inst_e_nxy), .A0_f (new_AGEMA_signal_4455), .A1_t (new_AGEMA_signal_4456), .A1_f (new_AGEMA_signal_4457), .B0_t (StateFromRhoPi[166]), .B0_f (new_AGEMA_signal_3611), .B1_t (new_AGEMA_signal_3612), .B1_f (new_AGEMA_signal_3613), .Z0_t (StateFromChi[166]), .Z0_f (new_AGEMA_signal_5061), .Z1_t (new_AGEMA_signal_5062), .Z1_f (new_AGEMA_signal_5063) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_1__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[54]), .A0_f (new_AGEMA_signal_3950), .A1_t (new_AGEMA_signal_3951), .A1_f (new_AGEMA_signal_3952), .B0_t (StateFromRhoPi[94]), .B0_f (new_AGEMA_signal_3902), .B1_t (new_AGEMA_signal_3903), .B1_f (new_AGEMA_signal_3904), .Z0_t (CHI_GEN_SLICES_6__GEN_ROWS_1__sbox_and_xor_inst_a_nxy), .Z0_f (new_AGEMA_signal_4458), .Z1_t (new_AGEMA_signal_4459), .Z1_f (new_AGEMA_signal_4460) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_1__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_6__GEN_ROWS_1__sbox_and_xor_inst_a_nxy), .A0_f (new_AGEMA_signal_4458), .A1_t (new_AGEMA_signal_4459), .A1_f (new_AGEMA_signal_4460), .B0_t (StateFromRhoPi[14]), .B0_f (new_AGEMA_signal_3533), .B1_t (new_AGEMA_signal_3534), .B1_f (new_AGEMA_signal_3535), .Z0_t (StateFromChi[14]), .Z0_f (new_AGEMA_signal_5064), .Z1_t (new_AGEMA_signal_5065), .Z1_f (new_AGEMA_signal_5066) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_1__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[94]), .A0_f (new_AGEMA_signal_3902), .A1_t (new_AGEMA_signal_3903), .A1_f (new_AGEMA_signal_3904), .B0_t (StateFromRhoPi[134]), .B0_f (new_AGEMA_signal_3674), .B1_t (new_AGEMA_signal_3675), .B1_f (new_AGEMA_signal_3676), .Z0_t (CHI_GEN_SLICES_6__GEN_ROWS_1__sbox_and_xor_inst_b_nxy), .Z0_f (new_AGEMA_signal_4461), .Z1_t (new_AGEMA_signal_4462), .Z1_f (new_AGEMA_signal_4463) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_1__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_6__GEN_ROWS_1__sbox_and_xor_inst_b_nxy), .A0_f (new_AGEMA_signal_4461), .A1_t (new_AGEMA_signal_4462), .A1_f (new_AGEMA_signal_4463), .B0_t (StateFromRhoPi[54]), .B0_f (new_AGEMA_signal_3950), .B1_t (new_AGEMA_signal_3951), .B1_f (new_AGEMA_signal_3952), .Z0_t (StateFromChi[54]), .Z0_f (new_AGEMA_signal_5067), .Z1_t (new_AGEMA_signal_5068), .Z1_f (new_AGEMA_signal_5069) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_1__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[134]), .A0_f (new_AGEMA_signal_3674), .A1_t (new_AGEMA_signal_3675), .A1_f (new_AGEMA_signal_3676), .B0_t (StateFromRhoPi[174]), .B0_f (new_AGEMA_signal_3686), .B1_t (new_AGEMA_signal_3687), .B1_f (new_AGEMA_signal_3688), .Z0_t (CHI_GEN_SLICES_6__GEN_ROWS_1__sbox_and_xor_inst_c_nxy), .Z0_f (new_AGEMA_signal_4464), .Z1_t (new_AGEMA_signal_4465), .Z1_f (new_AGEMA_signal_4466) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_1__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_6__GEN_ROWS_1__sbox_and_xor_inst_c_nxy), .A0_f (new_AGEMA_signal_4464), .A1_t (new_AGEMA_signal_4465), .A1_f (new_AGEMA_signal_4466), .B0_t (StateFromRhoPi[94]), .B0_f (new_AGEMA_signal_3902), .B1_t (new_AGEMA_signal_3903), .B1_f (new_AGEMA_signal_3904), .Z0_t (StateFromChi[94]), .Z0_f (new_AGEMA_signal_5070), .Z1_t (new_AGEMA_signal_5071), .Z1_f (new_AGEMA_signal_5072) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_1__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[174]), .A0_f (new_AGEMA_signal_3686), .A1_t (new_AGEMA_signal_3687), .A1_f (new_AGEMA_signal_3688), .B0_t (StateFromRhoPi[14]), .B0_f (new_AGEMA_signal_3533), .B1_t (new_AGEMA_signal_3534), .B1_f (new_AGEMA_signal_3535), .Z0_t (CHI_GEN_SLICES_6__GEN_ROWS_1__sbox_and_xor_inst_d_nxy), .Z0_f (new_AGEMA_signal_4467), .Z1_t (new_AGEMA_signal_4468), .Z1_f (new_AGEMA_signal_4469) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_1__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_6__GEN_ROWS_1__sbox_and_xor_inst_d_nxy), .A0_f (new_AGEMA_signal_4467), .A1_t (new_AGEMA_signal_4468), .A1_f (new_AGEMA_signal_4469), .B0_t (StateFromRhoPi[134]), .B0_f (new_AGEMA_signal_3674), .B1_t (new_AGEMA_signal_3675), .B1_f (new_AGEMA_signal_3676), .Z0_t (StateFromChi[134]), .Z0_f (new_AGEMA_signal_5073), .Z1_t (new_AGEMA_signal_5074), .Z1_f (new_AGEMA_signal_5075) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_1__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[14]), .A0_f (new_AGEMA_signal_3533), .A1_t (new_AGEMA_signal_3534), .A1_f (new_AGEMA_signal_3535), .B0_t (StateFromRhoPi[54]), .B0_f (new_AGEMA_signal_3950), .B1_t (new_AGEMA_signal_3951), .B1_f (new_AGEMA_signal_3952), .Z0_t (CHI_GEN_SLICES_6__GEN_ROWS_1__sbox_and_xor_inst_e_nxy), .Z0_f (new_AGEMA_signal_4470), .Z1_t (new_AGEMA_signal_4471), .Z1_f (new_AGEMA_signal_4472) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_1__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_6__GEN_ROWS_1__sbox_and_xor_inst_e_nxy), .A0_f (new_AGEMA_signal_4470), .A1_t (new_AGEMA_signal_4471), .A1_f (new_AGEMA_signal_4472), .B0_t (StateFromRhoPi[174]), .B0_f (new_AGEMA_signal_3686), .B1_t (new_AGEMA_signal_3687), .B1_f (new_AGEMA_signal_3688), .Z0_t (StateFromChi[174]), .Z0_f (new_AGEMA_signal_5076), .Z1_t (new_AGEMA_signal_5077), .Z1_f (new_AGEMA_signal_5078) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_2__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[62]), .A0_f (new_AGEMA_signal_3425), .A1_t (new_AGEMA_signal_3426), .A1_f (new_AGEMA_signal_3427), .B0_t (StateFromRhoPi[102]), .B0_f (new_AGEMA_signal_3932), .B1_t (new_AGEMA_signal_3933), .B1_f (new_AGEMA_signal_3934), .Z0_t (CHI_GEN_SLICES_6__GEN_ROWS_2__sbox_and_xor_inst_a_nxy), .Z0_f (new_AGEMA_signal_4473), .Z1_t (new_AGEMA_signal_4474), .Z1_f (new_AGEMA_signal_4475) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_2__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_6__GEN_ROWS_2__sbox_and_xor_inst_a_nxy), .A0_f (new_AGEMA_signal_4473), .A1_t (new_AGEMA_signal_4474), .A1_f (new_AGEMA_signal_4475), .B0_t (StateFromRhoPi[22]), .B0_f (new_AGEMA_signal_3893), .B1_t (new_AGEMA_signal_3894), .B1_f (new_AGEMA_signal_3895), .Z0_t (StateFromChi[22]), .Z0_f (new_AGEMA_signal_5079), .Z1_t (new_AGEMA_signal_5080), .Z1_f (new_AGEMA_signal_5081) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_2__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[102]), .A0_f (new_AGEMA_signal_3932), .A1_t (new_AGEMA_signal_3933), .A1_f (new_AGEMA_signal_3934), .B0_t (StateFromRhoPi[142]), .B0_f (new_AGEMA_signal_3434), .B1_t (new_AGEMA_signal_3435), .B1_f (new_AGEMA_signal_3436), .Z0_t (CHI_GEN_SLICES_6__GEN_ROWS_2__sbox_and_xor_inst_b_nxy), .Z0_f (new_AGEMA_signal_4476), .Z1_t (new_AGEMA_signal_4477), .Z1_f (new_AGEMA_signal_4478) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_2__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_6__GEN_ROWS_2__sbox_and_xor_inst_b_nxy), .A0_f (new_AGEMA_signal_4476), .A1_t (new_AGEMA_signal_4477), .A1_f (new_AGEMA_signal_4478), .B0_t (StateFromRhoPi[62]), .B0_f (new_AGEMA_signal_3425), .B1_t (new_AGEMA_signal_3426), .B1_f (new_AGEMA_signal_3427), .Z0_t (StateFromChi[62]), .Z0_f (new_AGEMA_signal_5082), .Z1_t (new_AGEMA_signal_5083), .Z1_f (new_AGEMA_signal_5084) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_2__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[142]), .A0_f (new_AGEMA_signal_3434), .A1_t (new_AGEMA_signal_3435), .A1_f (new_AGEMA_signal_3436), .B0_t (StateFromRhoPi[182]), .B0_f (new_AGEMA_signal_3866), .B1_t (new_AGEMA_signal_3867), .B1_f (new_AGEMA_signal_3868), .Z0_t (CHI_GEN_SLICES_6__GEN_ROWS_2__sbox_and_xor_inst_c_nxy), .Z0_f (new_AGEMA_signal_4479), .Z1_t (new_AGEMA_signal_4480), .Z1_f (new_AGEMA_signal_4481) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_2__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_6__GEN_ROWS_2__sbox_and_xor_inst_c_nxy), .A0_f (new_AGEMA_signal_4479), .A1_t (new_AGEMA_signal_4480), .A1_f (new_AGEMA_signal_4481), .B0_t (StateFromRhoPi[102]), .B0_f (new_AGEMA_signal_3932), .B1_t (new_AGEMA_signal_3933), .B1_f (new_AGEMA_signal_3934), .Z0_t (StateFromChi[102]), .Z0_f (new_AGEMA_signal_5085), .Z1_t (new_AGEMA_signal_5086), .Z1_f (new_AGEMA_signal_5087) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_2__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[182]), .A0_f (new_AGEMA_signal_3866), .A1_t (new_AGEMA_signal_3867), .A1_f (new_AGEMA_signal_3868), .B0_t (StateFromRhoPi[22]), .B0_f (new_AGEMA_signal_3893), .B1_t (new_AGEMA_signal_3894), .B1_f (new_AGEMA_signal_3895), .Z0_t (CHI_GEN_SLICES_6__GEN_ROWS_2__sbox_and_xor_inst_d_nxy), .Z0_f (new_AGEMA_signal_4482), .Z1_t (new_AGEMA_signal_4483), .Z1_f (new_AGEMA_signal_4484) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_2__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_6__GEN_ROWS_2__sbox_and_xor_inst_d_nxy), .A0_f (new_AGEMA_signal_4482), .A1_t (new_AGEMA_signal_4483), .A1_f (new_AGEMA_signal_4484), .B0_t (StateFromRhoPi[142]), .B0_f (new_AGEMA_signal_3434), .B1_t (new_AGEMA_signal_3435), .B1_f (new_AGEMA_signal_3436), .Z0_t (StateFromChi[142]), .Z0_f (new_AGEMA_signal_5088), .Z1_t (new_AGEMA_signal_5089), .Z1_f (new_AGEMA_signal_5090) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_2__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[22]), .A0_f (new_AGEMA_signal_3893), .A1_t (new_AGEMA_signal_3894), .A1_f (new_AGEMA_signal_3895), .B0_t (StateFromRhoPi[62]), .B0_f (new_AGEMA_signal_3425), .B1_t (new_AGEMA_signal_3426), .B1_f (new_AGEMA_signal_3427), .Z0_t (CHI_GEN_SLICES_6__GEN_ROWS_2__sbox_and_xor_inst_e_nxy), .Z0_f (new_AGEMA_signal_4485), .Z1_t (new_AGEMA_signal_4486), .Z1_f (new_AGEMA_signal_4487) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_2__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_6__GEN_ROWS_2__sbox_and_xor_inst_e_nxy), .A0_f (new_AGEMA_signal_4485), .A1_t (new_AGEMA_signal_4486), .A1_f (new_AGEMA_signal_4487), .B0_t (StateFromRhoPi[182]), .B0_f (new_AGEMA_signal_3866), .B1_t (new_AGEMA_signal_3867), .B1_f (new_AGEMA_signal_3868), .Z0_t (StateFromChi[182]), .Z0_f (new_AGEMA_signal_5091), .Z1_t (new_AGEMA_signal_5092), .Z1_f (new_AGEMA_signal_5093) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_3__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[70]), .A0_f (new_AGEMA_signal_3710), .A1_t (new_AGEMA_signal_3711), .A1_f (new_AGEMA_signal_3712), .B0_t (StateFromRhoPi[110]), .B0_f (new_AGEMA_signal_3812), .B1_t (new_AGEMA_signal_3813), .B1_f (new_AGEMA_signal_3814), .Z0_t (CHI_GEN_SLICES_6__GEN_ROWS_3__sbox_and_xor_inst_a_nxy), .Z0_f (new_AGEMA_signal_4488), .Z1_t (new_AGEMA_signal_4489), .Z1_f (new_AGEMA_signal_4490) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_3__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_6__GEN_ROWS_3__sbox_and_xor_inst_a_nxy), .A0_f (new_AGEMA_signal_4488), .A1_t (new_AGEMA_signal_4489), .A1_f (new_AGEMA_signal_4490), .B0_t (StateFromRhoPi[30]), .B0_f (new_AGEMA_signal_3788), .B1_t (new_AGEMA_signal_3789), .B1_f (new_AGEMA_signal_3790), .Z0_t (StateFromChi[30]), .Z0_f (new_AGEMA_signal_5094), .Z1_t (new_AGEMA_signal_5095), .Z1_f (new_AGEMA_signal_5096) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_3__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[110]), .A0_f (new_AGEMA_signal_3812), .A1_t (new_AGEMA_signal_3813), .A1_f (new_AGEMA_signal_3814), .B0_t (StateFromRhoPi[150]), .B0_f (new_AGEMA_signal_3449), .B1_t (new_AGEMA_signal_3450), .B1_f (new_AGEMA_signal_3451), .Z0_t (CHI_GEN_SLICES_6__GEN_ROWS_3__sbox_and_xor_inst_b_nxy), .Z0_f (new_AGEMA_signal_4491), .Z1_t (new_AGEMA_signal_4492), .Z1_f (new_AGEMA_signal_4493) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_3__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_6__GEN_ROWS_3__sbox_and_xor_inst_b_nxy), .A0_f (new_AGEMA_signal_4491), .A1_t (new_AGEMA_signal_4492), .A1_f (new_AGEMA_signal_4493), .B0_t (StateFromRhoPi[70]), .B0_f (new_AGEMA_signal_3710), .B1_t (new_AGEMA_signal_3711), .B1_f (new_AGEMA_signal_3712), .Z0_t (StateFromChi[70]), .Z0_f (new_AGEMA_signal_5097), .Z1_t (new_AGEMA_signal_5098), .Z1_f (new_AGEMA_signal_5099) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_3__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[150]), .A0_f (new_AGEMA_signal_3449), .A1_t (new_AGEMA_signal_3450), .A1_f (new_AGEMA_signal_3451), .B0_t (StateFromRhoPi[190]), .B0_f (new_AGEMA_signal_3911), .B1_t (new_AGEMA_signal_3912), .B1_f (new_AGEMA_signal_3913), .Z0_t (CHI_GEN_SLICES_6__GEN_ROWS_3__sbox_and_xor_inst_c_nxy), .Z0_f (new_AGEMA_signal_4494), .Z1_t (new_AGEMA_signal_4495), .Z1_f (new_AGEMA_signal_4496) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_3__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_6__GEN_ROWS_3__sbox_and_xor_inst_c_nxy), .A0_f (new_AGEMA_signal_4494), .A1_t (new_AGEMA_signal_4495), .A1_f (new_AGEMA_signal_4496), .B0_t (StateFromRhoPi[110]), .B0_f (new_AGEMA_signal_3812), .B1_t (new_AGEMA_signal_3813), .B1_f (new_AGEMA_signal_3814), .Z0_t (StateFromChi[110]), .Z0_f (new_AGEMA_signal_5100), .Z1_t (new_AGEMA_signal_5101), .Z1_f (new_AGEMA_signal_5102) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_3__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[190]), .A0_f (new_AGEMA_signal_3911), .A1_t (new_AGEMA_signal_3912), .A1_f (new_AGEMA_signal_3913), .B0_t (StateFromRhoPi[30]), .B0_f (new_AGEMA_signal_3788), .B1_t (new_AGEMA_signal_3789), .B1_f (new_AGEMA_signal_3790), .Z0_t (CHI_GEN_SLICES_6__GEN_ROWS_3__sbox_and_xor_inst_d_nxy), .Z0_f (new_AGEMA_signal_4497), .Z1_t (new_AGEMA_signal_4498), .Z1_f (new_AGEMA_signal_4499) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_3__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_6__GEN_ROWS_3__sbox_and_xor_inst_d_nxy), .A0_f (new_AGEMA_signal_4497), .A1_t (new_AGEMA_signal_4498), .A1_f (new_AGEMA_signal_4499), .B0_t (StateFromRhoPi[150]), .B0_f (new_AGEMA_signal_3449), .B1_t (new_AGEMA_signal_3450), .B1_f (new_AGEMA_signal_3451), .Z0_t (StateFromChi[150]), .Z0_f (new_AGEMA_signal_5103), .Z1_t (new_AGEMA_signal_5104), .Z1_f (new_AGEMA_signal_5105) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_3__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[30]), .A0_f (new_AGEMA_signal_3788), .A1_t (new_AGEMA_signal_3789), .A1_f (new_AGEMA_signal_3790), .B0_t (StateFromRhoPi[70]), .B0_f (new_AGEMA_signal_3710), .B1_t (new_AGEMA_signal_3711), .B1_f (new_AGEMA_signal_3712), .Z0_t (CHI_GEN_SLICES_6__GEN_ROWS_3__sbox_and_xor_inst_e_nxy), .Z0_f (new_AGEMA_signal_4500), .Z1_t (new_AGEMA_signal_4501), .Z1_f (new_AGEMA_signal_4502) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_3__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_6__GEN_ROWS_3__sbox_and_xor_inst_e_nxy), .A0_f (new_AGEMA_signal_4500), .A1_t (new_AGEMA_signal_4501), .A1_f (new_AGEMA_signal_4502), .B0_t (StateFromRhoPi[190]), .B0_f (new_AGEMA_signal_3911), .B1_t (new_AGEMA_signal_3912), .B1_f (new_AGEMA_signal_3913), .Z0_t (StateFromChi[190]), .Z0_f (new_AGEMA_signal_5106), .Z1_t (new_AGEMA_signal_5107), .Z1_f (new_AGEMA_signal_5108) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_4__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[78]), .A0_f (new_AGEMA_signal_3755), .A1_t (new_AGEMA_signal_3756), .A1_f (new_AGEMA_signal_3757), .B0_t (StateFromRhoPi[118]), .B0_f (new_AGEMA_signal_3392), .B1_t (new_AGEMA_signal_3393), .B1_f (new_AGEMA_signal_3394), .Z0_t (CHI_GEN_SLICES_6__GEN_ROWS_4__sbox_and_xor_inst_a_nxy), .Z0_f (new_AGEMA_signal_4503), .Z1_t (new_AGEMA_signal_4504), .Z1_f (new_AGEMA_signal_4505) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_4__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_6__GEN_ROWS_4__sbox_and_xor_inst_a_nxy), .A0_f (new_AGEMA_signal_4503), .A1_t (new_AGEMA_signal_4504), .A1_f (new_AGEMA_signal_4505), .B0_t (StateFromRhoPi[38]), .B0_f (new_AGEMA_signal_3428), .B1_t (new_AGEMA_signal_3429), .B1_f (new_AGEMA_signal_3430), .Z0_t (StateFromChi[38]), .Z0_f (new_AGEMA_signal_5109), .Z1_t (new_AGEMA_signal_5110), .Z1_f (new_AGEMA_signal_5111) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_4__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[118]), .A0_f (new_AGEMA_signal_3392), .A1_t (new_AGEMA_signal_3393), .A1_f (new_AGEMA_signal_3394), .B0_t (StateFromRhoPi[158]), .B0_f (new_AGEMA_signal_3839), .B1_t (new_AGEMA_signal_3840), .B1_f (new_AGEMA_signal_3841), .Z0_t (CHI_GEN_SLICES_6__GEN_ROWS_4__sbox_and_xor_inst_b_nxy), .Z0_f (new_AGEMA_signal_4506), .Z1_t (new_AGEMA_signal_4507), .Z1_f (new_AGEMA_signal_4508) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_4__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_6__GEN_ROWS_4__sbox_and_xor_inst_b_nxy), .A0_f (new_AGEMA_signal_4506), .A1_t (new_AGEMA_signal_4507), .A1_f (new_AGEMA_signal_4508), .B0_t (StateFromRhoPi[78]), .B0_f (new_AGEMA_signal_3755), .B1_t (new_AGEMA_signal_3756), .B1_f (new_AGEMA_signal_3757), .Z0_t (StateFromChi[78]), .Z0_f (new_AGEMA_signal_5112), .Z1_t (new_AGEMA_signal_5113), .Z1_f (new_AGEMA_signal_5114) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_4__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[158]), .A0_f (new_AGEMA_signal_3839), .A1_t (new_AGEMA_signal_3840), .A1_f (new_AGEMA_signal_3841), .B0_t (StateFromRhoPi[198]), .B0_f (new_AGEMA_signal_3806), .B1_t (new_AGEMA_signal_3807), .B1_f (new_AGEMA_signal_3808), .Z0_t (CHI_GEN_SLICES_6__GEN_ROWS_4__sbox_and_xor_inst_c_nxy), .Z0_f (new_AGEMA_signal_4509), .Z1_t (new_AGEMA_signal_4510), .Z1_f (new_AGEMA_signal_4511) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_4__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_6__GEN_ROWS_4__sbox_and_xor_inst_c_nxy), .A0_f (new_AGEMA_signal_4509), .A1_t (new_AGEMA_signal_4510), .A1_f (new_AGEMA_signal_4511), .B0_t (StateFromRhoPi[118]), .B0_f (new_AGEMA_signal_3392), .B1_t (new_AGEMA_signal_3393), .B1_f (new_AGEMA_signal_3394), .Z0_t (StateFromChi[118]), .Z0_f (new_AGEMA_signal_5115), .Z1_t (new_AGEMA_signal_5116), .Z1_f (new_AGEMA_signal_5117) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_4__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[198]), .A0_f (new_AGEMA_signal_3806), .A1_t (new_AGEMA_signal_3807), .A1_f (new_AGEMA_signal_3808), .B0_t (StateFromRhoPi[38]), .B0_f (new_AGEMA_signal_3428), .B1_t (new_AGEMA_signal_3429), .B1_f (new_AGEMA_signal_3430), .Z0_t (CHI_GEN_SLICES_6__GEN_ROWS_4__sbox_and_xor_inst_d_nxy), .Z0_f (new_AGEMA_signal_4512), .Z1_t (new_AGEMA_signal_4513), .Z1_f (new_AGEMA_signal_4514) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_4__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_6__GEN_ROWS_4__sbox_and_xor_inst_d_nxy), .A0_f (new_AGEMA_signal_4512), .A1_t (new_AGEMA_signal_4513), .A1_f (new_AGEMA_signal_4514), .B0_t (StateFromRhoPi[158]), .B0_f (new_AGEMA_signal_3839), .B1_t (new_AGEMA_signal_3840), .B1_f (new_AGEMA_signal_3841), .Z0_t (StateFromChi[158]), .Z0_f (new_AGEMA_signal_5118), .Z1_t (new_AGEMA_signal_5119), .Z1_f (new_AGEMA_signal_5120) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_4__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[38]), .A0_f (new_AGEMA_signal_3428), .A1_t (new_AGEMA_signal_3429), .A1_f (new_AGEMA_signal_3430), .B0_t (StateFromRhoPi[78]), .B0_f (new_AGEMA_signal_3755), .B1_t (new_AGEMA_signal_3756), .B1_f (new_AGEMA_signal_3757), .Z0_t (CHI_GEN_SLICES_6__GEN_ROWS_4__sbox_and_xor_inst_e_nxy), .Z0_f (new_AGEMA_signal_4515), .Z1_t (new_AGEMA_signal_4516), .Z1_f (new_AGEMA_signal_4517) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_4__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_6__GEN_ROWS_4__sbox_and_xor_inst_e_nxy), .A0_f (new_AGEMA_signal_4515), .A1_t (new_AGEMA_signal_4516), .A1_f (new_AGEMA_signal_4517), .B0_t (StateFromRhoPi[198]), .B0_f (new_AGEMA_signal_3806), .B1_t (new_AGEMA_signal_3807), .B1_f (new_AGEMA_signal_3808), .Z0_t (StateFromChi[198]), .Z0_f (new_AGEMA_signal_5121), .Z1_t (new_AGEMA_signal_5122), .Z1_f (new_AGEMA_signal_5123) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_0__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[47]), .A0_f (new_AGEMA_signal_3485), .A1_t (new_AGEMA_signal_3486), .A1_f (new_AGEMA_signal_3487), .B0_t (StateFromRhoPi[87]), .B0_f (new_AGEMA_signal_3827), .B1_t (new_AGEMA_signal_3828), .B1_f (new_AGEMA_signal_3829), .Z0_t (CHI_GEN_SLICES_7__GEN_ROWS_0__sbox_and_xor_inst_a_nxy), .Z0_f (new_AGEMA_signal_4518), .Z1_t (new_AGEMA_signal_4519), .Z1_f (new_AGEMA_signal_4520) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_0__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_7__GEN_ROWS_0__sbox_and_xor_inst_a_nxy), .A0_f (new_AGEMA_signal_4518), .A1_t (new_AGEMA_signal_4519), .A1_f (new_AGEMA_signal_4520), .B0_t (StateFromRhoPi[7]), .B0_f (new_AGEMA_signal_3728), .B1_t (new_AGEMA_signal_3729), .B1_f (new_AGEMA_signal_3730), .Z0_t (CHI_ChiOut_7), .Z0_f (new_AGEMA_signal_5124), .Z1_t (new_AGEMA_signal_5125), .Z1_f (new_AGEMA_signal_5126) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_0__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[87]), .A0_f (new_AGEMA_signal_3827), .A1_t (new_AGEMA_signal_3828), .A1_f (new_AGEMA_signal_3829), .B0_t (StateFromRhoPi[127]), .B0_f (new_AGEMA_signal_3524), .B1_t (new_AGEMA_signal_3525), .B1_f (new_AGEMA_signal_3526), .Z0_t (CHI_GEN_SLICES_7__GEN_ROWS_0__sbox_and_xor_inst_b_nxy), .Z0_f (new_AGEMA_signal_4521), .Z1_t (new_AGEMA_signal_4522), .Z1_f (new_AGEMA_signal_4523) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_0__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_7__GEN_ROWS_0__sbox_and_xor_inst_b_nxy), .A0_f (new_AGEMA_signal_4521), .A1_t (new_AGEMA_signal_4522), .A1_f (new_AGEMA_signal_4523), .B0_t (StateFromRhoPi[47]), .B0_f (new_AGEMA_signal_3485), .B1_t (new_AGEMA_signal_3486), .B1_f (new_AGEMA_signal_3487), .Z0_t (StateFromChi[47]), .Z0_f (new_AGEMA_signal_5127), .Z1_t (new_AGEMA_signal_5128), .Z1_f (new_AGEMA_signal_5129) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_0__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[127]), .A0_f (new_AGEMA_signal_3524), .A1_t (new_AGEMA_signal_3525), .A1_f (new_AGEMA_signal_3526), .B0_t (StateFromRhoPi[167]), .B0_f (new_AGEMA_signal_3491), .B1_t (new_AGEMA_signal_3492), .B1_f (new_AGEMA_signal_3493), .Z0_t (CHI_GEN_SLICES_7__GEN_ROWS_0__sbox_and_xor_inst_c_nxy), .Z0_f (new_AGEMA_signal_4524), .Z1_t (new_AGEMA_signal_4525), .Z1_f (new_AGEMA_signal_4526) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_0__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_7__GEN_ROWS_0__sbox_and_xor_inst_c_nxy), .A0_f (new_AGEMA_signal_4524), .A1_t (new_AGEMA_signal_4525), .A1_f (new_AGEMA_signal_4526), .B0_t (StateFromRhoPi[87]), .B0_f (new_AGEMA_signal_3827), .B1_t (new_AGEMA_signal_3828), .B1_f (new_AGEMA_signal_3829), .Z0_t (StateFromChi[87]), .Z0_f (new_AGEMA_signal_5130), .Z1_t (new_AGEMA_signal_5131), .Z1_f (new_AGEMA_signal_5132) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_0__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[167]), .A0_f (new_AGEMA_signal_3491), .A1_t (new_AGEMA_signal_3492), .A1_f (new_AGEMA_signal_3493), .B0_t (StateFromRhoPi[7]), .B0_f (new_AGEMA_signal_3728), .B1_t (new_AGEMA_signal_3729), .B1_f (new_AGEMA_signal_3730), .Z0_t (CHI_GEN_SLICES_7__GEN_ROWS_0__sbox_and_xor_inst_d_nxy), .Z0_f (new_AGEMA_signal_4527), .Z1_t (new_AGEMA_signal_4528), .Z1_f (new_AGEMA_signal_4529) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_0__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_7__GEN_ROWS_0__sbox_and_xor_inst_d_nxy), .A0_f (new_AGEMA_signal_4527), .A1_t (new_AGEMA_signal_4528), .A1_f (new_AGEMA_signal_4529), .B0_t (StateFromRhoPi[127]), .B0_f (new_AGEMA_signal_3524), .B1_t (new_AGEMA_signal_3525), .B1_f (new_AGEMA_signal_3526), .Z0_t (StateFromChi[127]), .Z0_f (new_AGEMA_signal_5133), .Z1_t (new_AGEMA_signal_5134), .Z1_f (new_AGEMA_signal_5135) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_0__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[7]), .A0_f (new_AGEMA_signal_3728), .A1_t (new_AGEMA_signal_3729), .A1_f (new_AGEMA_signal_3730), .B0_t (StateFromRhoPi[47]), .B0_f (new_AGEMA_signal_3485), .B1_t (new_AGEMA_signal_3486), .B1_f (new_AGEMA_signal_3487), .Z0_t (CHI_GEN_SLICES_7__GEN_ROWS_0__sbox_and_xor_inst_e_nxy), .Z0_f (new_AGEMA_signal_4530), .Z1_t (new_AGEMA_signal_4531), .Z1_f (new_AGEMA_signal_4532) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_0__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_7__GEN_ROWS_0__sbox_and_xor_inst_e_nxy), .A0_f (new_AGEMA_signal_4530), .A1_t (new_AGEMA_signal_4531), .A1_f (new_AGEMA_signal_4532), .B0_t (StateFromRhoPi[167]), .B0_f (new_AGEMA_signal_3491), .B1_t (new_AGEMA_signal_3492), .B1_f (new_AGEMA_signal_3493), .Z0_t (StateFromChi[167]), .Z0_f (new_AGEMA_signal_5136), .Z1_t (new_AGEMA_signal_5137), .Z1_f (new_AGEMA_signal_5138) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_1__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[55]), .A0_f (new_AGEMA_signal_3785), .A1_t (new_AGEMA_signal_3786), .A1_f (new_AGEMA_signal_3787), .B0_t (StateFromRhoPi[95]), .B0_f (new_AGEMA_signal_3872), .B1_t (new_AGEMA_signal_3873), .B1_f (new_AGEMA_signal_3874), .Z0_t (CHI_GEN_SLICES_7__GEN_ROWS_1__sbox_and_xor_inst_a_nxy), .Z0_f (new_AGEMA_signal_4533), .Z1_t (new_AGEMA_signal_4534), .Z1_f (new_AGEMA_signal_4535) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_1__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_7__GEN_ROWS_1__sbox_and_xor_inst_a_nxy), .A0_f (new_AGEMA_signal_4533), .A1_t (new_AGEMA_signal_4534), .A1_f (new_AGEMA_signal_4535), .B0_t (StateFromRhoPi[15]), .B0_f (new_AGEMA_signal_3983), .B1_t (new_AGEMA_signal_3984), .B1_f (new_AGEMA_signal_3985), .Z0_t (StateFromChi[15]), .Z0_f (new_AGEMA_signal_5139), .Z1_t (new_AGEMA_signal_5140), .Z1_f (new_AGEMA_signal_5141) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_1__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[95]), .A0_f (new_AGEMA_signal_3872), .A1_t (new_AGEMA_signal_3873), .A1_f (new_AGEMA_signal_3874), .B0_t (StateFromRhoPi[135]), .B0_f (new_AGEMA_signal_3584), .B1_t (new_AGEMA_signal_3585), .B1_f (new_AGEMA_signal_3586), .Z0_t (CHI_GEN_SLICES_7__GEN_ROWS_1__sbox_and_xor_inst_b_nxy), .Z0_f (new_AGEMA_signal_4536), .Z1_t (new_AGEMA_signal_4537), .Z1_f (new_AGEMA_signal_4538) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_1__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_7__GEN_ROWS_1__sbox_and_xor_inst_b_nxy), .A0_f (new_AGEMA_signal_4536), .A1_t (new_AGEMA_signal_4537), .A1_f (new_AGEMA_signal_4538), .B0_t (StateFromRhoPi[55]), .B0_f (new_AGEMA_signal_3785), .B1_t (new_AGEMA_signal_3786), .B1_f (new_AGEMA_signal_3787), .Z0_t (StateFromChi[55]), .Z0_f (new_AGEMA_signal_5142), .Z1_t (new_AGEMA_signal_5143), .Z1_f (new_AGEMA_signal_5144) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_1__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[135]), .A0_f (new_AGEMA_signal_3584), .A1_t (new_AGEMA_signal_3585), .A1_f (new_AGEMA_signal_3586), .B0_t (StateFromRhoPi[175]), .B0_f (new_AGEMA_signal_3551), .B1_t (new_AGEMA_signal_3552), .B1_f (new_AGEMA_signal_3553), .Z0_t (CHI_GEN_SLICES_7__GEN_ROWS_1__sbox_and_xor_inst_c_nxy), .Z0_f (new_AGEMA_signal_4539), .Z1_t (new_AGEMA_signal_4540), .Z1_f (new_AGEMA_signal_4541) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_1__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_7__GEN_ROWS_1__sbox_and_xor_inst_c_nxy), .A0_f (new_AGEMA_signal_4539), .A1_t (new_AGEMA_signal_4540), .A1_f (new_AGEMA_signal_4541), .B0_t (StateFromRhoPi[95]), .B0_f (new_AGEMA_signal_3872), .B1_t (new_AGEMA_signal_3873), .B1_f (new_AGEMA_signal_3874), .Z0_t (StateFromChi[95]), .Z0_f (new_AGEMA_signal_5145), .Z1_t (new_AGEMA_signal_5146), .Z1_f (new_AGEMA_signal_5147) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_1__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[175]), .A0_f (new_AGEMA_signal_3551), .A1_t (new_AGEMA_signal_3552), .A1_f (new_AGEMA_signal_3553), .B0_t (StateFromRhoPi[15]), .B0_f (new_AGEMA_signal_3983), .B1_t (new_AGEMA_signal_3984), .B1_f (new_AGEMA_signal_3985), .Z0_t (CHI_GEN_SLICES_7__GEN_ROWS_1__sbox_and_xor_inst_d_nxy), .Z0_f (new_AGEMA_signal_4542), .Z1_t (new_AGEMA_signal_4543), .Z1_f (new_AGEMA_signal_4544) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_1__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_7__GEN_ROWS_1__sbox_and_xor_inst_d_nxy), .A0_f (new_AGEMA_signal_4542), .A1_t (new_AGEMA_signal_4543), .A1_f (new_AGEMA_signal_4544), .B0_t (StateFromRhoPi[135]), .B0_f (new_AGEMA_signal_3584), .B1_t (new_AGEMA_signal_3585), .B1_f (new_AGEMA_signal_3586), .Z0_t (StateFromChi[135]), .Z0_f (new_AGEMA_signal_5148), .Z1_t (new_AGEMA_signal_5149), .Z1_f (new_AGEMA_signal_5150) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_1__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[15]), .A0_f (new_AGEMA_signal_3983), .A1_t (new_AGEMA_signal_3984), .A1_f (new_AGEMA_signal_3985), .B0_t (StateFromRhoPi[55]), .B0_f (new_AGEMA_signal_3785), .B1_t (new_AGEMA_signal_3786), .B1_f (new_AGEMA_signal_3787), .Z0_t (CHI_GEN_SLICES_7__GEN_ROWS_1__sbox_and_xor_inst_e_nxy), .Z0_f (new_AGEMA_signal_4545), .Z1_t (new_AGEMA_signal_4546), .Z1_f (new_AGEMA_signal_4547) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_1__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_7__GEN_ROWS_1__sbox_and_xor_inst_e_nxy), .A0_f (new_AGEMA_signal_4545), .A1_t (new_AGEMA_signal_4546), .A1_f (new_AGEMA_signal_4547), .B0_t (StateFromRhoPi[175]), .B0_f (new_AGEMA_signal_3551), .B1_t (new_AGEMA_signal_3552), .B1_f (new_AGEMA_signal_3553), .Z0_t (StateFromChi[175]), .Z0_f (new_AGEMA_signal_5151), .Z1_t (new_AGEMA_signal_5152), .Z1_f (new_AGEMA_signal_5153) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_2__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[63]), .A0_f (new_AGEMA_signal_3695), .A1_t (new_AGEMA_signal_3696), .A1_f (new_AGEMA_signal_3697), .B0_t (StateFromRhoPi[103]), .B0_f (new_AGEMA_signal_3917), .B1_t (new_AGEMA_signal_3918), .B1_f (new_AGEMA_signal_3919), .Z0_t (CHI_GEN_SLICES_7__GEN_ROWS_2__sbox_and_xor_inst_a_nxy), .Z0_f (new_AGEMA_signal_4548), .Z1_t (new_AGEMA_signal_4549), .Z1_f (new_AGEMA_signal_4550) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_2__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_7__GEN_ROWS_2__sbox_and_xor_inst_a_nxy), .A0_f (new_AGEMA_signal_4548), .A1_t (new_AGEMA_signal_4549), .A1_f (new_AGEMA_signal_4550), .B0_t (StateFromRhoPi[23]), .B0_f (new_AGEMA_signal_3413), .B1_t (new_AGEMA_signal_3414), .B1_f (new_AGEMA_signal_3415), .Z0_t (StateFromChi[23]), .Z0_f (new_AGEMA_signal_5154), .Z1_t (new_AGEMA_signal_5155), .Z1_f (new_AGEMA_signal_5156) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_2__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[103]), .A0_f (new_AGEMA_signal_3917), .A1_t (new_AGEMA_signal_3918), .A1_f (new_AGEMA_signal_3919), .B0_t (StateFromRhoPi[143]), .B0_f (new_AGEMA_signal_3389), .B1_t (new_AGEMA_signal_3390), .B1_f (new_AGEMA_signal_3391), .Z0_t (CHI_GEN_SLICES_7__GEN_ROWS_2__sbox_and_xor_inst_b_nxy), .Z0_f (new_AGEMA_signal_4551), .Z1_t (new_AGEMA_signal_4552), .Z1_f (new_AGEMA_signal_4553) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_2__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_7__GEN_ROWS_2__sbox_and_xor_inst_b_nxy), .A0_f (new_AGEMA_signal_4551), .A1_t (new_AGEMA_signal_4552), .A1_f (new_AGEMA_signal_4553), .B0_t (StateFromRhoPi[63]), .B0_f (new_AGEMA_signal_3695), .B1_t (new_AGEMA_signal_3696), .B1_f (new_AGEMA_signal_3697), .Z0_t (StateFromChi[63]), .Z0_f (new_AGEMA_signal_5157), .Z1_t (new_AGEMA_signal_5158), .Z1_f (new_AGEMA_signal_5159) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_2__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[143]), .A0_f (new_AGEMA_signal_3389), .A1_t (new_AGEMA_signal_3390), .A1_f (new_AGEMA_signal_3391), .B0_t (StateFromRhoPi[183]), .B0_f (new_AGEMA_signal_3836), .B1_t (new_AGEMA_signal_3837), .B1_f (new_AGEMA_signal_3838), .Z0_t (CHI_GEN_SLICES_7__GEN_ROWS_2__sbox_and_xor_inst_c_nxy), .Z0_f (new_AGEMA_signal_4554), .Z1_t (new_AGEMA_signal_4555), .Z1_f (new_AGEMA_signal_4556) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_2__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_7__GEN_ROWS_2__sbox_and_xor_inst_c_nxy), .A0_f (new_AGEMA_signal_4554), .A1_t (new_AGEMA_signal_4555), .A1_f (new_AGEMA_signal_4556), .B0_t (StateFromRhoPi[103]), .B0_f (new_AGEMA_signal_3917), .B1_t (new_AGEMA_signal_3918), .B1_f (new_AGEMA_signal_3919), .Z0_t (StateFromChi[103]), .Z0_f (new_AGEMA_signal_5160), .Z1_t (new_AGEMA_signal_5161), .Z1_f (new_AGEMA_signal_5162) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_2__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[183]), .A0_f (new_AGEMA_signal_3836), .A1_t (new_AGEMA_signal_3837), .A1_f (new_AGEMA_signal_3838), .B0_t (StateFromRhoPi[23]), .B0_f (new_AGEMA_signal_3413), .B1_t (new_AGEMA_signal_3414), .B1_f (new_AGEMA_signal_3415), .Z0_t (CHI_GEN_SLICES_7__GEN_ROWS_2__sbox_and_xor_inst_d_nxy), .Z0_f (new_AGEMA_signal_4557), .Z1_t (new_AGEMA_signal_4558), .Z1_f (new_AGEMA_signal_4559) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_2__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_7__GEN_ROWS_2__sbox_and_xor_inst_d_nxy), .A0_f (new_AGEMA_signal_4557), .A1_t (new_AGEMA_signal_4558), .A1_f (new_AGEMA_signal_4559), .B0_t (StateFromRhoPi[143]), .B0_f (new_AGEMA_signal_3389), .B1_t (new_AGEMA_signal_3390), .B1_f (new_AGEMA_signal_3391), .Z0_t (StateFromChi[143]), .Z0_f (new_AGEMA_signal_5163), .Z1_t (new_AGEMA_signal_5164), .Z1_f (new_AGEMA_signal_5165) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_2__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[23]), .A0_f (new_AGEMA_signal_3413), .A1_t (new_AGEMA_signal_3414), .A1_f (new_AGEMA_signal_3415), .B0_t (StateFromRhoPi[63]), .B0_f (new_AGEMA_signal_3695), .B1_t (new_AGEMA_signal_3696), .B1_f (new_AGEMA_signal_3697), .Z0_t (CHI_GEN_SLICES_7__GEN_ROWS_2__sbox_and_xor_inst_e_nxy), .Z0_f (new_AGEMA_signal_4560), .Z1_t (new_AGEMA_signal_4561), .Z1_f (new_AGEMA_signal_4562) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_2__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_7__GEN_ROWS_2__sbox_and_xor_inst_e_nxy), .A0_f (new_AGEMA_signal_4560), .A1_t (new_AGEMA_signal_4561), .A1_f (new_AGEMA_signal_4562), .B0_t (StateFromRhoPi[183]), .B0_f (new_AGEMA_signal_3836), .B1_t (new_AGEMA_signal_3837), .B1_f (new_AGEMA_signal_3838), .Z0_t (StateFromChi[183]), .Z0_f (new_AGEMA_signal_5166), .Z1_t (new_AGEMA_signal_5167), .Z1_f (new_AGEMA_signal_5168) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_3__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[71]), .A0_f (new_AGEMA_signal_3905), .A1_t (new_AGEMA_signal_3906), .A1_f (new_AGEMA_signal_3907), .B0_t (StateFromRhoPi[111]), .B0_f (new_AGEMA_signal_3887), .B1_t (new_AGEMA_signal_3888), .B1_f (new_AGEMA_signal_3889), .Z0_t (CHI_GEN_SLICES_7__GEN_ROWS_3__sbox_and_xor_inst_a_nxy), .Z0_f (new_AGEMA_signal_4563), .Z1_t (new_AGEMA_signal_4564), .Z1_f (new_AGEMA_signal_4565) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_3__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_7__GEN_ROWS_3__sbox_and_xor_inst_a_nxy), .A0_f (new_AGEMA_signal_4563), .A1_t (new_AGEMA_signal_4564), .A1_f (new_AGEMA_signal_4565), .B0_t (StateFromRhoPi[31]), .B0_f (new_AGEMA_signal_3473), .B1_t (new_AGEMA_signal_3474), .B1_f (new_AGEMA_signal_3475), .Z0_t (StateFromChi[31]), .Z0_f (new_AGEMA_signal_5169), .Z1_t (new_AGEMA_signal_5170), .Z1_f (new_AGEMA_signal_5171) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_3__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[111]), .A0_f (new_AGEMA_signal_3887), .A1_t (new_AGEMA_signal_3888), .A1_f (new_AGEMA_signal_3889), .B0_t (StateFromRhoPi[151]), .B0_f (new_AGEMA_signal_3419), .B1_t (new_AGEMA_signal_3420), .B1_f (new_AGEMA_signal_3421), .Z0_t (CHI_GEN_SLICES_7__GEN_ROWS_3__sbox_and_xor_inst_b_nxy), .Z0_f (new_AGEMA_signal_4566), .Z1_t (new_AGEMA_signal_4567), .Z1_f (new_AGEMA_signal_4568) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_3__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_7__GEN_ROWS_3__sbox_and_xor_inst_b_nxy), .A0_f (new_AGEMA_signal_4566), .A1_t (new_AGEMA_signal_4567), .A1_f (new_AGEMA_signal_4568), .B0_t (StateFromRhoPi[71]), .B0_f (new_AGEMA_signal_3905), .B1_t (new_AGEMA_signal_3906), .B1_f (new_AGEMA_signal_3907), .Z0_t (StateFromChi[71]), .Z0_f (new_AGEMA_signal_5172), .Z1_t (new_AGEMA_signal_5173), .Z1_f (new_AGEMA_signal_5174) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_3__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[151]), .A0_f (new_AGEMA_signal_3419), .A1_t (new_AGEMA_signal_3420), .A1_f (new_AGEMA_signal_3421), .B0_t (StateFromRhoPi[191]), .B0_f (new_AGEMA_signal_3746), .B1_t (new_AGEMA_signal_3747), .B1_f (new_AGEMA_signal_3748), .Z0_t (CHI_GEN_SLICES_7__GEN_ROWS_3__sbox_and_xor_inst_c_nxy), .Z0_f (new_AGEMA_signal_4569), .Z1_t (new_AGEMA_signal_4570), .Z1_f (new_AGEMA_signal_4571) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_3__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_7__GEN_ROWS_3__sbox_and_xor_inst_c_nxy), .A0_f (new_AGEMA_signal_4569), .A1_t (new_AGEMA_signal_4570), .A1_f (new_AGEMA_signal_4571), .B0_t (StateFromRhoPi[111]), .B0_f (new_AGEMA_signal_3887), .B1_t (new_AGEMA_signal_3888), .B1_f (new_AGEMA_signal_3889), .Z0_t (StateFromChi[111]), .Z0_f (new_AGEMA_signal_5175), .Z1_t (new_AGEMA_signal_5176), .Z1_f (new_AGEMA_signal_5177) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_3__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[191]), .A0_f (new_AGEMA_signal_3746), .A1_t (new_AGEMA_signal_3747), .A1_f (new_AGEMA_signal_3748), .B0_t (StateFromRhoPi[31]), .B0_f (new_AGEMA_signal_3473), .B1_t (new_AGEMA_signal_3474), .B1_f (new_AGEMA_signal_3475), .Z0_t (CHI_GEN_SLICES_7__GEN_ROWS_3__sbox_and_xor_inst_d_nxy), .Z0_f (new_AGEMA_signal_4572), .Z1_t (new_AGEMA_signal_4573), .Z1_f (new_AGEMA_signal_4574) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_3__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_7__GEN_ROWS_3__sbox_and_xor_inst_d_nxy), .A0_f (new_AGEMA_signal_4572), .A1_t (new_AGEMA_signal_4573), .A1_f (new_AGEMA_signal_4574), .B0_t (StateFromRhoPi[151]), .B0_f (new_AGEMA_signal_3419), .B1_t (new_AGEMA_signal_3420), .B1_f (new_AGEMA_signal_3421), .Z0_t (StateFromChi[151]), .Z0_f (new_AGEMA_signal_5178), .Z1_t (new_AGEMA_signal_5179), .Z1_f (new_AGEMA_signal_5180) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_3__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[31]), .A0_f (new_AGEMA_signal_3473), .A1_t (new_AGEMA_signal_3474), .A1_f (new_AGEMA_signal_3475), .B0_t (StateFromRhoPi[71]), .B0_f (new_AGEMA_signal_3905), .B1_t (new_AGEMA_signal_3906), .B1_f (new_AGEMA_signal_3907), .Z0_t (CHI_GEN_SLICES_7__GEN_ROWS_3__sbox_and_xor_inst_e_nxy), .Z0_f (new_AGEMA_signal_4575), .Z1_t (new_AGEMA_signal_4576), .Z1_f (new_AGEMA_signal_4577) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_3__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_7__GEN_ROWS_3__sbox_and_xor_inst_e_nxy), .A0_f (new_AGEMA_signal_4575), .A1_t (new_AGEMA_signal_4576), .A1_f (new_AGEMA_signal_4577), .B0_t (StateFromRhoPi[191]), .B0_f (new_AGEMA_signal_3746), .B1_t (new_AGEMA_signal_3747), .B1_f (new_AGEMA_signal_3748), .Z0_t (StateFromChi[191]), .Z0_f (new_AGEMA_signal_5181), .Z1_t (new_AGEMA_signal_5182), .Z1_f (new_AGEMA_signal_5183) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_4__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[79]), .A0_f (new_AGEMA_signal_3665), .A1_t (new_AGEMA_signal_3666), .A1_f (new_AGEMA_signal_3667), .B0_t (StateFromRhoPi[119]), .B0_f (new_AGEMA_signal_3617), .B1_t (new_AGEMA_signal_3618), .B1_f (new_AGEMA_signal_3619), .Z0_t (CHI_GEN_SLICES_7__GEN_ROWS_4__sbox_and_xor_inst_a_nxy), .Z0_f (new_AGEMA_signal_4578), .Z1_t (new_AGEMA_signal_4579), .Z1_f (new_AGEMA_signal_4580) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_4__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_7__GEN_ROWS_4__sbox_and_xor_inst_a_nxy), .A0_f (new_AGEMA_signal_4578), .A1_t (new_AGEMA_signal_4579), .A1_f (new_AGEMA_signal_4580), .B0_t (StateFromRhoPi[39]), .B0_f (new_AGEMA_signal_3698), .B1_t (new_AGEMA_signal_3699), .B1_f (new_AGEMA_signal_3700), .Z0_t (StateFromChi[39]), .Z0_f (new_AGEMA_signal_5184), .Z1_t (new_AGEMA_signal_5185), .Z1_f (new_AGEMA_signal_5186) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_4__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[119]), .A0_f (new_AGEMA_signal_3617), .A1_t (new_AGEMA_signal_3618), .A1_f (new_AGEMA_signal_3619), .B0_t (StateFromRhoPi[159]), .B0_f (new_AGEMA_signal_3764), .B1_t (new_AGEMA_signal_3765), .B1_f (new_AGEMA_signal_3766), .Z0_t (CHI_GEN_SLICES_7__GEN_ROWS_4__sbox_and_xor_inst_b_nxy), .Z0_f (new_AGEMA_signal_4581), .Z1_t (new_AGEMA_signal_4582), .Z1_f (new_AGEMA_signal_4583) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_4__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_7__GEN_ROWS_4__sbox_and_xor_inst_b_nxy), .A0_f (new_AGEMA_signal_4581), .A1_t (new_AGEMA_signal_4582), .A1_f (new_AGEMA_signal_4583), .B0_t (StateFromRhoPi[79]), .B0_f (new_AGEMA_signal_3665), .B1_t (new_AGEMA_signal_3666), .B1_f (new_AGEMA_signal_3667), .Z0_t (StateFromChi[79]), .Z0_f (new_AGEMA_signal_5187), .Z1_t (new_AGEMA_signal_5188), .Z1_f (new_AGEMA_signal_5189) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_4__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[159]), .A0_f (new_AGEMA_signal_3764), .A1_t (new_AGEMA_signal_3765), .A1_f (new_AGEMA_signal_3766), .B0_t (StateFromRhoPi[199]), .B0_f (new_AGEMA_signal_3881), .B1_t (new_AGEMA_signal_3882), .B1_f (new_AGEMA_signal_3883), .Z0_t (CHI_GEN_SLICES_7__GEN_ROWS_4__sbox_and_xor_inst_c_nxy), .Z0_f (new_AGEMA_signal_4584), .Z1_t (new_AGEMA_signal_4585), .Z1_f (new_AGEMA_signal_4586) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_4__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_7__GEN_ROWS_4__sbox_and_xor_inst_c_nxy), .A0_f (new_AGEMA_signal_4584), .A1_t (new_AGEMA_signal_4585), .A1_f (new_AGEMA_signal_4586), .B0_t (StateFromRhoPi[119]), .B0_f (new_AGEMA_signal_3617), .B1_t (new_AGEMA_signal_3618), .B1_f (new_AGEMA_signal_3619), .Z0_t (StateFromChi[119]), .Z0_f (new_AGEMA_signal_5190), .Z1_t (new_AGEMA_signal_5191), .Z1_f (new_AGEMA_signal_5192) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_4__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[199]), .A0_f (new_AGEMA_signal_3881), .A1_t (new_AGEMA_signal_3882), .A1_f (new_AGEMA_signal_3883), .B0_t (StateFromRhoPi[39]), .B0_f (new_AGEMA_signal_3698), .B1_t (new_AGEMA_signal_3699), .B1_f (new_AGEMA_signal_3700), .Z0_t (CHI_GEN_SLICES_7__GEN_ROWS_4__sbox_and_xor_inst_d_nxy), .Z0_f (new_AGEMA_signal_4587), .Z1_t (new_AGEMA_signal_4588), .Z1_f (new_AGEMA_signal_4589) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_4__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_7__GEN_ROWS_4__sbox_and_xor_inst_d_nxy), .A0_f (new_AGEMA_signal_4587), .A1_t (new_AGEMA_signal_4588), .A1_f (new_AGEMA_signal_4589), .B0_t (StateFromRhoPi[159]), .B0_f (new_AGEMA_signal_3764), .B1_t (new_AGEMA_signal_3765), .B1_f (new_AGEMA_signal_3766), .Z0_t (StateFromChi[159]), .Z0_f (new_AGEMA_signal_5193), .Z1_t (new_AGEMA_signal_5194), .Z1_f (new_AGEMA_signal_5195) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_4__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[39]), .A0_f (new_AGEMA_signal_3698), .A1_t (new_AGEMA_signal_3699), .A1_f (new_AGEMA_signal_3700), .B0_t (StateFromRhoPi[79]), .B0_f (new_AGEMA_signal_3665), .B1_t (new_AGEMA_signal_3666), .B1_f (new_AGEMA_signal_3667), .Z0_t (CHI_GEN_SLICES_7__GEN_ROWS_4__sbox_and_xor_inst_e_nxy), .Z0_f (new_AGEMA_signal_4590), .Z1_t (new_AGEMA_signal_4591), .Z1_f (new_AGEMA_signal_4592) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_4__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_7__GEN_ROWS_4__sbox_and_xor_inst_e_nxy), .A0_f (new_AGEMA_signal_4590), .A1_t (new_AGEMA_signal_4591), .A1_f (new_AGEMA_signal_4592), .B0_t (StateFromRhoPi[199]), .B0_f (new_AGEMA_signal_3881), .B1_t (new_AGEMA_signal_3882), .B1_f (new_AGEMA_signal_3883), .Z0_t (StateFromChi[199]), .Z0_f (new_AGEMA_signal_5196), .Z1_t (new_AGEMA_signal_5197), .Z1_f (new_AGEMA_signal_5198) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b1), .NL(1'b1)) KECCAK_CONTROL_U42 ( .A0_t (KECCAK_CONTROL_n47), .A0_f (new_AGEMA_signal_2988), .B0_t (Reset_t), .B0_f (Reset_f), .Z0_t (KECCAK_CONTROL_CtrlStatexDP[0]), .Z0_f (new_AGEMA_signal_2853) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_U41 ( .A0_t (KECCAK_CONTROL_n45), .A0_f (new_AGEMA_signal_2852), .B0_t (KECCAK_CONTROL_CtrlStatexDP[0]), .B0_f (new_AGEMA_signal_2853), .Z0_t (KECCAK_CONTROL_n47), .Z0_f (new_AGEMA_signal_2988) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_U40 ( .A0_t (KECCAK_CONTROL_CtrlStatexDP_reg_1__Q), .A0_f (new_AGEMA_signal_2850), .B0_t (KECCAK_CONTROL_CtrlStatexDP[2]), .B0_f (new_AGEMA_signal_2851), .Z0_t (KECCAK_CONTROL_n45), .Z0_f (new_AGEMA_signal_2852) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) KECCAK_CONTROL_U39 ( .A0_t (Reset_t), .A0_f (Reset_f), .B0_t (KECCAK_CONTROL_n44), .B0_f (new_AGEMA_signal_4593), .Z0_t (KECCAK_CONTROL_RoundCountxDP[4]), .Z0_f (new_AGEMA_signal_2998) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b0)) KECCAK_CONTROL_U38 ( .A0_t (KECCAK_CONTROL_RoundCountxDP[4]), .A0_f (new_AGEMA_signal_2998), .B0_t (KECCAK_CONTROL_n43), .B0_f (new_AGEMA_signal_3988), .Z0_t (KECCAK_CONTROL_n44), .Z0_f (new_AGEMA_signal_4593) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) KECCAK_CONTROL_U37 ( .A0_t (KECCAK_CONTROL_RoundCountxDP[4]), .A0_f (new_AGEMA_signal_2998), .B0_t (KECCAK_CONTROL_n34), .B0_f (new_AGEMA_signal_3378), .Z0_t (KECCAK_CONTROL_RoundCountLastxDP_reg_Q), .Z0_f (new_AGEMA_signal_2856) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_U36 ( .A0_t (Reset_t), .A0_f (Reset_f), .B0_t (KECCAK_CONTROL_n33), .B0_f (new_AGEMA_signal_3246), .Z0_t (KECCAK_CONTROL_n34), .Z0_f (new_AGEMA_signal_3378) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_U35 ( .A0_t (KECCAK_CONTROL_n32), .A0_f (new_AGEMA_signal_2990), .B0_t (KECCAK_CONTROL_RoundCountxDP[1]), .B0_f (new_AGEMA_signal_2863), .Z0_t (KECCAK_CONTROL_n33), .Z0_f (new_AGEMA_signal_3246) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_U34 ( .A0_t (KECCAK_CONTROL_RoundCountxDP[0]), .A0_f (new_AGEMA_signal_2989), .B0_t (KECCAK_CONTROL_n30), .B0_f (new_AGEMA_signal_2860), .Z0_t (KECCAK_CONTROL_n32), .Z0_f (new_AGEMA_signal_2990) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) KECCAK_CONTROL_U33 ( .A0_t (Reset_t), .A0_f (Reset_f), .B0_t (KECCAK_CONTROL_n29), .B0_f (new_AGEMA_signal_3247), .Z0_t (KECCAK_CONTROL_CtrlStatexDP[2]), .Z0_f (new_AGEMA_signal_2851) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_U32 ( .A0_t (KECCAK_CONTROL_CtrlStatexDP[2]), .A0_f (new_AGEMA_signal_2851), .B0_t (KECCAK_CONTROL_n28), .B0_f (new_AGEMA_signal_2991), .Z0_t (KECCAK_CONTROL_n29), .Z0_f (new_AGEMA_signal_3247) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_U31 ( .A0_t (KECCAK_CONTROL_n27), .A0_f (new_AGEMA_signal_2854), .B0_t (KECCAK_CONTROL_RoundCountLastxDP_reg_Q), .B0_f (new_AGEMA_signal_2856), .Z0_t (KECCAK_CONTROL_n28), .Z0_f (new_AGEMA_signal_2991) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_U30 ( .A0_t (KECCAK_CONTROL_CtrlStatexDP[0]), .A0_f (new_AGEMA_signal_2853), .B0_t (KECCAK_CONTROL_CtrlStatexDP_reg_1__Q), .B0_f (new_AGEMA_signal_2850), .Z0_t (KECCAK_CONTROL_n27), .Z0_f (new_AGEMA_signal_2854) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) KECCAK_CONTROL_U29 ( .A0_t (Reset_t), .A0_f (Reset_f), .B0_t (KECCAK_CONTROL_n25), .B0_f (new_AGEMA_signal_3986), .Z0_t (KECCAK_CONTROL_RoundCountxDP[2]), .Z0_f (new_AGEMA_signal_2859) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b0)) KECCAK_CONTROL_U28 ( .A0_t (KECCAK_CONTROL_RoundCountxDP[2]), .A0_f (new_AGEMA_signal_2859), .B0_t (KECCAK_CONTROL_n23), .B0_f (new_AGEMA_signal_3380), .Z0_t (KECCAK_CONTROL_n25), .Z0_f (new_AGEMA_signal_3986) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) KECCAK_CONTROL_U27 ( .A0_t (Reset_t), .A0_f (Reset_f), .B0_t (KECCAK_CONTROL_n22), .B0_f (new_AGEMA_signal_3248), .Z0_t (KECCAK_CONTROL_CtrlStatexDP_reg_1__Q), .Z0_f (new_AGEMA_signal_2850) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_U26 ( .A0_t (KECCAK_CONTROL_n21), .A0_f (new_AGEMA_signal_2992), .B0_t (KECCAK_CONTROL_n20), .B0_f (new_AGEMA_signal_2855), .Z0_t (KECCAK_CONTROL_n22), .Z0_f (new_AGEMA_signal_3248) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_U25 ( .A0_t (KECCAK_CONTROL_CtrlStatexDP[2]), .A0_f (new_AGEMA_signal_2851), .B0_t (KECCAK_CONTROL_CtrlStatexDP[0]), .B0_f (new_AGEMA_signal_2853), .Z0_t (KECCAK_CONTROL_n20), .Z0_f (new_AGEMA_signal_2855) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_U24 ( .A0_t (KECCAK_CONTROL_CtrlStatexDP_reg_1__Q), .A0_f (new_AGEMA_signal_2850), .B0_t (KECCAK_CONTROL_n19), .B0_f (new_AGEMA_signal_2857), .Z0_t (KECCAK_CONTROL_n21), .Z0_f (new_AGEMA_signal_2992) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_U23 ( .A0_t (KECCAK_CONTROL_CtrlStatexDP[2]), .A0_f (new_AGEMA_signal_2851), .B0_t (KECCAK_CONTROL_RoundCountLastxDP_reg_Q), .B0_f (new_AGEMA_signal_2856), .Z0_t (KECCAK_CONTROL_n19), .Z0_f (new_AGEMA_signal_2857) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) KECCAK_CONTROL_U22 ( .A0_t (Reset_t), .A0_f (Reset_f), .B0_t (KECCAK_CONTROL_n18), .B0_f (new_AGEMA_signal_3379), .Z0_t (KECCAK_CONTROL_RoundCountxDP[1]), .Z0_f (new_AGEMA_signal_2863) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) KECCAK_CONTROL_U21 ( .A0_t (KECCAK_CONTROL_n17), .A0_f (new_AGEMA_signal_3249), .B0_t (KECCAK_CONTROL_RoundCountxDP[1]), .B0_f (new_AGEMA_signal_2863), .Z0_t (KECCAK_CONTROL_n18), .Z0_f (new_AGEMA_signal_3379) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) KECCAK_CONTROL_U20 ( .A0_t (KECCAK_CONTROL_n16), .A0_f (new_AGEMA_signal_4595), .B0_t (KECCAK_CONTROL_n15), .B0_f (new_AGEMA_signal_4594), .Z0_t (KECCAK_CONTROL_RoundCountxDP[3]), .Z0_f (new_AGEMA_signal_2858) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_U19 ( .A0_t (KECCAK_CONTROL_RoundCountxDP[3]), .A0_f (new_AGEMA_signal_2858), .B0_t (KECCAK_CONTROL_n14), .B0_f (new_AGEMA_signal_3987), .Z0_t (KECCAK_CONTROL_n15), .Z0_f (new_AGEMA_signal_4594) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_U18 ( .A0_t (KECCAK_CONTROL_RoundCountxDP[2]), .A0_f (new_AGEMA_signal_2859), .B0_t (KECCAK_CONTROL_n23), .B0_f (new_AGEMA_signal_3380), .Z0_t (KECCAK_CONTROL_n14), .Z0_f (new_AGEMA_signal_3987) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_U16 ( .A0_t (Reset_t), .A0_f (Reset_f), .B0_t (KECCAK_CONTROL_n43), .B0_f (new_AGEMA_signal_3988), .Z0_t (KECCAK_CONTROL_n16), .Z0_f (new_AGEMA_signal_4595) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_U15 ( .A0_t (KECCAK_CONTROL_n30), .A0_f (new_AGEMA_signal_2860), .B0_t (KECCAK_CONTROL_n23), .B0_f (new_AGEMA_signal_3380), .Z0_t (KECCAK_CONTROL_n43), .Z0_f (new_AGEMA_signal_3988) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_U14 ( .A0_t (KECCAK_CONTROL_n17), .A0_f (new_AGEMA_signal_3249), .B0_t (KECCAK_CONTROL_RoundCountxDP[1]), .B0_f (new_AGEMA_signal_2863), .Z0_t (KECCAK_CONTROL_n23), .Z0_f (new_AGEMA_signal_3380) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_U12 ( .A0_t (KECCAK_CONTROL_n13), .A0_f (new_AGEMA_signal_2993), .B0_t (KECCAK_CONTROL_RoundCountxDP[0]), .B0_f (new_AGEMA_signal_2989), .Z0_t (KECCAK_CONTROL_n17), .Z0_f (new_AGEMA_signal_3249) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_U11 ( .A0_t (KECCAK_CONTROL_RoundCountxDP[3]), .A0_f (new_AGEMA_signal_2858), .B0_t (KECCAK_CONTROL_RoundCountxDP[2]), .B0_f (new_AGEMA_signal_2859), .Z0_t (KECCAK_CONTROL_n30), .Z0_f (new_AGEMA_signal_2860) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) KECCAK_CONTROL_U9 ( .A0_t (Reset_t), .A0_f (Reset_f), .B0_t (KECCAK_CONTROL_n11), .B0_f (new_AGEMA_signal_3250), .Z0_t (KECCAK_CONTROL_RoundCountxDP[0]), .Z0_f (new_AGEMA_signal_2989) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b0)) KECCAK_CONTROL_U8 ( .A0_t (KECCAK_CONTROL_RoundCountxDP[0]), .A0_f (new_AGEMA_signal_2989), .B0_t (KECCAK_CONTROL_n13), .B0_f (new_AGEMA_signal_2993), .Z0_t (KECCAK_CONTROL_n11), .Z0_f (new_AGEMA_signal_3250) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_U7 ( .A0_t (KECCAK_CONTROL_n10), .A0_f (new_AGEMA_signal_2861), .B0_t (KECCAK_CONTROL_CtrlStatexDP[2]), .B0_f (new_AGEMA_signal_2851), .Z0_t (KECCAK_CONTROL_n13), .Z0_f (new_AGEMA_signal_2993) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b0)) KECCAK_CONTROL_U5 ( .A0_t (KECCAK_CONTROL_CtrlStatexDP[0]), .A0_f (new_AGEMA_signal_2853), .B0_t (KECCAK_CONTROL_CtrlStatexDP_reg_1__Q), .B0_f (new_AGEMA_signal_2850), .Z0_t (KECCAK_CONTROL_n10), .Z0_f (new_AGEMA_signal_2861) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_U2 ( .A0_t (KECCAK_CONTROL_CtrlStatexDP[2]), .A0_f (new_AGEMA_signal_2851), .B0_t (KECCAK_CONTROL_n8), .B0_f (new_AGEMA_signal_2862), .Z0_t (Ready_t), .Z0_f (Ready_f) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_U1 ( .A0_t (KECCAK_CONTROL_CtrlStatexDP_reg_1__Q), .A0_f (new_AGEMA_signal_2850), .B0_t (KECCAK_CONTROL_CtrlStatexDP[0]), .B0_f (new_AGEMA_signal_2853), .Z0_t (KECCAK_CONTROL_n8), .Z0_f (new_AGEMA_signal_2862) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_RC_GEN_U35 ( .A0_t (KECCAK_CONTROL_RC_GEN_n3), .A0_f (new_AGEMA_signal_2865), .B0_t (KECCAK_CONTROL_RC_GEN_n28), .B0_f (new_AGEMA_signal_3251), .Z0_t (KECCAK_CONTROL_RC_GEN_n24), .Z0_f (new_AGEMA_signal_3381) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_RC_GEN_U34 ( .A0_t (KECCAK_CONTROL_RC_GEN_n27), .A0_f (new_AGEMA_signal_2864), .B0_t (KECCAK_CONTROL_RC_GEN_n26), .B0_f (new_AGEMA_signal_3002), .Z0_t (KECCAK_CONTROL_RC_GEN_n28), .Z0_f (new_AGEMA_signal_3251) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_RC_GEN_U33 ( .A0_t (KECCAK_CONTROL_RoundCountxDP[4]), .A0_f (new_AGEMA_signal_2998), .B0_t (KECCAK_CONTROL_RC_GEN_n25), .B0_f (new_AGEMA_signal_3989), .Z0_t (IotaRC_3), .Z0_f (new_AGEMA_signal_4596) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_RC_GEN_U31 ( .A0_t (KECCAK_CONTROL_RC_GEN_n22), .A0_f (new_AGEMA_signal_3383), .B0_t (KECCAK_CONTROL_RC_GEN_n19), .B0_f (new_AGEMA_signal_3382), .Z0_t (KECCAK_CONTROL_RC_GEN_n25), .Z0_f (new_AGEMA_signal_3989) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_RC_GEN_U30 ( .A0_t (KECCAK_CONTROL_RoundCountxDP[0]), .A0_f (new_AGEMA_signal_2989), .B0_t (KECCAK_CONTROL_RC_GEN_n18), .B0_f (new_AGEMA_signal_3252), .Z0_t (KECCAK_CONTROL_RC_GEN_n19), .Z0_f (new_AGEMA_signal_3382) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_RC_GEN_U29 ( .A0_t (KECCAK_CONTROL_RoundCountxDP[3]), .A0_f (new_AGEMA_signal_2858), .B0_t (KECCAK_CONTROL_RC_GEN_n17), .B0_f (new_AGEMA_signal_2995), .Z0_t (KECCAK_CONTROL_RC_GEN_n18), .Z0_f (new_AGEMA_signal_3252) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_RC_GEN_U27 ( .A0_t (KECCAK_CONTROL_RC_GEN_n27), .A0_f (new_AGEMA_signal_2864), .B0_t (KECCAK_CONTROL_RC_GEN_n15), .B0_f (new_AGEMA_signal_2867), .Z0_t (KECCAK_CONTROL_RC_GEN_n17), .Z0_f (new_AGEMA_signal_2995) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_RC_GEN_U24 ( .A0_t (KECCAK_CONTROL_RC_GEN_n14), .A0_f (new_AGEMA_signal_3253), .B0_t (KECCAK_CONTROL_RC_GEN_n13), .B0_f (new_AGEMA_signal_2996), .Z0_t (KECCAK_CONTROL_RC_GEN_n22), .Z0_f (new_AGEMA_signal_3383) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_RC_GEN_U23 ( .A0_t (KECCAK_CONTROL_RoundCountxDP[3]), .A0_f (new_AGEMA_signal_2858), .B0_t (KECCAK_CONTROL_RC_GEN_n27), .B0_f (new_AGEMA_signal_2864), .Z0_t (KECCAK_CONTROL_RC_GEN_n13), .Z0_f (new_AGEMA_signal_2996) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_RC_GEN_U22 ( .A0_t (KECCAK_CONTROL_RoundCountxDP[2]), .A0_f (new_AGEMA_signal_2859), .B0_t (KECCAK_CONTROL_RoundCountxDP[1]), .B0_f (new_AGEMA_signal_2863), .Z0_t (KECCAK_CONTROL_RC_GEN_n27), .Z0_f (new_AGEMA_signal_2864) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_RC_GEN_U21 ( .A0_t (KECCAK_CONTROL_RoundCountxDP[2]), .A0_f (new_AGEMA_signal_2859), .B0_t (KECCAK_CONTROL_RC_GEN_n12), .B0_f (new_AGEMA_signal_2997), .Z0_t (KECCAK_CONTROL_RC_GEN_n14), .Z0_f (new_AGEMA_signal_3253) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_RC_GEN_U20 ( .A0_t (KECCAK_CONTROL_RC_GEN_n11), .A0_f (new_AGEMA_signal_2866), .B0_t (KECCAK_CONTROL_RoundCountxDP[0]), .B0_f (new_AGEMA_signal_2989), .Z0_t (KECCAK_CONTROL_RC_GEN_n12), .Z0_f (new_AGEMA_signal_2997) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_RC_GEN_U18 ( .A0_t (KECCAK_CONTROL_RoundCountxDP[0]), .A0_f (new_AGEMA_signal_2989), .B0_t (KECCAK_CONTROL_RC_GEN_n9), .B0_f (new_AGEMA_signal_3000), .Z0_t (KECCAK_CONTROL_RC_GEN_n30), .Z0_f (new_AGEMA_signal_3254) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_RC_GEN_U17 ( .A0_t (KECCAK_CONTROL_RC_GEN_n9), .A0_f (new_AGEMA_signal_3000), .B0_t (KECCAK_CONTROL_RC_GEN_n8), .B0_f (new_AGEMA_signal_2999), .Z0_t (KECCAK_CONTROL_RC_GEN_n20), .Z0_f (new_AGEMA_signal_3255) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_RC_GEN_U16 ( .A0_t (KECCAK_CONTROL_RC_GEN_n3), .A0_f (new_AGEMA_signal_2865), .B0_t (KECCAK_CONTROL_RoundCountxDP[4]), .B0_f (new_AGEMA_signal_2998), .Z0_t (KECCAK_CONTROL_RC_GEN_n8), .Z0_f (new_AGEMA_signal_2999) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_RC_GEN_U15 ( .A0_t (KECCAK_CONTROL_RC_GEN_n15), .A0_f (new_AGEMA_signal_2867), .B0_t (KECCAK_CONTROL_RoundCountxDP[3]), .B0_f (new_AGEMA_signal_2858), .Z0_t (KECCAK_CONTROL_RC_GEN_n9), .Z0_f (new_AGEMA_signal_3000) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_RC_GEN_U14 ( .A0_t (KECCAK_CONTROL_RoundCountxDP[4]), .A0_f (new_AGEMA_signal_2998), .B0_t (KECCAK_CONTROL_RC_GEN_n6), .B0_f (new_AGEMA_signal_3384), .Z0_t (IotaRC[0]), .Z0_f (new_AGEMA_signal_3990) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_RC_GEN_U13 ( .A0_t (KECCAK_CONTROL_RoundCountxDP[2]), .A0_f (new_AGEMA_signal_2859), .B0_t (KECCAK_CONTROL_RC_GEN_n5), .B0_f (new_AGEMA_signal_3256), .Z0_t (KECCAK_CONTROL_RC_GEN_n6), .Z0_f (new_AGEMA_signal_3384) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_RC_GEN_U12 ( .A0_t (KECCAK_CONTROL_RC_GEN_n4), .A0_f (new_AGEMA_signal_3001), .B0_t (KECCAK_CONTROL_RoundCountxDP[0]), .B0_f (new_AGEMA_signal_2989), .Z0_t (KECCAK_CONTROL_RC_GEN_n5), .Z0_f (new_AGEMA_signal_3256) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_RC_GEN_U11 ( .A0_t (KECCAK_CONTROL_RC_GEN_n11), .A0_f (new_AGEMA_signal_2866), .B0_t (KECCAK_CONTROL_RC_GEN_n3), .B0_f (new_AGEMA_signal_2865), .Z0_t (KECCAK_CONTROL_RC_GEN_n4), .Z0_f (new_AGEMA_signal_3001) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_RC_GEN_U9 ( .A0_t (KECCAK_CONTROL_RoundCountxDP[4]), .A0_f (new_AGEMA_signal_2998), .B0_t (KECCAK_CONTROL_RC_GEN_n2), .B0_f (new_AGEMA_signal_3257), .Z0_t (KECCAK_CONTROL_RC_GEN_n21), .Z0_f (new_AGEMA_signal_3385) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_RC_GEN_U8 ( .A0_t (KECCAK_CONTROL_RC_GEN_n26), .A0_f (new_AGEMA_signal_3002), .B0_t (KECCAK_CONTROL_RC_GEN_n3), .B0_f (new_AGEMA_signal_2865), .Z0_t (KECCAK_CONTROL_RC_GEN_n2), .Z0_f (new_AGEMA_signal_3257) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_RC_GEN_U7 ( .A0_t (KECCAK_CONTROL_RoundCountxDP[3]), .A0_f (new_AGEMA_signal_2858), .B0_t (KECCAK_CONTROL_RoundCountxDP[1]), .B0_f (new_AGEMA_signal_2863), .Z0_t (KECCAK_CONTROL_RC_GEN_n3), .Z0_f (new_AGEMA_signal_2865) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_RC_GEN_U6 ( .A0_t (KECCAK_CONTROL_RoundCountxDP[2]), .A0_f (new_AGEMA_signal_2859), .B0_t (KECCAK_CONTROL_RC_GEN_n11), .B0_f (new_AGEMA_signal_2866), .Z0_t (KECCAK_CONTROL_RC_GEN_n26), .Z0_f (new_AGEMA_signal_3002) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_RC_GEN_U5 ( .A0_t (KECCAK_CONTROL_RoundCountxDP[1]), .A0_f (new_AGEMA_signal_2863), .B0_t (KECCAK_CONTROL_RoundCountxDP[3]), .B0_f (new_AGEMA_signal_2858), .Z0_t (KECCAK_CONTROL_RC_GEN_n11), .Z0_f (new_AGEMA_signal_2866) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) KECCAK_CONTROL_RC_GEN_U2 ( .A0_t (KECCAK_CONTROL_RC_GEN_n15), .A0_f (new_AGEMA_signal_2867), .B0_t (KECCAK_CONTROL_RoundCountxDP[3]), .B0_f (new_AGEMA_signal_2858), .Z0_t (KECCAK_CONTROL_RC_GEN_n23), .Z0_f (new_AGEMA_signal_3003) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_RC_GEN_U1 ( .A0_t (KECCAK_CONTROL_RoundCountxDP[2]), .A0_f (new_AGEMA_signal_2859), .B0_t (KECCAK_CONTROL_RoundCountxDP[1]), .B0_f (new_AGEMA_signal_2863), .Z0_t (KECCAK_CONTROL_RC_GEN_n15), .Z0_f (new_AGEMA_signal_2867) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) KECCAK_CONTROL_RC_GEN_U25_XOR1_U1 ( .A0_t (KECCAK_CONTROL_RC_GEN_n21), .A0_f (new_AGEMA_signal_3385), .B0_t (KECCAK_CONTROL_RC_GEN_n20), .B0_f (new_AGEMA_signal_3255), .Z0_t (KECCAK_CONTROL_RC_GEN_U25_X), .Z0_f (new_AGEMA_signal_3991) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_RC_GEN_U25_AND1_U1 ( .A0_t (KECCAK_CONTROL_RoundCountxDP[0]), .A0_f (new_AGEMA_signal_2989), .B0_t (KECCAK_CONTROL_RC_GEN_U25_X), .B0_f (new_AGEMA_signal_3991), .Z0_t (KECCAK_CONTROL_RC_GEN_U25_Y), .Z0_f (new_AGEMA_signal_4597) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) KECCAK_CONTROL_RC_GEN_U25_XOR2_U1 ( .A0_t (KECCAK_CONTROL_RC_GEN_U25_Y), .A0_f (new_AGEMA_signal_4597), .B0_t (KECCAK_CONTROL_RC_GEN_n21), .B0_f (new_AGEMA_signal_3385), .Z0_t (IotaRC_7), .Z0_f (new_AGEMA_signal_5199) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) KECCAK_CONTROL_RC_GEN_U28_XOR1_U1 ( .A0_t (KECCAK_CONTROL_RC_GEN_n24), .A0_f (new_AGEMA_signal_3381), .B0_t (KECCAK_CONTROL_RC_GEN_n23), .B0_f (new_AGEMA_signal_3003), .Z0_t (KECCAK_CONTROL_RC_GEN_U28_X), .Z0_f (new_AGEMA_signal_3992) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_RC_GEN_U28_AND1_U1 ( .A0_t (KECCAK_CONTROL_RoundCountxDP[0]), .A0_f (new_AGEMA_signal_2989), .B0_t (KECCAK_CONTROL_RC_GEN_U28_X), .B0_f (new_AGEMA_signal_3992), .Z0_t (KECCAK_CONTROL_RC_GEN_U28_Y), .Z0_f (new_AGEMA_signal_4598) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) KECCAK_CONTROL_RC_GEN_U28_XOR2_U1 ( .A0_t (KECCAK_CONTROL_RC_GEN_U28_Y), .A0_f (new_AGEMA_signal_4598), .B0_t (KECCAK_CONTROL_RC_GEN_n24), .B0_f (new_AGEMA_signal_3381), .Z0_t (KECCAK_CONTROL_RC_GEN_n31), .Z0_f (new_AGEMA_signal_5200) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) KECCAK_CONTROL_RC_GEN_U32_XOR1_U1 ( .A0_t (KECCAK_CONTROL_RC_GEN_n31), .A0_f (new_AGEMA_signal_5200), .B0_t (KECCAK_CONTROL_RC_GEN_n30), .B0_f (new_AGEMA_signal_3254), .Z0_t (KECCAK_CONTROL_RC_GEN_U32_X), .Z0_f (new_AGEMA_signal_5210) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_RC_GEN_U32_AND1_U1 ( .A0_t (KECCAK_CONTROL_RoundCountxDP[4]), .A0_f (new_AGEMA_signal_2998), .B0_t (KECCAK_CONTROL_RC_GEN_U32_X), .B0_f (new_AGEMA_signal_5210), .Z0_t (KECCAK_CONTROL_RC_GEN_U32_Y), .Z0_f (new_AGEMA_signal_5823) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) KECCAK_CONTROL_RC_GEN_U32_XOR2_U1 ( .A0_t (KECCAK_CONTROL_RC_GEN_U32_Y), .A0_f (new_AGEMA_signal_5823), .B0_t (KECCAK_CONTROL_RC_GEN_n31), .B0_f (new_AGEMA_signal_5200), .Z0_t (IotaRC[1]), .Z0_f (new_AGEMA_signal_6421) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U810_XOR1_U1 ( .A0_t (StateOut[11]), .A0_f (new_AGEMA_signal_2184), .A1_t (new_AGEMA_signal_2185), .A1_f (new_AGEMA_signal_2186), .B0_t (StateFromChi[3]), .B0_f (new_AGEMA_signal_5207), .B1_t (new_AGEMA_signal_5208), .B1_f (new_AGEMA_signal_5209), .Z0_t (U810_X), .Z0_f (new_AGEMA_signal_5824), .Z1_t (new_AGEMA_signal_5825), .Z1_f (new_AGEMA_signal_5826) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U810_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U810_X), .B0_f (new_AGEMA_signal_5824), .B1_t (new_AGEMA_signal_5825), .B1_f (new_AGEMA_signal_5826), .Z0_t (U810_Y), .Z0_f (new_AGEMA_signal_6422), .Z1_t (new_AGEMA_signal_6423), .Z1_f (new_AGEMA_signal_6424) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U810_XOR2_U1 ( .A0_t (U810_Y), .A0_f (new_AGEMA_signal_6422), .A1_t (new_AGEMA_signal_6423), .A1_f (new_AGEMA_signal_6424), .B0_t (StateOut[11]), .B0_f (new_AGEMA_signal_2184), .B1_t (new_AGEMA_signal_2185), .B1_f (new_AGEMA_signal_2186), .Z0_t (OutData_s0_t[3]), .Z0_f (OutData_s0_f[3]), .Z1_t (OutData_s1_t[3]), .Z1_f (OutData_s1_f[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U812_XOR1_U1 ( .A0_t (StateOut[15]), .A0_f (new_AGEMA_signal_2346), .A1_t (new_AGEMA_signal_2347), .A1_f (new_AGEMA_signal_2348), .B0_t (StateFromChi[7]), .B0_f (new_AGEMA_signal_5204), .B1_t (new_AGEMA_signal_5205), .B1_f (new_AGEMA_signal_5206), .Z0_t (U812_X), .Z0_f (new_AGEMA_signal_5827), .Z1_t (new_AGEMA_signal_5828), .Z1_f (new_AGEMA_signal_5829) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U812_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U812_X), .B0_f (new_AGEMA_signal_5827), .B1_t (new_AGEMA_signal_5828), .B1_f (new_AGEMA_signal_5829), .Z0_t (U812_Y), .Z0_f (new_AGEMA_signal_6425), .Z1_t (new_AGEMA_signal_6426), .Z1_f (new_AGEMA_signal_6427) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U812_XOR2_U1 ( .A0_t (U812_Y), .A0_f (new_AGEMA_signal_6425), .A1_t (new_AGEMA_signal_6426), .A1_f (new_AGEMA_signal_6427), .B0_t (StateOut[15]), .B0_f (new_AGEMA_signal_2346), .B1_t (new_AGEMA_signal_2347), .B1_f (new_AGEMA_signal_2348), .Z0_t (OutData_s0_t[7]), .Z0_f (OutData_s0_f[7]), .Z1_t (OutData_s1_t[7]), .Z1_f (OutData_s1_f[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U814_XOR1_U1 ( .A0_t (StateOut[8]), .A0_f (new_AGEMA_signal_2202), .A1_t (new_AGEMA_signal_2203), .A1_f (new_AGEMA_signal_2204), .B0_t (StateFromChi[0]), .B0_f (new_AGEMA_signal_5201), .B1_t (new_AGEMA_signal_5202), .B1_f (new_AGEMA_signal_5203), .Z0_t (U814_X), .Z0_f (new_AGEMA_signal_5830), .Z1_t (new_AGEMA_signal_5831), .Z1_f (new_AGEMA_signal_5832) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U814_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U814_X), .B0_f (new_AGEMA_signal_5830), .B1_t (new_AGEMA_signal_5831), .B1_f (new_AGEMA_signal_5832), .Z0_t (U814_Y), .Z0_f (new_AGEMA_signal_6428), .Z1_t (new_AGEMA_signal_6429), .Z1_f (new_AGEMA_signal_6430) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U814_XOR2_U1 ( .A0_t (U814_Y), .A0_f (new_AGEMA_signal_6428), .A1_t (new_AGEMA_signal_6429), .A1_f (new_AGEMA_signal_6430), .B0_t (StateOut[8]), .B0_f (new_AGEMA_signal_2202), .B1_t (new_AGEMA_signal_2203), .B1_f (new_AGEMA_signal_2204), .Z0_t (OutData_s0_t[0]), .Z0_f (OutData_s0_f[0]), .Z1_t (OutData_s1_t[0]), .Z1_f (OutData_s1_f[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U816_XOR1_U1 ( .A0_t (StateOut[9]), .A0_f (new_AGEMA_signal_2760), .A1_t (new_AGEMA_signal_2761), .A1_f (new_AGEMA_signal_2762), .B0_t (StateFromChi[1]), .B0_f (new_AGEMA_signal_6431), .B1_t (new_AGEMA_signal_6432), .B1_f (new_AGEMA_signal_6433), .Z0_t (U816_X), .Z0_f (new_AGEMA_signal_6434), .Z1_t (new_AGEMA_signal_6435), .Z1_f (new_AGEMA_signal_6436) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U816_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U816_X), .B0_f (new_AGEMA_signal_6434), .B1_t (new_AGEMA_signal_6435), .B1_f (new_AGEMA_signal_6436), .Z0_t (U816_Y), .Z0_f (new_AGEMA_signal_6437), .Z1_t (new_AGEMA_signal_6438), .Z1_f (new_AGEMA_signal_6439) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U816_XOR2_U1 ( .A0_t (U816_Y), .A0_f (new_AGEMA_signal_6437), .A1_t (new_AGEMA_signal_6438), .A1_f (new_AGEMA_signal_6439), .B0_t (StateOut[9]), .B0_f (new_AGEMA_signal_2760), .B1_t (new_AGEMA_signal_2761), .B1_f (new_AGEMA_signal_2762), .Z0_t (OutData_s0_t[1]), .Z0_f (OutData_s0_f[1]), .Z1_t (OutData_s1_t[1]), .Z1_f (OutData_s1_f[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U817_XOR1_U1 ( .A0_t (StateOut[47]), .A0_f (new_AGEMA_signal_3072), .A1_t (new_AGEMA_signal_3073), .A1_f (new_AGEMA_signal_3074), .B0_t (StateFromChi[39]), .B0_f (new_AGEMA_signal_5184), .B1_t (new_AGEMA_signal_5185), .B1_f (new_AGEMA_signal_5186), .Z0_t (U817_X), .Z0_f (new_AGEMA_signal_5211), .Z1_t (new_AGEMA_signal_5212), .Z1_f (new_AGEMA_signal_5213) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U817_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U817_X), .B0_f (new_AGEMA_signal_5211), .B1_t (new_AGEMA_signal_5212), .B1_f (new_AGEMA_signal_5213), .Z0_t (U817_Y), .Z0_f (new_AGEMA_signal_5833), .Z1_t (new_AGEMA_signal_5834), .Z1_f (new_AGEMA_signal_5835) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U817_XOR2_U1 ( .A0_t (U817_Y), .A0_f (new_AGEMA_signal_5833), .A1_t (new_AGEMA_signal_5834), .A1_f (new_AGEMA_signal_5835), .B0_t (StateOut[47]), .B0_f (new_AGEMA_signal_3072), .B1_t (new_AGEMA_signal_3073), .B1_f (new_AGEMA_signal_3074), .Z0_t (StateOut[39]), .Z0_f (new_AGEMA_signal_2355), .Z1_t (new_AGEMA_signal_2356), .Z1_f (new_AGEMA_signal_2357) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U818_XOR1_U1 ( .A0_t (StateOut[71]), .A0_f (new_AGEMA_signal_2340), .A1_t (new_AGEMA_signal_2341), .A1_f (new_AGEMA_signal_2342), .B0_t (StateFromChi[63]), .B0_f (new_AGEMA_signal_5157), .B1_t (new_AGEMA_signal_5158), .B1_f (new_AGEMA_signal_5159), .Z0_t (U818_X), .Z0_f (new_AGEMA_signal_5214), .Z1_t (new_AGEMA_signal_5215), .Z1_f (new_AGEMA_signal_5216) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U818_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U818_X), .B0_f (new_AGEMA_signal_5214), .B1_t (new_AGEMA_signal_5215), .B1_f (new_AGEMA_signal_5216), .Z0_t (U818_Y), .Z0_f (new_AGEMA_signal_5836), .Z1_t (new_AGEMA_signal_5837), .Z1_f (new_AGEMA_signal_5838) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U818_XOR2_U1 ( .A0_t (U818_Y), .A0_f (new_AGEMA_signal_5836), .A1_t (new_AGEMA_signal_5837), .A1_f (new_AGEMA_signal_5838), .B0_t (StateOut[71]), .B0_f (new_AGEMA_signal_2340), .B1_t (new_AGEMA_signal_2341), .B1_f (new_AGEMA_signal_2342), .Z0_t (StateOut[63]), .Z0_f (new_AGEMA_signal_2331), .Z1_t (new_AGEMA_signal_2332), .Z1_f (new_AGEMA_signal_2333) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U820_XOR1_U1 ( .A0_t (StateOut[95]), .A0_f (new_AGEMA_signal_2472), .A1_t (new_AGEMA_signal_2473), .A1_f (new_AGEMA_signal_2474), .B0_t (StateFromChi[87]), .B0_f (new_AGEMA_signal_5130), .B1_t (new_AGEMA_signal_5131), .B1_f (new_AGEMA_signal_5132), .Z0_t (U820_X), .Z0_f (new_AGEMA_signal_5217), .Z1_t (new_AGEMA_signal_5218), .Z1_f (new_AGEMA_signal_5219) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U820_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U820_X), .B0_f (new_AGEMA_signal_5217), .B1_t (new_AGEMA_signal_5218), .B1_f (new_AGEMA_signal_5219), .Z0_t (U820_Y), .Z0_f (new_AGEMA_signal_5839), .Z1_t (new_AGEMA_signal_5840), .Z1_f (new_AGEMA_signal_5841) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U820_XOR2_U1 ( .A0_t (U820_Y), .A0_f (new_AGEMA_signal_5839), .A1_t (new_AGEMA_signal_5840), .A1_f (new_AGEMA_signal_5841), .B0_t (StateOut[95]), .B0_f (new_AGEMA_signal_2472), .B1_t (new_AGEMA_signal_2473), .B1_f (new_AGEMA_signal_2474), .Z0_t (StateOut[87]), .Z0_f (new_AGEMA_signal_2475), .Z1_t (new_AGEMA_signal_2476), .Z1_f (new_AGEMA_signal_2477) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U821_XOR1_U1 ( .A0_t (StateOut[127]), .A0_f (new_AGEMA_signal_3012), .A1_t (new_AGEMA_signal_3013), .A1_f (new_AGEMA_signal_3014), .B0_t (StateFromChi[119]), .B0_f (new_AGEMA_signal_5190), .B1_t (new_AGEMA_signal_5191), .B1_f (new_AGEMA_signal_5192), .Z0_t (U821_X), .Z0_f (new_AGEMA_signal_5220), .Z1_t (new_AGEMA_signal_5221), .Z1_f (new_AGEMA_signal_5222) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U821_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U821_X), .B0_f (new_AGEMA_signal_5220), .B1_t (new_AGEMA_signal_5221), .B1_f (new_AGEMA_signal_5222), .Z0_t (U821_Y), .Z0_f (new_AGEMA_signal_5842), .Z1_t (new_AGEMA_signal_5843), .Z1_f (new_AGEMA_signal_5844) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U821_XOR2_U1 ( .A0_t (U821_Y), .A0_f (new_AGEMA_signal_5842), .A1_t (new_AGEMA_signal_5843), .A1_f (new_AGEMA_signal_5844), .B0_t (StateOut[127]), .B0_f (new_AGEMA_signal_3012), .B1_t (new_AGEMA_signal_3013), .B1_f (new_AGEMA_signal_3014), .Z0_t (StateOut[119]), .Z0_f (new_AGEMA_signal_2484), .Z1_t (new_AGEMA_signal_2485), .Z1_f (new_AGEMA_signal_2486) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U822_XOR1_U1 ( .A0_t (StateOut[151]), .A0_f (new_AGEMA_signal_2160), .A1_t (new_AGEMA_signal_2161), .A1_f (new_AGEMA_signal_2162), .B0_t (StateFromChi[143]), .B0_f (new_AGEMA_signal_5163), .B1_t (new_AGEMA_signal_5164), .B1_f (new_AGEMA_signal_5165), .Z0_t (U822_X), .Z0_f (new_AGEMA_signal_5223), .Z1_t (new_AGEMA_signal_5224), .Z1_f (new_AGEMA_signal_5225) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U822_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U822_X), .B0_f (new_AGEMA_signal_5223), .B1_t (new_AGEMA_signal_5224), .B1_f (new_AGEMA_signal_5225), .Z0_t (U822_Y), .Z0_f (new_AGEMA_signal_5845), .Z1_t (new_AGEMA_signal_5846), .Z1_f (new_AGEMA_signal_5847) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U822_XOR2_U1 ( .A0_t (U822_Y), .A0_f (new_AGEMA_signal_5845), .A1_t (new_AGEMA_signal_5846), .A1_f (new_AGEMA_signal_5847), .B0_t (StateOut[151]), .B0_f (new_AGEMA_signal_2160), .B1_t (new_AGEMA_signal_2161), .B1_f (new_AGEMA_signal_2162), .Z0_t (StateOut[143]), .Z0_f (new_AGEMA_signal_2151), .Z1_t (new_AGEMA_signal_2152), .Z1_f (new_AGEMA_signal_2153) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U823_XOR1_U1 ( .A0_t (StateOut[159]), .A0_f (new_AGEMA_signal_2157), .A1_t (new_AGEMA_signal_2158), .A1_f (new_AGEMA_signal_2159), .B0_t (StateFromChi[151]), .B0_f (new_AGEMA_signal_5178), .B1_t (new_AGEMA_signal_5179), .B1_f (new_AGEMA_signal_5180), .Z0_t (U823_X), .Z0_f (new_AGEMA_signal_5226), .Z1_t (new_AGEMA_signal_5227), .Z1_f (new_AGEMA_signal_5228) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U823_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U823_X), .B0_f (new_AGEMA_signal_5226), .B1_t (new_AGEMA_signal_5227), .B1_f (new_AGEMA_signal_5228), .Z0_t (U823_Y), .Z0_f (new_AGEMA_signal_5848), .Z1_t (new_AGEMA_signal_5849), .Z1_f (new_AGEMA_signal_5850) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U823_XOR2_U1 ( .A0_t (U823_Y), .A0_f (new_AGEMA_signal_5848), .A1_t (new_AGEMA_signal_5849), .A1_f (new_AGEMA_signal_5850), .B0_t (StateOut[159]), .B0_f (new_AGEMA_signal_2157), .B1_t (new_AGEMA_signal_2158), .B1_f (new_AGEMA_signal_2159), .Z0_t (StateOut[151]), .Z0_f (new_AGEMA_signal_2160), .Z1_t (new_AGEMA_signal_2161), .Z1_f (new_AGEMA_signal_2162) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U824_XOR1_U1 ( .A0_t (StateOut[175]), .A0_f (new_AGEMA_signal_2436), .A1_t (new_AGEMA_signal_2437), .A1_f (new_AGEMA_signal_2438), .B0_t (StateFromChi[167]), .B0_f (new_AGEMA_signal_5136), .B1_t (new_AGEMA_signal_5137), .B1_f (new_AGEMA_signal_5138), .Z0_t (U824_X), .Z0_f (new_AGEMA_signal_5229), .Z1_t (new_AGEMA_signal_5230), .Z1_f (new_AGEMA_signal_5231) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U824_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U824_X), .B0_f (new_AGEMA_signal_5229), .B1_t (new_AGEMA_signal_5230), .B1_f (new_AGEMA_signal_5231), .Z0_t (U824_Y), .Z0_f (new_AGEMA_signal_5851), .Z1_t (new_AGEMA_signal_5852), .Z1_f (new_AGEMA_signal_5853) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U824_XOR2_U1 ( .A0_t (U824_Y), .A0_f (new_AGEMA_signal_5851), .A1_t (new_AGEMA_signal_5852), .A1_f (new_AGEMA_signal_5853), .B0_t (StateOut[175]), .B0_f (new_AGEMA_signal_2436), .B1_t (new_AGEMA_signal_2437), .B1_f (new_AGEMA_signal_2438), .Z0_t (StateOut[167]), .Z0_f (new_AGEMA_signal_2439), .Z1_t (new_AGEMA_signal_2440), .Z1_f (new_AGEMA_signal_2441) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U825_XOR1_U1 ( .A0_t (StateOut[46]), .A0_f (new_AGEMA_signal_2457), .A1_t (new_AGEMA_signal_2458), .A1_f (new_AGEMA_signal_2459), .B0_t (StateFromChi[38]), .B0_f (new_AGEMA_signal_5109), .B1_t (new_AGEMA_signal_5110), .B1_f (new_AGEMA_signal_5111), .Z0_t (U825_X), .Z0_f (new_AGEMA_signal_5232), .Z1_t (new_AGEMA_signal_5233), .Z1_f (new_AGEMA_signal_5234) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U825_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U825_X), .B0_f (new_AGEMA_signal_5232), .B1_t (new_AGEMA_signal_5233), .B1_f (new_AGEMA_signal_5234), .Z0_t (U825_Y), .Z0_f (new_AGEMA_signal_5854), .Z1_t (new_AGEMA_signal_5855), .Z1_f (new_AGEMA_signal_5856) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U825_XOR2_U1 ( .A0_t (U825_Y), .A0_f (new_AGEMA_signal_5854), .A1_t (new_AGEMA_signal_5855), .A1_f (new_AGEMA_signal_5856), .B0_t (StateOut[46]), .B0_f (new_AGEMA_signal_2457), .B1_t (new_AGEMA_signal_2458), .B1_f (new_AGEMA_signal_2459), .Z0_t (StateOut[38]), .Z0_f (new_AGEMA_signal_2139), .Z1_t (new_AGEMA_signal_2140), .Z1_f (new_AGEMA_signal_2141) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U827_XOR1_U1 ( .A0_t (StateOut[70]), .A0_f (new_AGEMA_signal_2463), .A1_t (new_AGEMA_signal_2464), .A1_f (new_AGEMA_signal_2465), .B0_t (StateFromChi[62]), .B0_f (new_AGEMA_signal_5082), .B1_t (new_AGEMA_signal_5083), .B1_f (new_AGEMA_signal_5084), .Z0_t (U827_X), .Z0_f (new_AGEMA_signal_5235), .Z1_t (new_AGEMA_signal_5236), .Z1_f (new_AGEMA_signal_5237) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U827_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U827_X), .B0_f (new_AGEMA_signal_5235), .B1_t (new_AGEMA_signal_5236), .B1_f (new_AGEMA_signal_5237), .Z0_t (U827_Y), .Z0_f (new_AGEMA_signal_5857), .Z1_t (new_AGEMA_signal_5858), .Z1_f (new_AGEMA_signal_5859) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U827_XOR2_U1 ( .A0_t (U827_Y), .A0_f (new_AGEMA_signal_5857), .A1_t (new_AGEMA_signal_5858), .A1_f (new_AGEMA_signal_5859), .B0_t (StateOut[70]), .B0_f (new_AGEMA_signal_2463), .B1_t (new_AGEMA_signal_2464), .B1_f (new_AGEMA_signal_2465), .Z0_t (StateOut[62]), .Z0_f (new_AGEMA_signal_3114), .Z1_t (new_AGEMA_signal_3115), .Z1_f (new_AGEMA_signal_3116) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U828_XOR1_U1 ( .A0_t (StateOut[126]), .A0_f (new_AGEMA_signal_3018), .A1_t (new_AGEMA_signal_3019), .A1_f (new_AGEMA_signal_3020), .B0_t (StateFromChi[118]), .B0_f (new_AGEMA_signal_5115), .B1_t (new_AGEMA_signal_5116), .B1_f (new_AGEMA_signal_5117), .Z0_t (U828_X), .Z0_f (new_AGEMA_signal_5238), .Z1_t (new_AGEMA_signal_5239), .Z1_f (new_AGEMA_signal_5240) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U828_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U828_X), .B0_f (new_AGEMA_signal_5238), .B1_t (new_AGEMA_signal_5239), .B1_f (new_AGEMA_signal_5240), .Z0_t (U828_Y), .Z0_f (new_AGEMA_signal_5860), .Z1_t (new_AGEMA_signal_5861), .Z1_f (new_AGEMA_signal_5862) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U828_XOR2_U1 ( .A0_t (U828_Y), .A0_f (new_AGEMA_signal_5860), .A1_t (new_AGEMA_signal_5861), .A1_f (new_AGEMA_signal_5862), .B0_t (StateOut[126]), .B0_f (new_AGEMA_signal_3018), .B1_t (new_AGEMA_signal_3019), .B1_f (new_AGEMA_signal_3020), .Z0_t (StateOut[118]), .Z0_f (new_AGEMA_signal_2697), .Z1_t (new_AGEMA_signal_2698), .Z1_f (new_AGEMA_signal_2699) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U830_XOR1_U1 ( .A0_t (StateOut[150]), .A0_f (new_AGEMA_signal_2178), .A1_t (new_AGEMA_signal_2179), .A1_f (new_AGEMA_signal_2180), .B0_t (StateFromChi[142]), .B0_f (new_AGEMA_signal_5088), .B1_t (new_AGEMA_signal_5089), .B1_f (new_AGEMA_signal_5090), .Z0_t (U830_X), .Z0_f (new_AGEMA_signal_5241), .Z1_t (new_AGEMA_signal_5242), .Z1_f (new_AGEMA_signal_5243) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U830_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U830_X), .B0_f (new_AGEMA_signal_5241), .B1_t (new_AGEMA_signal_5242), .B1_f (new_AGEMA_signal_5243), .Z0_t (U830_Y), .Z0_f (new_AGEMA_signal_5863), .Z1_t (new_AGEMA_signal_5864), .Z1_f (new_AGEMA_signal_5865) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U830_XOR2_U1 ( .A0_t (U830_Y), .A0_f (new_AGEMA_signal_5863), .A1_t (new_AGEMA_signal_5864), .A1_f (new_AGEMA_signal_5865), .B0_t (StateOut[150]), .B0_f (new_AGEMA_signal_2178), .B1_t (new_AGEMA_signal_2179), .B1_f (new_AGEMA_signal_2180), .Z0_t (StateOut[142]), .Z0_f (new_AGEMA_signal_2169), .Z1_t (new_AGEMA_signal_2170), .Z1_f (new_AGEMA_signal_2171) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U831_XOR1_U1 ( .A0_t (StateOut[158]), .A0_f (new_AGEMA_signal_2175), .A1_t (new_AGEMA_signal_2176), .A1_f (new_AGEMA_signal_2177), .B0_t (StateFromChi[150]), .B0_f (new_AGEMA_signal_5103), .B1_t (new_AGEMA_signal_5104), .B1_f (new_AGEMA_signal_5105), .Z0_t (U831_X), .Z0_f (new_AGEMA_signal_5244), .Z1_t (new_AGEMA_signal_5245), .Z1_f (new_AGEMA_signal_5246) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U831_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U831_X), .B0_f (new_AGEMA_signal_5244), .B1_t (new_AGEMA_signal_5245), .B1_f (new_AGEMA_signal_5246), .Z0_t (U831_Y), .Z0_f (new_AGEMA_signal_5866), .Z1_t (new_AGEMA_signal_5867), .Z1_f (new_AGEMA_signal_5868) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U831_XOR2_U1 ( .A0_t (U831_Y), .A0_f (new_AGEMA_signal_5866), .A1_t (new_AGEMA_signal_5867), .A1_f (new_AGEMA_signal_5868), .B0_t (StateOut[158]), .B0_f (new_AGEMA_signal_2175), .B1_t (new_AGEMA_signal_2176), .B1_f (new_AGEMA_signal_2177), .Z0_t (StateOut[150]), .Z0_f (new_AGEMA_signal_2178), .Z1_t (new_AGEMA_signal_2179), .Z1_f (new_AGEMA_signal_2180) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U832_XOR1_U1 ( .A0_t (StateOut[174]), .A0_f (new_AGEMA_signal_2490), .A1_t (new_AGEMA_signal_2491), .A1_f (new_AGEMA_signal_2492), .B0_t (StateFromChi[166]), .B0_f (new_AGEMA_signal_5061), .B1_t (new_AGEMA_signal_5062), .B1_f (new_AGEMA_signal_5063), .Z0_t (U832_X), .Z0_f (new_AGEMA_signal_5247), .Z1_t (new_AGEMA_signal_5248), .Z1_f (new_AGEMA_signal_5249) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U832_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U832_X), .B0_f (new_AGEMA_signal_5247), .B1_t (new_AGEMA_signal_5248), .B1_f (new_AGEMA_signal_5249), .Z0_t (U832_Y), .Z0_f (new_AGEMA_signal_5869), .Z1_t (new_AGEMA_signal_5870), .Z1_f (new_AGEMA_signal_5871) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U832_XOR2_U1 ( .A0_t (U832_Y), .A0_f (new_AGEMA_signal_5869), .A1_t (new_AGEMA_signal_5870), .A1_f (new_AGEMA_signal_5871), .B0_t (StateOut[174]), .B0_f (new_AGEMA_signal_2490), .B1_t (new_AGEMA_signal_2491), .B1_f (new_AGEMA_signal_2492), .Z0_t (StateOut[166]), .Z0_f (new_AGEMA_signal_2493), .Z1_t (new_AGEMA_signal_2494), .Z1_f (new_AGEMA_signal_2495) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U833_XOR1_U1 ( .A0_t (StateOut[182]), .A0_f (new_AGEMA_signal_3126), .A1_t (new_AGEMA_signal_3127), .A1_f (new_AGEMA_signal_3128), .B0_t (StateFromChi[174]), .B0_f (new_AGEMA_signal_5076), .B1_t (new_AGEMA_signal_5077), .B1_f (new_AGEMA_signal_5078), .Z0_t (U833_X), .Z0_f (new_AGEMA_signal_5250), .Z1_t (new_AGEMA_signal_5251), .Z1_f (new_AGEMA_signal_5252) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U833_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U833_X), .B0_f (new_AGEMA_signal_5250), .B1_t (new_AGEMA_signal_5251), .B1_f (new_AGEMA_signal_5252), .Z0_t (U833_Y), .Z0_f (new_AGEMA_signal_5872), .Z1_t (new_AGEMA_signal_5873), .Z1_f (new_AGEMA_signal_5874) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U833_XOR2_U1 ( .A0_t (U833_Y), .A0_f (new_AGEMA_signal_5872), .A1_t (new_AGEMA_signal_5873), .A1_f (new_AGEMA_signal_5874), .B0_t (StateOut[182]), .B0_f (new_AGEMA_signal_3126), .B1_t (new_AGEMA_signal_3127), .B1_f (new_AGEMA_signal_3128), .Z0_t (StateOut[174]), .Z0_f (new_AGEMA_signal_2490), .Z1_t (new_AGEMA_signal_2491), .Z1_f (new_AGEMA_signal_2492) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U834_XOR1_U1 ( .A0_t (StateOut[45]), .A0_f (new_AGEMA_signal_3132), .A1_t (new_AGEMA_signal_3133), .A1_f (new_AGEMA_signal_3134), .B0_t (StateFromChi[37]), .B0_f (new_AGEMA_signal_5034), .B1_t (new_AGEMA_signal_5035), .B1_f (new_AGEMA_signal_5036), .Z0_t (U834_X), .Z0_f (new_AGEMA_signal_5253), .Z1_t (new_AGEMA_signal_5254), .Z1_f (new_AGEMA_signal_5255) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U834_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U834_X), .B0_f (new_AGEMA_signal_5253), .B1_t (new_AGEMA_signal_5254), .B1_f (new_AGEMA_signal_5255), .Z0_t (U834_Y), .Z0_f (new_AGEMA_signal_5875), .Z1_t (new_AGEMA_signal_5876), .Z1_f (new_AGEMA_signal_5877) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U834_XOR2_U1 ( .A0_t (U834_Y), .A0_f (new_AGEMA_signal_5875), .A1_t (new_AGEMA_signal_5876), .A1_f (new_AGEMA_signal_5877), .B0_t (StateOut[45]), .B0_f (new_AGEMA_signal_3132), .B1_t (new_AGEMA_signal_3133), .B1_f (new_AGEMA_signal_3134), .Z0_t (StateOut[37]), .Z0_f (new_AGEMA_signal_2643), .Z1_t (new_AGEMA_signal_2644), .Z1_f (new_AGEMA_signal_2645) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U835_XOR1_U1 ( .A0_t (StateOut[61]), .A0_f (new_AGEMA_signal_2511), .A1_t (new_AGEMA_signal_2512), .A1_f (new_AGEMA_signal_2513), .B0_t (StateFromChi[53]), .B0_f (new_AGEMA_signal_4992), .B1_t (new_AGEMA_signal_4993), .B1_f (new_AGEMA_signal_4994), .Z0_t (U835_X), .Z0_f (new_AGEMA_signal_5256), .Z1_t (new_AGEMA_signal_5257), .Z1_f (new_AGEMA_signal_5258) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U835_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U835_X), .B0_f (new_AGEMA_signal_5256), .B1_t (new_AGEMA_signal_5257), .B1_f (new_AGEMA_signal_5258), .Z0_t (U835_Y), .Z0_f (new_AGEMA_signal_5878), .Z1_t (new_AGEMA_signal_5879), .Z1_f (new_AGEMA_signal_5880) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U835_XOR2_U1 ( .A0_t (U835_Y), .A0_f (new_AGEMA_signal_5878), .A1_t (new_AGEMA_signal_5879), .A1_f (new_AGEMA_signal_5880), .B0_t (StateOut[61]), .B0_f (new_AGEMA_signal_2511), .B1_t (new_AGEMA_signal_2512), .B1_f (new_AGEMA_signal_2513), .Z0_t (StateOut[53]), .Z0_f (new_AGEMA_signal_2508), .Z1_t (new_AGEMA_signal_2509), .Z1_f (new_AGEMA_signal_2510) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U836_XOR1_U1 ( .A0_t (StateOut[69]), .A0_f (new_AGEMA_signal_2520), .A1_t (new_AGEMA_signal_2521), .A1_f (new_AGEMA_signal_2522), .B0_t (StateFromChi[61]), .B0_f (new_AGEMA_signal_5007), .B1_t (new_AGEMA_signal_5008), .B1_f (new_AGEMA_signal_5009), .Z0_t (U836_X), .Z0_f (new_AGEMA_signal_5259), .Z1_t (new_AGEMA_signal_5260), .Z1_f (new_AGEMA_signal_5261) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U836_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U836_X), .B0_f (new_AGEMA_signal_5259), .B1_t (new_AGEMA_signal_5260), .B1_f (new_AGEMA_signal_5261), .Z0_t (U836_Y), .Z0_f (new_AGEMA_signal_5881), .Z1_t (new_AGEMA_signal_5882), .Z1_f (new_AGEMA_signal_5883) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U836_XOR2_U1 ( .A0_t (U836_Y), .A0_f (new_AGEMA_signal_5881), .A1_t (new_AGEMA_signal_5882), .A1_f (new_AGEMA_signal_5883), .B0_t (StateOut[69]), .B0_f (new_AGEMA_signal_2520), .B1_t (new_AGEMA_signal_2521), .B1_f (new_AGEMA_signal_2522), .Z0_t (StateOut[61]), .Z0_f (new_AGEMA_signal_2511), .Z1_t (new_AGEMA_signal_2512), .Z1_f (new_AGEMA_signal_2513) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U837_XOR1_U1 ( .A0_t (StateOut[77]), .A0_f (new_AGEMA_signal_2517), .A1_t (new_AGEMA_signal_2518), .A1_f (new_AGEMA_signal_2519), .B0_t (StateFromChi[69]), .B0_f (new_AGEMA_signal_5022), .B1_t (new_AGEMA_signal_5023), .B1_f (new_AGEMA_signal_5024), .Z0_t (U837_X), .Z0_f (new_AGEMA_signal_5262), .Z1_t (new_AGEMA_signal_5263), .Z1_f (new_AGEMA_signal_5264) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U837_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U837_X), .B0_f (new_AGEMA_signal_5262), .B1_t (new_AGEMA_signal_5263), .B1_f (new_AGEMA_signal_5264), .Z0_t (U837_Y), .Z0_f (new_AGEMA_signal_5884), .Z1_t (new_AGEMA_signal_5885), .Z1_f (new_AGEMA_signal_5886) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U837_XOR2_U1 ( .A0_t (U837_Y), .A0_f (new_AGEMA_signal_5884), .A1_t (new_AGEMA_signal_5885), .A1_f (new_AGEMA_signal_5886), .B0_t (StateOut[77]), .B0_f (new_AGEMA_signal_2517), .B1_t (new_AGEMA_signal_2518), .B1_f (new_AGEMA_signal_2519), .Z0_t (StateOut[69]), .Z0_f (new_AGEMA_signal_2520), .Z1_t (new_AGEMA_signal_2521), .Z1_f (new_AGEMA_signal_2522) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U838_XOR1_U1 ( .A0_t (StateOut[125]), .A0_f (new_AGEMA_signal_3144), .A1_t (new_AGEMA_signal_3145), .A1_f (new_AGEMA_signal_3146), .B0_t (StateFromChi[117]), .B0_f (new_AGEMA_signal_5040), .B1_t (new_AGEMA_signal_5041), .B1_f (new_AGEMA_signal_5042), .Z0_t (U838_X), .Z0_f (new_AGEMA_signal_5265), .Z1_t (new_AGEMA_signal_5266), .Z1_f (new_AGEMA_signal_5267) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U838_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U838_X), .B0_f (new_AGEMA_signal_5265), .B1_t (new_AGEMA_signal_5266), .B1_f (new_AGEMA_signal_5267), .Z0_t (U838_Y), .Z0_f (new_AGEMA_signal_5887), .Z1_t (new_AGEMA_signal_5888), .Z1_f (new_AGEMA_signal_5889) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U838_XOR2_U1 ( .A0_t (U838_Y), .A0_f (new_AGEMA_signal_5887), .A1_t (new_AGEMA_signal_5888), .A1_f (new_AGEMA_signal_5889), .B0_t (StateOut[125]), .B0_f (new_AGEMA_signal_3144), .B1_t (new_AGEMA_signal_3145), .B1_f (new_AGEMA_signal_3146), .Z0_t (StateOut[117]), .Z0_f (new_AGEMA_signal_2733), .Z1_t (new_AGEMA_signal_2734), .Z1_f (new_AGEMA_signal_2735) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U839_XOR1_U1 ( .A0_t (StateOut[149]), .A0_f (new_AGEMA_signal_2556), .A1_t (new_AGEMA_signal_2557), .A1_f (new_AGEMA_signal_2558), .B0_t (StateFromChi[141]), .B0_f (new_AGEMA_signal_5013), .B1_t (new_AGEMA_signal_5014), .B1_f (new_AGEMA_signal_5015), .Z0_t (U839_X), .Z0_f (new_AGEMA_signal_5268), .Z1_t (new_AGEMA_signal_5269), .Z1_f (new_AGEMA_signal_5270) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U839_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U839_X), .B0_f (new_AGEMA_signal_5268), .B1_t (new_AGEMA_signal_5269), .B1_f (new_AGEMA_signal_5270), .Z0_t (U839_Y), .Z0_f (new_AGEMA_signal_5890), .Z1_t (new_AGEMA_signal_5891), .Z1_f (new_AGEMA_signal_5892) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U839_XOR2_U1 ( .A0_t (U839_Y), .A0_f (new_AGEMA_signal_5890), .A1_t (new_AGEMA_signal_5891), .A1_f (new_AGEMA_signal_5892), .B0_t (StateOut[149]), .B0_f (new_AGEMA_signal_2556), .B1_t (new_AGEMA_signal_2557), .B1_f (new_AGEMA_signal_2558), .Z0_t (StateOut[141]), .Z0_f (new_AGEMA_signal_2547), .Z1_t (new_AGEMA_signal_2548), .Z1_f (new_AGEMA_signal_2549) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U841_XOR1_U1 ( .A0_t (StateOut[157]), .A0_f (new_AGEMA_signal_2553), .A1_t (new_AGEMA_signal_2554), .A1_f (new_AGEMA_signal_2555), .B0_t (StateFromChi[149]), .B0_f (new_AGEMA_signal_5028), .B1_t (new_AGEMA_signal_5029), .B1_f (new_AGEMA_signal_5030), .Z0_t (U841_X), .Z0_f (new_AGEMA_signal_5271), .Z1_t (new_AGEMA_signal_5272), .Z1_f (new_AGEMA_signal_5273) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U841_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U841_X), .B0_f (new_AGEMA_signal_5271), .B1_t (new_AGEMA_signal_5272), .B1_f (new_AGEMA_signal_5273), .Z0_t (U841_Y), .Z0_f (new_AGEMA_signal_5893), .Z1_t (new_AGEMA_signal_5894), .Z1_f (new_AGEMA_signal_5895) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U841_XOR2_U1 ( .A0_t (U841_Y), .A0_f (new_AGEMA_signal_5893), .A1_t (new_AGEMA_signal_5894), .A1_f (new_AGEMA_signal_5895), .B0_t (StateOut[157]), .B0_f (new_AGEMA_signal_2553), .B1_t (new_AGEMA_signal_2554), .B1_f (new_AGEMA_signal_2555), .Z0_t (StateOut[149]), .Z0_f (new_AGEMA_signal_2556), .Z1_t (new_AGEMA_signal_2557), .Z1_f (new_AGEMA_signal_2558) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U842_XOR1_U1 ( .A0_t (StateOut[173]), .A0_f (new_AGEMA_signal_2670), .A1_t (new_AGEMA_signal_2671), .A1_f (new_AGEMA_signal_2672), .B0_t (StateFromChi[165]), .B0_f (new_AGEMA_signal_4986), .B1_t (new_AGEMA_signal_4987), .B1_f (new_AGEMA_signal_4988), .Z0_t (U842_X), .Z0_f (new_AGEMA_signal_5274), .Z1_t (new_AGEMA_signal_5275), .Z1_f (new_AGEMA_signal_5276) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U842_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U842_X), .B0_f (new_AGEMA_signal_5274), .B1_t (new_AGEMA_signal_5275), .B1_f (new_AGEMA_signal_5276), .Z0_t (U842_Y), .Z0_f (new_AGEMA_signal_5896), .Z1_t (new_AGEMA_signal_5897), .Z1_f (new_AGEMA_signal_5898) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U842_XOR2_U1 ( .A0_t (U842_Y), .A0_f (new_AGEMA_signal_5896), .A1_t (new_AGEMA_signal_5897), .A1_f (new_AGEMA_signal_5898), .B0_t (StateOut[173]), .B0_f (new_AGEMA_signal_2670), .B1_t (new_AGEMA_signal_2671), .B1_f (new_AGEMA_signal_2672), .Z0_t (StateOut[165]), .Z0_f (new_AGEMA_signal_2673), .Z1_t (new_AGEMA_signal_2674), .Z1_f (new_AGEMA_signal_2675) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U843_XOR1_U1 ( .A0_t (StateOut[181]), .A0_f (new_AGEMA_signal_3186), .A1_t (new_AGEMA_signal_3187), .A1_f (new_AGEMA_signal_3188), .B0_t (StateFromChi[173]), .B0_f (new_AGEMA_signal_5001), .B1_t (new_AGEMA_signal_5002), .B1_f (new_AGEMA_signal_5003), .Z0_t (U843_X), .Z0_f (new_AGEMA_signal_5277), .Z1_t (new_AGEMA_signal_5278), .Z1_f (new_AGEMA_signal_5279) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U843_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U843_X), .B0_f (new_AGEMA_signal_5277), .B1_t (new_AGEMA_signal_5278), .B1_f (new_AGEMA_signal_5279), .Z0_t (U843_Y), .Z0_f (new_AGEMA_signal_5899), .Z1_t (new_AGEMA_signal_5900), .Z1_f (new_AGEMA_signal_5901) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U843_XOR2_U1 ( .A0_t (U843_Y), .A0_f (new_AGEMA_signal_5899), .A1_t (new_AGEMA_signal_5900), .A1_f (new_AGEMA_signal_5901), .B0_t (StateOut[181]), .B0_f (new_AGEMA_signal_3186), .B1_t (new_AGEMA_signal_3187), .B1_f (new_AGEMA_signal_3188), .Z0_t (StateOut[173]), .Z0_f (new_AGEMA_signal_2670), .Z1_t (new_AGEMA_signal_2671), .Z1_f (new_AGEMA_signal_2672) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U844_XOR1_U1 ( .A0_t (StateOut[36]), .A0_f (new_AGEMA_signal_2571), .A1_t (new_AGEMA_signal_2572), .A1_f (new_AGEMA_signal_2573), .B0_t (StateFromChi[28]), .B0_f (new_AGEMA_signal_4944), .B1_t (new_AGEMA_signal_4945), .B1_f (new_AGEMA_signal_4946), .Z0_t (U844_X), .Z0_f (new_AGEMA_signal_5280), .Z1_t (new_AGEMA_signal_5281), .Z1_f (new_AGEMA_signal_5282) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U844_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U844_X), .B0_f (new_AGEMA_signal_5280), .B1_t (new_AGEMA_signal_5281), .B1_f (new_AGEMA_signal_5282), .Z0_t (U844_Y), .Z0_f (new_AGEMA_signal_5902), .Z1_t (new_AGEMA_signal_5903), .Z1_f (new_AGEMA_signal_5904) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U844_XOR2_U1 ( .A0_t (U844_Y), .A0_f (new_AGEMA_signal_5902), .A1_t (new_AGEMA_signal_5903), .A1_f (new_AGEMA_signal_5904), .B0_t (StateOut[36]), .B0_f (new_AGEMA_signal_2571), .B1_t (new_AGEMA_signal_2572), .B1_f (new_AGEMA_signal_2573), .Z0_t (StateOut[28]), .Z0_f (new_AGEMA_signal_2574), .Z1_t (new_AGEMA_signal_2575), .Z1_f (new_AGEMA_signal_2576) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U845_XOR1_U1 ( .A0_t (StateOut[44]), .A0_f (new_AGEMA_signal_2601), .A1_t (new_AGEMA_signal_2602), .A1_f (new_AGEMA_signal_2603), .B0_t (StateFromChi[36]), .B0_f (new_AGEMA_signal_4959), .B1_t (new_AGEMA_signal_4960), .B1_f (new_AGEMA_signal_4961), .Z0_t (U845_X), .Z0_f (new_AGEMA_signal_5283), .Z1_t (new_AGEMA_signal_5284), .Z1_f (new_AGEMA_signal_5285) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U845_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U845_X), .B0_f (new_AGEMA_signal_5283), .B1_t (new_AGEMA_signal_5284), .B1_f (new_AGEMA_signal_5285), .Z0_t (U845_Y), .Z0_f (new_AGEMA_signal_5905), .Z1_t (new_AGEMA_signal_5906), .Z1_f (new_AGEMA_signal_5907) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U845_XOR2_U1 ( .A0_t (U845_Y), .A0_f (new_AGEMA_signal_5905), .A1_t (new_AGEMA_signal_5906), .A1_f (new_AGEMA_signal_5907), .B0_t (StateOut[44]), .B0_f (new_AGEMA_signal_2601), .B1_t (new_AGEMA_signal_2602), .B1_f (new_AGEMA_signal_2603), .Z0_t (StateOut[36]), .Z0_f (new_AGEMA_signal_2571), .Z1_t (new_AGEMA_signal_2572), .Z1_f (new_AGEMA_signal_2573) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U846_XOR1_U1 ( .A0_t (StateOut[60]), .A0_f (new_AGEMA_signal_3162), .A1_t (new_AGEMA_signal_3163), .A1_f (new_AGEMA_signal_3164), .B0_t (StateFromChi[52]), .B0_f (new_AGEMA_signal_4917), .B1_t (new_AGEMA_signal_4918), .B1_f (new_AGEMA_signal_4919), .Z0_t (U846_X), .Z0_f (new_AGEMA_signal_5286), .Z1_t (new_AGEMA_signal_5287), .Z1_f (new_AGEMA_signal_5288) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U846_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U846_X), .B0_f (new_AGEMA_signal_5286), .B1_t (new_AGEMA_signal_5287), .B1_f (new_AGEMA_signal_5288), .Z0_t (U846_Y), .Z0_f (new_AGEMA_signal_5908), .Z1_t (new_AGEMA_signal_5909), .Z1_f (new_AGEMA_signal_5910) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U846_XOR2_U1 ( .A0_t (U846_Y), .A0_f (new_AGEMA_signal_5908), .A1_t (new_AGEMA_signal_5909), .A1_f (new_AGEMA_signal_5910), .B0_t (StateOut[60]), .B0_f (new_AGEMA_signal_3162), .B1_t (new_AGEMA_signal_3163), .B1_f (new_AGEMA_signal_3164), .Z0_t (StateOut[52]), .Z0_f (new_AGEMA_signal_2598), .Z1_t (new_AGEMA_signal_2599), .Z1_f (new_AGEMA_signal_2600) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U847_XOR1_U1 ( .A0_t (StateOut[68]), .A0_f (new_AGEMA_signal_2607), .A1_t (new_AGEMA_signal_2608), .A1_f (new_AGEMA_signal_2609), .B0_t (StateFromChi[60]), .B0_f (new_AGEMA_signal_4932), .B1_t (new_AGEMA_signal_4933), .B1_f (new_AGEMA_signal_4934), .Z0_t (U847_X), .Z0_f (new_AGEMA_signal_5289), .Z1_t (new_AGEMA_signal_5290), .Z1_f (new_AGEMA_signal_5291) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U847_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U847_X), .B0_f (new_AGEMA_signal_5289), .B1_t (new_AGEMA_signal_5290), .B1_f (new_AGEMA_signal_5291), .Z0_t (U847_Y), .Z0_f (new_AGEMA_signal_5911), .Z1_t (new_AGEMA_signal_5912), .Z1_f (new_AGEMA_signal_5913) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U847_XOR2_U1 ( .A0_t (U847_Y), .A0_f (new_AGEMA_signal_5911), .A1_t (new_AGEMA_signal_5912), .A1_f (new_AGEMA_signal_5913), .B0_t (StateOut[68]), .B0_f (new_AGEMA_signal_2607), .B1_t (new_AGEMA_signal_2608), .B1_f (new_AGEMA_signal_2609), .Z0_t (StateOut[60]), .Z0_f (new_AGEMA_signal_3162), .Z1_t (new_AGEMA_signal_3163), .Z1_f (new_AGEMA_signal_3164) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U848_XOR1_U1 ( .A0_t (StateOut[92]), .A0_f (new_AGEMA_signal_2796), .A1_t (new_AGEMA_signal_2797), .A1_f (new_AGEMA_signal_2798), .B0_t (StateFromChi[84]), .B0_f (new_AGEMA_signal_4905), .B1_t (new_AGEMA_signal_4906), .B1_f (new_AGEMA_signal_4907), .Z0_t (U848_X), .Z0_f (new_AGEMA_signal_5292), .Z1_t (new_AGEMA_signal_5293), .Z1_f (new_AGEMA_signal_5294) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U848_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U848_X), .B0_f (new_AGEMA_signal_5292), .B1_t (new_AGEMA_signal_5293), .B1_f (new_AGEMA_signal_5294), .Z0_t (U848_Y), .Z0_f (new_AGEMA_signal_5914), .Z1_t (new_AGEMA_signal_5915), .Z1_f (new_AGEMA_signal_5916) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U848_XOR2_U1 ( .A0_t (U848_Y), .A0_f (new_AGEMA_signal_5914), .A1_t (new_AGEMA_signal_5915), .A1_f (new_AGEMA_signal_5916), .B0_t (StateOut[92]), .B0_f (new_AGEMA_signal_2796), .B1_t (new_AGEMA_signal_2797), .B1_f (new_AGEMA_signal_2798), .Z0_t (StateOut[84]), .Z0_f (new_AGEMA_signal_2799), .Z1_t (new_AGEMA_signal_2800), .Z1_f (new_AGEMA_signal_2801) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U849_XOR1_U1 ( .A0_t (StateOut[100]), .A0_f (new_AGEMA_signal_3228), .A1_t (new_AGEMA_signal_3229), .A1_f (new_AGEMA_signal_3230), .B0_t (StateFromChi[92]), .B0_f (new_AGEMA_signal_4920), .B1_t (new_AGEMA_signal_4921), .B1_f (new_AGEMA_signal_4922), .Z0_t (U849_X), .Z0_f (new_AGEMA_signal_5295), .Z1_t (new_AGEMA_signal_5296), .Z1_f (new_AGEMA_signal_5297) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U849_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U849_X), .B0_f (new_AGEMA_signal_5295), .B1_t (new_AGEMA_signal_5296), .B1_f (new_AGEMA_signal_5297), .Z0_t (U849_Y), .Z0_f (new_AGEMA_signal_5917), .Z1_t (new_AGEMA_signal_5918), .Z1_f (new_AGEMA_signal_5919) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U849_XOR2_U1 ( .A0_t (U849_Y), .A0_f (new_AGEMA_signal_5917), .A1_t (new_AGEMA_signal_5918), .A1_f (new_AGEMA_signal_5919), .B0_t (StateOut[100]), .B0_f (new_AGEMA_signal_3228), .B1_t (new_AGEMA_signal_3229), .B1_f (new_AGEMA_signal_3230), .Z0_t (StateOut[92]), .Z0_f (new_AGEMA_signal_2796), .Z1_t (new_AGEMA_signal_2797), .Z1_f (new_AGEMA_signal_2798) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U850_XOR1_U1 ( .A0_t (StateOut[124]), .A0_f (new_AGEMA_signal_3084), .A1_t (new_AGEMA_signal_3085), .A1_f (new_AGEMA_signal_3086), .B0_t (StateFromChi[116]), .B0_f (new_AGEMA_signal_4965), .B1_t (new_AGEMA_signal_4966), .B1_f (new_AGEMA_signal_4967), .Z0_t (U850_X), .Z0_f (new_AGEMA_signal_5298), .Z1_t (new_AGEMA_signal_5299), .Z1_f (new_AGEMA_signal_5300) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U850_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U850_X), .B0_f (new_AGEMA_signal_5298), .B1_t (new_AGEMA_signal_5299), .B1_f (new_AGEMA_signal_5300), .Z0_t (U850_Y), .Z0_f (new_AGEMA_signal_5920), .Z1_t (new_AGEMA_signal_5921), .Z1_f (new_AGEMA_signal_5922) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U850_XOR2_U1 ( .A0_t (U850_Y), .A0_f (new_AGEMA_signal_5920), .A1_t (new_AGEMA_signal_5921), .A1_f (new_AGEMA_signal_5922), .B0_t (StateOut[124]), .B0_f (new_AGEMA_signal_3084), .B1_t (new_AGEMA_signal_3085), .B1_f (new_AGEMA_signal_3086), .Z0_t (StateOut[116]), .Z0_f (new_AGEMA_signal_2808), .Z1_t (new_AGEMA_signal_2809), .Z1_f (new_AGEMA_signal_2810) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U851_XOR1_U1 ( .A0_t (StateOut[172]), .A0_f (new_AGEMA_signal_2706), .A1_t (new_AGEMA_signal_2707), .A1_f (new_AGEMA_signal_2708), .B0_t (StateFromChi[164]), .B0_f (new_AGEMA_signal_4911), .B1_t (new_AGEMA_signal_4912), .B1_f (new_AGEMA_signal_4913), .Z0_t (U851_X), .Z0_f (new_AGEMA_signal_5301), .Z1_t (new_AGEMA_signal_5302), .Z1_f (new_AGEMA_signal_5303) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U851_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U851_X), .B0_f (new_AGEMA_signal_5301), .B1_t (new_AGEMA_signal_5302), .B1_f (new_AGEMA_signal_5303), .Z0_t (U851_Y), .Z0_f (new_AGEMA_signal_5923), .Z1_t (new_AGEMA_signal_5924), .Z1_f (new_AGEMA_signal_5925) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U851_XOR2_U1 ( .A0_t (U851_Y), .A0_f (new_AGEMA_signal_5923), .A1_t (new_AGEMA_signal_5924), .A1_f (new_AGEMA_signal_5925), .B0_t (StateOut[172]), .B0_f (new_AGEMA_signal_2706), .B1_t (new_AGEMA_signal_2707), .B1_f (new_AGEMA_signal_2708), .Z0_t (StateOut[164]), .Z0_f (new_AGEMA_signal_2709), .Z1_t (new_AGEMA_signal_2710), .Z1_f (new_AGEMA_signal_2711) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U852_XOR1_U1 ( .A0_t (StateOut[180]), .A0_f (new_AGEMA_signal_3198), .A1_t (new_AGEMA_signal_3199), .A1_f (new_AGEMA_signal_3200), .B0_t (StateFromChi[172]), .B0_f (new_AGEMA_signal_4926), .B1_t (new_AGEMA_signal_4927), .B1_f (new_AGEMA_signal_4928), .Z0_t (U852_X), .Z0_f (new_AGEMA_signal_5304), .Z1_t (new_AGEMA_signal_5305), .Z1_f (new_AGEMA_signal_5306) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U852_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U852_X), .B0_f (new_AGEMA_signal_5304), .B1_t (new_AGEMA_signal_5305), .B1_f (new_AGEMA_signal_5306), .Z0_t (U852_Y), .Z0_f (new_AGEMA_signal_5926), .Z1_t (new_AGEMA_signal_5927), .Z1_f (new_AGEMA_signal_5928) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U852_XOR2_U1 ( .A0_t (U852_Y), .A0_f (new_AGEMA_signal_5926), .A1_t (new_AGEMA_signal_5927), .A1_f (new_AGEMA_signal_5928), .B0_t (StateOut[180]), .B0_f (new_AGEMA_signal_3198), .B1_t (new_AGEMA_signal_3199), .B1_f (new_AGEMA_signal_3200), .Z0_t (StateOut[172]), .Z0_f (new_AGEMA_signal_2706), .Z1_t (new_AGEMA_signal_2707), .Z1_f (new_AGEMA_signal_2708) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U853_XOR1_U1 ( .A0_t (StateOut[35]), .A0_f (new_AGEMA_signal_2193), .A1_t (new_AGEMA_signal_2194), .A1_f (new_AGEMA_signal_2195), .B0_t (StateFromChi[27]), .B0_f (new_AGEMA_signal_4869), .B1_t (new_AGEMA_signal_4870), .B1_f (new_AGEMA_signal_4871), .Z0_t (U853_X), .Z0_f (new_AGEMA_signal_5307), .Z1_t (new_AGEMA_signal_5308), .Z1_f (new_AGEMA_signal_5309) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U853_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U853_X), .B0_f (new_AGEMA_signal_5307), .B1_t (new_AGEMA_signal_5308), .B1_f (new_AGEMA_signal_5309), .Z0_t (U853_Y), .Z0_f (new_AGEMA_signal_5929), .Z1_t (new_AGEMA_signal_5930), .Z1_f (new_AGEMA_signal_5931) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U853_XOR2_U1 ( .A0_t (U853_Y), .A0_f (new_AGEMA_signal_5929), .A1_t (new_AGEMA_signal_5930), .A1_f (new_AGEMA_signal_5931), .B0_t (StateOut[35]), .B0_f (new_AGEMA_signal_2193), .B1_t (new_AGEMA_signal_2194), .B1_f (new_AGEMA_signal_2195), .Z0_t (StateOut[27]), .Z0_f (new_AGEMA_signal_2196), .Z1_t (new_AGEMA_signal_2197), .Z1_f (new_AGEMA_signal_2198) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U854_XOR1_U1 ( .A0_t (StateOut[59]), .A0_f (new_AGEMA_signal_3168), .A1_t (new_AGEMA_signal_3169), .A1_f (new_AGEMA_signal_3170), .B0_t (StateFromChi[51]), .B0_f (new_AGEMA_signal_4842), .B1_t (new_AGEMA_signal_4843), .B1_f (new_AGEMA_signal_4844), .Z0_t (U854_X), .Z0_f (new_AGEMA_signal_5310), .Z1_t (new_AGEMA_signal_5311), .Z1_f (new_AGEMA_signal_5312) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U854_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U854_X), .B0_f (new_AGEMA_signal_5310), .B1_t (new_AGEMA_signal_5311), .B1_f (new_AGEMA_signal_5312), .Z0_t (U854_Y), .Z0_f (new_AGEMA_signal_5932), .Z1_t (new_AGEMA_signal_5933), .Z1_f (new_AGEMA_signal_5934) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U854_XOR2_U1 ( .A0_t (U854_Y), .A0_f (new_AGEMA_signal_5932), .A1_t (new_AGEMA_signal_5933), .A1_f (new_AGEMA_signal_5934), .B0_t (StateOut[59]), .B0_f (new_AGEMA_signal_3168), .B1_t (new_AGEMA_signal_3169), .B1_f (new_AGEMA_signal_3170), .Z0_t (StateOut[51]), .Z0_f (new_AGEMA_signal_2616), .Z1_t (new_AGEMA_signal_2617), .Z1_f (new_AGEMA_signal_2618) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U855_XOR1_U1 ( .A0_t (StateOut[91]), .A0_f (new_AGEMA_signal_2814), .A1_t (new_AGEMA_signal_2815), .A1_f (new_AGEMA_signal_2816), .B0_t (StateFromChi[83]), .B0_f (new_AGEMA_signal_4830), .B1_t (new_AGEMA_signal_4831), .B1_f (new_AGEMA_signal_4832), .Z0_t (U855_X), .Z0_f (new_AGEMA_signal_5313), .Z1_t (new_AGEMA_signal_5314), .Z1_f (new_AGEMA_signal_5315) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U855_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U855_X), .B0_f (new_AGEMA_signal_5313), .B1_t (new_AGEMA_signal_5314), .B1_f (new_AGEMA_signal_5315), .Z0_t (U855_Y), .Z0_f (new_AGEMA_signal_5935), .Z1_t (new_AGEMA_signal_5936), .Z1_f (new_AGEMA_signal_5937) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U855_XOR2_U1 ( .A0_t (U855_Y), .A0_f (new_AGEMA_signal_5935), .A1_t (new_AGEMA_signal_5936), .A1_f (new_AGEMA_signal_5937), .B0_t (StateOut[91]), .B0_f (new_AGEMA_signal_2814), .B1_t (new_AGEMA_signal_2815), .B1_f (new_AGEMA_signal_2816), .Z0_t (StateOut[83]), .Z0_f (new_AGEMA_signal_2817), .Z1_t (new_AGEMA_signal_2818), .Z1_f (new_AGEMA_signal_2819) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U856_XOR1_U1 ( .A0_t (StateOut[155]), .A0_f (new_AGEMA_signal_2589), .A1_t (new_AGEMA_signal_2590), .A1_f (new_AGEMA_signal_2591), .B0_t (StateFromChi[147]), .B0_f (new_AGEMA_signal_4878), .B1_t (new_AGEMA_signal_4879), .B1_f (new_AGEMA_signal_4880), .Z0_t (U856_X), .Z0_f (new_AGEMA_signal_5316), .Z1_t (new_AGEMA_signal_5317), .Z1_f (new_AGEMA_signal_5318) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U856_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U856_X), .B0_f (new_AGEMA_signal_5316), .B1_t (new_AGEMA_signal_5317), .B1_f (new_AGEMA_signal_5318), .Z0_t (U856_Y), .Z0_f (new_AGEMA_signal_5938), .Z1_t (new_AGEMA_signal_5939), .Z1_f (new_AGEMA_signal_5940) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U856_XOR2_U1 ( .A0_t (U856_Y), .A0_f (new_AGEMA_signal_5938), .A1_t (new_AGEMA_signal_5939), .A1_f (new_AGEMA_signal_5940), .B0_t (StateOut[155]), .B0_f (new_AGEMA_signal_2589), .B1_t (new_AGEMA_signal_2590), .B1_f (new_AGEMA_signal_2591), .Z0_t (StateOut[147]), .Z0_f (new_AGEMA_signal_2592), .Z1_t (new_AGEMA_signal_2593), .Z1_f (new_AGEMA_signal_2594) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U857_XOR1_U1 ( .A0_t (StateOut[171]), .A0_f (new_AGEMA_signal_2778), .A1_t (new_AGEMA_signal_2779), .A1_f (new_AGEMA_signal_2780), .B0_t (StateFromChi[163]), .B0_f (new_AGEMA_signal_4836), .B1_t (new_AGEMA_signal_4837), .B1_f (new_AGEMA_signal_4838), .Z0_t (U857_X), .Z0_f (new_AGEMA_signal_5319), .Z1_t (new_AGEMA_signal_5320), .Z1_f (new_AGEMA_signal_5321) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U857_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U857_X), .B0_f (new_AGEMA_signal_5319), .B1_t (new_AGEMA_signal_5320), .B1_f (new_AGEMA_signal_5321), .Z0_t (U857_Y), .Z0_f (new_AGEMA_signal_5941), .Z1_t (new_AGEMA_signal_5942), .Z1_f (new_AGEMA_signal_5943) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U857_XOR2_U1 ( .A0_t (U857_Y), .A0_f (new_AGEMA_signal_5941), .A1_t (new_AGEMA_signal_5942), .A1_f (new_AGEMA_signal_5943), .B0_t (StateOut[171]), .B0_f (new_AGEMA_signal_2778), .B1_t (new_AGEMA_signal_2779), .B1_f (new_AGEMA_signal_2780), .Z0_t (StateOut[163]), .Z0_f (new_AGEMA_signal_2781), .Z1_t (new_AGEMA_signal_2782), .Z1_f (new_AGEMA_signal_2783) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U858_XOR1_U1 ( .A0_t (StateOut[179]), .A0_f (new_AGEMA_signal_3222), .A1_t (new_AGEMA_signal_3223), .A1_f (new_AGEMA_signal_3224), .B0_t (StateFromChi[171]), .B0_f (new_AGEMA_signal_4851), .B1_t (new_AGEMA_signal_4852), .B1_f (new_AGEMA_signal_4853), .Z0_t (U858_X), .Z0_f (new_AGEMA_signal_5322), .Z1_t (new_AGEMA_signal_5323), .Z1_f (new_AGEMA_signal_5324) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U858_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U858_X), .B0_f (new_AGEMA_signal_5322), .B1_t (new_AGEMA_signal_5323), .B1_f (new_AGEMA_signal_5324), .Z0_t (U858_Y), .Z0_f (new_AGEMA_signal_5944), .Z1_t (new_AGEMA_signal_5945), .Z1_f (new_AGEMA_signal_5946) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U858_XOR2_U1 ( .A0_t (U858_Y), .A0_f (new_AGEMA_signal_5944), .A1_t (new_AGEMA_signal_5945), .A1_f (new_AGEMA_signal_5946), .B0_t (StateOut[179]), .B0_f (new_AGEMA_signal_3222), .B1_t (new_AGEMA_signal_3223), .B1_f (new_AGEMA_signal_3224), .Z0_t (StateOut[171]), .Z0_f (new_AGEMA_signal_2778), .Z1_t (new_AGEMA_signal_2779), .Z1_f (new_AGEMA_signal_2780) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U859_XOR1_U1 ( .A0_t (StateOut[187]), .A0_f (new_AGEMA_signal_2787), .A1_t (new_AGEMA_signal_2788), .A1_f (new_AGEMA_signal_2789), .B0_t (StateFromChi[179]), .B0_f (new_AGEMA_signal_4866), .B1_t (new_AGEMA_signal_4867), .B1_f (new_AGEMA_signal_4868), .Z0_t (U859_X), .Z0_f (new_AGEMA_signal_5325), .Z1_t (new_AGEMA_signal_5326), .Z1_f (new_AGEMA_signal_5327) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U859_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U859_X), .B0_f (new_AGEMA_signal_5325), .B1_t (new_AGEMA_signal_5326), .B1_f (new_AGEMA_signal_5327), .Z0_t (U859_Y), .Z0_f (new_AGEMA_signal_5947), .Z1_t (new_AGEMA_signal_5948), .Z1_f (new_AGEMA_signal_5949) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U859_XOR2_U1 ( .A0_t (U859_Y), .A0_f (new_AGEMA_signal_5947), .A1_t (new_AGEMA_signal_5948), .A1_f (new_AGEMA_signal_5949), .B0_t (StateOut[187]), .B0_f (new_AGEMA_signal_2787), .B1_t (new_AGEMA_signal_2788), .B1_f (new_AGEMA_signal_2789), .Z0_t (StateOut[179]), .Z0_f (new_AGEMA_signal_3222), .Z1_t (new_AGEMA_signal_3223), .Z1_f (new_AGEMA_signal_3224) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U860_XOR1_U1 ( .A0_t (StateOut[34]), .A0_f (new_AGEMA_signal_2535), .A1_t (new_AGEMA_signal_2536), .A1_f (new_AGEMA_signal_2537), .B0_t (StateFromChi[26]), .B0_f (new_AGEMA_signal_4794), .B1_t (new_AGEMA_signal_4795), .B1_f (new_AGEMA_signal_4796), .Z0_t (U860_X), .Z0_f (new_AGEMA_signal_5328), .Z1_t (new_AGEMA_signal_5329), .Z1_f (new_AGEMA_signal_5330) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U860_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U860_X), .B0_f (new_AGEMA_signal_5328), .B1_t (new_AGEMA_signal_5329), .B1_f (new_AGEMA_signal_5330), .Z0_t (U860_Y), .Z0_f (new_AGEMA_signal_5950), .Z1_t (new_AGEMA_signal_5951), .Z1_f (new_AGEMA_signal_5952) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U860_XOR2_U1 ( .A0_t (U860_Y), .A0_f (new_AGEMA_signal_5950), .A1_t (new_AGEMA_signal_5951), .A1_f (new_AGEMA_signal_5952), .B0_t (StateOut[34]), .B0_f (new_AGEMA_signal_2535), .B1_t (new_AGEMA_signal_2536), .B1_f (new_AGEMA_signal_2537), .Z0_t (StateOut[26]), .Z0_f (new_AGEMA_signal_3138), .Z1_t (new_AGEMA_signal_3139), .Z1_f (new_AGEMA_signal_3140) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U861_XOR1_U1 ( .A0_t (StateOut[42]), .A0_f (new_AGEMA_signal_2655), .A1_t (new_AGEMA_signal_2656), .A1_f (new_AGEMA_signal_2657), .B0_t (StateFromChi[34]), .B0_f (new_AGEMA_signal_4809), .B1_t (new_AGEMA_signal_4810), .B1_f (new_AGEMA_signal_4811), .Z0_t (U861_X), .Z0_f (new_AGEMA_signal_5331), .Z1_t (new_AGEMA_signal_5332), .Z1_f (new_AGEMA_signal_5333) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U861_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U861_X), .B0_f (new_AGEMA_signal_5331), .B1_t (new_AGEMA_signal_5332), .B1_f (new_AGEMA_signal_5333), .Z0_t (U861_Y), .Z0_f (new_AGEMA_signal_5953), .Z1_t (new_AGEMA_signal_5954), .Z1_f (new_AGEMA_signal_5955) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U861_XOR2_U1 ( .A0_t (U861_Y), .A0_f (new_AGEMA_signal_5953), .A1_t (new_AGEMA_signal_5954), .A1_f (new_AGEMA_signal_5955), .B0_t (StateOut[42]), .B0_f (new_AGEMA_signal_2655), .B1_t (new_AGEMA_signal_2656), .B1_f (new_AGEMA_signal_2657), .Z0_t (StateOut[34]), .Z0_f (new_AGEMA_signal_2535), .Z1_t (new_AGEMA_signal_2536), .Z1_f (new_AGEMA_signal_2537) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U862_XOR1_U1 ( .A0_t (StateOut[58]), .A0_f (new_AGEMA_signal_2664), .A1_t (new_AGEMA_signal_2665), .A1_f (new_AGEMA_signal_2666), .B0_t (StateFromChi[50]), .B0_f (new_AGEMA_signal_4767), .B1_t (new_AGEMA_signal_4768), .B1_f (new_AGEMA_signal_4769), .Z0_t (U862_X), .Z0_f (new_AGEMA_signal_5334), .Z1_t (new_AGEMA_signal_5335), .Z1_f (new_AGEMA_signal_5336) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U862_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U862_X), .B0_f (new_AGEMA_signal_5334), .B1_t (new_AGEMA_signal_5335), .B1_f (new_AGEMA_signal_5336), .Z0_t (U862_Y), .Z0_f (new_AGEMA_signal_5956), .Z1_t (new_AGEMA_signal_5957), .Z1_f (new_AGEMA_signal_5958) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U862_XOR2_U1 ( .A0_t (U862_Y), .A0_f (new_AGEMA_signal_5956), .A1_t (new_AGEMA_signal_5957), .A1_f (new_AGEMA_signal_5958), .B0_t (StateOut[58]), .B0_f (new_AGEMA_signal_2664), .B1_t (new_AGEMA_signal_2665), .B1_f (new_AGEMA_signal_2666), .Z0_t (StateOut[50]), .Z0_f (new_AGEMA_signal_2652), .Z1_t (new_AGEMA_signal_2653), .Z1_f (new_AGEMA_signal_2654) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U863_XOR1_U1 ( .A0_t (StateOut[66]), .A0_f (new_AGEMA_signal_3180), .A1_t (new_AGEMA_signal_3181), .A1_f (new_AGEMA_signal_3182), .B0_t (StateFromChi[58]), .B0_f (new_AGEMA_signal_4782), .B1_t (new_AGEMA_signal_4783), .B1_f (new_AGEMA_signal_4784), .Z0_t (U863_X), .Z0_f (new_AGEMA_signal_5337), .Z1_t (new_AGEMA_signal_5338), .Z1_f (new_AGEMA_signal_5339) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U863_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U863_X), .B0_f (new_AGEMA_signal_5337), .B1_t (new_AGEMA_signal_5338), .B1_f (new_AGEMA_signal_5339), .Z0_t (U863_Y), .Z0_f (new_AGEMA_signal_5959), .Z1_t (new_AGEMA_signal_5960), .Z1_f (new_AGEMA_signal_5961) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U863_XOR2_U1 ( .A0_t (U863_Y), .A0_f (new_AGEMA_signal_5959), .A1_t (new_AGEMA_signal_5960), .A1_f (new_AGEMA_signal_5961), .B0_t (StateOut[66]), .B0_f (new_AGEMA_signal_3180), .B1_t (new_AGEMA_signal_3181), .B1_f (new_AGEMA_signal_3182), .Z0_t (StateOut[58]), .Z0_f (new_AGEMA_signal_2664), .Z1_t (new_AGEMA_signal_2665), .Z1_f (new_AGEMA_signal_2666) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U864_XOR1_U1 ( .A0_t (StateOut[90]), .A0_f (new_AGEMA_signal_2220), .A1_t (new_AGEMA_signal_2221), .A1_f (new_AGEMA_signal_2222), .B0_t (StateFromChi[82]), .B0_f (new_AGEMA_signal_4755), .B1_t (new_AGEMA_signal_4756), .B1_f (new_AGEMA_signal_4757), .Z0_t (U864_X), .Z0_f (new_AGEMA_signal_5340), .Z1_t (new_AGEMA_signal_5341), .Z1_f (new_AGEMA_signal_5342) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U864_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U864_X), .B0_f (new_AGEMA_signal_5340), .B1_t (new_AGEMA_signal_5341), .B1_f (new_AGEMA_signal_5342), .Z0_t (U864_Y), .Z0_f (new_AGEMA_signal_5962), .Z1_t (new_AGEMA_signal_5963), .Z1_f (new_AGEMA_signal_5964) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U864_XOR2_U1 ( .A0_t (U864_Y), .A0_f (new_AGEMA_signal_5962), .A1_t (new_AGEMA_signal_5963), .A1_f (new_AGEMA_signal_5964), .B0_t (StateOut[90]), .B0_f (new_AGEMA_signal_2220), .B1_t (new_AGEMA_signal_2221), .B1_f (new_AGEMA_signal_2222), .Z0_t (StateOut[82]), .Z0_f (new_AGEMA_signal_3036), .Z1_t (new_AGEMA_signal_3037), .Z1_f (new_AGEMA_signal_3038) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U865_XOR1_U1 ( .A0_t (StateOut[162]), .A0_f (new_AGEMA_signal_2835), .A1_t (new_AGEMA_signal_2836), .A1_f (new_AGEMA_signal_2837), .B0_t (StateFromChi[154]), .B0_f (new_AGEMA_signal_4818), .B1_t (new_AGEMA_signal_4819), .B1_f (new_AGEMA_signal_4820), .Z0_t (U865_X), .Z0_f (new_AGEMA_signal_5343), .Z1_t (new_AGEMA_signal_5344), .Z1_f (new_AGEMA_signal_5345) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U865_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U865_X), .B0_f (new_AGEMA_signal_5343), .B1_t (new_AGEMA_signal_5344), .B1_f (new_AGEMA_signal_5345), .Z0_t (U865_Y), .Z0_f (new_AGEMA_signal_5965), .Z1_t (new_AGEMA_signal_5966), .Z1_f (new_AGEMA_signal_5967) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U865_XOR2_U1 ( .A0_t (U865_Y), .A0_f (new_AGEMA_signal_5965), .A1_t (new_AGEMA_signal_5966), .A1_f (new_AGEMA_signal_5967), .B0_t (StateOut[162]), .B0_f (new_AGEMA_signal_2835), .B1_t (new_AGEMA_signal_2836), .B1_f (new_AGEMA_signal_2837), .Z0_t (StateOut[154]), .Z0_f (new_AGEMA_signal_2754), .Z1_t (new_AGEMA_signal_2755), .Z1_f (new_AGEMA_signal_2756) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U866_XOR1_U1 ( .A0_t (StateOut[33]), .A0_f (new_AGEMA_signal_2772), .A1_t (new_AGEMA_signal_2773), .A1_f (new_AGEMA_signal_2774), .B0_t (StateFromChi[25]), .B0_f (new_AGEMA_signal_4719), .B1_t (new_AGEMA_signal_4720), .B1_f (new_AGEMA_signal_4721), .Z0_t (U866_X), .Z0_f (new_AGEMA_signal_5346), .Z1_t (new_AGEMA_signal_5347), .Z1_f (new_AGEMA_signal_5348) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U866_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U866_X), .B0_f (new_AGEMA_signal_5346), .B1_t (new_AGEMA_signal_5347), .B1_f (new_AGEMA_signal_5348), .Z0_t (U866_Y), .Z0_f (new_AGEMA_signal_5968), .Z1_t (new_AGEMA_signal_5969), .Z1_f (new_AGEMA_signal_5970) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U866_XOR2_U1 ( .A0_t (U866_Y), .A0_f (new_AGEMA_signal_5968), .A1_t (new_AGEMA_signal_5969), .A1_f (new_AGEMA_signal_5970), .B0_t (StateOut[33]), .B0_f (new_AGEMA_signal_2772), .B1_t (new_AGEMA_signal_2773), .B1_f (new_AGEMA_signal_2774), .Z0_t (StateOut[25]), .Z0_f (new_AGEMA_signal_2769), .Z1_t (new_AGEMA_signal_2770), .Z1_f (new_AGEMA_signal_2771) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U867_XOR1_U1 ( .A0_t (StateOut[57]), .A0_f (new_AGEMA_signal_3102), .A1_t (new_AGEMA_signal_3103), .A1_f (new_AGEMA_signal_3104), .B0_t (StateFromChi[49]), .B0_f (new_AGEMA_signal_4692), .B1_t (new_AGEMA_signal_4693), .B1_f (new_AGEMA_signal_4694), .Z0_t (U867_X), .Z0_f (new_AGEMA_signal_5349), .Z1_t (new_AGEMA_signal_5350), .Z1_f (new_AGEMA_signal_5351) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U867_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U867_X), .B0_f (new_AGEMA_signal_5349), .B1_t (new_AGEMA_signal_5350), .B1_f (new_AGEMA_signal_5351), .Z0_t (U867_Y), .Z0_f (new_AGEMA_signal_5971), .Z1_t (new_AGEMA_signal_5972), .Z1_f (new_AGEMA_signal_5973) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U867_XOR2_U1 ( .A0_t (U867_Y), .A0_f (new_AGEMA_signal_5971), .A1_t (new_AGEMA_signal_5972), .A1_f (new_AGEMA_signal_5973), .B0_t (StateOut[57]), .B0_f (new_AGEMA_signal_3102), .B1_t (new_AGEMA_signal_3103), .B1_f (new_AGEMA_signal_3104), .Z0_t (StateOut[49]), .Z0_f (new_AGEMA_signal_2418), .Z1_t (new_AGEMA_signal_2419), .Z1_f (new_AGEMA_signal_2420) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U868_XOR1_U1 ( .A0_t (StateOut[89]), .A0_f (new_AGEMA_signal_2292), .A1_t (new_AGEMA_signal_2293), .A1_f (new_AGEMA_signal_2294), .B0_t (StateFromChi[81]), .B0_f (new_AGEMA_signal_4680), .B1_t (new_AGEMA_signal_4681), .B1_f (new_AGEMA_signal_4682), .Z0_t (U868_X), .Z0_f (new_AGEMA_signal_5352), .Z1_t (new_AGEMA_signal_5353), .Z1_f (new_AGEMA_signal_5354) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U868_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U868_X), .B0_f (new_AGEMA_signal_5352), .B1_t (new_AGEMA_signal_5353), .B1_f (new_AGEMA_signal_5354), .Z0_t (U868_Y), .Z0_f (new_AGEMA_signal_5974), .Z1_t (new_AGEMA_signal_5975), .Z1_f (new_AGEMA_signal_5976) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U868_XOR2_U1 ( .A0_t (U868_Y), .A0_f (new_AGEMA_signal_5974), .A1_t (new_AGEMA_signal_5975), .A1_f (new_AGEMA_signal_5976), .B0_t (StateOut[89]), .B0_f (new_AGEMA_signal_2292), .B1_t (new_AGEMA_signal_2293), .B1_f (new_AGEMA_signal_2294), .Z0_t (StateOut[81]), .Z0_f (new_AGEMA_signal_3060), .Z1_t (new_AGEMA_signal_3061), .Z1_f (new_AGEMA_signal_3062) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U869_XOR1_U1 ( .A0_t (StateOut[145]), .A0_f (new_AGEMA_signal_2286), .A1_t (new_AGEMA_signal_2287), .A1_f (new_AGEMA_signal_2288), .B0_t (StateFromChi[137]), .B0_f (new_AGEMA_signal_4713), .B1_t (new_AGEMA_signal_4714), .B1_f (new_AGEMA_signal_4715), .Z0_t (U869_X), .Z0_f (new_AGEMA_signal_5355), .Z1_t (new_AGEMA_signal_5356), .Z1_f (new_AGEMA_signal_5357) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U869_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U869_X), .B0_f (new_AGEMA_signal_5355), .B1_t (new_AGEMA_signal_5356), .B1_f (new_AGEMA_signal_5357), .Z0_t (U869_Y), .Z0_f (new_AGEMA_signal_5977), .Z1_t (new_AGEMA_signal_5978), .Z1_f (new_AGEMA_signal_5979) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U869_XOR2_U1 ( .A0_t (U869_Y), .A0_f (new_AGEMA_signal_5977), .A1_t (new_AGEMA_signal_5978), .A1_f (new_AGEMA_signal_5979), .B0_t (StateOut[145]), .B0_f (new_AGEMA_signal_2286), .B1_t (new_AGEMA_signal_2287), .B1_f (new_AGEMA_signal_2288), .Z0_t (StateOut[137]), .Z0_f (new_AGEMA_signal_2277), .Z1_t (new_AGEMA_signal_2278), .Z1_f (new_AGEMA_signal_2279) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U870_XOR1_U1 ( .A0_t (StateOut[177]), .A0_f (new_AGEMA_signal_3042), .A1_t (new_AGEMA_signal_3043), .A1_f (new_AGEMA_signal_3044), .B0_t (StateFromChi[169]), .B0_f (new_AGEMA_signal_4701), .B1_t (new_AGEMA_signal_4702), .B1_f (new_AGEMA_signal_4703), .Z0_t (U870_X), .Z0_f (new_AGEMA_signal_5358), .Z1_t (new_AGEMA_signal_5359), .Z1_f (new_AGEMA_signal_5360) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U870_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U870_X), .B0_f (new_AGEMA_signal_5358), .B1_t (new_AGEMA_signal_5359), .B1_f (new_AGEMA_signal_5360), .Z0_t (U870_Y), .Z0_f (new_AGEMA_signal_5980), .Z1_t (new_AGEMA_signal_5981), .Z1_f (new_AGEMA_signal_5982) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U870_XOR2_U1 ( .A0_t (U870_Y), .A0_f (new_AGEMA_signal_5980), .A1_t (new_AGEMA_signal_5981), .A1_f (new_AGEMA_signal_5982), .B0_t (StateOut[177]), .B0_f (new_AGEMA_signal_3042), .B1_t (new_AGEMA_signal_3043), .B1_f (new_AGEMA_signal_3044), .Z0_t (StateOut[169]), .Z0_f (new_AGEMA_signal_2238), .Z1_t (new_AGEMA_signal_2239), .Z1_f (new_AGEMA_signal_2240) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U871_XOR1_U1 ( .A0_t (StateOut[32]), .A0_f (new_AGEMA_signal_2211), .A1_t (new_AGEMA_signal_2212), .A1_f (new_AGEMA_signal_2213), .B0_t (StateFromChi[24]), .B0_f (new_AGEMA_signal_4644), .B1_t (new_AGEMA_signal_4645), .B1_f (new_AGEMA_signal_4646), .Z0_t (U871_X), .Z0_f (new_AGEMA_signal_5361), .Z1_t (new_AGEMA_signal_5362), .Z1_f (new_AGEMA_signal_5363) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U871_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U871_X), .B0_f (new_AGEMA_signal_5361), .B1_t (new_AGEMA_signal_5362), .B1_f (new_AGEMA_signal_5363), .Z0_t (U871_Y), .Z0_f (new_AGEMA_signal_5983), .Z1_t (new_AGEMA_signal_5984), .Z1_f (new_AGEMA_signal_5985) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U871_XOR2_U1 ( .A0_t (U871_Y), .A0_f (new_AGEMA_signal_5983), .A1_t (new_AGEMA_signal_5984), .A1_f (new_AGEMA_signal_5985), .B0_t (StateOut[32]), .B0_f (new_AGEMA_signal_2211), .B1_t (new_AGEMA_signal_2212), .B1_f (new_AGEMA_signal_2213), .Z0_t (StateOut[24]), .Z0_f (new_AGEMA_signal_2214), .Z1_t (new_AGEMA_signal_2215), .Z1_f (new_AGEMA_signal_2216) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U872_XOR1_U1 ( .A0_t (StateOut[120]), .A0_f (new_AGEMA_signal_2403), .A1_t (new_AGEMA_signal_2404), .A1_f (new_AGEMA_signal_2405), .B0_t (StateFromChi[112]), .B0_f (new_AGEMA_signal_4665), .B1_t (new_AGEMA_signal_4666), .B1_f (new_AGEMA_signal_4667), .Z0_t (U872_X), .Z0_f (new_AGEMA_signal_5364), .Z1_t (new_AGEMA_signal_5365), .Z1_f (new_AGEMA_signal_5366) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U872_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U872_X), .B0_f (new_AGEMA_signal_5364), .B1_t (new_AGEMA_signal_5365), .B1_f (new_AGEMA_signal_5366), .Z0_t (U872_Y), .Z0_f (new_AGEMA_signal_5986), .Z1_t (new_AGEMA_signal_5987), .Z1_f (new_AGEMA_signal_5988) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U872_XOR2_U1 ( .A0_t (U872_Y), .A0_f (new_AGEMA_signal_5986), .A1_t (new_AGEMA_signal_5987), .A1_f (new_AGEMA_signal_5988), .B0_t (StateOut[120]), .B0_f (new_AGEMA_signal_2403), .B1_t (new_AGEMA_signal_2404), .B1_f (new_AGEMA_signal_2405), .Z0_t (StateOut[112]), .Z0_f (new_AGEMA_signal_2394), .Z1_t (new_AGEMA_signal_2395), .Z1_f (new_AGEMA_signal_2396) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U873_XOR1_U1 ( .A0_t (StateOut[144]), .A0_f (new_AGEMA_signal_3096), .A1_t (new_AGEMA_signal_3097), .A1_f (new_AGEMA_signal_3098), .B0_t (StateFromChi[136]), .B0_f (new_AGEMA_signal_4638), .B1_t (new_AGEMA_signal_4639), .B1_f (new_AGEMA_signal_4640), .Z0_t (U873_X), .Z0_f (new_AGEMA_signal_5367), .Z1_t (new_AGEMA_signal_5368), .Z1_f (new_AGEMA_signal_5369) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U873_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U873_X), .B0_f (new_AGEMA_signal_5367), .B1_t (new_AGEMA_signal_5368), .B1_f (new_AGEMA_signal_5369), .Z0_t (U873_Y), .Z0_f (new_AGEMA_signal_5989), .Z1_t (new_AGEMA_signal_5990), .Z1_f (new_AGEMA_signal_5991) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U873_XOR2_U1 ( .A0_t (U873_Y), .A0_f (new_AGEMA_signal_5989), .A1_t (new_AGEMA_signal_5990), .A1_f (new_AGEMA_signal_5991), .B0_t (StateOut[144]), .B0_f (new_AGEMA_signal_3096), .B1_t (new_AGEMA_signal_3097), .B1_f (new_AGEMA_signal_3098), .Z0_t (StateOut[136]), .Z0_f (new_AGEMA_signal_2412), .Z1_t (new_AGEMA_signal_2413), .Z1_f (new_AGEMA_signal_2414) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U874_XOR1_U1 ( .A0_t (StateOut[152]), .A0_f (new_AGEMA_signal_2409), .A1_t (new_AGEMA_signal_2410), .A1_f (new_AGEMA_signal_2411), .B0_t (StateFromChi[144]), .B0_f (new_AGEMA_signal_4653), .B1_t (new_AGEMA_signal_4654), .B1_f (new_AGEMA_signal_4655), .Z0_t (U874_X), .Z0_f (new_AGEMA_signal_5370), .Z1_t (new_AGEMA_signal_5371), .Z1_f (new_AGEMA_signal_5372) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U874_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U874_X), .B0_f (new_AGEMA_signal_5370), .B1_t (new_AGEMA_signal_5371), .B1_f (new_AGEMA_signal_5372), .Z0_t (U874_Y), .Z0_f (new_AGEMA_signal_5992), .Z1_t (new_AGEMA_signal_5993), .Z1_f (new_AGEMA_signal_5994) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U874_XOR2_U1 ( .A0_t (U874_Y), .A0_f (new_AGEMA_signal_5992), .A1_t (new_AGEMA_signal_5993), .A1_f (new_AGEMA_signal_5994), .B0_t (StateOut[152]), .B0_f (new_AGEMA_signal_2409), .B1_t (new_AGEMA_signal_2410), .B1_f (new_AGEMA_signal_2411), .Z0_t (StateOut[144]), .Z0_f (new_AGEMA_signal_3096), .Z1_t (new_AGEMA_signal_3097), .Z1_f (new_AGEMA_signal_3098) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U875_XOR1_U1 ( .A0_t (StateOut[31]), .A0_f (new_AGEMA_signal_2358), .A1_t (new_AGEMA_signal_2359), .A1_f (new_AGEMA_signal_2360), .B0_t (StateFromChi[23]), .B0_f (new_AGEMA_signal_5154), .B1_t (new_AGEMA_signal_5155), .B1_f (new_AGEMA_signal_5156), .Z0_t (U875_X), .Z0_f (new_AGEMA_signal_5373), .Z1_t (new_AGEMA_signal_5374), .Z1_f (new_AGEMA_signal_5375) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U875_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U875_X), .B0_f (new_AGEMA_signal_5373), .B1_t (new_AGEMA_signal_5374), .B1_f (new_AGEMA_signal_5375), .Z0_t (U875_Y), .Z0_f (new_AGEMA_signal_5995), .Z1_t (new_AGEMA_signal_5996), .Z1_f (new_AGEMA_signal_5997) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U875_XOR2_U1 ( .A0_t (U875_Y), .A0_f (new_AGEMA_signal_5995), .A1_t (new_AGEMA_signal_5996), .A1_f (new_AGEMA_signal_5997), .B0_t (StateOut[31]), .B0_f (new_AGEMA_signal_2358), .B1_t (new_AGEMA_signal_2359), .B1_f (new_AGEMA_signal_2360), .Z0_t (StateOut[23]), .Z0_f (new_AGEMA_signal_2349), .Z1_t (new_AGEMA_signal_2350), .Z1_f (new_AGEMA_signal_2351) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U876_XOR1_U1 ( .A0_t (StateOut[39]), .A0_f (new_AGEMA_signal_2355), .A1_t (new_AGEMA_signal_2356), .A1_f (new_AGEMA_signal_2357), .B0_t (StateFromChi[31]), .B0_f (new_AGEMA_signal_5169), .B1_t (new_AGEMA_signal_5170), .B1_f (new_AGEMA_signal_5171), .Z0_t (U876_X), .Z0_f (new_AGEMA_signal_5376), .Z1_t (new_AGEMA_signal_5377), .Z1_f (new_AGEMA_signal_5378) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U876_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U876_X), .B0_f (new_AGEMA_signal_5376), .B1_t (new_AGEMA_signal_5377), .B1_f (new_AGEMA_signal_5378), .Z0_t (U876_Y), .Z0_f (new_AGEMA_signal_5998), .Z1_t (new_AGEMA_signal_5999), .Z1_f (new_AGEMA_signal_6000) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U876_XOR2_U1 ( .A0_t (U876_Y), .A0_f (new_AGEMA_signal_5998), .A1_t (new_AGEMA_signal_5999), .A1_f (new_AGEMA_signal_6000), .B0_t (StateOut[39]), .B0_f (new_AGEMA_signal_2355), .B1_t (new_AGEMA_signal_2356), .B1_f (new_AGEMA_signal_2357), .Z0_t (StateOut[31]), .Z0_f (new_AGEMA_signal_2358), .Z1_t (new_AGEMA_signal_2359), .Z1_f (new_AGEMA_signal_2360) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U877_XOR1_U1 ( .A0_t (StateOut[63]), .A0_f (new_AGEMA_signal_2331), .A1_t (new_AGEMA_signal_2332), .A1_f (new_AGEMA_signal_2333), .B0_t (StateFromChi[55]), .B0_f (new_AGEMA_signal_5142), .B1_t (new_AGEMA_signal_5143), .B1_f (new_AGEMA_signal_5144), .Z0_t (U877_X), .Z0_f (new_AGEMA_signal_5379), .Z1_t (new_AGEMA_signal_5380), .Z1_f (new_AGEMA_signal_5381) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U877_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U877_X), .B0_f (new_AGEMA_signal_5379), .B1_t (new_AGEMA_signal_5380), .B1_f (new_AGEMA_signal_5381), .Z0_t (U877_Y), .Z0_f (new_AGEMA_signal_6001), .Z1_t (new_AGEMA_signal_6002), .Z1_f (new_AGEMA_signal_6003) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U877_XOR2_U1 ( .A0_t (U877_Y), .A0_f (new_AGEMA_signal_6001), .A1_t (new_AGEMA_signal_6002), .A1_f (new_AGEMA_signal_6003), .B0_t (StateOut[63]), .B0_f (new_AGEMA_signal_2331), .B1_t (new_AGEMA_signal_2332), .B1_f (new_AGEMA_signal_2333), .Z0_t (StateOut[55]), .Z0_f (new_AGEMA_signal_2328), .Z1_t (new_AGEMA_signal_2329), .Z1_f (new_AGEMA_signal_2330) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U878_XOR1_U1 ( .A0_t (StateOut[119]), .A0_f (new_AGEMA_signal_2484), .A1_t (new_AGEMA_signal_2485), .A1_f (new_AGEMA_signal_2486), .B0_t (StateFromChi[111]), .B0_f (new_AGEMA_signal_5175), .B1_t (new_AGEMA_signal_5176), .B1_f (new_AGEMA_signal_5177), .Z0_t (U878_X), .Z0_f (new_AGEMA_signal_5382), .Z1_t (new_AGEMA_signal_5383), .Z1_f (new_AGEMA_signal_5384) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U878_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U878_X), .B0_f (new_AGEMA_signal_5382), .B1_t (new_AGEMA_signal_5383), .B1_f (new_AGEMA_signal_5384), .Z0_t (U878_Y), .Z0_f (new_AGEMA_signal_6004), .Z1_t (new_AGEMA_signal_6005), .Z1_f (new_AGEMA_signal_6006) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U878_XOR2_U1 ( .A0_t (U878_Y), .A0_f (new_AGEMA_signal_6004), .A1_t (new_AGEMA_signal_6005), .A1_f (new_AGEMA_signal_6006), .B0_t (StateOut[119]), .B0_f (new_AGEMA_signal_2484), .B1_t (new_AGEMA_signal_2485), .B1_f (new_AGEMA_signal_2486), .Z0_t (StateOut[111]), .Z0_f (new_AGEMA_signal_2481), .Z1_t (new_AGEMA_signal_2482), .Z1_f (new_AGEMA_signal_2483) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U879_XOR1_U1 ( .A0_t (StateOut[183]), .A0_f (new_AGEMA_signal_3108), .A1_t (new_AGEMA_signal_3109), .A1_f (new_AGEMA_signal_3110), .B0_t (StateFromChi[175]), .B0_f (new_AGEMA_signal_5151), .B1_t (new_AGEMA_signal_5152), .B1_f (new_AGEMA_signal_5153), .Z0_t (U879_X), .Z0_f (new_AGEMA_signal_5385), .Z1_t (new_AGEMA_signal_5386), .Z1_f (new_AGEMA_signal_5387) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U879_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U879_X), .B0_f (new_AGEMA_signal_5385), .B1_t (new_AGEMA_signal_5386), .B1_f (new_AGEMA_signal_5387), .Z0_t (U879_Y), .Z0_f (new_AGEMA_signal_6007), .Z1_t (new_AGEMA_signal_6008), .Z1_f (new_AGEMA_signal_6009) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U879_XOR2_U1 ( .A0_t (U879_Y), .A0_f (new_AGEMA_signal_6007), .A1_t (new_AGEMA_signal_6008), .A1_f (new_AGEMA_signal_6009), .B0_t (StateOut[183]), .B0_f (new_AGEMA_signal_3108), .B1_t (new_AGEMA_signal_3109), .B1_f (new_AGEMA_signal_3110), .Z0_t (StateOut[175]), .Z0_f (new_AGEMA_signal_2436), .Z1_t (new_AGEMA_signal_2437), .Z1_f (new_AGEMA_signal_2438) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U880_XOR1_U1 ( .A0_t (InData_s0_t[7]), .A0_f (InData_s0_f[7]), .A1_t (InData_s1_t[7]), .A1_f (InData_s1_f[7]), .B0_t (StateFromChi[199]), .B0_f (new_AGEMA_signal_5196), .B1_t (new_AGEMA_signal_5197), .B1_f (new_AGEMA_signal_5198), .Z0_t (U880_X), .Z0_f (new_AGEMA_signal_5391), .Z1_t (new_AGEMA_signal_5392), .Z1_f (new_AGEMA_signal_5393) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U880_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U880_X), .B0_f (new_AGEMA_signal_5391), .B1_t (new_AGEMA_signal_5392), .B1_f (new_AGEMA_signal_5393), .Z0_t (U880_Y), .Z0_f (new_AGEMA_signal_6010), .Z1_t (new_AGEMA_signal_6011), .Z1_f (new_AGEMA_signal_6012) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U880_XOR2_U1 ( .A0_t (U880_Y), .A0_f (new_AGEMA_signal_6010), .A1_t (new_AGEMA_signal_6011), .A1_f (new_AGEMA_signal_6012), .B0_t (InData_s0_t[7]), .B0_f (InData_s0_f[7]), .B1_t (InData_s1_t[7]), .B1_f (InData_s1_f[7]), .Z0_t (StateOut[199]), .Z0_f (new_AGEMA_signal_2448), .Z1_t (new_AGEMA_signal_2449), .Z1_f (new_AGEMA_signal_2450) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U881_XOR1_U1 ( .A0_t (StateOut[30]), .A0_f (new_AGEMA_signal_2142), .A1_t (new_AGEMA_signal_2143), .A1_f (new_AGEMA_signal_2144), .B0_t (StateFromChi[22]), .B0_f (new_AGEMA_signal_5079), .B1_t (new_AGEMA_signal_5080), .B1_f (new_AGEMA_signal_5081), .Z0_t (U881_X), .Z0_f (new_AGEMA_signal_5394), .Z1_t (new_AGEMA_signal_5395), .Z1_f (new_AGEMA_signal_5396) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U881_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U881_X), .B0_f (new_AGEMA_signal_5394), .B1_t (new_AGEMA_signal_5395), .B1_f (new_AGEMA_signal_5396), .Z0_t (U881_Y), .Z0_f (new_AGEMA_signal_6013), .Z1_t (new_AGEMA_signal_6014), .Z1_f (new_AGEMA_signal_6015) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U881_XOR2_U1 ( .A0_t (U881_Y), .A0_f (new_AGEMA_signal_6013), .A1_t (new_AGEMA_signal_6014), .A1_f (new_AGEMA_signal_6015), .B0_t (StateOut[30]), .B0_f (new_AGEMA_signal_2142), .B1_t (new_AGEMA_signal_2143), .B1_f (new_AGEMA_signal_2144), .Z0_t (StateOut[22]), .Z0_f (new_AGEMA_signal_2133), .Z1_t (new_AGEMA_signal_2134), .Z1_f (new_AGEMA_signal_2135) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U882_XOR1_U1 ( .A0_t (StateOut[38]), .A0_f (new_AGEMA_signal_2139), .A1_t (new_AGEMA_signal_2140), .A1_f (new_AGEMA_signal_2141), .B0_t (StateFromChi[30]), .B0_f (new_AGEMA_signal_5094), .B1_t (new_AGEMA_signal_5095), .B1_f (new_AGEMA_signal_5096), .Z0_t (U882_X), .Z0_f (new_AGEMA_signal_5397), .Z1_t (new_AGEMA_signal_5398), .Z1_f (new_AGEMA_signal_5399) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U882_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U882_X), .B0_f (new_AGEMA_signal_5397), .B1_t (new_AGEMA_signal_5398), .B1_f (new_AGEMA_signal_5399), .Z0_t (U882_Y), .Z0_f (new_AGEMA_signal_6016), .Z1_t (new_AGEMA_signal_6017), .Z1_f (new_AGEMA_signal_6018) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U882_XOR2_U1 ( .A0_t (U882_Y), .A0_f (new_AGEMA_signal_6016), .A1_t (new_AGEMA_signal_6017), .A1_f (new_AGEMA_signal_6018), .B0_t (StateOut[38]), .B0_f (new_AGEMA_signal_2139), .B1_t (new_AGEMA_signal_2140), .B1_f (new_AGEMA_signal_2141), .Z0_t (StateOut[30]), .Z0_f (new_AGEMA_signal_2142), .Z1_t (new_AGEMA_signal_2143), .Z1_f (new_AGEMA_signal_2144) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U883_XOR1_U1 ( .A0_t (StateOut[62]), .A0_f (new_AGEMA_signal_3114), .A1_t (new_AGEMA_signal_3115), .A1_f (new_AGEMA_signal_3116), .B0_t (StateFromChi[54]), .B0_f (new_AGEMA_signal_5067), .B1_t (new_AGEMA_signal_5068), .B1_f (new_AGEMA_signal_5069), .Z0_t (U883_X), .Z0_f (new_AGEMA_signal_5400), .Z1_t (new_AGEMA_signal_5401), .Z1_f (new_AGEMA_signal_5402) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U883_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U883_X), .B0_f (new_AGEMA_signal_5400), .B1_t (new_AGEMA_signal_5401), .B1_f (new_AGEMA_signal_5402), .Z0_t (U883_Y), .Z0_f (new_AGEMA_signal_6019), .Z1_t (new_AGEMA_signal_6020), .Z1_f (new_AGEMA_signal_6021) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U883_XOR2_U1 ( .A0_t (U883_Y), .A0_f (new_AGEMA_signal_6019), .A1_t (new_AGEMA_signal_6020), .A1_f (new_AGEMA_signal_6021), .B0_t (StateOut[62]), .B0_f (new_AGEMA_signal_3114), .B1_t (new_AGEMA_signal_3115), .B1_f (new_AGEMA_signal_3116), .Z0_t (StateOut[54]), .Z0_f (new_AGEMA_signal_2454), .Z1_t (new_AGEMA_signal_2455), .Z1_f (new_AGEMA_signal_2456) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U884_XOR1_U1 ( .A0_t (StateOut[94]), .A0_f (new_AGEMA_signal_2688), .A1_t (new_AGEMA_signal_2689), .A1_f (new_AGEMA_signal_2690), .B0_t (StateFromChi[86]), .B0_f (new_AGEMA_signal_5055), .B1_t (new_AGEMA_signal_5056), .B1_f (new_AGEMA_signal_5057), .Z0_t (U884_X), .Z0_f (new_AGEMA_signal_5403), .Z1_t (new_AGEMA_signal_5404), .Z1_f (new_AGEMA_signal_5405) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U884_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U884_X), .B0_f (new_AGEMA_signal_5403), .B1_t (new_AGEMA_signal_5404), .B1_f (new_AGEMA_signal_5405), .Z0_t (U884_Y), .Z0_f (new_AGEMA_signal_6022), .Z1_t (new_AGEMA_signal_6023), .Z1_f (new_AGEMA_signal_6024) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U884_XOR2_U1 ( .A0_t (U884_Y), .A0_f (new_AGEMA_signal_6022), .A1_t (new_AGEMA_signal_6023), .A1_f (new_AGEMA_signal_6024), .B0_t (StateOut[94]), .B0_f (new_AGEMA_signal_2688), .B1_t (new_AGEMA_signal_2689), .B1_f (new_AGEMA_signal_2690), .Z0_t (StateOut[86]), .Z0_f (new_AGEMA_signal_2691), .Z1_t (new_AGEMA_signal_2692), .Z1_f (new_AGEMA_signal_2693) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U885_XOR1_U1 ( .A0_t (StateOut[118]), .A0_f (new_AGEMA_signal_2697), .A1_t (new_AGEMA_signal_2698), .A1_f (new_AGEMA_signal_2699), .B0_t (StateFromChi[110]), .B0_f (new_AGEMA_signal_5100), .B1_t (new_AGEMA_signal_5101), .B1_f (new_AGEMA_signal_5102), .Z0_t (U885_X), .Z0_f (new_AGEMA_signal_5406), .Z1_t (new_AGEMA_signal_5407), .Z1_f (new_AGEMA_signal_5408) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U885_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U885_X), .B0_f (new_AGEMA_signal_5406), .B1_t (new_AGEMA_signal_5407), .B1_f (new_AGEMA_signal_5408), .Z0_t (U885_Y), .Z0_f (new_AGEMA_signal_6025), .Z1_t (new_AGEMA_signal_6026), .Z1_f (new_AGEMA_signal_6027) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U885_XOR2_U1 ( .A0_t (U885_Y), .A0_f (new_AGEMA_signal_6025), .A1_t (new_AGEMA_signal_6026), .A1_f (new_AGEMA_signal_6027), .B0_t (StateOut[118]), .B0_f (new_AGEMA_signal_2697), .B1_t (new_AGEMA_signal_2698), .B1_f (new_AGEMA_signal_2699), .Z0_t (StateOut[110]), .Z0_f (new_AGEMA_signal_3192), .Z1_t (new_AGEMA_signal_3193), .Z1_f (new_AGEMA_signal_3194) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U886_XOR1_U1 ( .A0_t (InData_s0_t[6]), .A0_f (InData_s0_f[6]), .A1_t (InData_s1_t[6]), .A1_f (InData_s1_f[6]), .B0_t (StateFromChi[198]), .B0_f (new_AGEMA_signal_5121), .B1_t (new_AGEMA_signal_5122), .B1_f (new_AGEMA_signal_5123), .Z0_t (U886_X), .Z0_f (new_AGEMA_signal_5412), .Z1_t (new_AGEMA_signal_5413), .Z1_f (new_AGEMA_signal_5414) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U886_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U886_X), .B0_f (new_AGEMA_signal_5412), .B1_t (new_AGEMA_signal_5413), .B1_f (new_AGEMA_signal_5414), .Z0_t (U886_Y), .Z0_f (new_AGEMA_signal_6028), .Z1_t (new_AGEMA_signal_6029), .Z1_f (new_AGEMA_signal_6030) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U886_XOR2_U1 ( .A0_t (U886_Y), .A0_f (new_AGEMA_signal_6028), .A1_t (new_AGEMA_signal_6029), .A1_f (new_AGEMA_signal_6030), .B0_t (InData_s0_t[6]), .B0_f (InData_s0_f[6]), .B1_t (InData_s1_t[6]), .B1_f (InData_s1_f[6]), .Z0_t (StateOut[198]), .Z0_f (new_AGEMA_signal_2502), .Z1_t (new_AGEMA_signal_2503), .Z1_f (new_AGEMA_signal_2504) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U887_XOR1_U1 ( .A0_t (StateOut[29]), .A0_f (new_AGEMA_signal_3174), .A1_t (new_AGEMA_signal_3175), .A1_f (new_AGEMA_signal_3176), .B0_t (StateFromChi[21]), .B0_f (new_AGEMA_signal_5004), .B1_t (new_AGEMA_signal_5005), .B1_f (new_AGEMA_signal_5006), .Z0_t (U887_X), .Z0_f (new_AGEMA_signal_5415), .Z1_t (new_AGEMA_signal_5416), .Z1_f (new_AGEMA_signal_5417) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U887_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U887_X), .B0_f (new_AGEMA_signal_5415), .B1_t (new_AGEMA_signal_5416), .B1_f (new_AGEMA_signal_5417), .Z0_t (U887_Y), .Z0_f (new_AGEMA_signal_6031), .Z1_t (new_AGEMA_signal_6032), .Z1_f (new_AGEMA_signal_6033) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U887_XOR2_U1 ( .A0_t (U887_Y), .A0_f (new_AGEMA_signal_6031), .A1_t (new_AGEMA_signal_6032), .A1_f (new_AGEMA_signal_6033), .B0_t (StateOut[29]), .B0_f (new_AGEMA_signal_3174), .B1_t (new_AGEMA_signal_3175), .B1_f (new_AGEMA_signal_3176), .Z0_t (StateOut[21]), .Z0_f (new_AGEMA_signal_2646), .Z1_t (new_AGEMA_signal_2647), .Z1_f (new_AGEMA_signal_2648) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U888_XOR1_U1 ( .A0_t (StateOut[37]), .A0_f (new_AGEMA_signal_2643), .A1_t (new_AGEMA_signal_2644), .A1_f (new_AGEMA_signal_2645), .B0_t (StateFromChi[29]), .B0_f (new_AGEMA_signal_5019), .B1_t (new_AGEMA_signal_5020), .B1_f (new_AGEMA_signal_5021), .Z0_t (U888_X), .Z0_f (new_AGEMA_signal_5418), .Z1_t (new_AGEMA_signal_5419), .Z1_f (new_AGEMA_signal_5420) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U888_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U888_X), .B0_f (new_AGEMA_signal_5418), .B1_t (new_AGEMA_signal_5419), .B1_f (new_AGEMA_signal_5420), .Z0_t (U888_Y), .Z0_f (new_AGEMA_signal_6034), .Z1_t (new_AGEMA_signal_6035), .Z1_f (new_AGEMA_signal_6036) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U888_XOR2_U1 ( .A0_t (U888_Y), .A0_f (new_AGEMA_signal_6034), .A1_t (new_AGEMA_signal_6035), .A1_f (new_AGEMA_signal_6036), .B0_t (StateOut[37]), .B0_f (new_AGEMA_signal_2643), .B1_t (new_AGEMA_signal_2644), .B1_f (new_AGEMA_signal_2645), .Z0_t (StateOut[29]), .Z0_f (new_AGEMA_signal_3174), .Z1_t (new_AGEMA_signal_3175), .Z1_f (new_AGEMA_signal_3176) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U889_XOR1_U1 ( .A0_t (StateOut[93]), .A0_f (new_AGEMA_signal_2724), .A1_t (new_AGEMA_signal_2725), .A1_f (new_AGEMA_signal_2726), .B0_t (StateFromChi[85]), .B0_f (new_AGEMA_signal_4980), .B1_t (new_AGEMA_signal_4981), .B1_f (new_AGEMA_signal_4982), .Z0_t (U889_X), .Z0_f (new_AGEMA_signal_5421), .Z1_t (new_AGEMA_signal_5422), .Z1_f (new_AGEMA_signal_5423) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U889_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U889_X), .B0_f (new_AGEMA_signal_5421), .B1_t (new_AGEMA_signal_5422), .B1_f (new_AGEMA_signal_5423), .Z0_t (U889_Y), .Z0_f (new_AGEMA_signal_6037), .Z1_t (new_AGEMA_signal_6038), .Z1_f (new_AGEMA_signal_6039) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U889_XOR2_U1 ( .A0_t (U889_Y), .A0_f (new_AGEMA_signal_6037), .A1_t (new_AGEMA_signal_6038), .A1_f (new_AGEMA_signal_6039), .B0_t (StateOut[93]), .B0_f (new_AGEMA_signal_2724), .B1_t (new_AGEMA_signal_2725), .B1_f (new_AGEMA_signal_2726), .Z0_t (StateOut[85]), .Z0_f (new_AGEMA_signal_2727), .Z1_t (new_AGEMA_signal_2728), .Z1_f (new_AGEMA_signal_2729) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U890_XOR1_U1 ( .A0_t (StateOut[141]), .A0_f (new_AGEMA_signal_2547), .A1_t (new_AGEMA_signal_2548), .A1_f (new_AGEMA_signal_2549), .B0_t (StateFromChi[133]), .B0_f (new_AGEMA_signal_4998), .B1_t (new_AGEMA_signal_4999), .B1_f (new_AGEMA_signal_5000), .Z0_t (U890_X), .Z0_f (new_AGEMA_signal_5424), .Z1_t (new_AGEMA_signal_5425), .Z1_f (new_AGEMA_signal_5426) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U890_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U890_X), .B0_f (new_AGEMA_signal_5424), .B1_t (new_AGEMA_signal_5425), .B1_f (new_AGEMA_signal_5426), .Z0_t (U890_Y), .Z0_f (new_AGEMA_signal_6040), .Z1_t (new_AGEMA_signal_6041), .Z1_f (new_AGEMA_signal_6042) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U890_XOR2_U1 ( .A0_t (U890_Y), .A0_f (new_AGEMA_signal_6040), .A1_t (new_AGEMA_signal_6041), .A1_f (new_AGEMA_signal_6042), .B0_t (StateOut[141]), .B0_f (new_AGEMA_signal_2547), .B1_t (new_AGEMA_signal_2548), .B1_f (new_AGEMA_signal_2549), .Z0_t (StateOut[133]), .Z0_f (new_AGEMA_signal_2544), .Z1_t (new_AGEMA_signal_2545), .Z1_f (new_AGEMA_signal_2546) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U891_XOR1_U1 ( .A0_t (StateOut[52]), .A0_f (new_AGEMA_signal_2598), .A1_t (new_AGEMA_signal_2599), .A1_f (new_AGEMA_signal_2600), .B0_t (StateFromChi[44]), .B0_f (new_AGEMA_signal_4902), .B1_t (new_AGEMA_signal_4903), .B1_f (new_AGEMA_signal_4904), .Z0_t (U891_X), .Z0_f (new_AGEMA_signal_5427), .Z1_t (new_AGEMA_signal_5428), .Z1_f (new_AGEMA_signal_5429) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U891_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U891_X), .B0_f (new_AGEMA_signal_5427), .B1_t (new_AGEMA_signal_5428), .B1_f (new_AGEMA_signal_5429), .Z0_t (U891_Y), .Z0_f (new_AGEMA_signal_6043), .Z1_t (new_AGEMA_signal_6044), .Z1_f (new_AGEMA_signal_6045) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U891_XOR2_U1 ( .A0_t (U891_Y), .A0_f (new_AGEMA_signal_6043), .A1_t (new_AGEMA_signal_6044), .A1_f (new_AGEMA_signal_6045), .B0_t (StateOut[52]), .B0_f (new_AGEMA_signal_2598), .B1_t (new_AGEMA_signal_2599), .B1_f (new_AGEMA_signal_2600), .Z0_t (StateOut[44]), .Z0_f (new_AGEMA_signal_2601), .Z1_t (new_AGEMA_signal_2602), .Z1_f (new_AGEMA_signal_2603) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U892_XOR1_U1 ( .A0_t (StateOut[76]), .A0_f (new_AGEMA_signal_2610), .A1_t (new_AGEMA_signal_2611), .A1_f (new_AGEMA_signal_2612), .B0_t (StateFromChi[68]), .B0_f (new_AGEMA_signal_4947), .B1_t (new_AGEMA_signal_4948), .B1_f (new_AGEMA_signal_4949), .Z0_t (U892_X), .Z0_f (new_AGEMA_signal_5430), .Z1_t (new_AGEMA_signal_5431), .Z1_f (new_AGEMA_signal_5432) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U892_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U892_X), .B0_f (new_AGEMA_signal_5430), .B1_t (new_AGEMA_signal_5431), .B1_f (new_AGEMA_signal_5432), .Z0_t (U892_Y), .Z0_f (new_AGEMA_signal_6046), .Z1_t (new_AGEMA_signal_6047), .Z1_f (new_AGEMA_signal_6048) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U892_XOR2_U1 ( .A0_t (U892_Y), .A0_f (new_AGEMA_signal_6046), .A1_t (new_AGEMA_signal_6047), .A1_f (new_AGEMA_signal_6048), .B0_t (StateOut[76]), .B0_f (new_AGEMA_signal_2610), .B1_t (new_AGEMA_signal_2611), .B1_f (new_AGEMA_signal_2612), .Z0_t (StateOut[68]), .Z0_f (new_AGEMA_signal_2607), .Z1_t (new_AGEMA_signal_2608), .Z1_f (new_AGEMA_signal_2609) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U893_XOR1_U1 ( .A0_t (StateOut[140]), .A0_f (new_AGEMA_signal_2367), .A1_t (new_AGEMA_signal_2368), .A1_f (new_AGEMA_signal_2369), .B0_t (StateFromChi[132]), .B0_f (new_AGEMA_signal_4923), .B1_t (new_AGEMA_signal_4924), .B1_f (new_AGEMA_signal_4925), .Z0_t (U893_X), .Z0_f (new_AGEMA_signal_5433), .Z1_t (new_AGEMA_signal_5434), .Z1_f (new_AGEMA_signal_5435) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U893_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U893_X), .B0_f (new_AGEMA_signal_5433), .B1_t (new_AGEMA_signal_5434), .B1_f (new_AGEMA_signal_5435), .Z0_t (U893_Y), .Z0_f (new_AGEMA_signal_6049), .Z1_t (new_AGEMA_signal_6050), .Z1_f (new_AGEMA_signal_6051) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U893_XOR2_U1 ( .A0_t (U893_Y), .A0_f (new_AGEMA_signal_6049), .A1_t (new_AGEMA_signal_6050), .A1_f (new_AGEMA_signal_6051), .B0_t (StateOut[140]), .B0_f (new_AGEMA_signal_2367), .B1_t (new_AGEMA_signal_2368), .B1_f (new_AGEMA_signal_2369), .Z0_t (StateOut[132]), .Z0_f (new_AGEMA_signal_2364), .Z1_t (new_AGEMA_signal_2365), .Z1_f (new_AGEMA_signal_2366) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U894_XOR1_U1 ( .A0_t (StateOut[148]), .A0_f (new_AGEMA_signal_2376), .A1_t (new_AGEMA_signal_2377), .A1_f (new_AGEMA_signal_2378), .B0_t (StateFromChi[140]), .B0_f (new_AGEMA_signal_4938), .B1_t (new_AGEMA_signal_4939), .B1_f (new_AGEMA_signal_4940), .Z0_t (U894_X), .Z0_f (new_AGEMA_signal_5436), .Z1_t (new_AGEMA_signal_5437), .Z1_f (new_AGEMA_signal_5438) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U894_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U894_X), .B0_f (new_AGEMA_signal_5436), .B1_t (new_AGEMA_signal_5437), .B1_f (new_AGEMA_signal_5438), .Z0_t (U894_Y), .Z0_f (new_AGEMA_signal_6052), .Z1_t (new_AGEMA_signal_6053), .Z1_f (new_AGEMA_signal_6054) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U894_XOR2_U1 ( .A0_t (U894_Y), .A0_f (new_AGEMA_signal_6052), .A1_t (new_AGEMA_signal_6053), .A1_f (new_AGEMA_signal_6054), .B0_t (StateOut[148]), .B0_f (new_AGEMA_signal_2376), .B1_t (new_AGEMA_signal_2377), .B1_f (new_AGEMA_signal_2378), .Z0_t (StateOut[140]), .Z0_f (new_AGEMA_signal_2367), .Z1_t (new_AGEMA_signal_2368), .Z1_f (new_AGEMA_signal_2369) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U895_XOR1_U1 ( .A0_t (StateOut[156]), .A0_f (new_AGEMA_signal_2373), .A1_t (new_AGEMA_signal_2374), .A1_f (new_AGEMA_signal_2375), .B0_t (StateFromChi[148]), .B0_f (new_AGEMA_signal_4953), .B1_t (new_AGEMA_signal_4954), .B1_f (new_AGEMA_signal_4955), .Z0_t (U895_X), .Z0_f (new_AGEMA_signal_5439), .Z1_t (new_AGEMA_signal_5440), .Z1_f (new_AGEMA_signal_5441) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U895_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U895_X), .B0_f (new_AGEMA_signal_5439), .B1_t (new_AGEMA_signal_5440), .B1_f (new_AGEMA_signal_5441), .Z0_t (U895_Y), .Z0_f (new_AGEMA_signal_6055), .Z1_t (new_AGEMA_signal_6056), .Z1_f (new_AGEMA_signal_6057) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U895_XOR2_U1 ( .A0_t (U895_Y), .A0_f (new_AGEMA_signal_6055), .A1_t (new_AGEMA_signal_6056), .A1_f (new_AGEMA_signal_6057), .B0_t (StateOut[156]), .B0_f (new_AGEMA_signal_2373), .B1_t (new_AGEMA_signal_2374), .B1_f (new_AGEMA_signal_2375), .Z0_t (StateOut[148]), .Z0_f (new_AGEMA_signal_2376), .Z1_t (new_AGEMA_signal_2377), .Z1_f (new_AGEMA_signal_2378) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U896_XOR1_U1 ( .A0_t (StateOut[43]), .A0_f (new_AGEMA_signal_2619), .A1_t (new_AGEMA_signal_2620), .A1_f (new_AGEMA_signal_2621), .B0_t (StateFromChi[35]), .B0_f (new_AGEMA_signal_4884), .B1_t (new_AGEMA_signal_4885), .B1_f (new_AGEMA_signal_4886), .Z0_t (U896_X), .Z0_f (new_AGEMA_signal_5442), .Z1_t (new_AGEMA_signal_5443), .Z1_f (new_AGEMA_signal_5444) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U896_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U896_X), .B0_f (new_AGEMA_signal_5442), .B1_t (new_AGEMA_signal_5443), .B1_f (new_AGEMA_signal_5444), .Z0_t (U896_Y), .Z0_f (new_AGEMA_signal_6058), .Z1_t (new_AGEMA_signal_6059), .Z1_f (new_AGEMA_signal_6060) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U896_XOR2_U1 ( .A0_t (U896_Y), .A0_f (new_AGEMA_signal_6058), .A1_t (new_AGEMA_signal_6059), .A1_f (new_AGEMA_signal_6060), .B0_t (StateOut[43]), .B0_f (new_AGEMA_signal_2619), .B1_t (new_AGEMA_signal_2620), .B1_f (new_AGEMA_signal_2621), .Z0_t (StateOut[35]), .Z0_f (new_AGEMA_signal_2193), .Z1_t (new_AGEMA_signal_2194), .Z1_f (new_AGEMA_signal_2195) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U897_XOR1_U1 ( .A0_t (StateOut[51]), .A0_f (new_AGEMA_signal_2616), .A1_t (new_AGEMA_signal_2617), .A1_f (new_AGEMA_signal_2618), .B0_t (StateFromChi[43]), .B0_f (new_AGEMA_signal_4827), .B1_t (new_AGEMA_signal_4828), .B1_f (new_AGEMA_signal_4829), .Z0_t (U897_X), .Z0_f (new_AGEMA_signal_5445), .Z1_t (new_AGEMA_signal_5446), .Z1_f (new_AGEMA_signal_5447) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U897_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U897_X), .B0_f (new_AGEMA_signal_5445), .B1_t (new_AGEMA_signal_5446), .B1_f (new_AGEMA_signal_5447), .Z0_t (U897_Y), .Z0_f (new_AGEMA_signal_6061), .Z1_t (new_AGEMA_signal_6062), .Z1_f (new_AGEMA_signal_6063) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U897_XOR2_U1 ( .A0_t (U897_Y), .A0_f (new_AGEMA_signal_6061), .A1_t (new_AGEMA_signal_6062), .A1_f (new_AGEMA_signal_6063), .B0_t (StateOut[51]), .B0_f (new_AGEMA_signal_2616), .B1_t (new_AGEMA_signal_2617), .B1_f (new_AGEMA_signal_2618), .Z0_t (StateOut[43]), .Z0_f (new_AGEMA_signal_2619), .Z1_t (new_AGEMA_signal_2620), .Z1_f (new_AGEMA_signal_2621) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U898_XOR1_U1 ( .A0_t (StateOut[67]), .A0_f (new_AGEMA_signal_2625), .A1_t (new_AGEMA_signal_2626), .A1_f (new_AGEMA_signal_2627), .B0_t (StateFromChi[59]), .B0_f (new_AGEMA_signal_4857), .B1_t (new_AGEMA_signal_4858), .B1_f (new_AGEMA_signal_4859), .Z0_t (U898_X), .Z0_f (new_AGEMA_signal_5448), .Z1_t (new_AGEMA_signal_5449), .Z1_f (new_AGEMA_signal_5450) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U898_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U898_X), .B0_f (new_AGEMA_signal_5448), .B1_t (new_AGEMA_signal_5449), .B1_f (new_AGEMA_signal_5450), .Z0_t (U898_Y), .Z0_f (new_AGEMA_signal_6064), .Z1_t (new_AGEMA_signal_6065), .Z1_f (new_AGEMA_signal_6066) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U898_XOR2_U1 ( .A0_t (U898_Y), .A0_f (new_AGEMA_signal_6064), .A1_t (new_AGEMA_signal_6065), .A1_f (new_AGEMA_signal_6066), .B0_t (StateOut[67]), .B0_f (new_AGEMA_signal_2625), .B1_t (new_AGEMA_signal_2626), .B1_f (new_AGEMA_signal_2627), .Z0_t (StateOut[59]), .Z0_f (new_AGEMA_signal_3168), .Z1_t (new_AGEMA_signal_3169), .Z1_f (new_AGEMA_signal_3170) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U899_XOR1_U1 ( .A0_t (StateOut[75]), .A0_f (new_AGEMA_signal_2628), .A1_t (new_AGEMA_signal_2629), .A1_f (new_AGEMA_signal_2630), .B0_t (StateFromChi[67]), .B0_f (new_AGEMA_signal_4872), .B1_t (new_AGEMA_signal_4873), .B1_f (new_AGEMA_signal_4874), .Z0_t (U899_X), .Z0_f (new_AGEMA_signal_5451), .Z1_t (new_AGEMA_signal_5452), .Z1_f (new_AGEMA_signal_5453) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U899_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U899_X), .B0_f (new_AGEMA_signal_5451), .B1_t (new_AGEMA_signal_5452), .B1_f (new_AGEMA_signal_5453), .Z0_t (U899_Y), .Z0_f (new_AGEMA_signal_6067), .Z1_t (new_AGEMA_signal_6068), .Z1_f (new_AGEMA_signal_6069) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U899_XOR2_U1 ( .A0_t (U899_Y), .A0_f (new_AGEMA_signal_6067), .A1_t (new_AGEMA_signal_6068), .A1_f (new_AGEMA_signal_6069), .B0_t (StateOut[75]), .B0_f (new_AGEMA_signal_2628), .B1_t (new_AGEMA_signal_2629), .B1_f (new_AGEMA_signal_2630), .Z0_t (StateOut[67]), .Z0_f (new_AGEMA_signal_2625), .Z1_t (new_AGEMA_signal_2626), .Z1_f (new_AGEMA_signal_2627) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U900_XOR1_U1 ( .A0_t (StateOut[99]), .A0_f (new_AGEMA_signal_2826), .A1_t (new_AGEMA_signal_2827), .A1_f (new_AGEMA_signal_2828), .B0_t (StateFromChi[91]), .B0_f (new_AGEMA_signal_4845), .B1_t (new_AGEMA_signal_4846), .B1_f (new_AGEMA_signal_4847), .Z0_t (U900_X), .Z0_f (new_AGEMA_signal_5454), .Z1_t (new_AGEMA_signal_5455), .Z1_f (new_AGEMA_signal_5456) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U900_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U900_X), .B0_f (new_AGEMA_signal_5454), .B1_t (new_AGEMA_signal_5455), .B1_f (new_AGEMA_signal_5456), .Z0_t (U900_Y), .Z0_f (new_AGEMA_signal_6070), .Z1_t (new_AGEMA_signal_6071), .Z1_f (new_AGEMA_signal_6072) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U900_XOR2_U1 ( .A0_t (U900_Y), .A0_f (new_AGEMA_signal_6070), .A1_t (new_AGEMA_signal_6071), .A1_f (new_AGEMA_signal_6072), .B0_t (StateOut[99]), .B0_f (new_AGEMA_signal_2826), .B1_t (new_AGEMA_signal_2827), .B1_f (new_AGEMA_signal_2828), .Z0_t (StateOut[91]), .Z0_f (new_AGEMA_signal_2814), .Z1_t (new_AGEMA_signal_2815), .Z1_f (new_AGEMA_signal_2816) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U901_XOR1_U1 ( .A0_t (StateOut[123]), .A0_f (new_AGEMA_signal_3156), .A1_t (new_AGEMA_signal_3157), .A1_f (new_AGEMA_signal_3158), .B0_t (StateFromChi[115]), .B0_f (new_AGEMA_signal_4890), .B1_t (new_AGEMA_signal_4891), .B1_f (new_AGEMA_signal_4892), .Z0_t (U901_X), .Z0_f (new_AGEMA_signal_5457), .Z1_t (new_AGEMA_signal_5458), .Z1_f (new_AGEMA_signal_5459) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U901_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U901_X), .B0_f (new_AGEMA_signal_5457), .B1_t (new_AGEMA_signal_5458), .B1_f (new_AGEMA_signal_5459), .Z0_t (U901_Y), .Z0_f (new_AGEMA_signal_6073), .Z1_t (new_AGEMA_signal_6074), .Z1_f (new_AGEMA_signal_6075) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U901_XOR2_U1 ( .A0_t (U901_Y), .A0_f (new_AGEMA_signal_6073), .A1_t (new_AGEMA_signal_6074), .A1_f (new_AGEMA_signal_6075), .B0_t (StateOut[123]), .B0_f (new_AGEMA_signal_3156), .B1_t (new_AGEMA_signal_3157), .B1_f (new_AGEMA_signal_3158), .Z0_t (StateOut[115]), .Z0_f (new_AGEMA_signal_2823), .Z1_t (new_AGEMA_signal_2824), .Z1_f (new_AGEMA_signal_2825) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U902_XOR1_U1 ( .A0_t (StateOut[139]), .A0_f (new_AGEMA_signal_2583), .A1_t (new_AGEMA_signal_2584), .A1_f (new_AGEMA_signal_2585), .B0_t (StateFromChi[131]), .B0_f (new_AGEMA_signal_4848), .B1_t (new_AGEMA_signal_4849), .B1_f (new_AGEMA_signal_4850), .Z0_t (U902_X), .Z0_f (new_AGEMA_signal_5460), .Z1_t (new_AGEMA_signal_5461), .Z1_f (new_AGEMA_signal_5462) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U902_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U902_X), .B0_f (new_AGEMA_signal_5460), .B1_t (new_AGEMA_signal_5461), .B1_f (new_AGEMA_signal_5462), .Z0_t (U902_Y), .Z0_f (new_AGEMA_signal_6076), .Z1_t (new_AGEMA_signal_6077), .Z1_f (new_AGEMA_signal_6078) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U902_XOR2_U1 ( .A0_t (U902_Y), .A0_f (new_AGEMA_signal_6076), .A1_t (new_AGEMA_signal_6077), .A1_f (new_AGEMA_signal_6078), .B0_t (StateOut[139]), .B0_f (new_AGEMA_signal_2583), .B1_t (new_AGEMA_signal_2584), .B1_f (new_AGEMA_signal_2585), .Z0_t (StateOut[131]), .Z0_f (new_AGEMA_signal_2580), .Z1_t (new_AGEMA_signal_2581), .Z1_f (new_AGEMA_signal_2582) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U903_XOR1_U1 ( .A0_t (StateOut[147]), .A0_f (new_AGEMA_signal_2592), .A1_t (new_AGEMA_signal_2593), .A1_f (new_AGEMA_signal_2594), .B0_t (StateFromChi[139]), .B0_f (new_AGEMA_signal_4863), .B1_t (new_AGEMA_signal_4864), .B1_f (new_AGEMA_signal_4865), .Z0_t (U903_X), .Z0_f (new_AGEMA_signal_5463), .Z1_t (new_AGEMA_signal_5464), .Z1_f (new_AGEMA_signal_5465) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U903_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U903_X), .B0_f (new_AGEMA_signal_5463), .B1_t (new_AGEMA_signal_5464), .B1_f (new_AGEMA_signal_5465), .Z0_t (U903_Y), .Z0_f (new_AGEMA_signal_6079), .Z1_t (new_AGEMA_signal_6080), .Z1_f (new_AGEMA_signal_6081) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U903_XOR2_U1 ( .A0_t (U903_Y), .A0_f (new_AGEMA_signal_6079), .A1_t (new_AGEMA_signal_6080), .A1_f (new_AGEMA_signal_6081), .B0_t (StateOut[147]), .B0_f (new_AGEMA_signal_2592), .B1_t (new_AGEMA_signal_2593), .B1_f (new_AGEMA_signal_2594), .Z0_t (StateOut[139]), .Z0_f (new_AGEMA_signal_2583), .Z1_t (new_AGEMA_signal_2584), .Z1_f (new_AGEMA_signal_2585) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U904_XOR1_U1 ( .A0_t (StateOut[50]), .A0_f (new_AGEMA_signal_2652), .A1_t (new_AGEMA_signal_2653), .A1_f (new_AGEMA_signal_2654), .B0_t (StateFromChi[42]), .B0_f (new_AGEMA_signal_4752), .B1_t (new_AGEMA_signal_4753), .B1_f (new_AGEMA_signal_4754), .Z0_t (U904_X), .Z0_f (new_AGEMA_signal_5466), .Z1_t (new_AGEMA_signal_5467), .Z1_f (new_AGEMA_signal_5468) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U904_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U904_X), .B0_f (new_AGEMA_signal_5466), .B1_t (new_AGEMA_signal_5467), .B1_f (new_AGEMA_signal_5468), .Z0_t (U904_Y), .Z0_f (new_AGEMA_signal_6082), .Z1_t (new_AGEMA_signal_6083), .Z1_f (new_AGEMA_signal_6084) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U904_XOR2_U1 ( .A0_t (U904_Y), .A0_f (new_AGEMA_signal_6082), .A1_t (new_AGEMA_signal_6083), .A1_f (new_AGEMA_signal_6084), .B0_t (StateOut[50]), .B0_f (new_AGEMA_signal_2652), .B1_t (new_AGEMA_signal_2653), .B1_f (new_AGEMA_signal_2654), .Z0_t (StateOut[42]), .Z0_f (new_AGEMA_signal_2655), .Z1_t (new_AGEMA_signal_2656), .Z1_f (new_AGEMA_signal_2657) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U905_XOR1_U1 ( .A0_t (StateOut[98]), .A0_f (new_AGEMA_signal_2223), .A1_t (new_AGEMA_signal_2224), .A1_f (new_AGEMA_signal_2225), .B0_t (StateFromChi[90]), .B0_f (new_AGEMA_signal_4770), .B1_t (new_AGEMA_signal_4771), .B1_f (new_AGEMA_signal_4772), .Z0_t (U905_X), .Z0_f (new_AGEMA_signal_5469), .Z1_t (new_AGEMA_signal_5470), .Z1_f (new_AGEMA_signal_5471) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U905_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U905_X), .B0_f (new_AGEMA_signal_5469), .B1_t (new_AGEMA_signal_5470), .B1_f (new_AGEMA_signal_5471), .Z0_t (U905_Y), .Z0_f (new_AGEMA_signal_6085), .Z1_t (new_AGEMA_signal_6086), .Z1_f (new_AGEMA_signal_6087) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U905_XOR2_U1 ( .A0_t (U905_Y), .A0_f (new_AGEMA_signal_6085), .A1_t (new_AGEMA_signal_6086), .A1_f (new_AGEMA_signal_6087), .B0_t (StateOut[98]), .B0_f (new_AGEMA_signal_2223), .B1_t (new_AGEMA_signal_2224), .B1_f (new_AGEMA_signal_2225), .Z0_t (StateOut[90]), .Z0_f (new_AGEMA_signal_2220), .Z1_t (new_AGEMA_signal_2221), .Z1_f (new_AGEMA_signal_2222) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U906_XOR1_U1 ( .A0_t (StateOut[114]), .A0_f (new_AGEMA_signal_2229), .A1_t (new_AGEMA_signal_2230), .A1_f (new_AGEMA_signal_2231), .B0_t (StateFromChi[106]), .B0_f (new_AGEMA_signal_4800), .B1_t (new_AGEMA_signal_4801), .B1_f (new_AGEMA_signal_4802), .Z0_t (U906_X), .Z0_f (new_AGEMA_signal_5472), .Z1_t (new_AGEMA_signal_5473), .Z1_f (new_AGEMA_signal_5474) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U906_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U906_X), .B0_f (new_AGEMA_signal_5472), .B1_t (new_AGEMA_signal_5473), .B1_f (new_AGEMA_signal_5474), .Z0_t (U906_Y), .Z0_f (new_AGEMA_signal_6088), .Z1_t (new_AGEMA_signal_6089), .Z1_f (new_AGEMA_signal_6090) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U906_XOR2_U1 ( .A0_t (U906_Y), .A0_f (new_AGEMA_signal_6088), .A1_t (new_AGEMA_signal_6089), .A1_f (new_AGEMA_signal_6090), .B0_t (StateOut[114]), .B0_f (new_AGEMA_signal_2229), .B1_t (new_AGEMA_signal_2230), .B1_f (new_AGEMA_signal_2231), .Z0_t (StateOut[106]), .Z0_f (new_AGEMA_signal_2232), .Z1_t (new_AGEMA_signal_2233), .Z1_f (new_AGEMA_signal_2234) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U907_XOR1_U1 ( .A0_t (StateOut[122]), .A0_f (new_AGEMA_signal_2745), .A1_t (new_AGEMA_signal_2746), .A1_f (new_AGEMA_signal_2747), .B0_t (StateFromChi[114]), .B0_f (new_AGEMA_signal_4815), .B1_t (new_AGEMA_signal_4816), .B1_f (new_AGEMA_signal_4817), .Z0_t (U907_X), .Z0_f (new_AGEMA_signal_5475), .Z1_t (new_AGEMA_signal_5476), .Z1_f (new_AGEMA_signal_5477) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U907_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U907_X), .B0_f (new_AGEMA_signal_5475), .B1_t (new_AGEMA_signal_5476), .B1_f (new_AGEMA_signal_5477), .Z0_t (U907_Y), .Z0_f (new_AGEMA_signal_6091), .Z1_t (new_AGEMA_signal_6092), .Z1_f (new_AGEMA_signal_6093) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U907_XOR2_U1 ( .A0_t (U907_Y), .A0_f (new_AGEMA_signal_6091), .A1_t (new_AGEMA_signal_6092), .A1_f (new_AGEMA_signal_6093), .B0_t (StateOut[122]), .B0_f (new_AGEMA_signal_2745), .B1_t (new_AGEMA_signal_2746), .B1_f (new_AGEMA_signal_2747), .Z0_t (StateOut[114]), .Z0_f (new_AGEMA_signal_2229), .Z1_t (new_AGEMA_signal_2230), .Z1_f (new_AGEMA_signal_2231) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U908_XOR1_U1 ( .A0_t (StateOut[138]), .A0_f (new_AGEMA_signal_3210), .A1_t (new_AGEMA_signal_3211), .A1_f (new_AGEMA_signal_3212), .B0_t (StateFromChi[130]), .B0_f (new_AGEMA_signal_4773), .B1_t (new_AGEMA_signal_4774), .B1_f (new_AGEMA_signal_4775), .Z0_t (U908_X), .Z0_f (new_AGEMA_signal_5478), .Z1_t (new_AGEMA_signal_5479), .Z1_f (new_AGEMA_signal_5480) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U908_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U908_X), .B0_f (new_AGEMA_signal_5478), .B1_t (new_AGEMA_signal_5479), .B1_f (new_AGEMA_signal_5480), .Z0_t (U908_Y), .Z0_f (new_AGEMA_signal_6094), .Z1_t (new_AGEMA_signal_6095), .Z1_f (new_AGEMA_signal_6096) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U908_XOR2_U1 ( .A0_t (U908_Y), .A0_f (new_AGEMA_signal_6094), .A1_t (new_AGEMA_signal_6095), .A1_f (new_AGEMA_signal_6096), .B0_t (StateOut[138]), .B0_f (new_AGEMA_signal_3210), .B1_t (new_AGEMA_signal_3211), .B1_f (new_AGEMA_signal_3212), .Z0_t (StateOut[130]), .Z0_f (new_AGEMA_signal_2742), .Z1_t (new_AGEMA_signal_2743), .Z1_f (new_AGEMA_signal_2744) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U909_XOR1_U1 ( .A0_t (StateOut[146]), .A0_f (new_AGEMA_signal_2751), .A1_t (new_AGEMA_signal_2752), .A1_f (new_AGEMA_signal_2753), .B0_t (StateFromChi[138]), .B0_f (new_AGEMA_signal_4788), .B1_t (new_AGEMA_signal_4789), .B1_f (new_AGEMA_signal_4790), .Z0_t (U909_X), .Z0_f (new_AGEMA_signal_5481), .Z1_t (new_AGEMA_signal_5482), .Z1_f (new_AGEMA_signal_5483) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U909_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U909_X), .B0_f (new_AGEMA_signal_5481), .B1_t (new_AGEMA_signal_5482), .B1_f (new_AGEMA_signal_5483), .Z0_t (U909_Y), .Z0_f (new_AGEMA_signal_6097), .Z1_t (new_AGEMA_signal_6098), .Z1_f (new_AGEMA_signal_6099) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U909_XOR2_U1 ( .A0_t (U909_Y), .A0_f (new_AGEMA_signal_6097), .A1_t (new_AGEMA_signal_6098), .A1_f (new_AGEMA_signal_6099), .B0_t (StateOut[146]), .B0_f (new_AGEMA_signal_2751), .B1_t (new_AGEMA_signal_2752), .B1_f (new_AGEMA_signal_2753), .Z0_t (StateOut[138]), .Z0_f (new_AGEMA_signal_3210), .Z1_t (new_AGEMA_signal_3211), .Z1_f (new_AGEMA_signal_3212) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U910_XOR1_U1 ( .A0_t (StateOut[154]), .A0_f (new_AGEMA_signal_2754), .A1_t (new_AGEMA_signal_2755), .A1_f (new_AGEMA_signal_2756), .B0_t (StateFromChi[146]), .B0_f (new_AGEMA_signal_4803), .B1_t (new_AGEMA_signal_4804), .B1_f (new_AGEMA_signal_4805), .Z0_t (U910_X), .Z0_f (new_AGEMA_signal_5484), .Z1_t (new_AGEMA_signal_5485), .Z1_f (new_AGEMA_signal_5486) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U910_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U910_X), .B0_f (new_AGEMA_signal_5484), .B1_t (new_AGEMA_signal_5485), .B1_f (new_AGEMA_signal_5486), .Z0_t (U910_Y), .Z0_f (new_AGEMA_signal_6100), .Z1_t (new_AGEMA_signal_6101), .Z1_f (new_AGEMA_signal_6102) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U910_XOR2_U1 ( .A0_t (U910_Y), .A0_f (new_AGEMA_signal_6100), .A1_t (new_AGEMA_signal_6101), .A1_f (new_AGEMA_signal_6102), .B0_t (StateOut[154]), .B0_f (new_AGEMA_signal_2754), .B1_t (new_AGEMA_signal_2755), .B1_f (new_AGEMA_signal_2756), .Z0_t (StateOut[146]), .Z0_f (new_AGEMA_signal_2751), .Z1_t (new_AGEMA_signal_2752), .Z1_f (new_AGEMA_signal_2753) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U911_XOR1_U1 ( .A0_t (StateOut[170]), .A0_f (new_AGEMA_signal_2832), .A1_t (new_AGEMA_signal_2833), .A1_f (new_AGEMA_signal_2834), .B0_t (StateFromChi[162]), .B0_f (new_AGEMA_signal_4761), .B1_t (new_AGEMA_signal_4762), .B1_f (new_AGEMA_signal_4763), .Z0_t (U911_X), .Z0_f (new_AGEMA_signal_5487), .Z1_t (new_AGEMA_signal_5488), .Z1_f (new_AGEMA_signal_5489) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U911_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U911_X), .B0_f (new_AGEMA_signal_5487), .B1_t (new_AGEMA_signal_5488), .B1_f (new_AGEMA_signal_5489), .Z0_t (U911_Y), .Z0_f (new_AGEMA_signal_6103), .Z1_t (new_AGEMA_signal_6104), .Z1_f (new_AGEMA_signal_6105) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U911_XOR2_U1 ( .A0_t (U911_Y), .A0_f (new_AGEMA_signal_6103), .A1_t (new_AGEMA_signal_6104), .A1_f (new_AGEMA_signal_6105), .B0_t (StateOut[170]), .B0_f (new_AGEMA_signal_2832), .B1_t (new_AGEMA_signal_2833), .B1_f (new_AGEMA_signal_2834), .Z0_t (StateOut[162]), .Z0_f (new_AGEMA_signal_2835), .Z1_t (new_AGEMA_signal_2836), .Z1_f (new_AGEMA_signal_2837) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U912_XOR1_U1 ( .A0_t (StateOut[178]), .A0_f (new_AGEMA_signal_2844), .A1_t (new_AGEMA_signal_2845), .A1_f (new_AGEMA_signal_2846), .B0_t (StateFromChi[170]), .B0_f (new_AGEMA_signal_4776), .B1_t (new_AGEMA_signal_4777), .B1_f (new_AGEMA_signal_4778), .Z0_t (U912_X), .Z0_f (new_AGEMA_signal_5490), .Z1_t (new_AGEMA_signal_5491), .Z1_f (new_AGEMA_signal_5492) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U912_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U912_X), .B0_f (new_AGEMA_signal_5490), .B1_t (new_AGEMA_signal_5491), .B1_f (new_AGEMA_signal_5492), .Z0_t (U912_Y), .Z0_f (new_AGEMA_signal_6106), .Z1_t (new_AGEMA_signal_6107), .Z1_f (new_AGEMA_signal_6108) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U912_XOR2_U1 ( .A0_t (U912_Y), .A0_f (new_AGEMA_signal_6106), .A1_t (new_AGEMA_signal_6107), .A1_f (new_AGEMA_signal_6108), .B0_t (StateOut[178]), .B0_f (new_AGEMA_signal_2844), .B1_t (new_AGEMA_signal_2845), .B1_f (new_AGEMA_signal_2846), .Z0_t (StateOut[170]), .Z0_f (new_AGEMA_signal_2832), .Z1_t (new_AGEMA_signal_2833), .Z1_f (new_AGEMA_signal_2834) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U913_XOR1_U1 ( .A0_t (StateOut[186]), .A0_f (new_AGEMA_signal_3240), .A1_t (new_AGEMA_signal_3241), .A1_f (new_AGEMA_signal_3242), .B0_t (StateFromChi[178]), .B0_f (new_AGEMA_signal_4791), .B1_t (new_AGEMA_signal_4792), .B1_f (new_AGEMA_signal_4793), .Z0_t (U913_X), .Z0_f (new_AGEMA_signal_5493), .Z1_t (new_AGEMA_signal_5494), .Z1_f (new_AGEMA_signal_5495) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U913_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U913_X), .B0_f (new_AGEMA_signal_5493), .B1_t (new_AGEMA_signal_5494), .B1_f (new_AGEMA_signal_5495), .Z0_t (U913_Y), .Z0_f (new_AGEMA_signal_6109), .Z1_t (new_AGEMA_signal_6110), .Z1_f (new_AGEMA_signal_6111) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U913_XOR2_U1 ( .A0_t (U913_Y), .A0_f (new_AGEMA_signal_6109), .A1_t (new_AGEMA_signal_6110), .A1_f (new_AGEMA_signal_6111), .B0_t (StateOut[186]), .B0_f (new_AGEMA_signal_3240), .B1_t (new_AGEMA_signal_3241), .B1_f (new_AGEMA_signal_3242), .Z0_t (StateOut[178]), .Z0_f (new_AGEMA_signal_2844), .Z1_t (new_AGEMA_signal_2845), .Z1_f (new_AGEMA_signal_2846) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U914_XOR1_U1 ( .A0_t (InData_s0_t[2]), .A0_f (InData_s0_f[2]), .A1_t (InData_s1_t[2]), .A1_f (InData_s1_f[2]), .B0_t (StateFromChi[194]), .B0_f (new_AGEMA_signal_4821), .B1_t (new_AGEMA_signal_4822), .B1_f (new_AGEMA_signal_4823), .Z0_t (U914_X), .Z0_f (new_AGEMA_signal_5499), .Z1_t (new_AGEMA_signal_5500), .Z1_f (new_AGEMA_signal_5501) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U914_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U914_X), .B0_f (new_AGEMA_signal_5499), .B1_t (new_AGEMA_signal_5500), .B1_f (new_AGEMA_signal_5501), .Z0_t (U914_Y), .Z0_f (new_AGEMA_signal_6112), .Z1_t (new_AGEMA_signal_6113), .Z1_f (new_AGEMA_signal_6114) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U914_XOR2_U1 ( .A0_t (U914_Y), .A0_f (new_AGEMA_signal_6112), .A1_t (new_AGEMA_signal_6113), .A1_f (new_AGEMA_signal_6114), .B0_t (InData_s0_t[2]), .B0_f (InData_s0_f[2]), .B1_t (InData_s1_t[2]), .B1_f (InData_s1_f[2]), .Z0_t (StateOut[194]), .Z0_f (new_AGEMA_signal_2841), .Z1_t (new_AGEMA_signal_2842), .Z1_f (new_AGEMA_signal_2843) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U915_XOR1_U1 ( .A0_t (StateOut[25]), .A0_f (new_AGEMA_signal_2769), .A1_t (new_AGEMA_signal_2770), .A1_f (new_AGEMA_signal_2771), .B0_t (StateFromChi[17]), .B0_f (new_AGEMA_signal_4704), .B1_t (new_AGEMA_signal_4705), .B1_f (new_AGEMA_signal_4706), .Z0_t (U915_X), .Z0_f (new_AGEMA_signal_5502), .Z1_t (new_AGEMA_signal_5503), .Z1_f (new_AGEMA_signal_5504) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U915_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U915_X), .B0_f (new_AGEMA_signal_5502), .B1_t (new_AGEMA_signal_5503), .B1_f (new_AGEMA_signal_5504), .Z0_t (U915_Y), .Z0_f (new_AGEMA_signal_6115), .Z1_t (new_AGEMA_signal_6116), .Z1_f (new_AGEMA_signal_6117) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U915_XOR2_U1 ( .A0_t (U915_Y), .A0_f (new_AGEMA_signal_6115), .A1_t (new_AGEMA_signal_6116), .A1_f (new_AGEMA_signal_6117), .B0_t (StateOut[25]), .B0_f (new_AGEMA_signal_2769), .B1_t (new_AGEMA_signal_2770), .B1_f (new_AGEMA_signal_2771), .Z0_t (StateOut[17]), .Z0_f (new_AGEMA_signal_3216), .Z1_t (new_AGEMA_signal_3217), .Z1_f (new_AGEMA_signal_3218) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U916_XOR1_U1 ( .A0_t (StateOut[41]), .A0_f (new_AGEMA_signal_2421), .A1_t (new_AGEMA_signal_2422), .A1_f (new_AGEMA_signal_2423), .B0_t (StateFromChi[33]), .B0_f (new_AGEMA_signal_4734), .B1_t (new_AGEMA_signal_4735), .B1_f (new_AGEMA_signal_4736), .Z0_t (U916_X), .Z0_f (new_AGEMA_signal_5505), .Z1_t (new_AGEMA_signal_5506), .Z1_f (new_AGEMA_signal_5507) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U916_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U916_X), .B0_f (new_AGEMA_signal_5505), .B1_t (new_AGEMA_signal_5506), .B1_f (new_AGEMA_signal_5507), .Z0_t (U916_Y), .Z0_f (new_AGEMA_signal_6118), .Z1_t (new_AGEMA_signal_6119), .Z1_f (new_AGEMA_signal_6120) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U916_XOR2_U1 ( .A0_t (U916_Y), .A0_f (new_AGEMA_signal_6118), .A1_t (new_AGEMA_signal_6119), .A1_f (new_AGEMA_signal_6120), .B0_t (StateOut[41]), .B0_f (new_AGEMA_signal_2421), .B1_t (new_AGEMA_signal_2422), .B1_f (new_AGEMA_signal_2423), .Z0_t (StateOut[33]), .Z0_f (new_AGEMA_signal_2772), .Z1_t (new_AGEMA_signal_2773), .Z1_f (new_AGEMA_signal_2774) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U917_XOR1_U1 ( .A0_t (StateOut[49]), .A0_f (new_AGEMA_signal_2418), .A1_t (new_AGEMA_signal_2419), .A1_f (new_AGEMA_signal_2420), .B0_t (StateFromChi[41]), .B0_f (new_AGEMA_signal_4677), .B1_t (new_AGEMA_signal_4678), .B1_f (new_AGEMA_signal_4679), .Z0_t (U917_X), .Z0_f (new_AGEMA_signal_5508), .Z1_t (new_AGEMA_signal_5509), .Z1_f (new_AGEMA_signal_5510) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U917_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U917_X), .B0_f (new_AGEMA_signal_5508), .B1_t (new_AGEMA_signal_5509), .B1_f (new_AGEMA_signal_5510), .Z0_t (U917_Y), .Z0_f (new_AGEMA_signal_6121), .Z1_t (new_AGEMA_signal_6122), .Z1_f (new_AGEMA_signal_6123) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U917_XOR2_U1 ( .A0_t (U917_Y), .A0_f (new_AGEMA_signal_6121), .A1_t (new_AGEMA_signal_6122), .A1_f (new_AGEMA_signal_6123), .B0_t (StateOut[49]), .B0_f (new_AGEMA_signal_2418), .B1_t (new_AGEMA_signal_2419), .B1_f (new_AGEMA_signal_2420), .Z0_t (StateOut[41]), .Z0_f (new_AGEMA_signal_2421), .Z1_t (new_AGEMA_signal_2422), .Z1_f (new_AGEMA_signal_2423) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U918_XOR1_U1 ( .A0_t (StateOut[65]), .A0_f (new_AGEMA_signal_2427), .A1_t (new_AGEMA_signal_2428), .A1_f (new_AGEMA_signal_2429), .B0_t (StateFromChi[57]), .B0_f (new_AGEMA_signal_4707), .B1_t (new_AGEMA_signal_4708), .B1_f (new_AGEMA_signal_4709), .Z0_t (U918_X), .Z0_f (new_AGEMA_signal_5511), .Z1_t (new_AGEMA_signal_5512), .Z1_f (new_AGEMA_signal_5513) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U918_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U918_X), .B0_f (new_AGEMA_signal_5511), .B1_t (new_AGEMA_signal_5512), .B1_f (new_AGEMA_signal_5513), .Z0_t (U918_Y), .Z0_f (new_AGEMA_signal_6124), .Z1_t (new_AGEMA_signal_6125), .Z1_f (new_AGEMA_signal_6126) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U918_XOR2_U1 ( .A0_t (U918_Y), .A0_f (new_AGEMA_signal_6124), .A1_t (new_AGEMA_signal_6125), .A1_f (new_AGEMA_signal_6126), .B0_t (StateOut[65]), .B0_f (new_AGEMA_signal_2427), .B1_t (new_AGEMA_signal_2428), .B1_f (new_AGEMA_signal_2429), .Z0_t (StateOut[57]), .Z0_f (new_AGEMA_signal_3102), .Z1_t (new_AGEMA_signal_3103), .Z1_f (new_AGEMA_signal_3104) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U919_XOR1_U1 ( .A0_t (StateOut[113]), .A0_f (new_AGEMA_signal_2301), .A1_t (new_AGEMA_signal_2302), .A1_f (new_AGEMA_signal_2303), .B0_t (StateFromChi[105]), .B0_f (new_AGEMA_signal_4725), .B1_t (new_AGEMA_signal_4726), .B1_f (new_AGEMA_signal_4727), .Z0_t (U919_X), .Z0_f (new_AGEMA_signal_5514), .Z1_t (new_AGEMA_signal_5515), .Z1_f (new_AGEMA_signal_5516) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U919_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U919_X), .B0_f (new_AGEMA_signal_5514), .B1_t (new_AGEMA_signal_5515), .B1_f (new_AGEMA_signal_5516), .Z0_t (U919_Y), .Z0_f (new_AGEMA_signal_6127), .Z1_t (new_AGEMA_signal_6128), .Z1_f (new_AGEMA_signal_6129) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U919_XOR2_U1 ( .A0_t (U919_Y), .A0_f (new_AGEMA_signal_6127), .A1_t (new_AGEMA_signal_6128), .A1_f (new_AGEMA_signal_6129), .B0_t (StateOut[113]), .B0_f (new_AGEMA_signal_2301), .B1_t (new_AGEMA_signal_2302), .B1_f (new_AGEMA_signal_2303), .Z0_t (StateOut[105]), .Z0_f (new_AGEMA_signal_2304), .Z1_t (new_AGEMA_signal_2305), .Z1_f (new_AGEMA_signal_2306) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U920_XOR1_U1 ( .A0_t (StateOut[121]), .A0_f (new_AGEMA_signal_3054), .A1_t (new_AGEMA_signal_3055), .A1_f (new_AGEMA_signal_3056), .B0_t (StateFromChi[113]), .B0_f (new_AGEMA_signal_4740), .B1_t (new_AGEMA_signal_4741), .B1_f (new_AGEMA_signal_4742), .Z0_t (U920_X), .Z0_f (new_AGEMA_signal_5517), .Z1_t (new_AGEMA_signal_5518), .Z1_f (new_AGEMA_signal_5519) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U920_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U920_X), .B0_f (new_AGEMA_signal_5517), .B1_t (new_AGEMA_signal_5518), .B1_f (new_AGEMA_signal_5519), .Z0_t (U920_Y), .Z0_f (new_AGEMA_signal_6130), .Z1_t (new_AGEMA_signal_6131), .Z1_f (new_AGEMA_signal_6132) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U920_XOR2_U1 ( .A0_t (U920_Y), .A0_f (new_AGEMA_signal_6130), .A1_t (new_AGEMA_signal_6131), .A1_f (new_AGEMA_signal_6132), .B0_t (StateOut[121]), .B0_f (new_AGEMA_signal_3054), .B1_t (new_AGEMA_signal_3055), .B1_f (new_AGEMA_signal_3056), .Z0_t (StateOut[113]), .Z0_f (new_AGEMA_signal_2301), .Z1_t (new_AGEMA_signal_2302), .Z1_f (new_AGEMA_signal_2303) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U921_XOR1_U1 ( .A0_t (StateOut[137]), .A0_f (new_AGEMA_signal_2277), .A1_t (new_AGEMA_signal_2278), .A1_f (new_AGEMA_signal_2279), .B0_t (StateFromChi[129]), .B0_f (new_AGEMA_signal_4698), .B1_t (new_AGEMA_signal_4699), .B1_f (new_AGEMA_signal_4700), .Z0_t (U921_X), .Z0_f (new_AGEMA_signal_5520), .Z1_t (new_AGEMA_signal_5521), .Z1_f (new_AGEMA_signal_5522) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U921_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U921_X), .B0_f (new_AGEMA_signal_5520), .B1_t (new_AGEMA_signal_5521), .B1_f (new_AGEMA_signal_5522), .Z0_t (U921_Y), .Z0_f (new_AGEMA_signal_6133), .Z1_t (new_AGEMA_signal_6134), .Z1_f (new_AGEMA_signal_6135) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U921_XOR2_U1 ( .A0_t (U921_Y), .A0_f (new_AGEMA_signal_6133), .A1_t (new_AGEMA_signal_6134), .A1_f (new_AGEMA_signal_6135), .B0_t (StateOut[137]), .B0_f (new_AGEMA_signal_2277), .B1_t (new_AGEMA_signal_2278), .B1_f (new_AGEMA_signal_2279), .Z0_t (StateOut[129]), .Z0_f (new_AGEMA_signal_2274), .Z1_t (new_AGEMA_signal_2275), .Z1_f (new_AGEMA_signal_2276) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U922_XOR1_U1 ( .A0_t (StateOut[153]), .A0_f (new_AGEMA_signal_2283), .A1_t (new_AGEMA_signal_2284), .A1_f (new_AGEMA_signal_2285), .B0_t (StateFromChi[145]), .B0_f (new_AGEMA_signal_4728), .B1_t (new_AGEMA_signal_4729), .B1_f (new_AGEMA_signal_4730), .Z0_t (U922_X), .Z0_f (new_AGEMA_signal_5523), .Z1_t (new_AGEMA_signal_5524), .Z1_f (new_AGEMA_signal_5525) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U922_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U922_X), .B0_f (new_AGEMA_signal_5523), .B1_t (new_AGEMA_signal_5524), .B1_f (new_AGEMA_signal_5525), .Z0_t (U922_Y), .Z0_f (new_AGEMA_signal_6136), .Z1_t (new_AGEMA_signal_6137), .Z1_f (new_AGEMA_signal_6138) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U922_XOR2_U1 ( .A0_t (U922_Y), .A0_f (new_AGEMA_signal_6136), .A1_t (new_AGEMA_signal_6137), .A1_f (new_AGEMA_signal_6138), .B0_t (StateOut[153]), .B0_f (new_AGEMA_signal_2283), .B1_t (new_AGEMA_signal_2284), .B1_f (new_AGEMA_signal_2285), .Z0_t (StateOut[145]), .Z0_f (new_AGEMA_signal_2286), .Z1_t (new_AGEMA_signal_2287), .Z1_f (new_AGEMA_signal_2288) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U923_XOR1_U1 ( .A0_t (StateOut[161]), .A0_f (new_AGEMA_signal_2241), .A1_t (new_AGEMA_signal_2242), .A1_f (new_AGEMA_signal_2243), .B0_t (StateFromChi[153]), .B0_f (new_AGEMA_signal_4743), .B1_t (new_AGEMA_signal_4744), .B1_f (new_AGEMA_signal_4745), .Z0_t (U923_X), .Z0_f (new_AGEMA_signal_5526), .Z1_t (new_AGEMA_signal_5527), .Z1_f (new_AGEMA_signal_5528) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U923_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U923_X), .B0_f (new_AGEMA_signal_5526), .B1_t (new_AGEMA_signal_5527), .B1_f (new_AGEMA_signal_5528), .Z0_t (U923_Y), .Z0_f (new_AGEMA_signal_6139), .Z1_t (new_AGEMA_signal_6140), .Z1_f (new_AGEMA_signal_6141) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U923_XOR2_U1 ( .A0_t (U923_Y), .A0_f (new_AGEMA_signal_6139), .A1_t (new_AGEMA_signal_6140), .A1_f (new_AGEMA_signal_6141), .B0_t (StateOut[161]), .B0_f (new_AGEMA_signal_2241), .B1_t (new_AGEMA_signal_2242), .B1_f (new_AGEMA_signal_2243), .Z0_t (StateOut[153]), .Z0_f (new_AGEMA_signal_2283), .Z1_t (new_AGEMA_signal_2284), .Z1_f (new_AGEMA_signal_2285) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U924_XOR1_U1 ( .A0_t (StateOut[169]), .A0_f (new_AGEMA_signal_2238), .A1_t (new_AGEMA_signal_2239), .A1_f (new_AGEMA_signal_2240), .B0_t (StateFromChi[161]), .B0_f (new_AGEMA_signal_4686), .B1_t (new_AGEMA_signal_4687), .B1_f (new_AGEMA_signal_4688), .Z0_t (U924_X), .Z0_f (new_AGEMA_signal_5529), .Z1_t (new_AGEMA_signal_5530), .Z1_f (new_AGEMA_signal_5531) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U924_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U924_X), .B0_f (new_AGEMA_signal_5529), .B1_t (new_AGEMA_signal_5530), .B1_f (new_AGEMA_signal_5531), .Z0_t (U924_Y), .Z0_f (new_AGEMA_signal_6142), .Z1_t (new_AGEMA_signal_6143), .Z1_f (new_AGEMA_signal_6144) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U924_XOR2_U1 ( .A0_t (U924_Y), .A0_f (new_AGEMA_signal_6142), .A1_t (new_AGEMA_signal_6143), .A1_f (new_AGEMA_signal_6144), .B0_t (StateOut[169]), .B0_f (new_AGEMA_signal_2238), .B1_t (new_AGEMA_signal_2239), .B1_f (new_AGEMA_signal_2240), .Z0_t (StateOut[161]), .Z0_f (new_AGEMA_signal_2241), .Z1_t (new_AGEMA_signal_2242), .Z1_f (new_AGEMA_signal_2243) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U925_XOR1_U1 ( .A0_t (StateOut[185]), .A0_f (new_AGEMA_signal_2247), .A1_t (new_AGEMA_signal_2248), .A1_f (new_AGEMA_signal_2249), .B0_t (StateFromChi[177]), .B0_f (new_AGEMA_signal_4716), .B1_t (new_AGEMA_signal_4717), .B1_f (new_AGEMA_signal_4718), .Z0_t (U925_X), .Z0_f (new_AGEMA_signal_5532), .Z1_t (new_AGEMA_signal_5533), .Z1_f (new_AGEMA_signal_5534) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U925_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U925_X), .B0_f (new_AGEMA_signal_5532), .B1_t (new_AGEMA_signal_5533), .B1_f (new_AGEMA_signal_5534), .Z0_t (U925_Y), .Z0_f (new_AGEMA_signal_6145), .Z1_t (new_AGEMA_signal_6146), .Z1_f (new_AGEMA_signal_6147) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U925_XOR2_U1 ( .A0_t (U925_Y), .A0_f (new_AGEMA_signal_6145), .A1_t (new_AGEMA_signal_6146), .A1_f (new_AGEMA_signal_6147), .B0_t (StateOut[185]), .B0_f (new_AGEMA_signal_2247), .B1_t (new_AGEMA_signal_2248), .B1_f (new_AGEMA_signal_2249), .Z0_t (StateOut[177]), .Z0_f (new_AGEMA_signal_3042), .Z1_t (new_AGEMA_signal_3043), .Z1_f (new_AGEMA_signal_3044) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U926_XOR1_U1 ( .A0_t (InData_s0_t[1]), .A0_f (InData_s0_f[1]), .A1_t (InData_s1_t[1]), .A1_f (InData_s1_f[1]), .B0_t (StateFromChi[193]), .B0_f (new_AGEMA_signal_4746), .B1_t (new_AGEMA_signal_4747), .B1_f (new_AGEMA_signal_4748), .Z0_t (U926_X), .Z0_f (new_AGEMA_signal_5538), .Z1_t (new_AGEMA_signal_5539), .Z1_f (new_AGEMA_signal_5540) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U926_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U926_X), .B0_f (new_AGEMA_signal_5538), .B1_t (new_AGEMA_signal_5539), .B1_f (new_AGEMA_signal_5540), .Z0_t (U926_Y), .Z0_f (new_AGEMA_signal_6148), .Z1_t (new_AGEMA_signal_6149), .Z1_f (new_AGEMA_signal_6150) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U926_XOR2_U1 ( .A0_t (U926_Y), .A0_f (new_AGEMA_signal_6148), .A1_t (new_AGEMA_signal_6149), .A1_f (new_AGEMA_signal_6150), .B0_t (InData_s0_t[1]), .B0_f (InData_s0_f[1]), .B1_t (InData_s1_t[1]), .B1_f (InData_s1_f[1]), .Z0_t (StateOut[193]), .Z0_f (new_AGEMA_signal_2250), .Z1_t (new_AGEMA_signal_2251), .Z1_f (new_AGEMA_signal_2252) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U927_XOR1_U1 ( .A0_t (StateOut[24]), .A0_f (new_AGEMA_signal_2214), .A1_t (new_AGEMA_signal_2215), .A1_f (new_AGEMA_signal_2216), .B0_t (StateFromChi[16]), .B0_f (new_AGEMA_signal_4629), .B1_t (new_AGEMA_signal_4630), .B1_f (new_AGEMA_signal_4631), .Z0_t (U927_X), .Z0_f (new_AGEMA_signal_5541), .Z1_t (new_AGEMA_signal_5542), .Z1_f (new_AGEMA_signal_5543) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U927_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U927_X), .B0_f (new_AGEMA_signal_5541), .B1_t (new_AGEMA_signal_5542), .B1_f (new_AGEMA_signal_5543), .Z0_t (U927_Y), .Z0_f (new_AGEMA_signal_6151), .Z1_t (new_AGEMA_signal_6152), .Z1_f (new_AGEMA_signal_6153) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U927_XOR2_U1 ( .A0_t (U927_Y), .A0_f (new_AGEMA_signal_6151), .A1_t (new_AGEMA_signal_6152), .A1_f (new_AGEMA_signal_6153), .B0_t (StateOut[24]), .B0_f (new_AGEMA_signal_2214), .B1_t (new_AGEMA_signal_2215), .B1_f (new_AGEMA_signal_2216), .Z0_t (StateOut[16]), .Z0_f (new_AGEMA_signal_2205), .Z1_t (new_AGEMA_signal_2206), .Z1_f (new_AGEMA_signal_2207) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U928_XOR1_U1 ( .A0_t (StateOut[40]), .A0_f (new_AGEMA_signal_2259), .A1_t (new_AGEMA_signal_2260), .A1_f (new_AGEMA_signal_2261), .B0_t (StateFromChi[32]), .B0_f (new_AGEMA_signal_4659), .B1_t (new_AGEMA_signal_4660), .B1_f (new_AGEMA_signal_4661), .Z0_t (U928_X), .Z0_f (new_AGEMA_signal_5544), .Z1_t (new_AGEMA_signal_5545), .Z1_f (new_AGEMA_signal_5546) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U928_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U928_X), .B0_f (new_AGEMA_signal_5544), .B1_t (new_AGEMA_signal_5545), .B1_f (new_AGEMA_signal_5546), .Z0_t (U928_Y), .Z0_f (new_AGEMA_signal_6154), .Z1_t (new_AGEMA_signal_6155), .Z1_f (new_AGEMA_signal_6156) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U928_XOR2_U1 ( .A0_t (U928_Y), .A0_f (new_AGEMA_signal_6154), .A1_t (new_AGEMA_signal_6155), .A1_f (new_AGEMA_signal_6156), .B0_t (StateOut[40]), .B0_f (new_AGEMA_signal_2259), .B1_t (new_AGEMA_signal_2260), .B1_f (new_AGEMA_signal_2261), .Z0_t (StateOut[32]), .Z0_f (new_AGEMA_signal_2211), .Z1_t (new_AGEMA_signal_2212), .Z1_f (new_AGEMA_signal_2213) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U929_XOR1_U1 ( .A0_t (StateOut[48]), .A0_f (new_AGEMA_signal_2256), .A1_t (new_AGEMA_signal_2257), .A1_f (new_AGEMA_signal_2258), .B0_t (StateFromChi[40]), .B0_f (new_AGEMA_signal_4602), .B1_t (new_AGEMA_signal_4603), .B1_f (new_AGEMA_signal_4604), .Z0_t (U929_X), .Z0_f (new_AGEMA_signal_5547), .Z1_t (new_AGEMA_signal_5548), .Z1_f (new_AGEMA_signal_5549) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U929_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U929_X), .B0_f (new_AGEMA_signal_5547), .B1_t (new_AGEMA_signal_5548), .B1_f (new_AGEMA_signal_5549), .Z0_t (U929_Y), .Z0_f (new_AGEMA_signal_6157), .Z1_t (new_AGEMA_signal_6158), .Z1_f (new_AGEMA_signal_6159) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U929_XOR2_U1 ( .A0_t (U929_Y), .A0_f (new_AGEMA_signal_6157), .A1_t (new_AGEMA_signal_6158), .A1_f (new_AGEMA_signal_6159), .B0_t (StateOut[48]), .B0_f (new_AGEMA_signal_2256), .B1_t (new_AGEMA_signal_2257), .B1_f (new_AGEMA_signal_2258), .Z0_t (StateOut[40]), .Z0_f (new_AGEMA_signal_2259), .Z1_t (new_AGEMA_signal_2260), .Z1_f (new_AGEMA_signal_2261) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U930_XOR1_U1 ( .A0_t (StateOut[56]), .A0_f (new_AGEMA_signal_2268), .A1_t (new_AGEMA_signal_2269), .A1_f (new_AGEMA_signal_2270), .B0_t (StateFromChi[48]), .B0_f (new_AGEMA_signal_4617), .B1_t (new_AGEMA_signal_4618), .B1_f (new_AGEMA_signal_4619), .Z0_t (U930_X), .Z0_f (new_AGEMA_signal_5550), .Z1_t (new_AGEMA_signal_5551), .Z1_f (new_AGEMA_signal_5552) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U930_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U930_X), .B0_f (new_AGEMA_signal_5550), .B1_t (new_AGEMA_signal_5551), .B1_f (new_AGEMA_signal_5552), .Z0_t (U930_Y), .Z0_f (new_AGEMA_signal_6160), .Z1_t (new_AGEMA_signal_6161), .Z1_f (new_AGEMA_signal_6162) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U930_XOR2_U1 ( .A0_t (U930_Y), .A0_f (new_AGEMA_signal_6160), .A1_t (new_AGEMA_signal_6161), .A1_f (new_AGEMA_signal_6162), .B0_t (StateOut[56]), .B0_f (new_AGEMA_signal_2268), .B1_t (new_AGEMA_signal_2269), .B1_f (new_AGEMA_signal_2270), .Z0_t (StateOut[48]), .Z0_f (new_AGEMA_signal_2256), .Z1_t (new_AGEMA_signal_2257), .Z1_f (new_AGEMA_signal_2258) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U931_XOR1_U1 ( .A0_t (StateOut[64]), .A0_f (new_AGEMA_signal_3048), .A1_t (new_AGEMA_signal_3049), .A1_f (new_AGEMA_signal_3050), .B0_t (StateFromChi[56]), .B0_f (new_AGEMA_signal_4632), .B1_t (new_AGEMA_signal_4633), .B1_f (new_AGEMA_signal_4634), .Z0_t (U931_X), .Z0_f (new_AGEMA_signal_5553), .Z1_t (new_AGEMA_signal_5554), .Z1_f (new_AGEMA_signal_5555) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U931_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U931_X), .B0_f (new_AGEMA_signal_5553), .B1_t (new_AGEMA_signal_5554), .B1_f (new_AGEMA_signal_5555), .Z0_t (U931_Y), .Z0_f (new_AGEMA_signal_6163), .Z1_t (new_AGEMA_signal_6164), .Z1_f (new_AGEMA_signal_6165) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U931_XOR2_U1 ( .A0_t (U931_Y), .A0_f (new_AGEMA_signal_6163), .A1_t (new_AGEMA_signal_6164), .A1_f (new_AGEMA_signal_6165), .B0_t (StateOut[64]), .B0_f (new_AGEMA_signal_3048), .B1_t (new_AGEMA_signal_3049), .B1_f (new_AGEMA_signal_3050), .Z0_t (StateOut[56]), .Z0_f (new_AGEMA_signal_2268), .Z1_t (new_AGEMA_signal_2269), .Z1_f (new_AGEMA_signal_2270) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U932_XOR1_U1 ( .A0_t (StateOut[88]), .A0_f (new_AGEMA_signal_2382), .A1_t (new_AGEMA_signal_2383), .A1_f (new_AGEMA_signal_2384), .B0_t (StateFromChi[80]), .B0_f (new_AGEMA_signal_4605), .B1_t (new_AGEMA_signal_4606), .B1_f (new_AGEMA_signal_4607), .Z0_t (U932_X), .Z0_f (new_AGEMA_signal_5556), .Z1_t (new_AGEMA_signal_5557), .Z1_f (new_AGEMA_signal_5558) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U932_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U932_X), .B0_f (new_AGEMA_signal_5556), .B1_t (new_AGEMA_signal_5557), .B1_f (new_AGEMA_signal_5558), .Z0_t (U932_Y), .Z0_f (new_AGEMA_signal_6166), .Z1_t (new_AGEMA_signal_6167), .Z1_f (new_AGEMA_signal_6168) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U932_XOR2_U1 ( .A0_t (U932_Y), .A0_f (new_AGEMA_signal_6166), .A1_t (new_AGEMA_signal_6167), .A1_f (new_AGEMA_signal_6168), .B0_t (StateOut[88]), .B0_f (new_AGEMA_signal_2382), .B1_t (new_AGEMA_signal_2383), .B1_f (new_AGEMA_signal_2384), .Z0_t (StateOut[80]), .Z0_f (new_AGEMA_signal_2385), .Z1_t (new_AGEMA_signal_2386), .Z1_f (new_AGEMA_signal_2387) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U933_XOR1_U1 ( .A0_t (StateOut[112]), .A0_f (new_AGEMA_signal_2394), .A1_t (new_AGEMA_signal_2395), .A1_f (new_AGEMA_signal_2396), .B0_t (StateFromChi[104]), .B0_f (new_AGEMA_signal_4650), .B1_t (new_AGEMA_signal_4651), .B1_f (new_AGEMA_signal_4652), .Z0_t (U933_X), .Z0_f (new_AGEMA_signal_5559), .Z1_t (new_AGEMA_signal_5560), .Z1_f (new_AGEMA_signal_5561) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U933_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U933_X), .B0_f (new_AGEMA_signal_5559), .B1_t (new_AGEMA_signal_5560), .B1_f (new_AGEMA_signal_5561), .Z0_t (U933_Y), .Z0_f (new_AGEMA_signal_6169), .Z1_t (new_AGEMA_signal_6170), .Z1_f (new_AGEMA_signal_6171) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U933_XOR2_U1 ( .A0_t (U933_Y), .A0_f (new_AGEMA_signal_6169), .A1_t (new_AGEMA_signal_6170), .A1_f (new_AGEMA_signal_6171), .B0_t (StateOut[112]), .B0_f (new_AGEMA_signal_2394), .B1_t (new_AGEMA_signal_2395), .B1_f (new_AGEMA_signal_2396), .Z0_t (StateOut[104]), .Z0_f (new_AGEMA_signal_2391), .Z1_t (new_AGEMA_signal_2392), .Z1_f (new_AGEMA_signal_2393) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U934_XOR1_U1 ( .A0_t (StateOut[160]), .A0_f (new_AGEMA_signal_3066), .A1_t (new_AGEMA_signal_3067), .A1_f (new_AGEMA_signal_3068), .B0_t (StateFromChi[152]), .B0_f (new_AGEMA_signal_4668), .B1_t (new_AGEMA_signal_4669), .B1_f (new_AGEMA_signal_4670), .Z0_t (U934_X), .Z0_f (new_AGEMA_signal_5562), .Z1_t (new_AGEMA_signal_5563), .Z1_f (new_AGEMA_signal_5564) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U934_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U934_X), .B0_f (new_AGEMA_signal_5562), .B1_t (new_AGEMA_signal_5563), .B1_f (new_AGEMA_signal_5564), .Z0_t (U934_Y), .Z0_f (new_AGEMA_signal_6172), .Z1_t (new_AGEMA_signal_6173), .Z1_f (new_AGEMA_signal_6174) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U934_XOR2_U1 ( .A0_t (U934_Y), .A0_f (new_AGEMA_signal_6172), .A1_t (new_AGEMA_signal_6173), .A1_f (new_AGEMA_signal_6174), .B0_t (StateOut[160]), .B0_f (new_AGEMA_signal_3066), .B1_t (new_AGEMA_signal_3067), .B1_f (new_AGEMA_signal_3068), .Z0_t (StateOut[152]), .Z0_f (new_AGEMA_signal_2409), .Z1_t (new_AGEMA_signal_2410), .Z1_f (new_AGEMA_signal_2411) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U935_XOR1_U1 ( .A0_t (StateOut[168]), .A0_f (new_AGEMA_signal_2310), .A1_t (new_AGEMA_signal_2311), .A1_f (new_AGEMA_signal_2312), .B0_t (StateFromChi[160]), .B0_f (new_AGEMA_signal_4611), .B1_t (new_AGEMA_signal_4612), .B1_f (new_AGEMA_signal_4613), .Z0_t (U935_X), .Z0_f (new_AGEMA_signal_5565), .Z1_t (new_AGEMA_signal_5566), .Z1_f (new_AGEMA_signal_5567) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U935_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U935_X), .B0_f (new_AGEMA_signal_5565), .B1_t (new_AGEMA_signal_5566), .B1_f (new_AGEMA_signal_5567), .Z0_t (U935_Y), .Z0_f (new_AGEMA_signal_6175), .Z1_t (new_AGEMA_signal_6176), .Z1_f (new_AGEMA_signal_6177) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U935_XOR2_U1 ( .A0_t (U935_Y), .A0_f (new_AGEMA_signal_6175), .A1_t (new_AGEMA_signal_6176), .A1_f (new_AGEMA_signal_6177), .B0_t (StateOut[168]), .B0_f (new_AGEMA_signal_2310), .B1_t (new_AGEMA_signal_2311), .B1_f (new_AGEMA_signal_2312), .Z0_t (StateOut[160]), .Z0_f (new_AGEMA_signal_3066), .Z1_t (new_AGEMA_signal_3067), .Z1_f (new_AGEMA_signal_3068) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U936_XOR1_U1 ( .A0_t (StateOut[176]), .A0_f (new_AGEMA_signal_2313), .A1_t (new_AGEMA_signal_2314), .A1_f (new_AGEMA_signal_2315), .B0_t (StateFromChi[168]), .B0_f (new_AGEMA_signal_4626), .B1_t (new_AGEMA_signal_4627), .B1_f (new_AGEMA_signal_4628), .Z0_t (U936_X), .Z0_f (new_AGEMA_signal_5568), .Z1_t (new_AGEMA_signal_5569), .Z1_f (new_AGEMA_signal_5570) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U936_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U936_X), .B0_f (new_AGEMA_signal_5568), .B1_t (new_AGEMA_signal_5569), .B1_f (new_AGEMA_signal_5570), .Z0_t (U936_Y), .Z0_f (new_AGEMA_signal_6178), .Z1_t (new_AGEMA_signal_6179), .Z1_f (new_AGEMA_signal_6180) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U936_XOR2_U1 ( .A0_t (U936_Y), .A0_f (new_AGEMA_signal_6178), .A1_t (new_AGEMA_signal_6179), .A1_f (new_AGEMA_signal_6180), .B0_t (StateOut[176]), .B0_f (new_AGEMA_signal_2313), .B1_t (new_AGEMA_signal_2314), .B1_f (new_AGEMA_signal_2315), .Z0_t (StateOut[168]), .Z0_f (new_AGEMA_signal_2310), .Z1_t (new_AGEMA_signal_2311), .Z1_f (new_AGEMA_signal_2312) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U937_XOR1_U1 ( .A0_t (InData_s0_t[0]), .A0_f (InData_s0_f[0]), .A1_t (InData_s1_t[0]), .A1_f (InData_s1_f[0]), .B0_t (StateFromChi[192]), .B0_f (new_AGEMA_signal_4671), .B1_t (new_AGEMA_signal_4672), .B1_f (new_AGEMA_signal_4673), .Z0_t (U937_X), .Z0_f (new_AGEMA_signal_5574), .Z1_t (new_AGEMA_signal_5575), .Z1_f (new_AGEMA_signal_5576) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U937_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U937_X), .B0_f (new_AGEMA_signal_5574), .B1_t (new_AGEMA_signal_5575), .B1_f (new_AGEMA_signal_5576), .Z0_t (U937_Y), .Z0_f (new_AGEMA_signal_6181), .Z1_t (new_AGEMA_signal_6182), .Z1_f (new_AGEMA_signal_6183) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U937_XOR2_U1 ( .A0_t (U937_Y), .A0_f (new_AGEMA_signal_6181), .A1_t (new_AGEMA_signal_6182), .A1_f (new_AGEMA_signal_6183), .B0_t (InData_s0_t[0]), .B0_f (InData_s0_f[0]), .B1_t (InData_s1_t[0]), .B1_f (InData_s1_f[0]), .Z0_t (StateOut[192]), .Z0_f (new_AGEMA_signal_2319), .Z1_t (new_AGEMA_signal_2320), .Z1_f (new_AGEMA_signal_2321) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U938_XOR1_U1 ( .A0_t (StateOut[23]), .A0_f (new_AGEMA_signal_2349), .A1_t (new_AGEMA_signal_2350), .A1_f (new_AGEMA_signal_2351), .B0_t (StateFromChi[15]), .B0_f (new_AGEMA_signal_5139), .B1_t (new_AGEMA_signal_5140), .B1_f (new_AGEMA_signal_5141), .Z0_t (U938_X), .Z0_f (new_AGEMA_signal_5577), .Z1_t (new_AGEMA_signal_5578), .Z1_f (new_AGEMA_signal_5579) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U938_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U938_X), .B0_f (new_AGEMA_signal_5577), .B1_t (new_AGEMA_signal_5578), .B1_f (new_AGEMA_signal_5579), .Z0_t (U938_Y), .Z0_f (new_AGEMA_signal_6184), .Z1_t (new_AGEMA_signal_6185), .Z1_f (new_AGEMA_signal_6186) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U938_XOR2_U1 ( .A0_t (U938_Y), .A0_f (new_AGEMA_signal_6184), .A1_t (new_AGEMA_signal_6185), .A1_f (new_AGEMA_signal_6186), .B0_t (StateOut[23]), .B0_f (new_AGEMA_signal_2349), .B1_t (new_AGEMA_signal_2350), .B1_f (new_AGEMA_signal_2351), .Z0_t (StateOut[15]), .Z0_f (new_AGEMA_signal_2346), .Z1_t (new_AGEMA_signal_2347), .Z1_f (new_AGEMA_signal_2348) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U939_XOR1_U1 ( .A0_t (StateOut[55]), .A0_f (new_AGEMA_signal_2328), .A1_t (new_AGEMA_signal_2329), .A1_f (new_AGEMA_signal_2330), .B0_t (StateFromChi[47]), .B0_f (new_AGEMA_signal_5127), .B1_t (new_AGEMA_signal_5128), .B1_f (new_AGEMA_signal_5129), .Z0_t (U939_X), .Z0_f (new_AGEMA_signal_5580), .Z1_t (new_AGEMA_signal_5581), .Z1_f (new_AGEMA_signal_5582) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U939_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U939_X), .B0_f (new_AGEMA_signal_5580), .B1_t (new_AGEMA_signal_5581), .B1_f (new_AGEMA_signal_5582), .Z0_t (U939_Y), .Z0_f (new_AGEMA_signal_6187), .Z1_t (new_AGEMA_signal_6188), .Z1_f (new_AGEMA_signal_6189) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U939_XOR2_U1 ( .A0_t (U939_Y), .A0_f (new_AGEMA_signal_6187), .A1_t (new_AGEMA_signal_6188), .A1_f (new_AGEMA_signal_6189), .B0_t (StateOut[55]), .B0_f (new_AGEMA_signal_2328), .B1_t (new_AGEMA_signal_2329), .B1_f (new_AGEMA_signal_2330), .Z0_t (StateOut[47]), .Z0_f (new_AGEMA_signal_3072), .Z1_t (new_AGEMA_signal_3073), .Z1_f (new_AGEMA_signal_3074) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U940_XOR1_U1 ( .A0_t (StateOut[79]), .A0_f (new_AGEMA_signal_2337), .A1_t (new_AGEMA_signal_2338), .A1_f (new_AGEMA_signal_2339), .B0_t (StateFromChi[71]), .B0_f (new_AGEMA_signal_5172), .B1_t (new_AGEMA_signal_5173), .B1_f (new_AGEMA_signal_5174), .Z0_t (U940_X), .Z0_f (new_AGEMA_signal_5583), .Z1_t (new_AGEMA_signal_5584), .Z1_f (new_AGEMA_signal_5585) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U940_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U940_X), .B0_f (new_AGEMA_signal_5583), .B1_t (new_AGEMA_signal_5584), .B1_f (new_AGEMA_signal_5585), .Z0_t (U940_Y), .Z0_f (new_AGEMA_signal_6190), .Z1_t (new_AGEMA_signal_6191), .Z1_f (new_AGEMA_signal_6192) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U940_XOR2_U1 ( .A0_t (U940_Y), .A0_f (new_AGEMA_signal_6190), .A1_t (new_AGEMA_signal_6191), .A1_f (new_AGEMA_signal_6192), .B0_t (StateOut[79]), .B0_f (new_AGEMA_signal_2337), .B1_t (new_AGEMA_signal_2338), .B1_f (new_AGEMA_signal_2339), .Z0_t (StateOut[71]), .Z0_f (new_AGEMA_signal_2340), .Z1_t (new_AGEMA_signal_2341), .Z1_f (new_AGEMA_signal_2342) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U941_XOR1_U1 ( .A0_t (StateOut[87]), .A0_f (new_AGEMA_signal_2475), .A1_t (new_AGEMA_signal_2476), .A1_f (new_AGEMA_signal_2477), .B0_t (StateFromChi[79]), .B0_f (new_AGEMA_signal_5187), .B1_t (new_AGEMA_signal_5188), .B1_f (new_AGEMA_signal_5189), .Z0_t (U941_X), .Z0_f (new_AGEMA_signal_5586), .Z1_t (new_AGEMA_signal_5587), .Z1_f (new_AGEMA_signal_5588) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U941_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U941_X), .B0_f (new_AGEMA_signal_5586), .B1_t (new_AGEMA_signal_5587), .B1_f (new_AGEMA_signal_5588), .Z0_t (U941_Y), .Z0_f (new_AGEMA_signal_6193), .Z1_t (new_AGEMA_signal_6194), .Z1_f (new_AGEMA_signal_6195) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U941_XOR2_U1 ( .A0_t (U941_Y), .A0_f (new_AGEMA_signal_6193), .A1_t (new_AGEMA_signal_6194), .A1_f (new_AGEMA_signal_6195), .B0_t (StateOut[87]), .B0_f (new_AGEMA_signal_2475), .B1_t (new_AGEMA_signal_2476), .B1_f (new_AGEMA_signal_2477), .Z0_t (StateOut[79]), .Z0_f (new_AGEMA_signal_2337), .Z1_t (new_AGEMA_signal_2338), .Z1_f (new_AGEMA_signal_2339) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U942_XOR1_U1 ( .A0_t (StateOut[103]), .A0_f (new_AGEMA_signal_3120), .A1_t (new_AGEMA_signal_3121), .A1_f (new_AGEMA_signal_3122), .B0_t (StateFromChi[95]), .B0_f (new_AGEMA_signal_5145), .B1_t (new_AGEMA_signal_5146), .B1_f (new_AGEMA_signal_5147), .Z0_t (U942_X), .Z0_f (new_AGEMA_signal_5589), .Z1_t (new_AGEMA_signal_5590), .Z1_f (new_AGEMA_signal_5591) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U942_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U942_X), .B0_f (new_AGEMA_signal_5589), .B1_t (new_AGEMA_signal_5590), .B1_f (new_AGEMA_signal_5591), .Z0_t (U942_Y), .Z0_f (new_AGEMA_signal_6196), .Z1_t (new_AGEMA_signal_6197), .Z1_f (new_AGEMA_signal_6198) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U942_XOR2_U1 ( .A0_t (U942_Y), .A0_f (new_AGEMA_signal_6196), .A1_t (new_AGEMA_signal_6197), .A1_f (new_AGEMA_signal_6198), .B0_t (StateOut[103]), .B0_f (new_AGEMA_signal_3120), .B1_t (new_AGEMA_signal_3121), .B1_f (new_AGEMA_signal_3122), .Z0_t (StateOut[95]), .Z0_f (new_AGEMA_signal_2472), .Z1_t (new_AGEMA_signal_2473), .Z1_f (new_AGEMA_signal_2474) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U943_XOR1_U1 ( .A0_t (StateOut[111]), .A0_f (new_AGEMA_signal_2481), .A1_t (new_AGEMA_signal_2482), .A1_f (new_AGEMA_signal_2483), .B0_t (StateFromChi[103]), .B0_f (new_AGEMA_signal_5160), .B1_t (new_AGEMA_signal_5161), .B1_f (new_AGEMA_signal_5162), .Z0_t (U943_X), .Z0_f (new_AGEMA_signal_5592), .Z1_t (new_AGEMA_signal_5593), .Z1_f (new_AGEMA_signal_5594) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U943_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U943_X), .B0_f (new_AGEMA_signal_5592), .B1_t (new_AGEMA_signal_5593), .B1_f (new_AGEMA_signal_5594), .Z0_t (U943_Y), .Z0_f (new_AGEMA_signal_6199), .Z1_t (new_AGEMA_signal_6200), .Z1_f (new_AGEMA_signal_6201) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U943_XOR2_U1 ( .A0_t (U943_Y), .A0_f (new_AGEMA_signal_6199), .A1_t (new_AGEMA_signal_6200), .A1_f (new_AGEMA_signal_6201), .B0_t (StateOut[111]), .B0_f (new_AGEMA_signal_2481), .B1_t (new_AGEMA_signal_2482), .B1_f (new_AGEMA_signal_2483), .Z0_t (StateOut[103]), .Z0_f (new_AGEMA_signal_3120), .Z1_t (new_AGEMA_signal_3121), .Z1_f (new_AGEMA_signal_3122) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U944_XOR1_U1 ( .A0_t (StateOut[135]), .A0_f (new_AGEMA_signal_2148), .A1_t (new_AGEMA_signal_2149), .A1_f (new_AGEMA_signal_2150), .B0_t (StateFromChi[127]), .B0_f (new_AGEMA_signal_5133), .B1_t (new_AGEMA_signal_5134), .B1_f (new_AGEMA_signal_5135), .Z0_t (U944_X), .Z0_f (new_AGEMA_signal_5595), .Z1_t (new_AGEMA_signal_5596), .Z1_f (new_AGEMA_signal_5597) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U944_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U944_X), .B0_f (new_AGEMA_signal_5595), .B1_t (new_AGEMA_signal_5596), .B1_f (new_AGEMA_signal_5597), .Z0_t (U944_Y), .Z0_f (new_AGEMA_signal_6202), .Z1_t (new_AGEMA_signal_6203), .Z1_f (new_AGEMA_signal_6204) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U944_XOR2_U1 ( .A0_t (U944_Y), .A0_f (new_AGEMA_signal_6202), .A1_t (new_AGEMA_signal_6203), .A1_f (new_AGEMA_signal_6204), .B0_t (StateOut[135]), .B0_f (new_AGEMA_signal_2148), .B1_t (new_AGEMA_signal_2149), .B1_f (new_AGEMA_signal_2150), .Z0_t (StateOut[127]), .Z0_f (new_AGEMA_signal_3012), .Z1_t (new_AGEMA_signal_3013), .Z1_f (new_AGEMA_signal_3014) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U945_XOR1_U1 ( .A0_t (StateOut[143]), .A0_f (new_AGEMA_signal_2151), .A1_t (new_AGEMA_signal_2152), .A1_f (new_AGEMA_signal_2153), .B0_t (StateFromChi[135]), .B0_f (new_AGEMA_signal_5148), .B1_t (new_AGEMA_signal_5149), .B1_f (new_AGEMA_signal_5150), .Z0_t (U945_X), .Z0_f (new_AGEMA_signal_5598), .Z1_t (new_AGEMA_signal_5599), .Z1_f (new_AGEMA_signal_5600) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U945_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U945_X), .B0_f (new_AGEMA_signal_5598), .B1_t (new_AGEMA_signal_5599), .B1_f (new_AGEMA_signal_5600), .Z0_t (U945_Y), .Z0_f (new_AGEMA_signal_6205), .Z1_t (new_AGEMA_signal_6206), .Z1_f (new_AGEMA_signal_6207) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U945_XOR2_U1 ( .A0_t (U945_Y), .A0_f (new_AGEMA_signal_6205), .A1_t (new_AGEMA_signal_6206), .A1_f (new_AGEMA_signal_6207), .B0_t (StateOut[143]), .B0_f (new_AGEMA_signal_2151), .B1_t (new_AGEMA_signal_2152), .B1_f (new_AGEMA_signal_2153), .Z0_t (StateOut[135]), .Z0_f (new_AGEMA_signal_2148), .Z1_t (new_AGEMA_signal_2149), .Z1_f (new_AGEMA_signal_2150) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U946_XOR1_U1 ( .A0_t (StateOut[167]), .A0_f (new_AGEMA_signal_2439), .A1_t (new_AGEMA_signal_2440), .A1_f (new_AGEMA_signal_2441), .B0_t (StateFromChi[159]), .B0_f (new_AGEMA_signal_5193), .B1_t (new_AGEMA_signal_5194), .B1_f (new_AGEMA_signal_5195), .Z0_t (U946_X), .Z0_f (new_AGEMA_signal_5601), .Z1_t (new_AGEMA_signal_5602), .Z1_f (new_AGEMA_signal_5603) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U946_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U946_X), .B0_f (new_AGEMA_signal_5601), .B1_t (new_AGEMA_signal_5602), .B1_f (new_AGEMA_signal_5603), .Z0_t (U946_Y), .Z0_f (new_AGEMA_signal_6208), .Z1_t (new_AGEMA_signal_6209), .Z1_f (new_AGEMA_signal_6210) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U946_XOR2_U1 ( .A0_t (U946_Y), .A0_f (new_AGEMA_signal_6208), .A1_t (new_AGEMA_signal_6209), .A1_f (new_AGEMA_signal_6210), .B0_t (StateOut[167]), .B0_f (new_AGEMA_signal_2439), .B1_t (new_AGEMA_signal_2440), .B1_f (new_AGEMA_signal_2441), .Z0_t (StateOut[159]), .Z0_f (new_AGEMA_signal_2157), .Z1_t (new_AGEMA_signal_2158), .Z1_f (new_AGEMA_signal_2159) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U947_XOR1_U1 ( .A0_t (StateOut[191]), .A0_f (new_AGEMA_signal_2445), .A1_t (new_AGEMA_signal_2446), .A1_f (new_AGEMA_signal_2447), .B0_t (StateFromChi[183]), .B0_f (new_AGEMA_signal_5166), .B1_t (new_AGEMA_signal_5167), .B1_f (new_AGEMA_signal_5168), .Z0_t (U947_X), .Z0_f (new_AGEMA_signal_5604), .Z1_t (new_AGEMA_signal_5605), .Z1_f (new_AGEMA_signal_5606) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U947_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U947_X), .B0_f (new_AGEMA_signal_5604), .B1_t (new_AGEMA_signal_5605), .B1_f (new_AGEMA_signal_5606), .Z0_t (U947_Y), .Z0_f (new_AGEMA_signal_6211), .Z1_t (new_AGEMA_signal_6212), .Z1_f (new_AGEMA_signal_6213) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U947_XOR2_U1 ( .A0_t (U947_Y), .A0_f (new_AGEMA_signal_6211), .A1_t (new_AGEMA_signal_6212), .A1_f (new_AGEMA_signal_6213), .B0_t (StateOut[191]), .B0_f (new_AGEMA_signal_2445), .B1_t (new_AGEMA_signal_2446), .B1_f (new_AGEMA_signal_2447), .Z0_t (StateOut[183]), .Z0_f (new_AGEMA_signal_3108), .Z1_t (new_AGEMA_signal_3109), .Z1_f (new_AGEMA_signal_3110) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U948_XOR1_U1 ( .A0_t (StateOut[199]), .A0_f (new_AGEMA_signal_2448), .A1_t (new_AGEMA_signal_2449), .A1_f (new_AGEMA_signal_2450), .B0_t (StateFromChi[191]), .B0_f (new_AGEMA_signal_5181), .B1_t (new_AGEMA_signal_5182), .B1_f (new_AGEMA_signal_5183), .Z0_t (U948_X), .Z0_f (new_AGEMA_signal_5607), .Z1_t (new_AGEMA_signal_5608), .Z1_f (new_AGEMA_signal_5609) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U948_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U948_X), .B0_f (new_AGEMA_signal_5607), .B1_t (new_AGEMA_signal_5608), .B1_f (new_AGEMA_signal_5609), .Z0_t (U948_Y), .Z0_f (new_AGEMA_signal_6214), .Z1_t (new_AGEMA_signal_6215), .Z1_f (new_AGEMA_signal_6216) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U948_XOR2_U1 ( .A0_t (U948_Y), .A0_f (new_AGEMA_signal_6214), .A1_t (new_AGEMA_signal_6215), .A1_f (new_AGEMA_signal_6216), .B0_t (StateOut[199]), .B0_f (new_AGEMA_signal_2448), .B1_t (new_AGEMA_signal_2449), .B1_f (new_AGEMA_signal_2450), .Z0_t (StateOut[191]), .Z0_f (new_AGEMA_signal_2445), .Z1_t (new_AGEMA_signal_2446), .Z1_f (new_AGEMA_signal_2447) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U949_XOR1_U1 ( .A0_t (StateOut[22]), .A0_f (new_AGEMA_signal_2133), .A1_t (new_AGEMA_signal_2134), .A1_f (new_AGEMA_signal_2135), .B0_t (StateFromChi[14]), .B0_f (new_AGEMA_signal_5064), .B1_t (new_AGEMA_signal_5065), .B1_f (new_AGEMA_signal_5066), .Z0_t (U949_X), .Z0_f (new_AGEMA_signal_5610), .Z1_t (new_AGEMA_signal_5611), .Z1_f (new_AGEMA_signal_5612) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U949_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U949_X), .B0_f (new_AGEMA_signal_5610), .B1_t (new_AGEMA_signal_5611), .B1_f (new_AGEMA_signal_5612), .Z0_t (U949_Y), .Z0_f (new_AGEMA_signal_6217), .Z1_t (new_AGEMA_signal_6218), .Z1_f (new_AGEMA_signal_6219) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U949_XOR2_U1 ( .A0_t (U949_Y), .A0_f (new_AGEMA_signal_6217), .A1_t (new_AGEMA_signal_6218), .A1_f (new_AGEMA_signal_6219), .B0_t (StateOut[22]), .B0_f (new_AGEMA_signal_2133), .B1_t (new_AGEMA_signal_2134), .B1_f (new_AGEMA_signal_2135), .Z0_t (StateOut[14]), .Z0_f (new_AGEMA_signal_2130), .Z1_t (new_AGEMA_signal_2131), .Z1_f (new_AGEMA_signal_2132) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U950_XOR1_U1 ( .A0_t (StateOut[54]), .A0_f (new_AGEMA_signal_2454), .A1_t (new_AGEMA_signal_2455), .A1_f (new_AGEMA_signal_2456), .B0_t (StateFromChi[46]), .B0_f (new_AGEMA_signal_5052), .B1_t (new_AGEMA_signal_5053), .B1_f (new_AGEMA_signal_5054), .Z0_t (U950_X), .Z0_f (new_AGEMA_signal_5613), .Z1_t (new_AGEMA_signal_5614), .Z1_f (new_AGEMA_signal_5615) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U950_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U950_X), .B0_f (new_AGEMA_signal_5613), .B1_t (new_AGEMA_signal_5614), .B1_f (new_AGEMA_signal_5615), .Z0_t (U950_Y), .Z0_f (new_AGEMA_signal_6220), .Z1_t (new_AGEMA_signal_6221), .Z1_f (new_AGEMA_signal_6222) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U950_XOR2_U1 ( .A0_t (U950_Y), .A0_f (new_AGEMA_signal_6220), .A1_t (new_AGEMA_signal_6221), .A1_f (new_AGEMA_signal_6222), .B0_t (StateOut[54]), .B0_f (new_AGEMA_signal_2454), .B1_t (new_AGEMA_signal_2455), .B1_f (new_AGEMA_signal_2456), .Z0_t (StateOut[46]), .Z0_f (new_AGEMA_signal_2457), .Z1_t (new_AGEMA_signal_2458), .Z1_f (new_AGEMA_signal_2459) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U951_XOR1_U1 ( .A0_t (StateOut[78]), .A0_f (new_AGEMA_signal_2466), .A1_t (new_AGEMA_signal_2467), .A1_f (new_AGEMA_signal_2468), .B0_t (StateFromChi[70]), .B0_f (new_AGEMA_signal_5097), .B1_t (new_AGEMA_signal_5098), .B1_f (new_AGEMA_signal_5099), .Z0_t (U951_X), .Z0_f (new_AGEMA_signal_5616), .Z1_t (new_AGEMA_signal_5617), .Z1_f (new_AGEMA_signal_5618) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U951_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U951_X), .B0_f (new_AGEMA_signal_5616), .B1_t (new_AGEMA_signal_5617), .B1_f (new_AGEMA_signal_5618), .Z0_t (U951_Y), .Z0_f (new_AGEMA_signal_6223), .Z1_t (new_AGEMA_signal_6224), .Z1_f (new_AGEMA_signal_6225) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U951_XOR2_U1 ( .A0_t (U951_Y), .A0_f (new_AGEMA_signal_6223), .A1_t (new_AGEMA_signal_6224), .A1_f (new_AGEMA_signal_6225), .B0_t (StateOut[78]), .B0_f (new_AGEMA_signal_2466), .B1_t (new_AGEMA_signal_2467), .B1_f (new_AGEMA_signal_2468), .Z0_t (StateOut[70]), .Z0_f (new_AGEMA_signal_2463), .Z1_t (new_AGEMA_signal_2464), .Z1_f (new_AGEMA_signal_2465) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U952_XOR1_U1 ( .A0_t (StateOut[86]), .A0_f (new_AGEMA_signal_2691), .A1_t (new_AGEMA_signal_2692), .A1_f (new_AGEMA_signal_2693), .B0_t (StateFromChi[78]), .B0_f (new_AGEMA_signal_5112), .B1_t (new_AGEMA_signal_5113), .B1_f (new_AGEMA_signal_5114), .Z0_t (U952_X), .Z0_f (new_AGEMA_signal_5619), .Z1_t (new_AGEMA_signal_5620), .Z1_f (new_AGEMA_signal_5621) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U952_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U952_X), .B0_f (new_AGEMA_signal_5619), .B1_t (new_AGEMA_signal_5620), .B1_f (new_AGEMA_signal_5621), .Z0_t (U952_Y), .Z0_f (new_AGEMA_signal_6226), .Z1_t (new_AGEMA_signal_6227), .Z1_f (new_AGEMA_signal_6228) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U952_XOR2_U1 ( .A0_t (U952_Y), .A0_f (new_AGEMA_signal_6226), .A1_t (new_AGEMA_signal_6227), .A1_f (new_AGEMA_signal_6228), .B0_t (StateOut[86]), .B0_f (new_AGEMA_signal_2691), .B1_t (new_AGEMA_signal_2692), .B1_f (new_AGEMA_signal_2693), .Z0_t (StateOut[78]), .Z0_f (new_AGEMA_signal_2466), .Z1_t (new_AGEMA_signal_2467), .Z1_f (new_AGEMA_signal_2468) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U953_XOR1_U1 ( .A0_t (StateOut[102]), .A0_f (new_AGEMA_signal_2700), .A1_t (new_AGEMA_signal_2701), .A1_f (new_AGEMA_signal_2702), .B0_t (StateFromChi[94]), .B0_f (new_AGEMA_signal_5070), .B1_t (new_AGEMA_signal_5071), .B1_f (new_AGEMA_signal_5072), .Z0_t (U953_X), .Z0_f (new_AGEMA_signal_5622), .Z1_t (new_AGEMA_signal_5623), .Z1_f (new_AGEMA_signal_5624) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U953_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U953_X), .B0_f (new_AGEMA_signal_5622), .B1_t (new_AGEMA_signal_5623), .B1_f (new_AGEMA_signal_5624), .Z0_t (U953_Y), .Z0_f (new_AGEMA_signal_6229), .Z1_t (new_AGEMA_signal_6230), .Z1_f (new_AGEMA_signal_6231) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U953_XOR2_U1 ( .A0_t (U953_Y), .A0_f (new_AGEMA_signal_6229), .A1_t (new_AGEMA_signal_6230), .A1_f (new_AGEMA_signal_6231), .B0_t (StateOut[102]), .B0_f (new_AGEMA_signal_2700), .B1_t (new_AGEMA_signal_2701), .B1_f (new_AGEMA_signal_2702), .Z0_t (StateOut[94]), .Z0_f (new_AGEMA_signal_2688), .Z1_t (new_AGEMA_signal_2689), .Z1_f (new_AGEMA_signal_2690) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U954_XOR1_U1 ( .A0_t (StateOut[110]), .A0_f (new_AGEMA_signal_3192), .A1_t (new_AGEMA_signal_3193), .A1_f (new_AGEMA_signal_3194), .B0_t (StateFromChi[102]), .B0_f (new_AGEMA_signal_5085), .B1_t (new_AGEMA_signal_5086), .B1_f (new_AGEMA_signal_5087), .Z0_t (U954_X), .Z0_f (new_AGEMA_signal_5625), .Z1_t (new_AGEMA_signal_5626), .Z1_f (new_AGEMA_signal_5627) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U954_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U954_X), .B0_f (new_AGEMA_signal_5625), .B1_t (new_AGEMA_signal_5626), .B1_f (new_AGEMA_signal_5627), .Z0_t (U954_Y), .Z0_f (new_AGEMA_signal_6232), .Z1_t (new_AGEMA_signal_6233), .Z1_f (new_AGEMA_signal_6234) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U954_XOR2_U1 ( .A0_t (U954_Y), .A0_f (new_AGEMA_signal_6232), .A1_t (new_AGEMA_signal_6233), .A1_f (new_AGEMA_signal_6234), .B0_t (StateOut[110]), .B0_f (new_AGEMA_signal_3192), .B1_t (new_AGEMA_signal_3193), .B1_f (new_AGEMA_signal_3194), .Z0_t (StateOut[102]), .Z0_f (new_AGEMA_signal_2700), .Z1_t (new_AGEMA_signal_2701), .Z1_f (new_AGEMA_signal_2702) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U955_XOR1_U1 ( .A0_t (StateOut[134]), .A0_f (new_AGEMA_signal_2166), .A1_t (new_AGEMA_signal_2167), .A1_f (new_AGEMA_signal_2168), .B0_t (StateFromChi[126]), .B0_f (new_AGEMA_signal_5058), .B1_t (new_AGEMA_signal_5059), .B1_f (new_AGEMA_signal_5060), .Z0_t (U955_X), .Z0_f (new_AGEMA_signal_5628), .Z1_t (new_AGEMA_signal_5629), .Z1_f (new_AGEMA_signal_5630) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U955_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U955_X), .B0_f (new_AGEMA_signal_5628), .B1_t (new_AGEMA_signal_5629), .B1_f (new_AGEMA_signal_5630), .Z0_t (U955_Y), .Z0_f (new_AGEMA_signal_6235), .Z1_t (new_AGEMA_signal_6236), .Z1_f (new_AGEMA_signal_6237) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U955_XOR2_U1 ( .A0_t (U955_Y), .A0_f (new_AGEMA_signal_6235), .A1_t (new_AGEMA_signal_6236), .A1_f (new_AGEMA_signal_6237), .B0_t (StateOut[134]), .B0_f (new_AGEMA_signal_2166), .B1_t (new_AGEMA_signal_2167), .B1_f (new_AGEMA_signal_2168), .Z0_t (StateOut[126]), .Z0_f (new_AGEMA_signal_3018), .Z1_t (new_AGEMA_signal_3019), .Z1_f (new_AGEMA_signal_3020) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U956_XOR1_U1 ( .A0_t (StateOut[142]), .A0_f (new_AGEMA_signal_2169), .A1_t (new_AGEMA_signal_2170), .A1_f (new_AGEMA_signal_2171), .B0_t (StateFromChi[134]), .B0_f (new_AGEMA_signal_5073), .B1_t (new_AGEMA_signal_5074), .B1_f (new_AGEMA_signal_5075), .Z0_t (U956_X), .Z0_f (new_AGEMA_signal_5631), .Z1_t (new_AGEMA_signal_5632), .Z1_f (new_AGEMA_signal_5633) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U956_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U956_X), .B0_f (new_AGEMA_signal_5631), .B1_t (new_AGEMA_signal_5632), .B1_f (new_AGEMA_signal_5633), .Z0_t (U956_Y), .Z0_f (new_AGEMA_signal_6238), .Z1_t (new_AGEMA_signal_6239), .Z1_f (new_AGEMA_signal_6240) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U956_XOR2_U1 ( .A0_t (U956_Y), .A0_f (new_AGEMA_signal_6238), .A1_t (new_AGEMA_signal_6239), .A1_f (new_AGEMA_signal_6240), .B0_t (StateOut[142]), .B0_f (new_AGEMA_signal_2169), .B1_t (new_AGEMA_signal_2170), .B1_f (new_AGEMA_signal_2171), .Z0_t (StateOut[134]), .Z0_f (new_AGEMA_signal_2166), .Z1_t (new_AGEMA_signal_2167), .Z1_f (new_AGEMA_signal_2168) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U957_XOR1_U1 ( .A0_t (StateOut[166]), .A0_f (new_AGEMA_signal_2493), .A1_t (new_AGEMA_signal_2494), .A1_f (new_AGEMA_signal_2495), .B0_t (StateFromChi[158]), .B0_f (new_AGEMA_signal_5118), .B1_t (new_AGEMA_signal_5119), .B1_f (new_AGEMA_signal_5120), .Z0_t (U957_X), .Z0_f (new_AGEMA_signal_5634), .Z1_t (new_AGEMA_signal_5635), .Z1_f (new_AGEMA_signal_5636) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U957_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U957_X), .B0_f (new_AGEMA_signal_5634), .B1_t (new_AGEMA_signal_5635), .B1_f (new_AGEMA_signal_5636), .Z0_t (U957_Y), .Z0_f (new_AGEMA_signal_6241), .Z1_t (new_AGEMA_signal_6242), .Z1_f (new_AGEMA_signal_6243) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U957_XOR2_U1 ( .A0_t (U957_Y), .A0_f (new_AGEMA_signal_6241), .A1_t (new_AGEMA_signal_6242), .A1_f (new_AGEMA_signal_6243), .B0_t (StateOut[166]), .B0_f (new_AGEMA_signal_2493), .B1_t (new_AGEMA_signal_2494), .B1_f (new_AGEMA_signal_2495), .Z0_t (StateOut[158]), .Z0_f (new_AGEMA_signal_2175), .Z1_t (new_AGEMA_signal_2176), .Z1_f (new_AGEMA_signal_2177) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U958_XOR1_U1 ( .A0_t (StateOut[190]), .A0_f (new_AGEMA_signal_2499), .A1_t (new_AGEMA_signal_2500), .A1_f (new_AGEMA_signal_2501), .B0_t (StateFromChi[182]), .B0_f (new_AGEMA_signal_5091), .B1_t (new_AGEMA_signal_5092), .B1_f (new_AGEMA_signal_5093), .Z0_t (U958_X), .Z0_f (new_AGEMA_signal_5637), .Z1_t (new_AGEMA_signal_5638), .Z1_f (new_AGEMA_signal_5639) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U958_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U958_X), .B0_f (new_AGEMA_signal_5637), .B1_t (new_AGEMA_signal_5638), .B1_f (new_AGEMA_signal_5639), .Z0_t (U958_Y), .Z0_f (new_AGEMA_signal_6244), .Z1_t (new_AGEMA_signal_6245), .Z1_f (new_AGEMA_signal_6246) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U958_XOR2_U1 ( .A0_t (U958_Y), .A0_f (new_AGEMA_signal_6244), .A1_t (new_AGEMA_signal_6245), .A1_f (new_AGEMA_signal_6246), .B0_t (StateOut[190]), .B0_f (new_AGEMA_signal_2499), .B1_t (new_AGEMA_signal_2500), .B1_f (new_AGEMA_signal_2501), .Z0_t (StateOut[182]), .Z0_f (new_AGEMA_signal_3126), .Z1_t (new_AGEMA_signal_3127), .Z1_f (new_AGEMA_signal_3128) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U959_XOR1_U1 ( .A0_t (StateOut[198]), .A0_f (new_AGEMA_signal_2502), .A1_t (new_AGEMA_signal_2503), .A1_f (new_AGEMA_signal_2504), .B0_t (StateFromChi[190]), .B0_f (new_AGEMA_signal_5106), .B1_t (new_AGEMA_signal_5107), .B1_f (new_AGEMA_signal_5108), .Z0_t (U959_X), .Z0_f (new_AGEMA_signal_5640), .Z1_t (new_AGEMA_signal_5641), .Z1_f (new_AGEMA_signal_5642) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U959_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U959_X), .B0_f (new_AGEMA_signal_5640), .B1_t (new_AGEMA_signal_5641), .B1_f (new_AGEMA_signal_5642), .Z0_t (U959_Y), .Z0_f (new_AGEMA_signal_6247), .Z1_t (new_AGEMA_signal_6248), .Z1_f (new_AGEMA_signal_6249) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U959_XOR2_U1 ( .A0_t (U959_Y), .A0_f (new_AGEMA_signal_6247), .A1_t (new_AGEMA_signal_6248), .A1_f (new_AGEMA_signal_6249), .B0_t (StateOut[198]), .B0_f (new_AGEMA_signal_2502), .B1_t (new_AGEMA_signal_2503), .B1_f (new_AGEMA_signal_2504), .Z0_t (StateOut[190]), .Z0_f (new_AGEMA_signal_2499), .Z1_t (new_AGEMA_signal_2500), .Z1_f (new_AGEMA_signal_2501) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U960_XOR1_U1 ( .A0_t (StateOut[21]), .A0_f (new_AGEMA_signal_2646), .A1_t (new_AGEMA_signal_2647), .A1_f (new_AGEMA_signal_2648), .B0_t (StateFromChi[13]), .B0_f (new_AGEMA_signal_4989), .B1_t (new_AGEMA_signal_4990), .B1_f (new_AGEMA_signal_4991), .Z0_t (U960_X), .Z0_f (new_AGEMA_signal_5643), .Z1_t (new_AGEMA_signal_5644), .Z1_f (new_AGEMA_signal_5645) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U960_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U960_X), .B0_f (new_AGEMA_signal_5643), .B1_t (new_AGEMA_signal_5644), .B1_f (new_AGEMA_signal_5645), .Z0_t (U960_Y), .Z0_f (new_AGEMA_signal_6250), .Z1_t (new_AGEMA_signal_6251), .Z1_f (new_AGEMA_signal_6252) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U960_XOR2_U1 ( .A0_t (U960_Y), .A0_f (new_AGEMA_signal_6250), .A1_t (new_AGEMA_signal_6251), .A1_f (new_AGEMA_signal_6252), .B0_t (StateOut[21]), .B0_f (new_AGEMA_signal_2646), .B1_t (new_AGEMA_signal_2647), .B1_f (new_AGEMA_signal_2648), .Z0_t (StateOut[13]), .Z0_f (new_AGEMA_signal_2634), .Z1_t (new_AGEMA_signal_2635), .Z1_f (new_AGEMA_signal_2636) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U961_XOR1_U1 ( .A0_t (StateOut[53]), .A0_f (new_AGEMA_signal_2508), .A1_t (new_AGEMA_signal_2509), .A1_f (new_AGEMA_signal_2510), .B0_t (StateFromChi[45]), .B0_f (new_AGEMA_signal_4977), .B1_t (new_AGEMA_signal_4978), .B1_f (new_AGEMA_signal_4979), .Z0_t (U961_X), .Z0_f (new_AGEMA_signal_5646), .Z1_t (new_AGEMA_signal_5647), .Z1_f (new_AGEMA_signal_5648) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U961_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U961_X), .B0_f (new_AGEMA_signal_5646), .B1_t (new_AGEMA_signal_5647), .B1_f (new_AGEMA_signal_5648), .Z0_t (U961_Y), .Z0_f (new_AGEMA_signal_6253), .Z1_t (new_AGEMA_signal_6254), .Z1_f (new_AGEMA_signal_6255) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U961_XOR2_U1 ( .A0_t (U961_Y), .A0_f (new_AGEMA_signal_6253), .A1_t (new_AGEMA_signal_6254), .A1_f (new_AGEMA_signal_6255), .B0_t (StateOut[53]), .B0_f (new_AGEMA_signal_2508), .B1_t (new_AGEMA_signal_2509), .B1_f (new_AGEMA_signal_2510), .Z0_t (StateOut[45]), .Z0_f (new_AGEMA_signal_3132), .Z1_t (new_AGEMA_signal_3133), .Z1_f (new_AGEMA_signal_3134) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U962_XOR1_U1 ( .A0_t (StateOut[85]), .A0_f (new_AGEMA_signal_2727), .A1_t (new_AGEMA_signal_2728), .A1_f (new_AGEMA_signal_2729), .B0_t (StateFromChi[77]), .B0_f (new_AGEMA_signal_5037), .B1_t (new_AGEMA_signal_5038), .B1_f (new_AGEMA_signal_5039), .Z0_t (U962_X), .Z0_f (new_AGEMA_signal_5649), .Z1_t (new_AGEMA_signal_5650), .Z1_f (new_AGEMA_signal_5651) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U962_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U962_X), .B0_f (new_AGEMA_signal_5649), .B1_t (new_AGEMA_signal_5650), .B1_f (new_AGEMA_signal_5651), .Z0_t (U962_Y), .Z0_f (new_AGEMA_signal_6256), .Z1_t (new_AGEMA_signal_6257), .Z1_f (new_AGEMA_signal_6258) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U962_XOR2_U1 ( .A0_t (U962_Y), .A0_f (new_AGEMA_signal_6256), .A1_t (new_AGEMA_signal_6257), .A1_f (new_AGEMA_signal_6258), .B0_t (StateOut[85]), .B0_f (new_AGEMA_signal_2727), .B1_t (new_AGEMA_signal_2728), .B1_f (new_AGEMA_signal_2729), .Z0_t (StateOut[77]), .Z0_f (new_AGEMA_signal_2517), .Z1_t (new_AGEMA_signal_2518), .Z1_f (new_AGEMA_signal_2519) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U963_XOR1_U1 ( .A0_t (StateOut[101]), .A0_f (new_AGEMA_signal_2736), .A1_t (new_AGEMA_signal_2737), .A1_f (new_AGEMA_signal_2738), .B0_t (StateFromChi[93]), .B0_f (new_AGEMA_signal_4995), .B1_t (new_AGEMA_signal_4996), .B1_f (new_AGEMA_signal_4997), .Z0_t (U963_X), .Z0_f (new_AGEMA_signal_5652), .Z1_t (new_AGEMA_signal_5653), .Z1_f (new_AGEMA_signal_5654) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U963_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U963_X), .B0_f (new_AGEMA_signal_5652), .B1_t (new_AGEMA_signal_5653), .B1_f (new_AGEMA_signal_5654), .Z0_t (U963_Y), .Z0_f (new_AGEMA_signal_6259), .Z1_t (new_AGEMA_signal_6260), .Z1_f (new_AGEMA_signal_6261) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U963_XOR2_U1 ( .A0_t (U963_Y), .A0_f (new_AGEMA_signal_6259), .A1_t (new_AGEMA_signal_6260), .A1_f (new_AGEMA_signal_6261), .B0_t (StateOut[101]), .B0_f (new_AGEMA_signal_2736), .B1_t (new_AGEMA_signal_2737), .B1_f (new_AGEMA_signal_2738), .Z0_t (StateOut[93]), .Z0_f (new_AGEMA_signal_2724), .Z1_t (new_AGEMA_signal_2725), .Z1_f (new_AGEMA_signal_2726) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U964_XOR1_U1 ( .A0_t (StateOut[109]), .A0_f (new_AGEMA_signal_3204), .A1_t (new_AGEMA_signal_3205), .A1_f (new_AGEMA_signal_3206), .B0_t (StateFromChi[101]), .B0_f (new_AGEMA_signal_5010), .B1_t (new_AGEMA_signal_5011), .B1_f (new_AGEMA_signal_5012), .Z0_t (U964_X), .Z0_f (new_AGEMA_signal_5655), .Z1_t (new_AGEMA_signal_5656), .Z1_f (new_AGEMA_signal_5657) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U964_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U964_X), .B0_f (new_AGEMA_signal_5655), .B1_t (new_AGEMA_signal_5656), .B1_f (new_AGEMA_signal_5657), .Z0_t (U964_Y), .Z0_f (new_AGEMA_signal_6262), .Z1_t (new_AGEMA_signal_6263), .Z1_f (new_AGEMA_signal_6264) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U964_XOR2_U1 ( .A0_t (U964_Y), .A0_f (new_AGEMA_signal_6262), .A1_t (new_AGEMA_signal_6263), .A1_f (new_AGEMA_signal_6264), .B0_t (StateOut[109]), .B0_f (new_AGEMA_signal_3204), .B1_t (new_AGEMA_signal_3205), .B1_f (new_AGEMA_signal_3206), .Z0_t (StateOut[101]), .Z0_f (new_AGEMA_signal_2736), .Z1_t (new_AGEMA_signal_2737), .Z1_f (new_AGEMA_signal_2738) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U965_XOR1_U1 ( .A0_t (StateOut[117]), .A0_f (new_AGEMA_signal_2733), .A1_t (new_AGEMA_signal_2734), .A1_f (new_AGEMA_signal_2735), .B0_t (StateFromChi[109]), .B0_f (new_AGEMA_signal_5025), .B1_t (new_AGEMA_signal_5026), .B1_f (new_AGEMA_signal_5027), .Z0_t (U965_X), .Z0_f (new_AGEMA_signal_5658), .Z1_t (new_AGEMA_signal_5659), .Z1_f (new_AGEMA_signal_5660) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U965_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U965_X), .B0_f (new_AGEMA_signal_5658), .B1_t (new_AGEMA_signal_5659), .B1_f (new_AGEMA_signal_5660), .Z0_t (U965_Y), .Z0_f (new_AGEMA_signal_6265), .Z1_t (new_AGEMA_signal_6266), .Z1_f (new_AGEMA_signal_6267) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U965_XOR2_U1 ( .A0_t (U965_Y), .A0_f (new_AGEMA_signal_6265), .A1_t (new_AGEMA_signal_6266), .A1_f (new_AGEMA_signal_6267), .B0_t (StateOut[117]), .B0_f (new_AGEMA_signal_2733), .B1_t (new_AGEMA_signal_2734), .B1_f (new_AGEMA_signal_2735), .Z0_t (StateOut[109]), .Z0_f (new_AGEMA_signal_3204), .Z1_t (new_AGEMA_signal_3205), .Z1_f (new_AGEMA_signal_3206) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U966_XOR1_U1 ( .A0_t (StateOut[133]), .A0_f (new_AGEMA_signal_2544), .A1_t (new_AGEMA_signal_2545), .A1_f (new_AGEMA_signal_2546), .B0_t (StateFromChi[125]), .B0_f (new_AGEMA_signal_4983), .B1_t (new_AGEMA_signal_4984), .B1_f (new_AGEMA_signal_4985), .Z0_t (U966_X), .Z0_f (new_AGEMA_signal_5661), .Z1_t (new_AGEMA_signal_5662), .Z1_f (new_AGEMA_signal_5663) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U966_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U966_X), .B0_f (new_AGEMA_signal_5661), .B1_t (new_AGEMA_signal_5662), .B1_f (new_AGEMA_signal_5663), .Z0_t (U966_Y), .Z0_f (new_AGEMA_signal_6268), .Z1_t (new_AGEMA_signal_6269), .Z1_f (new_AGEMA_signal_6270) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U966_XOR2_U1 ( .A0_t (U966_Y), .A0_f (new_AGEMA_signal_6268), .A1_t (new_AGEMA_signal_6269), .A1_f (new_AGEMA_signal_6270), .B0_t (StateOut[133]), .B0_f (new_AGEMA_signal_2544), .B1_t (new_AGEMA_signal_2545), .B1_f (new_AGEMA_signal_2546), .Z0_t (StateOut[125]), .Z0_f (new_AGEMA_signal_3144), .Z1_t (new_AGEMA_signal_3145), .Z1_f (new_AGEMA_signal_3146) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U967_XOR1_U1 ( .A0_t (StateOut[165]), .A0_f (new_AGEMA_signal_2673), .A1_t (new_AGEMA_signal_2674), .A1_f (new_AGEMA_signal_2675), .B0_t (StateFromChi[157]), .B0_f (new_AGEMA_signal_5043), .B1_t (new_AGEMA_signal_5044), .B1_f (new_AGEMA_signal_5045), .Z0_t (U967_X), .Z0_f (new_AGEMA_signal_5664), .Z1_t (new_AGEMA_signal_5665), .Z1_f (new_AGEMA_signal_5666) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U967_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U967_X), .B0_f (new_AGEMA_signal_5664), .B1_t (new_AGEMA_signal_5665), .B1_f (new_AGEMA_signal_5666), .Z0_t (U967_Y), .Z0_f (new_AGEMA_signal_6271), .Z1_t (new_AGEMA_signal_6272), .Z1_f (new_AGEMA_signal_6273) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U967_XOR2_U1 ( .A0_t (U967_Y), .A0_f (new_AGEMA_signal_6271), .A1_t (new_AGEMA_signal_6272), .A1_f (new_AGEMA_signal_6273), .B0_t (StateOut[165]), .B0_f (new_AGEMA_signal_2673), .B1_t (new_AGEMA_signal_2674), .B1_f (new_AGEMA_signal_2675), .Z0_t (StateOut[157]), .Z0_f (new_AGEMA_signal_2553), .Z1_t (new_AGEMA_signal_2554), .Z1_f (new_AGEMA_signal_2555) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U968_XOR1_U1 ( .A0_t (StateOut[189]), .A0_f (new_AGEMA_signal_2679), .A1_t (new_AGEMA_signal_2680), .A1_f (new_AGEMA_signal_2681), .B0_t (StateFromChi[181]), .B0_f (new_AGEMA_signal_5016), .B1_t (new_AGEMA_signal_5017), .B1_f (new_AGEMA_signal_5018), .Z0_t (U968_X), .Z0_f (new_AGEMA_signal_5667), .Z1_t (new_AGEMA_signal_5668), .Z1_f (new_AGEMA_signal_5669) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U968_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U968_X), .B0_f (new_AGEMA_signal_5667), .B1_t (new_AGEMA_signal_5668), .B1_f (new_AGEMA_signal_5669), .Z0_t (U968_Y), .Z0_f (new_AGEMA_signal_6274), .Z1_t (new_AGEMA_signal_6275), .Z1_f (new_AGEMA_signal_6276) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U968_XOR2_U1 ( .A0_t (U968_Y), .A0_f (new_AGEMA_signal_6274), .A1_t (new_AGEMA_signal_6275), .A1_f (new_AGEMA_signal_6276), .B0_t (StateOut[189]), .B0_f (new_AGEMA_signal_2679), .B1_t (new_AGEMA_signal_2680), .B1_f (new_AGEMA_signal_2681), .Z0_t (StateOut[181]), .Z0_f (new_AGEMA_signal_3186), .Z1_t (new_AGEMA_signal_3187), .Z1_f (new_AGEMA_signal_3188) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U969_XOR1_U1 ( .A0_t (StateOut[197]), .A0_f (new_AGEMA_signal_2682), .A1_t (new_AGEMA_signal_2683), .A1_f (new_AGEMA_signal_2684), .B0_t (StateFromChi[189]), .B0_f (new_AGEMA_signal_5031), .B1_t (new_AGEMA_signal_5032), .B1_f (new_AGEMA_signal_5033), .Z0_t (U969_X), .Z0_f (new_AGEMA_signal_5670), .Z1_t (new_AGEMA_signal_5671), .Z1_f (new_AGEMA_signal_5672) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U969_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U969_X), .B0_f (new_AGEMA_signal_5670), .B1_t (new_AGEMA_signal_5671), .B1_f (new_AGEMA_signal_5672), .Z0_t (U969_Y), .Z0_f (new_AGEMA_signal_6277), .Z1_t (new_AGEMA_signal_6278), .Z1_f (new_AGEMA_signal_6279) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U969_XOR2_U1 ( .A0_t (U969_Y), .A0_f (new_AGEMA_signal_6277), .A1_t (new_AGEMA_signal_6278), .A1_f (new_AGEMA_signal_6279), .B0_t (StateOut[197]), .B0_f (new_AGEMA_signal_2682), .B1_t (new_AGEMA_signal_2683), .B1_f (new_AGEMA_signal_2684), .Z0_t (StateOut[189]), .Z0_f (new_AGEMA_signal_2679), .Z1_t (new_AGEMA_signal_2680), .Z1_f (new_AGEMA_signal_2681) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U970_XOR1_U1 ( .A0_t (InData_s0_t[5]), .A0_f (InData_s0_f[5]), .A1_t (InData_s1_t[5]), .A1_f (InData_s1_f[5]), .B0_t (StateFromChi[197]), .B0_f (new_AGEMA_signal_5046), .B1_t (new_AGEMA_signal_5047), .B1_f (new_AGEMA_signal_5048), .Z0_t (U970_X), .Z0_f (new_AGEMA_signal_5676), .Z1_t (new_AGEMA_signal_5677), .Z1_f (new_AGEMA_signal_5678) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U970_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U970_X), .B0_f (new_AGEMA_signal_5676), .B1_t (new_AGEMA_signal_5677), .B1_f (new_AGEMA_signal_5678), .Z0_t (U970_Y), .Z0_f (new_AGEMA_signal_6280), .Z1_t (new_AGEMA_signal_6281), .Z1_f (new_AGEMA_signal_6282) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U970_XOR2_U1 ( .A0_t (U970_Y), .A0_f (new_AGEMA_signal_6280), .A1_t (new_AGEMA_signal_6281), .A1_f (new_AGEMA_signal_6282), .B0_t (InData_s0_t[5]), .B0_f (InData_s0_f[5]), .B1_t (InData_s1_t[5]), .B1_f (InData_s1_f[5]), .Z0_t (StateOut[197]), .Z0_f (new_AGEMA_signal_2682), .Z1_t (new_AGEMA_signal_2683), .Z1_f (new_AGEMA_signal_2684) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U971_XOR1_U1 ( .A0_t (StateOut[20]), .A0_f (new_AGEMA_signal_2565), .A1_t (new_AGEMA_signal_2566), .A1_f (new_AGEMA_signal_2567), .B0_t (StateFromChi[12]), .B0_f (new_AGEMA_signal_4914), .B1_t (new_AGEMA_signal_4915), .B1_f (new_AGEMA_signal_4916), .Z0_t (U971_X), .Z0_f (new_AGEMA_signal_5679), .Z1_t (new_AGEMA_signal_5680), .Z1_f (new_AGEMA_signal_5681) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U971_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U971_X), .B0_f (new_AGEMA_signal_5679), .B1_t (new_AGEMA_signal_5680), .B1_f (new_AGEMA_signal_5681), .Z0_t (U971_Y), .Z0_f (new_AGEMA_signal_6283), .Z1_t (new_AGEMA_signal_6284), .Z1_f (new_AGEMA_signal_6285) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U971_XOR2_U1 ( .A0_t (U971_Y), .A0_f (new_AGEMA_signal_6283), .A1_t (new_AGEMA_signal_6284), .A1_f (new_AGEMA_signal_6285), .B0_t (StateOut[20]), .B0_f (new_AGEMA_signal_2565), .B1_t (new_AGEMA_signal_2566), .B1_f (new_AGEMA_signal_2567), .Z0_t (StateOut[12]), .Z0_f (new_AGEMA_signal_2562), .Z1_t (new_AGEMA_signal_2563), .Z1_f (new_AGEMA_signal_2564) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U972_XOR1_U1 ( .A0_t (StateOut[28]), .A0_f (new_AGEMA_signal_2574), .A1_t (new_AGEMA_signal_2575), .A1_f (new_AGEMA_signal_2576), .B0_t (StateFromChi[20]), .B0_f (new_AGEMA_signal_4929), .B1_t (new_AGEMA_signal_4930), .B1_f (new_AGEMA_signal_4931), .Z0_t (U972_X), .Z0_f (new_AGEMA_signal_5682), .Z1_t (new_AGEMA_signal_5683), .Z1_f (new_AGEMA_signal_5684) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U972_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U972_X), .B0_f (new_AGEMA_signal_5682), .B1_t (new_AGEMA_signal_5683), .B1_f (new_AGEMA_signal_5684), .Z0_t (U972_Y), .Z0_f (new_AGEMA_signal_6286), .Z1_t (new_AGEMA_signal_6287), .Z1_f (new_AGEMA_signal_6288) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U972_XOR2_U1 ( .A0_t (U972_Y), .A0_f (new_AGEMA_signal_6286), .A1_t (new_AGEMA_signal_6287), .A1_f (new_AGEMA_signal_6288), .B0_t (StateOut[28]), .B0_f (new_AGEMA_signal_2574), .B1_t (new_AGEMA_signal_2575), .B1_f (new_AGEMA_signal_2576), .Z0_t (StateOut[20]), .Z0_f (new_AGEMA_signal_2565), .Z1_t (new_AGEMA_signal_2566), .Z1_f (new_AGEMA_signal_2567) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U973_XOR1_U1 ( .A0_t (StateOut[84]), .A0_f (new_AGEMA_signal_2799), .A1_t (new_AGEMA_signal_2800), .A1_f (new_AGEMA_signal_2801), .B0_t (StateFromChi[76]), .B0_f (new_AGEMA_signal_4962), .B1_t (new_AGEMA_signal_4963), .B1_f (new_AGEMA_signal_4964), .Z0_t (U973_X), .Z0_f (new_AGEMA_signal_5685), .Z1_t (new_AGEMA_signal_5686), .Z1_f (new_AGEMA_signal_5687) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U973_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U973_X), .B0_f (new_AGEMA_signal_5685), .B1_t (new_AGEMA_signal_5686), .B1_f (new_AGEMA_signal_5687), .Z0_t (U973_Y), .Z0_f (new_AGEMA_signal_6289), .Z1_t (new_AGEMA_signal_6290), .Z1_f (new_AGEMA_signal_6291) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U973_XOR2_U1 ( .A0_t (U973_Y), .A0_f (new_AGEMA_signal_6289), .A1_t (new_AGEMA_signal_6290), .A1_f (new_AGEMA_signal_6291), .B0_t (StateOut[84]), .B0_f (new_AGEMA_signal_2799), .B1_t (new_AGEMA_signal_2800), .B1_f (new_AGEMA_signal_2801), .Z0_t (StateOut[76]), .Z0_f (new_AGEMA_signal_2610), .Z1_t (new_AGEMA_signal_2611), .Z1_f (new_AGEMA_signal_2612) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U974_XOR1_U1 ( .A0_t (StateOut[108]), .A0_f (new_AGEMA_signal_2805), .A1_t (new_AGEMA_signal_2806), .A1_f (new_AGEMA_signal_2807), .B0_t (StateFromChi[100]), .B0_f (new_AGEMA_signal_4935), .B1_t (new_AGEMA_signal_4936), .B1_f (new_AGEMA_signal_4937), .Z0_t (U974_X), .Z0_f (new_AGEMA_signal_5688), .Z1_t (new_AGEMA_signal_5689), .Z1_f (new_AGEMA_signal_5690) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U974_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U974_X), .B0_f (new_AGEMA_signal_5688), .B1_t (new_AGEMA_signal_5689), .B1_f (new_AGEMA_signal_5690), .Z0_t (U974_Y), .Z0_f (new_AGEMA_signal_6292), .Z1_t (new_AGEMA_signal_6293), .Z1_f (new_AGEMA_signal_6294) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U974_XOR2_U1 ( .A0_t (U974_Y), .A0_f (new_AGEMA_signal_6292), .A1_t (new_AGEMA_signal_6293), .A1_f (new_AGEMA_signal_6294), .B0_t (StateOut[108]), .B0_f (new_AGEMA_signal_2805), .B1_t (new_AGEMA_signal_2806), .B1_f (new_AGEMA_signal_2807), .Z0_t (StateOut[100]), .Z0_f (new_AGEMA_signal_3228), .Z1_t (new_AGEMA_signal_3229), .Z1_f (new_AGEMA_signal_3230) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U975_XOR1_U1 ( .A0_t (StateOut[116]), .A0_f (new_AGEMA_signal_2808), .A1_t (new_AGEMA_signal_2809), .A1_f (new_AGEMA_signal_2810), .B0_t (StateFromChi[108]), .B0_f (new_AGEMA_signal_4950), .B1_t (new_AGEMA_signal_4951), .B1_f (new_AGEMA_signal_4952), .Z0_t (U975_X), .Z0_f (new_AGEMA_signal_5691), .Z1_t (new_AGEMA_signal_5692), .Z1_f (new_AGEMA_signal_5693) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U975_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U975_X), .B0_f (new_AGEMA_signal_5691), .B1_t (new_AGEMA_signal_5692), .B1_f (new_AGEMA_signal_5693), .Z0_t (U975_Y), .Z0_f (new_AGEMA_signal_6295), .Z1_t (new_AGEMA_signal_6296), .Z1_f (new_AGEMA_signal_6297) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U975_XOR2_U1 ( .A0_t (U975_Y), .A0_f (new_AGEMA_signal_6295), .A1_t (new_AGEMA_signal_6296), .A1_f (new_AGEMA_signal_6297), .B0_t (StateOut[116]), .B0_f (new_AGEMA_signal_2808), .B1_t (new_AGEMA_signal_2809), .B1_f (new_AGEMA_signal_2810), .Z0_t (StateOut[108]), .Z0_f (new_AGEMA_signal_2805), .Z1_t (new_AGEMA_signal_2806), .Z1_f (new_AGEMA_signal_2807) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U976_XOR1_U1 ( .A0_t (StateOut[132]), .A0_f (new_AGEMA_signal_2364), .A1_t (new_AGEMA_signal_2365), .A1_f (new_AGEMA_signal_2366), .B0_t (StateFromChi[124]), .B0_f (new_AGEMA_signal_4908), .B1_t (new_AGEMA_signal_4909), .B1_f (new_AGEMA_signal_4910), .Z0_t (U976_X), .Z0_f (new_AGEMA_signal_5694), .Z1_t (new_AGEMA_signal_5695), .Z1_f (new_AGEMA_signal_5696) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U976_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U976_X), .B0_f (new_AGEMA_signal_5694), .B1_t (new_AGEMA_signal_5695), .B1_f (new_AGEMA_signal_5696), .Z0_t (U976_Y), .Z0_f (new_AGEMA_signal_6298), .Z1_t (new_AGEMA_signal_6299), .Z1_f (new_AGEMA_signal_6300) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U976_XOR2_U1 ( .A0_t (U976_Y), .A0_f (new_AGEMA_signal_6298), .A1_t (new_AGEMA_signal_6299), .A1_f (new_AGEMA_signal_6300), .B0_t (StateOut[132]), .B0_f (new_AGEMA_signal_2364), .B1_t (new_AGEMA_signal_2365), .B1_f (new_AGEMA_signal_2366), .Z0_t (StateOut[124]), .Z0_f (new_AGEMA_signal_3084), .Z1_t (new_AGEMA_signal_3085), .Z1_f (new_AGEMA_signal_3086) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U977_XOR1_U1 ( .A0_t (StateOut[164]), .A0_f (new_AGEMA_signal_2709), .A1_t (new_AGEMA_signal_2710), .A1_f (new_AGEMA_signal_2711), .B0_t (StateFromChi[156]), .B0_f (new_AGEMA_signal_4968), .B1_t (new_AGEMA_signal_4969), .B1_f (new_AGEMA_signal_4970), .Z0_t (U977_X), .Z0_f (new_AGEMA_signal_5697), .Z1_t (new_AGEMA_signal_5698), .Z1_f (new_AGEMA_signal_5699) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U977_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U977_X), .B0_f (new_AGEMA_signal_5697), .B1_t (new_AGEMA_signal_5698), .B1_f (new_AGEMA_signal_5699), .Z0_t (U977_Y), .Z0_f (new_AGEMA_signal_6301), .Z1_t (new_AGEMA_signal_6302), .Z1_f (new_AGEMA_signal_6303) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U977_XOR2_U1 ( .A0_t (U977_Y), .A0_f (new_AGEMA_signal_6301), .A1_t (new_AGEMA_signal_6302), .A1_f (new_AGEMA_signal_6303), .B0_t (StateOut[164]), .B0_f (new_AGEMA_signal_2709), .B1_t (new_AGEMA_signal_2710), .B1_f (new_AGEMA_signal_2711), .Z0_t (StateOut[156]), .Z0_f (new_AGEMA_signal_2373), .Z1_t (new_AGEMA_signal_2374), .Z1_f (new_AGEMA_signal_2375) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U978_XOR1_U1 ( .A0_t (StateOut[188]), .A0_f (new_AGEMA_signal_2715), .A1_t (new_AGEMA_signal_2716), .A1_f (new_AGEMA_signal_2717), .B0_t (StateFromChi[180]), .B0_f (new_AGEMA_signal_4941), .B1_t (new_AGEMA_signal_4942), .B1_f (new_AGEMA_signal_4943), .Z0_t (U978_X), .Z0_f (new_AGEMA_signal_5700), .Z1_t (new_AGEMA_signal_5701), .Z1_f (new_AGEMA_signal_5702) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U978_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U978_X), .B0_f (new_AGEMA_signal_5700), .B1_t (new_AGEMA_signal_5701), .B1_f (new_AGEMA_signal_5702), .Z0_t (U978_Y), .Z0_f (new_AGEMA_signal_6304), .Z1_t (new_AGEMA_signal_6305), .Z1_f (new_AGEMA_signal_6306) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U978_XOR2_U1 ( .A0_t (U978_Y), .A0_f (new_AGEMA_signal_6304), .A1_t (new_AGEMA_signal_6305), .A1_f (new_AGEMA_signal_6306), .B0_t (StateOut[188]), .B0_f (new_AGEMA_signal_2715), .B1_t (new_AGEMA_signal_2716), .B1_f (new_AGEMA_signal_2717), .Z0_t (StateOut[180]), .Z0_f (new_AGEMA_signal_3198), .Z1_t (new_AGEMA_signal_3199), .Z1_f (new_AGEMA_signal_3200) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U979_XOR1_U1 ( .A0_t (StateOut[196]), .A0_f (new_AGEMA_signal_2718), .A1_t (new_AGEMA_signal_2719), .A1_f (new_AGEMA_signal_2720), .B0_t (StateFromChi[188]), .B0_f (new_AGEMA_signal_4956), .B1_t (new_AGEMA_signal_4957), .B1_f (new_AGEMA_signal_4958), .Z0_t (U979_X), .Z0_f (new_AGEMA_signal_5703), .Z1_t (new_AGEMA_signal_5704), .Z1_f (new_AGEMA_signal_5705) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U979_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U979_X), .B0_f (new_AGEMA_signal_5703), .B1_t (new_AGEMA_signal_5704), .B1_f (new_AGEMA_signal_5705), .Z0_t (U979_Y), .Z0_f (new_AGEMA_signal_6307), .Z1_t (new_AGEMA_signal_6308), .Z1_f (new_AGEMA_signal_6309) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U979_XOR2_U1 ( .A0_t (U979_Y), .A0_f (new_AGEMA_signal_6307), .A1_t (new_AGEMA_signal_6308), .A1_f (new_AGEMA_signal_6309), .B0_t (StateOut[196]), .B0_f (new_AGEMA_signal_2718), .B1_t (new_AGEMA_signal_2719), .B1_f (new_AGEMA_signal_2720), .Z0_t (StateOut[188]), .Z0_f (new_AGEMA_signal_2715), .Z1_t (new_AGEMA_signal_2716), .Z1_f (new_AGEMA_signal_2717) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U980_XOR1_U1 ( .A0_t (InData_s0_t[4]), .A0_f (InData_s0_f[4]), .A1_t (InData_s1_t[4]), .A1_f (InData_s1_f[4]), .B0_t (StateFromChi[196]), .B0_f (new_AGEMA_signal_4971), .B1_t (new_AGEMA_signal_4972), .B1_f (new_AGEMA_signal_4973), .Z0_t (U980_X), .Z0_f (new_AGEMA_signal_5709), .Z1_t (new_AGEMA_signal_5710), .Z1_f (new_AGEMA_signal_5711) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U980_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U980_X), .B0_f (new_AGEMA_signal_5709), .B1_t (new_AGEMA_signal_5710), .B1_f (new_AGEMA_signal_5711), .Z0_t (U980_Y), .Z0_f (new_AGEMA_signal_6310), .Z1_t (new_AGEMA_signal_6311), .Z1_f (new_AGEMA_signal_6312) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U980_XOR2_U1 ( .A0_t (U980_Y), .A0_f (new_AGEMA_signal_6310), .A1_t (new_AGEMA_signal_6311), .A1_f (new_AGEMA_signal_6312), .B0_t (InData_s0_t[4]), .B0_f (InData_s0_f[4]), .B1_t (InData_s1_t[4]), .B1_f (InData_s1_f[4]), .Z0_t (StateOut[196]), .Z0_f (new_AGEMA_signal_2718), .Z1_t (new_AGEMA_signal_2719), .Z1_f (new_AGEMA_signal_2720) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U981_XOR1_U1 ( .A0_t (StateOut[19]), .A0_f (new_AGEMA_signal_2187), .A1_t (new_AGEMA_signal_2188), .A1_f (new_AGEMA_signal_2189), .B0_t (StateFromChi[11]), .B0_f (new_AGEMA_signal_4839), .B1_t (new_AGEMA_signal_4840), .B1_f (new_AGEMA_signal_4841), .Z0_t (U981_X), .Z0_f (new_AGEMA_signal_5712), .Z1_t (new_AGEMA_signal_5713), .Z1_f (new_AGEMA_signal_5714) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U981_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U981_X), .B0_f (new_AGEMA_signal_5712), .B1_t (new_AGEMA_signal_5713), .B1_f (new_AGEMA_signal_5714), .Z0_t (U981_Y), .Z0_f (new_AGEMA_signal_6313), .Z1_t (new_AGEMA_signal_6314), .Z1_f (new_AGEMA_signal_6315) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U981_XOR2_U1 ( .A0_t (U981_Y), .A0_f (new_AGEMA_signal_6313), .A1_t (new_AGEMA_signal_6314), .A1_f (new_AGEMA_signal_6315), .B0_t (StateOut[19]), .B0_f (new_AGEMA_signal_2187), .B1_t (new_AGEMA_signal_2188), .B1_f (new_AGEMA_signal_2189), .Z0_t (StateOut[11]), .Z0_f (new_AGEMA_signal_2184), .Z1_t (new_AGEMA_signal_2185), .Z1_f (new_AGEMA_signal_2186) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U982_XOR1_U1 ( .A0_t (StateOut[27]), .A0_f (new_AGEMA_signal_2196), .A1_t (new_AGEMA_signal_2197), .A1_f (new_AGEMA_signal_2198), .B0_t (StateFromChi[19]), .B0_f (new_AGEMA_signal_4854), .B1_t (new_AGEMA_signal_4855), .B1_f (new_AGEMA_signal_4856), .Z0_t (U982_X), .Z0_f (new_AGEMA_signal_5715), .Z1_t (new_AGEMA_signal_5716), .Z1_f (new_AGEMA_signal_5717) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U982_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U982_X), .B0_f (new_AGEMA_signal_5715), .B1_t (new_AGEMA_signal_5716), .B1_f (new_AGEMA_signal_5717), .Z0_t (U982_Y), .Z0_f (new_AGEMA_signal_6316), .Z1_t (new_AGEMA_signal_6317), .Z1_f (new_AGEMA_signal_6318) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U982_XOR2_U1 ( .A0_t (U982_Y), .A0_f (new_AGEMA_signal_6316), .A1_t (new_AGEMA_signal_6317), .A1_f (new_AGEMA_signal_6318), .B0_t (StateOut[27]), .B0_f (new_AGEMA_signal_2196), .B1_t (new_AGEMA_signal_2197), .B1_f (new_AGEMA_signal_2198), .Z0_t (StateOut[19]), .Z0_f (new_AGEMA_signal_2187), .Z1_t (new_AGEMA_signal_2188), .Z1_f (new_AGEMA_signal_2189) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U983_XOR1_U1 ( .A0_t (StateOut[83]), .A0_f (new_AGEMA_signal_2817), .A1_t (new_AGEMA_signal_2818), .A1_f (new_AGEMA_signal_2819), .B0_t (StateFromChi[75]), .B0_f (new_AGEMA_signal_4887), .B1_t (new_AGEMA_signal_4888), .B1_f (new_AGEMA_signal_4889), .Z0_t (U983_X), .Z0_f (new_AGEMA_signal_5718), .Z1_t (new_AGEMA_signal_5719), .Z1_f (new_AGEMA_signal_5720) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U983_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U983_X), .B0_f (new_AGEMA_signal_5718), .B1_t (new_AGEMA_signal_5719), .B1_f (new_AGEMA_signal_5720), .Z0_t (U983_Y), .Z0_f (new_AGEMA_signal_6319), .Z1_t (new_AGEMA_signal_6320), .Z1_f (new_AGEMA_signal_6321) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U983_XOR2_U1 ( .A0_t (U983_Y), .A0_f (new_AGEMA_signal_6319), .A1_t (new_AGEMA_signal_6320), .A1_f (new_AGEMA_signal_6321), .B0_t (StateOut[83]), .B0_f (new_AGEMA_signal_2817), .B1_t (new_AGEMA_signal_2818), .B1_f (new_AGEMA_signal_2819), .Z0_t (StateOut[75]), .Z0_f (new_AGEMA_signal_2628), .Z1_t (new_AGEMA_signal_2629), .Z1_f (new_AGEMA_signal_2630) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U984_XOR1_U1 ( .A0_t (StateOut[107]), .A0_f (new_AGEMA_signal_3234), .A1_t (new_AGEMA_signal_3235), .A1_f (new_AGEMA_signal_3236), .B0_t (StateFromChi[99]), .B0_f (new_AGEMA_signal_4860), .B1_t (new_AGEMA_signal_4861), .B1_f (new_AGEMA_signal_4862), .Z0_t (U984_X), .Z0_f (new_AGEMA_signal_5721), .Z1_t (new_AGEMA_signal_5722), .Z1_f (new_AGEMA_signal_5723) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U984_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U984_X), .B0_f (new_AGEMA_signal_5721), .B1_t (new_AGEMA_signal_5722), .B1_f (new_AGEMA_signal_5723), .Z0_t (U984_Y), .Z0_f (new_AGEMA_signal_6322), .Z1_t (new_AGEMA_signal_6323), .Z1_f (new_AGEMA_signal_6324) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U984_XOR2_U1 ( .A0_t (U984_Y), .A0_f (new_AGEMA_signal_6322), .A1_t (new_AGEMA_signal_6323), .A1_f (new_AGEMA_signal_6324), .B0_t (StateOut[107]), .B0_f (new_AGEMA_signal_3234), .B1_t (new_AGEMA_signal_3235), .B1_f (new_AGEMA_signal_3236), .Z0_t (StateOut[99]), .Z0_f (new_AGEMA_signal_2826), .Z1_t (new_AGEMA_signal_2827), .Z1_f (new_AGEMA_signal_2828) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U985_XOR1_U1 ( .A0_t (StateOut[115]), .A0_f (new_AGEMA_signal_2823), .A1_t (new_AGEMA_signal_2824), .A1_f (new_AGEMA_signal_2825), .B0_t (StateFromChi[107]), .B0_f (new_AGEMA_signal_4875), .B1_t (new_AGEMA_signal_4876), .B1_f (new_AGEMA_signal_4877), .Z0_t (U985_X), .Z0_f (new_AGEMA_signal_5724), .Z1_t (new_AGEMA_signal_5725), .Z1_f (new_AGEMA_signal_5726) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U985_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U985_X), .B0_f (new_AGEMA_signal_5724), .B1_t (new_AGEMA_signal_5725), .B1_f (new_AGEMA_signal_5726), .Z0_t (U985_Y), .Z0_f (new_AGEMA_signal_6325), .Z1_t (new_AGEMA_signal_6326), .Z1_f (new_AGEMA_signal_6327) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U985_XOR2_U1 ( .A0_t (U985_Y), .A0_f (new_AGEMA_signal_6325), .A1_t (new_AGEMA_signal_6326), .A1_f (new_AGEMA_signal_6327), .B0_t (StateOut[115]), .B0_f (new_AGEMA_signal_2823), .B1_t (new_AGEMA_signal_2824), .B1_f (new_AGEMA_signal_2825), .Z0_t (StateOut[107]), .Z0_f (new_AGEMA_signal_3234), .Z1_t (new_AGEMA_signal_3235), .Z1_f (new_AGEMA_signal_3236) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U986_XOR1_U1 ( .A0_t (StateOut[131]), .A0_f (new_AGEMA_signal_2580), .A1_t (new_AGEMA_signal_2581), .A1_f (new_AGEMA_signal_2582), .B0_t (StateFromChi[123]), .B0_f (new_AGEMA_signal_4833), .B1_t (new_AGEMA_signal_4834), .B1_f (new_AGEMA_signal_4835), .Z0_t (U986_X), .Z0_f (new_AGEMA_signal_5727), .Z1_t (new_AGEMA_signal_5728), .Z1_f (new_AGEMA_signal_5729) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U986_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U986_X), .B0_f (new_AGEMA_signal_5727), .B1_t (new_AGEMA_signal_5728), .B1_f (new_AGEMA_signal_5729), .Z0_t (U986_Y), .Z0_f (new_AGEMA_signal_6328), .Z1_t (new_AGEMA_signal_6329), .Z1_f (new_AGEMA_signal_6330) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U986_XOR2_U1 ( .A0_t (U986_Y), .A0_f (new_AGEMA_signal_6328), .A1_t (new_AGEMA_signal_6329), .A1_f (new_AGEMA_signal_6330), .B0_t (StateOut[131]), .B0_f (new_AGEMA_signal_2580), .B1_t (new_AGEMA_signal_2581), .B1_f (new_AGEMA_signal_2582), .Z0_t (StateOut[123]), .Z0_f (new_AGEMA_signal_3156), .Z1_t (new_AGEMA_signal_3157), .Z1_f (new_AGEMA_signal_3158) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U987_XOR1_U1 ( .A0_t (StateOut[163]), .A0_f (new_AGEMA_signal_2781), .A1_t (new_AGEMA_signal_2782), .A1_f (new_AGEMA_signal_2783), .B0_t (StateFromChi[155]), .B0_f (new_AGEMA_signal_4893), .B1_t (new_AGEMA_signal_4894), .B1_f (new_AGEMA_signal_4895), .Z0_t (U987_X), .Z0_f (new_AGEMA_signal_5730), .Z1_t (new_AGEMA_signal_5731), .Z1_f (new_AGEMA_signal_5732) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U987_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U987_X), .B0_f (new_AGEMA_signal_5730), .B1_t (new_AGEMA_signal_5731), .B1_f (new_AGEMA_signal_5732), .Z0_t (U987_Y), .Z0_f (new_AGEMA_signal_6331), .Z1_t (new_AGEMA_signal_6332), .Z1_f (new_AGEMA_signal_6333) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U987_XOR2_U1 ( .A0_t (U987_Y), .A0_f (new_AGEMA_signal_6331), .A1_t (new_AGEMA_signal_6332), .A1_f (new_AGEMA_signal_6333), .B0_t (StateOut[163]), .B0_f (new_AGEMA_signal_2781), .B1_t (new_AGEMA_signal_2782), .B1_f (new_AGEMA_signal_2783), .Z0_t (StateOut[155]), .Z0_f (new_AGEMA_signal_2589), .Z1_t (new_AGEMA_signal_2590), .Z1_f (new_AGEMA_signal_2591) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U988_XOR1_U1 ( .A0_t (StateOut[195]), .A0_f (new_AGEMA_signal_2790), .A1_t (new_AGEMA_signal_2791), .A1_f (new_AGEMA_signal_2792), .B0_t (StateFromChi[187]), .B0_f (new_AGEMA_signal_4881), .B1_t (new_AGEMA_signal_4882), .B1_f (new_AGEMA_signal_4883), .Z0_t (U988_X), .Z0_f (new_AGEMA_signal_5733), .Z1_t (new_AGEMA_signal_5734), .Z1_f (new_AGEMA_signal_5735) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U988_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U988_X), .B0_f (new_AGEMA_signal_5733), .B1_t (new_AGEMA_signal_5734), .B1_f (new_AGEMA_signal_5735), .Z0_t (U988_Y), .Z0_f (new_AGEMA_signal_6334), .Z1_t (new_AGEMA_signal_6335), .Z1_f (new_AGEMA_signal_6336) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U988_XOR2_U1 ( .A0_t (U988_Y), .A0_f (new_AGEMA_signal_6334), .A1_t (new_AGEMA_signal_6335), .A1_f (new_AGEMA_signal_6336), .B0_t (StateOut[195]), .B0_f (new_AGEMA_signal_2790), .B1_t (new_AGEMA_signal_2791), .B1_f (new_AGEMA_signal_2792), .Z0_t (StateOut[187]), .Z0_f (new_AGEMA_signal_2787), .Z1_t (new_AGEMA_signal_2788), .Z1_f (new_AGEMA_signal_2789) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U989_XOR1_U1 ( .A0_t (InData_s0_t[3]), .A0_f (InData_s0_f[3]), .A1_t (InData_s1_t[3]), .A1_f (InData_s1_f[3]), .B0_t (StateFromChi[195]), .B0_f (new_AGEMA_signal_4896), .B1_t (new_AGEMA_signal_4897), .B1_f (new_AGEMA_signal_4898), .Z0_t (U989_X), .Z0_f (new_AGEMA_signal_5739), .Z1_t (new_AGEMA_signal_5740), .Z1_f (new_AGEMA_signal_5741) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U989_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U989_X), .B0_f (new_AGEMA_signal_5739), .B1_t (new_AGEMA_signal_5740), .B1_f (new_AGEMA_signal_5741), .Z0_t (U989_Y), .Z0_f (new_AGEMA_signal_6337), .Z1_t (new_AGEMA_signal_6338), .Z1_f (new_AGEMA_signal_6339) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U989_XOR2_U1 ( .A0_t (U989_Y), .A0_f (new_AGEMA_signal_6337), .A1_t (new_AGEMA_signal_6338), .A1_f (new_AGEMA_signal_6339), .B0_t (InData_s0_t[3]), .B0_f (InData_s0_f[3]), .B1_t (InData_s1_t[3]), .B1_f (InData_s1_f[3]), .Z0_t (StateOut[195]), .Z0_f (new_AGEMA_signal_2790), .Z1_t (new_AGEMA_signal_2791), .Z1_f (new_AGEMA_signal_2792) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U990_XOR1_U1 ( .A0_t (StateOut[18]), .A0_f (new_AGEMA_signal_2538), .A1_t (new_AGEMA_signal_2539), .A1_f (new_AGEMA_signal_2540), .B0_t (StateFromChi[10]), .B0_f (new_AGEMA_signal_4764), .B1_t (new_AGEMA_signal_4765), .B1_f (new_AGEMA_signal_4766), .Z0_t (U990_X), .Z0_f (new_AGEMA_signal_5742), .Z1_t (new_AGEMA_signal_5743), .Z1_f (new_AGEMA_signal_5744) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U990_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U990_X), .B0_f (new_AGEMA_signal_5742), .B1_t (new_AGEMA_signal_5743), .B1_f (new_AGEMA_signal_5744), .Z0_t (U990_Y), .Z0_f (new_AGEMA_signal_6340), .Z1_t (new_AGEMA_signal_6341), .Z1_f (new_AGEMA_signal_6342) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U990_XOR2_U1 ( .A0_t (U990_Y), .A0_f (new_AGEMA_signal_6340), .A1_t (new_AGEMA_signal_6341), .A1_f (new_AGEMA_signal_6342), .B0_t (StateOut[18]), .B0_f (new_AGEMA_signal_2538), .B1_t (new_AGEMA_signal_2539), .B1_f (new_AGEMA_signal_2540), .Z0_t (StateOut[10]), .Z0_f (new_AGEMA_signal_2526), .Z1_t (new_AGEMA_signal_2527), .Z1_f (new_AGEMA_signal_2528) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U991_XOR1_U1 ( .A0_t (StateOut[26]), .A0_f (new_AGEMA_signal_3138), .A1_t (new_AGEMA_signal_3139), .A1_f (new_AGEMA_signal_3140), .B0_t (StateFromChi[18]), .B0_f (new_AGEMA_signal_4779), .B1_t (new_AGEMA_signal_4780), .B1_f (new_AGEMA_signal_4781), .Z0_t (U991_X), .Z0_f (new_AGEMA_signal_5745), .Z1_t (new_AGEMA_signal_5746), .Z1_f (new_AGEMA_signal_5747) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U991_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U991_X), .B0_f (new_AGEMA_signal_5745), .B1_t (new_AGEMA_signal_5746), .B1_f (new_AGEMA_signal_5747), .Z0_t (U991_Y), .Z0_f (new_AGEMA_signal_6343), .Z1_t (new_AGEMA_signal_6344), .Z1_f (new_AGEMA_signal_6345) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U991_XOR2_U1 ( .A0_t (U991_Y), .A0_f (new_AGEMA_signal_6343), .A1_t (new_AGEMA_signal_6344), .A1_f (new_AGEMA_signal_6345), .B0_t (StateOut[26]), .B0_f (new_AGEMA_signal_3138), .B1_t (new_AGEMA_signal_3139), .B1_f (new_AGEMA_signal_3140), .Z0_t (StateOut[18]), .Z0_f (new_AGEMA_signal_2538), .Z1_t (new_AGEMA_signal_2539), .Z1_f (new_AGEMA_signal_2540) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U992_XOR1_U1 ( .A0_t (StateOut[74]), .A0_f (new_AGEMA_signal_2661), .A1_t (new_AGEMA_signal_2662), .A1_f (new_AGEMA_signal_2663), .B0_t (StateFromChi[66]), .B0_f (new_AGEMA_signal_4797), .B1_t (new_AGEMA_signal_4798), .B1_f (new_AGEMA_signal_4799), .Z0_t (U992_X), .Z0_f (new_AGEMA_signal_5748), .Z1_t (new_AGEMA_signal_5749), .Z1_f (new_AGEMA_signal_5750) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U992_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U992_X), .B0_f (new_AGEMA_signal_5748), .B1_t (new_AGEMA_signal_5749), .B1_f (new_AGEMA_signal_5750), .Z0_t (U992_Y), .Z0_f (new_AGEMA_signal_6346), .Z1_t (new_AGEMA_signal_6347), .Z1_f (new_AGEMA_signal_6348) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U992_XOR2_U1 ( .A0_t (U992_Y), .A0_f (new_AGEMA_signal_6346), .A1_t (new_AGEMA_signal_6347), .A1_f (new_AGEMA_signal_6348), .B0_t (StateOut[74]), .B0_f (new_AGEMA_signal_2661), .B1_t (new_AGEMA_signal_2662), .B1_f (new_AGEMA_signal_2663), .Z0_t (StateOut[66]), .Z0_f (new_AGEMA_signal_3180), .Z1_t (new_AGEMA_signal_3181), .Z1_f (new_AGEMA_signal_3182) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U993_XOR1_U1 ( .A0_t (StateOut[82]), .A0_f (new_AGEMA_signal_3036), .A1_t (new_AGEMA_signal_3037), .A1_f (new_AGEMA_signal_3038), .B0_t (StateFromChi[74]), .B0_f (new_AGEMA_signal_4812), .B1_t (new_AGEMA_signal_4813), .B1_f (new_AGEMA_signal_4814), .Z0_t (U993_X), .Z0_f (new_AGEMA_signal_5751), .Z1_t (new_AGEMA_signal_5752), .Z1_f (new_AGEMA_signal_5753) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U993_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U993_X), .B0_f (new_AGEMA_signal_5751), .B1_t (new_AGEMA_signal_5752), .B1_f (new_AGEMA_signal_5753), .Z0_t (U993_Y), .Z0_f (new_AGEMA_signal_6349), .Z1_t (new_AGEMA_signal_6350), .Z1_f (new_AGEMA_signal_6351) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U993_XOR2_U1 ( .A0_t (U993_Y), .A0_f (new_AGEMA_signal_6349), .A1_t (new_AGEMA_signal_6350), .A1_f (new_AGEMA_signal_6351), .B0_t (StateOut[82]), .B0_f (new_AGEMA_signal_3036), .B1_t (new_AGEMA_signal_3037), .B1_f (new_AGEMA_signal_3038), .Z0_t (StateOut[74]), .Z0_f (new_AGEMA_signal_2661), .Z1_t (new_AGEMA_signal_2662), .Z1_f (new_AGEMA_signal_2663) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U994_XOR1_U1 ( .A0_t (StateOut[106]), .A0_f (new_AGEMA_signal_2232), .A1_t (new_AGEMA_signal_2233), .A1_f (new_AGEMA_signal_2234), .B0_t (StateFromChi[98]), .B0_f (new_AGEMA_signal_4785), .B1_t (new_AGEMA_signal_4786), .B1_f (new_AGEMA_signal_4787), .Z0_t (U994_X), .Z0_f (new_AGEMA_signal_5754), .Z1_t (new_AGEMA_signal_5755), .Z1_f (new_AGEMA_signal_5756) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U994_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U994_X), .B0_f (new_AGEMA_signal_5754), .B1_t (new_AGEMA_signal_5755), .B1_f (new_AGEMA_signal_5756), .Z0_t (U994_Y), .Z0_f (new_AGEMA_signal_6352), .Z1_t (new_AGEMA_signal_6353), .Z1_f (new_AGEMA_signal_6354) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U994_XOR2_U1 ( .A0_t (U994_Y), .A0_f (new_AGEMA_signal_6352), .A1_t (new_AGEMA_signal_6353), .A1_f (new_AGEMA_signal_6354), .B0_t (StateOut[106]), .B0_f (new_AGEMA_signal_2232), .B1_t (new_AGEMA_signal_2233), .B1_f (new_AGEMA_signal_2234), .Z0_t (StateOut[98]), .Z0_f (new_AGEMA_signal_2223), .Z1_t (new_AGEMA_signal_2224), .Z1_f (new_AGEMA_signal_2225) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U995_XOR1_U1 ( .A0_t (StateOut[130]), .A0_f (new_AGEMA_signal_2742), .A1_t (new_AGEMA_signal_2743), .A1_f (new_AGEMA_signal_2744), .B0_t (StateFromChi[122]), .B0_f (new_AGEMA_signal_4758), .B1_t (new_AGEMA_signal_4759), .B1_f (new_AGEMA_signal_4760), .Z0_t (U995_X), .Z0_f (new_AGEMA_signal_5757), .Z1_t (new_AGEMA_signal_5758), .Z1_f (new_AGEMA_signal_5759) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U995_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U995_X), .B0_f (new_AGEMA_signal_5757), .B1_t (new_AGEMA_signal_5758), .B1_f (new_AGEMA_signal_5759), .Z0_t (U995_Y), .Z0_f (new_AGEMA_signal_6355), .Z1_t (new_AGEMA_signal_6356), .Z1_f (new_AGEMA_signal_6357) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U995_XOR2_U1 ( .A0_t (U995_Y), .A0_f (new_AGEMA_signal_6355), .A1_t (new_AGEMA_signal_6356), .A1_f (new_AGEMA_signal_6357), .B0_t (StateOut[130]), .B0_f (new_AGEMA_signal_2742), .B1_t (new_AGEMA_signal_2743), .B1_f (new_AGEMA_signal_2744), .Z0_t (StateOut[122]), .Z0_f (new_AGEMA_signal_2745), .Z1_t (new_AGEMA_signal_2746), .Z1_f (new_AGEMA_signal_2747) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U996_XOR1_U1 ( .A0_t (StateOut[194]), .A0_f (new_AGEMA_signal_2841), .A1_t (new_AGEMA_signal_2842), .A1_f (new_AGEMA_signal_2843), .B0_t (StateFromChi[186]), .B0_f (new_AGEMA_signal_4806), .B1_t (new_AGEMA_signal_4807), .B1_f (new_AGEMA_signal_4808), .Z0_t (U996_X), .Z0_f (new_AGEMA_signal_5760), .Z1_t (new_AGEMA_signal_5761), .Z1_f (new_AGEMA_signal_5762) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U996_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U996_X), .B0_f (new_AGEMA_signal_5760), .B1_t (new_AGEMA_signal_5761), .B1_f (new_AGEMA_signal_5762), .Z0_t (U996_Y), .Z0_f (new_AGEMA_signal_6358), .Z1_t (new_AGEMA_signal_6359), .Z1_f (new_AGEMA_signal_6360) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U996_XOR2_U1 ( .A0_t (U996_Y), .A0_f (new_AGEMA_signal_6358), .A1_t (new_AGEMA_signal_6359), .A1_f (new_AGEMA_signal_6360), .B0_t (StateOut[194]), .B0_f (new_AGEMA_signal_2841), .B1_t (new_AGEMA_signal_2842), .B1_f (new_AGEMA_signal_2843), .Z0_t (StateOut[186]), .Z0_f (new_AGEMA_signal_3240), .Z1_t (new_AGEMA_signal_3241), .Z1_f (new_AGEMA_signal_3242) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U997_XOR1_U1 ( .A0_t (StateOut[17]), .A0_f (new_AGEMA_signal_3216), .A1_t (new_AGEMA_signal_3217), .A1_f (new_AGEMA_signal_3218), .B0_t (StateFromChi[9]), .B0_f (new_AGEMA_signal_4689), .B1_t (new_AGEMA_signal_4690), .B1_f (new_AGEMA_signal_4691), .Z0_t (U997_X), .Z0_f (new_AGEMA_signal_5763), .Z1_t (new_AGEMA_signal_5764), .Z1_f (new_AGEMA_signal_5765) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U997_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U997_X), .B0_f (new_AGEMA_signal_5763), .B1_t (new_AGEMA_signal_5764), .B1_f (new_AGEMA_signal_5765), .Z0_t (U997_Y), .Z0_f (new_AGEMA_signal_6361), .Z1_t (new_AGEMA_signal_6362), .Z1_f (new_AGEMA_signal_6363) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U997_XOR2_U1 ( .A0_t (U997_Y), .A0_f (new_AGEMA_signal_6361), .A1_t (new_AGEMA_signal_6362), .A1_f (new_AGEMA_signal_6363), .B0_t (StateOut[17]), .B0_f (new_AGEMA_signal_3216), .B1_t (new_AGEMA_signal_3217), .B1_f (new_AGEMA_signal_3218), .Z0_t (StateOut[9]), .Z0_f (new_AGEMA_signal_2760), .Z1_t (new_AGEMA_signal_2761), .Z1_f (new_AGEMA_signal_2762) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U998_XOR1_U1 ( .A0_t (StateOut[73]), .A0_f (new_AGEMA_signal_2430), .A1_t (new_AGEMA_signal_2431), .A1_f (new_AGEMA_signal_2432), .B0_t (StateFromChi[65]), .B0_f (new_AGEMA_signal_4722), .B1_t (new_AGEMA_signal_4723), .B1_f (new_AGEMA_signal_4724), .Z0_t (U998_X), .Z0_f (new_AGEMA_signal_5766), .Z1_t (new_AGEMA_signal_5767), .Z1_f (new_AGEMA_signal_5768) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U998_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U998_X), .B0_f (new_AGEMA_signal_5766), .B1_t (new_AGEMA_signal_5767), .B1_f (new_AGEMA_signal_5768), .Z0_t (U998_Y), .Z0_f (new_AGEMA_signal_6364), .Z1_t (new_AGEMA_signal_6365), .Z1_f (new_AGEMA_signal_6366) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U998_XOR2_U1 ( .A0_t (U998_Y), .A0_f (new_AGEMA_signal_6364), .A1_t (new_AGEMA_signal_6365), .A1_f (new_AGEMA_signal_6366), .B0_t (StateOut[73]), .B0_f (new_AGEMA_signal_2430), .B1_t (new_AGEMA_signal_2431), .B1_f (new_AGEMA_signal_2432), .Z0_t (StateOut[65]), .Z0_f (new_AGEMA_signal_2427), .Z1_t (new_AGEMA_signal_2428), .Z1_f (new_AGEMA_signal_2429) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U999_XOR1_U1 ( .A0_t (StateOut[81]), .A0_f (new_AGEMA_signal_3060), .A1_t (new_AGEMA_signal_3061), .A1_f (new_AGEMA_signal_3062), .B0_t (StateFromChi[73]), .B0_f (new_AGEMA_signal_4737), .B1_t (new_AGEMA_signal_4738), .B1_f (new_AGEMA_signal_4739), .Z0_t (U999_X), .Z0_f (new_AGEMA_signal_5769), .Z1_t (new_AGEMA_signal_5770), .Z1_f (new_AGEMA_signal_5771) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U999_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U999_X), .B0_f (new_AGEMA_signal_5769), .B1_t (new_AGEMA_signal_5770), .B1_f (new_AGEMA_signal_5771), .Z0_t (U999_Y), .Z0_f (new_AGEMA_signal_6367), .Z1_t (new_AGEMA_signal_6368), .Z1_f (new_AGEMA_signal_6369) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U999_XOR2_U1 ( .A0_t (U999_Y), .A0_f (new_AGEMA_signal_6367), .A1_t (new_AGEMA_signal_6368), .A1_f (new_AGEMA_signal_6369), .B0_t (StateOut[81]), .B0_f (new_AGEMA_signal_3060), .B1_t (new_AGEMA_signal_3061), .B1_f (new_AGEMA_signal_3062), .Z0_t (StateOut[73]), .Z0_f (new_AGEMA_signal_2430), .Z1_t (new_AGEMA_signal_2431), .Z1_f (new_AGEMA_signal_2432) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1000_XOR1_U1 ( .A0_t (StateOut[97]), .A0_f (new_AGEMA_signal_2295), .A1_t (new_AGEMA_signal_2296), .A1_f (new_AGEMA_signal_2297), .B0_t (StateFromChi[89]), .B0_f (new_AGEMA_signal_4695), .B1_t (new_AGEMA_signal_4696), .B1_f (new_AGEMA_signal_4697), .Z0_t (U1000_X), .Z0_f (new_AGEMA_signal_5772), .Z1_t (new_AGEMA_signal_5773), .Z1_f (new_AGEMA_signal_5774) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1000_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U1000_X), .B0_f (new_AGEMA_signal_5772), .B1_t (new_AGEMA_signal_5773), .B1_f (new_AGEMA_signal_5774), .Z0_t (U1000_Y), .Z0_f (new_AGEMA_signal_6370), .Z1_t (new_AGEMA_signal_6371), .Z1_f (new_AGEMA_signal_6372) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U1000_XOR2_U1 ( .A0_t (U1000_Y), .A0_f (new_AGEMA_signal_6370), .A1_t (new_AGEMA_signal_6371), .A1_f (new_AGEMA_signal_6372), .B0_t (StateOut[97]), .B0_f (new_AGEMA_signal_2295), .B1_t (new_AGEMA_signal_2296), .B1_f (new_AGEMA_signal_2297), .Z0_t (StateOut[89]), .Z0_f (new_AGEMA_signal_2292), .Z1_t (new_AGEMA_signal_2293), .Z1_f (new_AGEMA_signal_2294) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1001_XOR1_U1 ( .A0_t (StateOut[105]), .A0_f (new_AGEMA_signal_2304), .A1_t (new_AGEMA_signal_2305), .A1_f (new_AGEMA_signal_2306), .B0_t (StateFromChi[97]), .B0_f (new_AGEMA_signal_4710), .B1_t (new_AGEMA_signal_4711), .B1_f (new_AGEMA_signal_4712), .Z0_t (U1001_X), .Z0_f (new_AGEMA_signal_5775), .Z1_t (new_AGEMA_signal_5776), .Z1_f (new_AGEMA_signal_5777) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1001_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U1001_X), .B0_f (new_AGEMA_signal_5775), .B1_t (new_AGEMA_signal_5776), .B1_f (new_AGEMA_signal_5777), .Z0_t (U1001_Y), .Z0_f (new_AGEMA_signal_6373), .Z1_t (new_AGEMA_signal_6374), .Z1_f (new_AGEMA_signal_6375) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U1001_XOR2_U1 ( .A0_t (U1001_Y), .A0_f (new_AGEMA_signal_6373), .A1_t (new_AGEMA_signal_6374), .A1_f (new_AGEMA_signal_6375), .B0_t (StateOut[105]), .B0_f (new_AGEMA_signal_2304), .B1_t (new_AGEMA_signal_2305), .B1_f (new_AGEMA_signal_2306), .Z0_t (StateOut[97]), .Z0_f (new_AGEMA_signal_2295), .Z1_t (new_AGEMA_signal_2296), .Z1_f (new_AGEMA_signal_2297) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1002_XOR1_U1 ( .A0_t (StateOut[129]), .A0_f (new_AGEMA_signal_2274), .A1_t (new_AGEMA_signal_2275), .A1_f (new_AGEMA_signal_2276), .B0_t (StateFromChi[121]), .B0_f (new_AGEMA_signal_4683), .B1_t (new_AGEMA_signal_4684), .B1_f (new_AGEMA_signal_4685), .Z0_t (U1002_X), .Z0_f (new_AGEMA_signal_5778), .Z1_t (new_AGEMA_signal_5779), .Z1_f (new_AGEMA_signal_5780) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1002_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U1002_X), .B0_f (new_AGEMA_signal_5778), .B1_t (new_AGEMA_signal_5779), .B1_f (new_AGEMA_signal_5780), .Z0_t (U1002_Y), .Z0_f (new_AGEMA_signal_6376), .Z1_t (new_AGEMA_signal_6377), .Z1_f (new_AGEMA_signal_6378) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U1002_XOR2_U1 ( .A0_t (U1002_Y), .A0_f (new_AGEMA_signal_6376), .A1_t (new_AGEMA_signal_6377), .A1_f (new_AGEMA_signal_6378), .B0_t (StateOut[129]), .B0_f (new_AGEMA_signal_2274), .B1_t (new_AGEMA_signal_2275), .B1_f (new_AGEMA_signal_2276), .Z0_t (StateOut[121]), .Z0_f (new_AGEMA_signal_3054), .Z1_t (new_AGEMA_signal_3055), .Z1_f (new_AGEMA_signal_3056) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1003_XOR1_U1 ( .A0_t (StateOut[193]), .A0_f (new_AGEMA_signal_2250), .A1_t (new_AGEMA_signal_2251), .A1_f (new_AGEMA_signal_2252), .B0_t (StateFromChi[185]), .B0_f (new_AGEMA_signal_4731), .B1_t (new_AGEMA_signal_4732), .B1_f (new_AGEMA_signal_4733), .Z0_t (U1003_X), .Z0_f (new_AGEMA_signal_5781), .Z1_t (new_AGEMA_signal_5782), .Z1_f (new_AGEMA_signal_5783) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1003_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U1003_X), .B0_f (new_AGEMA_signal_5781), .B1_t (new_AGEMA_signal_5782), .B1_f (new_AGEMA_signal_5783), .Z0_t (U1003_Y), .Z0_f (new_AGEMA_signal_6379), .Z1_t (new_AGEMA_signal_6380), .Z1_f (new_AGEMA_signal_6381) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U1003_XOR2_U1 ( .A0_t (U1003_Y), .A0_f (new_AGEMA_signal_6379), .A1_t (new_AGEMA_signal_6380), .A1_f (new_AGEMA_signal_6381), .B0_t (StateOut[193]), .B0_f (new_AGEMA_signal_2250), .B1_t (new_AGEMA_signal_2251), .B1_f (new_AGEMA_signal_2252), .Z0_t (StateOut[185]), .Z0_f (new_AGEMA_signal_2247), .Z1_t (new_AGEMA_signal_2248), .Z1_f (new_AGEMA_signal_2249) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1004_XOR1_U1 ( .A0_t (StateOut[16]), .A0_f (new_AGEMA_signal_2205), .A1_t (new_AGEMA_signal_2206), .A1_f (new_AGEMA_signal_2207), .B0_t (StateFromChi[8]), .B0_f (new_AGEMA_signal_4614), .B1_t (new_AGEMA_signal_4615), .B1_f (new_AGEMA_signal_4616), .Z0_t (U1004_X), .Z0_f (new_AGEMA_signal_5784), .Z1_t (new_AGEMA_signal_5785), .Z1_f (new_AGEMA_signal_5786) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1004_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U1004_X), .B0_f (new_AGEMA_signal_5784), .B1_t (new_AGEMA_signal_5785), .B1_f (new_AGEMA_signal_5786), .Z0_t (U1004_Y), .Z0_f (new_AGEMA_signal_6382), .Z1_t (new_AGEMA_signal_6383), .Z1_f (new_AGEMA_signal_6384) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U1004_XOR2_U1 ( .A0_t (U1004_Y), .A0_f (new_AGEMA_signal_6382), .A1_t (new_AGEMA_signal_6383), .A1_f (new_AGEMA_signal_6384), .B0_t (StateOut[16]), .B0_f (new_AGEMA_signal_2205), .B1_t (new_AGEMA_signal_2206), .B1_f (new_AGEMA_signal_2207), .Z0_t (StateOut[8]), .Z0_f (new_AGEMA_signal_2202), .Z1_t (new_AGEMA_signal_2203), .Z1_f (new_AGEMA_signal_2204) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1005_XOR1_U1 ( .A0_t (StateOut[72]), .A0_f (new_AGEMA_signal_2265), .A1_t (new_AGEMA_signal_2266), .A1_f (new_AGEMA_signal_2267), .B0_t (StateFromChi[64]), .B0_f (new_AGEMA_signal_4647), .B1_t (new_AGEMA_signal_4648), .B1_f (new_AGEMA_signal_4649), .Z0_t (U1005_X), .Z0_f (new_AGEMA_signal_5787), .Z1_t (new_AGEMA_signal_5788), .Z1_f (new_AGEMA_signal_5789) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1005_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U1005_X), .B0_f (new_AGEMA_signal_5787), .B1_t (new_AGEMA_signal_5788), .B1_f (new_AGEMA_signal_5789), .Z0_t (U1005_Y), .Z0_f (new_AGEMA_signal_6385), .Z1_t (new_AGEMA_signal_6386), .Z1_f (new_AGEMA_signal_6387) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U1005_XOR2_U1 ( .A0_t (U1005_Y), .A0_f (new_AGEMA_signal_6385), .A1_t (new_AGEMA_signal_6386), .A1_f (new_AGEMA_signal_6387), .B0_t (StateOut[72]), .B0_f (new_AGEMA_signal_2265), .B1_t (new_AGEMA_signal_2266), .B1_f (new_AGEMA_signal_2267), .Z0_t (StateOut[64]), .Z0_f (new_AGEMA_signal_3048), .Z1_t (new_AGEMA_signal_3049), .Z1_f (new_AGEMA_signal_3050) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1006_XOR1_U1 ( .A0_t (StateOut[80]), .A0_f (new_AGEMA_signal_2385), .A1_t (new_AGEMA_signal_2386), .A1_f (new_AGEMA_signal_2387), .B0_t (StateFromChi[72]), .B0_f (new_AGEMA_signal_4662), .B1_t (new_AGEMA_signal_4663), .B1_f (new_AGEMA_signal_4664), .Z0_t (U1006_X), .Z0_f (new_AGEMA_signal_5790), .Z1_t (new_AGEMA_signal_5791), .Z1_f (new_AGEMA_signal_5792) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1006_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U1006_X), .B0_f (new_AGEMA_signal_5790), .B1_t (new_AGEMA_signal_5791), .B1_f (new_AGEMA_signal_5792), .Z0_t (U1006_Y), .Z0_f (new_AGEMA_signal_6388), .Z1_t (new_AGEMA_signal_6389), .Z1_f (new_AGEMA_signal_6390) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U1006_XOR2_U1 ( .A0_t (U1006_Y), .A0_f (new_AGEMA_signal_6388), .A1_t (new_AGEMA_signal_6389), .A1_f (new_AGEMA_signal_6390), .B0_t (StateOut[80]), .B0_f (new_AGEMA_signal_2385), .B1_t (new_AGEMA_signal_2386), .B1_f (new_AGEMA_signal_2387), .Z0_t (StateOut[72]), .Z0_f (new_AGEMA_signal_2265), .Z1_t (new_AGEMA_signal_2266), .Z1_f (new_AGEMA_signal_2267) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1007_XOR1_U1 ( .A0_t (StateOut[96]), .A0_f (new_AGEMA_signal_3090), .A1_t (new_AGEMA_signal_3091), .A1_f (new_AGEMA_signal_3092), .B0_t (StateFromChi[88]), .B0_f (new_AGEMA_signal_4620), .B1_t (new_AGEMA_signal_4621), .B1_f (new_AGEMA_signal_4622), .Z0_t (U1007_X), .Z0_f (new_AGEMA_signal_5793), .Z1_t (new_AGEMA_signal_5794), .Z1_f (new_AGEMA_signal_5795) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1007_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U1007_X), .B0_f (new_AGEMA_signal_5793), .B1_t (new_AGEMA_signal_5794), .B1_f (new_AGEMA_signal_5795), .Z0_t (U1007_Y), .Z0_f (new_AGEMA_signal_6391), .Z1_t (new_AGEMA_signal_6392), .Z1_f (new_AGEMA_signal_6393) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U1007_XOR2_U1 ( .A0_t (U1007_Y), .A0_f (new_AGEMA_signal_6391), .A1_t (new_AGEMA_signal_6392), .A1_f (new_AGEMA_signal_6393), .B0_t (StateOut[96]), .B0_f (new_AGEMA_signal_3090), .B1_t (new_AGEMA_signal_3091), .B1_f (new_AGEMA_signal_3092), .Z0_t (StateOut[88]), .Z0_f (new_AGEMA_signal_2382), .Z1_t (new_AGEMA_signal_2383), .Z1_f (new_AGEMA_signal_2384) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1008_XOR1_U1 ( .A0_t (StateOut[104]), .A0_f (new_AGEMA_signal_2391), .A1_t (new_AGEMA_signal_2392), .A1_f (new_AGEMA_signal_2393), .B0_t (StateFromChi[96]), .B0_f (new_AGEMA_signal_4635), .B1_t (new_AGEMA_signal_4636), .B1_f (new_AGEMA_signal_4637), .Z0_t (U1008_X), .Z0_f (new_AGEMA_signal_5796), .Z1_t (new_AGEMA_signal_5797), .Z1_f (new_AGEMA_signal_5798) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1008_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U1008_X), .B0_f (new_AGEMA_signal_5796), .B1_t (new_AGEMA_signal_5797), .B1_f (new_AGEMA_signal_5798), .Z0_t (U1008_Y), .Z0_f (new_AGEMA_signal_6394), .Z1_t (new_AGEMA_signal_6395), .Z1_f (new_AGEMA_signal_6396) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U1008_XOR2_U1 ( .A0_t (U1008_Y), .A0_f (new_AGEMA_signal_6394), .A1_t (new_AGEMA_signal_6395), .A1_f (new_AGEMA_signal_6396), .B0_t (StateOut[104]), .B0_f (new_AGEMA_signal_2391), .B1_t (new_AGEMA_signal_2392), .B1_f (new_AGEMA_signal_2393), .Z0_t (StateOut[96]), .Z0_f (new_AGEMA_signal_3090), .Z1_t (new_AGEMA_signal_3091), .Z1_f (new_AGEMA_signal_3092) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1009_XOR1_U1 ( .A0_t (StateOut[128]), .A0_f (new_AGEMA_signal_2400), .A1_t (new_AGEMA_signal_2401), .A1_f (new_AGEMA_signal_2402), .B0_t (StateFromChi[120]), .B0_f (new_AGEMA_signal_4608), .B1_t (new_AGEMA_signal_4609), .B1_f (new_AGEMA_signal_4610), .Z0_t (U1009_X), .Z0_f (new_AGEMA_signal_5799), .Z1_t (new_AGEMA_signal_5800), .Z1_f (new_AGEMA_signal_5801) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1009_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U1009_X), .B0_f (new_AGEMA_signal_5799), .B1_t (new_AGEMA_signal_5800), .B1_f (new_AGEMA_signal_5801), .Z0_t (U1009_Y), .Z0_f (new_AGEMA_signal_6397), .Z1_t (new_AGEMA_signal_6398), .Z1_f (new_AGEMA_signal_6399) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U1009_XOR2_U1 ( .A0_t (U1009_Y), .A0_f (new_AGEMA_signal_6397), .A1_t (new_AGEMA_signal_6398), .A1_f (new_AGEMA_signal_6399), .B0_t (StateOut[128]), .B0_f (new_AGEMA_signal_2400), .B1_t (new_AGEMA_signal_2401), .B1_f (new_AGEMA_signal_2402), .Z0_t (StateOut[120]), .Z0_f (new_AGEMA_signal_2403), .Z1_t (new_AGEMA_signal_2404), .Z1_f (new_AGEMA_signal_2405) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1010_XOR1_U1 ( .A0_t (StateOut[136]), .A0_f (new_AGEMA_signal_2412), .A1_t (new_AGEMA_signal_2413), .A1_f (new_AGEMA_signal_2414), .B0_t (StateFromChi[128]), .B0_f (new_AGEMA_signal_4623), .B1_t (new_AGEMA_signal_4624), .B1_f (new_AGEMA_signal_4625), .Z0_t (U1010_X), .Z0_f (new_AGEMA_signal_5802), .Z1_t (new_AGEMA_signal_5803), .Z1_f (new_AGEMA_signal_5804) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1010_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U1010_X), .B0_f (new_AGEMA_signal_5802), .B1_t (new_AGEMA_signal_5803), .B1_f (new_AGEMA_signal_5804), .Z0_t (U1010_Y), .Z0_f (new_AGEMA_signal_6400), .Z1_t (new_AGEMA_signal_6401), .Z1_f (new_AGEMA_signal_6402) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U1010_XOR2_U1 ( .A0_t (U1010_Y), .A0_f (new_AGEMA_signal_6400), .A1_t (new_AGEMA_signal_6401), .A1_f (new_AGEMA_signal_6402), .B0_t (StateOut[136]), .B0_f (new_AGEMA_signal_2412), .B1_t (new_AGEMA_signal_2413), .B1_f (new_AGEMA_signal_2414), .Z0_t (StateOut[128]), .Z0_f (new_AGEMA_signal_2400), .Z1_t (new_AGEMA_signal_2401), .Z1_f (new_AGEMA_signal_2402) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1011_XOR1_U1 ( .A0_t (StateOut[184]), .A0_f (new_AGEMA_signal_2322), .A1_t (new_AGEMA_signal_2323), .A1_f (new_AGEMA_signal_2324), .B0_t (StateFromChi[176]), .B0_f (new_AGEMA_signal_4641), .B1_t (new_AGEMA_signal_4642), .B1_f (new_AGEMA_signal_4643), .Z0_t (U1011_X), .Z0_f (new_AGEMA_signal_5805), .Z1_t (new_AGEMA_signal_5806), .Z1_f (new_AGEMA_signal_5807) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1011_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U1011_X), .B0_f (new_AGEMA_signal_5805), .B1_t (new_AGEMA_signal_5806), .B1_f (new_AGEMA_signal_5807), .Z0_t (U1011_Y), .Z0_f (new_AGEMA_signal_6403), .Z1_t (new_AGEMA_signal_6404), .Z1_f (new_AGEMA_signal_6405) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U1011_XOR2_U1 ( .A0_t (U1011_Y), .A0_f (new_AGEMA_signal_6403), .A1_t (new_AGEMA_signal_6404), .A1_f (new_AGEMA_signal_6405), .B0_t (StateOut[184]), .B0_f (new_AGEMA_signal_2322), .B1_t (new_AGEMA_signal_2323), .B1_f (new_AGEMA_signal_2324), .Z0_t (StateOut[176]), .Z0_f (new_AGEMA_signal_2313), .Z1_t (new_AGEMA_signal_2314), .Z1_f (new_AGEMA_signal_2315) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1012_XOR1_U1 ( .A0_t (StateOut[192]), .A0_f (new_AGEMA_signal_2319), .A1_t (new_AGEMA_signal_2320), .A1_f (new_AGEMA_signal_2321), .B0_t (StateFromChi[184]), .B0_f (new_AGEMA_signal_4656), .B1_t (new_AGEMA_signal_4657), .B1_f (new_AGEMA_signal_4658), .Z0_t (U1012_X), .Z0_f (new_AGEMA_signal_5808), .Z1_t (new_AGEMA_signal_5809), .Z1_f (new_AGEMA_signal_5810) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1012_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U1012_X), .B0_f (new_AGEMA_signal_5808), .B1_t (new_AGEMA_signal_5809), .B1_f (new_AGEMA_signal_5810), .Z0_t (U1012_Y), .Z0_f (new_AGEMA_signal_6406), .Z1_t (new_AGEMA_signal_6407), .Z1_f (new_AGEMA_signal_6408) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U1012_XOR2_U1 ( .A0_t (U1012_Y), .A0_f (new_AGEMA_signal_6406), .A1_t (new_AGEMA_signal_6407), .A1_f (new_AGEMA_signal_6408), .B0_t (StateOut[192]), .B0_f (new_AGEMA_signal_2319), .B1_t (new_AGEMA_signal_2320), .B1_f (new_AGEMA_signal_2321), .Z0_t (StateOut[184]), .Z0_f (new_AGEMA_signal_2322), .Z1_t (new_AGEMA_signal_2323), .Z1_f (new_AGEMA_signal_2324) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1013_XOR1_U1 ( .A0_t (StateOut[14]), .A0_f (new_AGEMA_signal_2130), .A1_t (new_AGEMA_signal_2131), .A1_f (new_AGEMA_signal_2132), .B0_t (StateFromChi[6]), .B0_f (new_AGEMA_signal_5049), .B1_t (new_AGEMA_signal_5050), .B1_f (new_AGEMA_signal_5051), .Z0_t (U1013_X), .Z0_f (new_AGEMA_signal_5811), .Z1_t (new_AGEMA_signal_5812), .Z1_f (new_AGEMA_signal_5813) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1013_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U1013_X), .B0_f (new_AGEMA_signal_5811), .B1_t (new_AGEMA_signal_5812), .B1_f (new_AGEMA_signal_5813), .Z0_t (U1013_Y), .Z0_f (new_AGEMA_signal_6409), .Z1_t (new_AGEMA_signal_6410), .Z1_f (new_AGEMA_signal_6411) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U1013_XOR2_U1 ( .A0_t (U1013_Y), .A0_f (new_AGEMA_signal_6409), .A1_t (new_AGEMA_signal_6410), .A1_f (new_AGEMA_signal_6411), .B0_t (StateOut[14]), .B0_f (new_AGEMA_signal_2130), .B1_t (new_AGEMA_signal_2131), .B1_f (new_AGEMA_signal_2132), .Z0_t (OutData_s0_t[6]), .Z0_f (OutData_s0_f[6]), .Z1_t (OutData_s1_t[6]), .Z1_f (OutData_s1_f[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1014_XOR1_U1 ( .A0_t (StateOut[13]), .A0_f (new_AGEMA_signal_2634), .A1_t (new_AGEMA_signal_2635), .A1_f (new_AGEMA_signal_2636), .B0_t (StateFromChi[5]), .B0_f (new_AGEMA_signal_4974), .B1_t (new_AGEMA_signal_4975), .B1_f (new_AGEMA_signal_4976), .Z0_t (U1014_X), .Z0_f (new_AGEMA_signal_5814), .Z1_t (new_AGEMA_signal_5815), .Z1_f (new_AGEMA_signal_5816) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1014_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U1014_X), .B0_f (new_AGEMA_signal_5814), .B1_t (new_AGEMA_signal_5815), .B1_f (new_AGEMA_signal_5816), .Z0_t (U1014_Y), .Z0_f (new_AGEMA_signal_6412), .Z1_t (new_AGEMA_signal_6413), .Z1_f (new_AGEMA_signal_6414) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U1014_XOR2_U1 ( .A0_t (U1014_Y), .A0_f (new_AGEMA_signal_6412), .A1_t (new_AGEMA_signal_6413), .A1_f (new_AGEMA_signal_6414), .B0_t (StateOut[13]), .B0_f (new_AGEMA_signal_2634), .B1_t (new_AGEMA_signal_2635), .B1_f (new_AGEMA_signal_2636), .Z0_t (OutData_s0_t[5]), .Z0_f (OutData_s0_f[5]), .Z1_t (OutData_s1_t[5]), .Z1_f (OutData_s1_f[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1015_XOR1_U1 ( .A0_t (StateOut[12]), .A0_f (new_AGEMA_signal_2562), .A1_t (new_AGEMA_signal_2563), .A1_f (new_AGEMA_signal_2564), .B0_t (StateFromChi[4]), .B0_f (new_AGEMA_signal_4899), .B1_t (new_AGEMA_signal_4900), .B1_f (new_AGEMA_signal_4901), .Z0_t (U1015_X), .Z0_f (new_AGEMA_signal_5817), .Z1_t (new_AGEMA_signal_5818), .Z1_f (new_AGEMA_signal_5819) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1015_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U1015_X), .B0_f (new_AGEMA_signal_5817), .B1_t (new_AGEMA_signal_5818), .B1_f (new_AGEMA_signal_5819), .Z0_t (U1015_Y), .Z0_f (new_AGEMA_signal_6415), .Z1_t (new_AGEMA_signal_6416), .Z1_f (new_AGEMA_signal_6417) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U1015_XOR2_U1 ( .A0_t (U1015_Y), .A0_f (new_AGEMA_signal_6415), .A1_t (new_AGEMA_signal_6416), .A1_f (new_AGEMA_signal_6417), .B0_t (StateOut[12]), .B0_f (new_AGEMA_signal_2562), .B1_t (new_AGEMA_signal_2563), .B1_f (new_AGEMA_signal_2564), .Z0_t (OutData_s0_t[4]), .Z0_f (OutData_s0_f[4]), .Z1_t (OutData_s1_t[4]), .Z1_f (OutData_s1_f[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1016_XOR1_U1 ( .A0_t (StateOut[10]), .A0_f (new_AGEMA_signal_2526), .A1_t (new_AGEMA_signal_2527), .A1_f (new_AGEMA_signal_2528), .B0_t (StateFromChi[2]), .B0_f (new_AGEMA_signal_4749), .B1_t (new_AGEMA_signal_4750), .B1_f (new_AGEMA_signal_4751), .Z0_t (U1016_X), .Z0_f (new_AGEMA_signal_5820), .Z1_t (new_AGEMA_signal_5821), .Z1_f (new_AGEMA_signal_5822) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1016_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (n9), .A1_f (new_AGEMA_signal_3005), .B0_t (U1016_X), .B0_f (new_AGEMA_signal_5820), .B1_t (new_AGEMA_signal_5821), .B1_f (new_AGEMA_signal_5822), .Z0_t (U1016_Y), .Z0_f (new_AGEMA_signal_6418), .Z1_t (new_AGEMA_signal_6419), .Z1_f (new_AGEMA_signal_6420) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U1016_XOR2_U1 ( .A0_t (U1016_Y), .A0_f (new_AGEMA_signal_6418), .A1_t (new_AGEMA_signal_6419), .A1_f (new_AGEMA_signal_6420), .B0_t (StateOut[10]), .B0_f (new_AGEMA_signal_2526), .B1_t (new_AGEMA_signal_2527), .B1_f (new_AGEMA_signal_2528), .Z0_t (OutData_s0_t[2]), .Z0_f (OutData_s0_f[2]), .Z1_t (OutData_s1_t[2]), .Z1_f (OutData_s1_f[2]) ) ;

    /* register cells */
endmodule
