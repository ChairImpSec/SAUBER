/* modified netlist. Source: module main in file /mnt/c/Users/amirm/Desktop/Papers_in_progress/SAUBER/Design for our FPGA/3-AES_Sbox_with_control_MUX/4-AGEMA/main.v */
/* 0 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 1 register stage(s) in total */

module main_SAUBER_Pipeline_d1 (value_in_s0_t, start_t, rst_t, value_in_s0_f, value_in_s1_t, value_in_s1_f, start_f, rst_f, value_out_s0_t, value_out_s0_f, value_out_s1_t, value_out_s1_f);
    input [7:0] value_in_s0_t ;
    input [3:0] start_t ;
    input rst_t ;
    input [7:0] value_in_s0_f ;
    input [7:0] value_in_s1_t ;
    input [7:0] value_in_s1_f ;
    input [3:0] start_f ;
    input rst_f ;
    output [7:0] value_out_s0_t ;
    output [7:0] value_out_s0_f ;
    output [7:0] value_out_s1_t ;
    output [7:0] value_out_s1_f ;
    wire n9 ;
    wire n10 ;
    wire [3:3] Inc_out ;
    wire [7:0] Sbox_in ;
    wire [3:0] Inc_Reg ;
    wire [3:0] Inc_in ;
    wire \M1.gen_loop_0__M.X ;
    wire \M1.gen_loop_0__M.Y ;
    wire \M1.gen_loop_1__M.X ;
    wire \M1.gen_loop_1__M.Y ;
    wire \M1.gen_loop_2__M.X ;
    wire \M1.gen_loop_2__M.Y ;
    wire \M1.gen_loop_3__M.X ;
    wire \M1.gen_loop_3__M.Y ;
    wire \M1.gen_loop_4__M.X ;
    wire \M1.gen_loop_4__M.Y ;
    wire \M1.gen_loop_5__M.X ;
    wire \M1.gen_loop_5__M.Y ;
    wire \M1.gen_loop_6__M.X ;
    wire \M1.gen_loop_6__M.Y ;
    wire \M1.gen_loop_7__M.X ;
    wire \M1.gen_loop_7__M.Y ;
    wire \SboxInst.T1 ;
    wire \SboxInst.T2 ;
    wire \SboxInst.T3 ;
    wire \SboxInst.T4 ;
    wire \SboxInst.T5 ;
    wire \SboxInst.T6 ;
    wire \SboxInst.T7 ;
    wire \SboxInst.T8 ;
    wire \SboxInst.T9 ;
    wire \SboxInst.T10 ;
    wire \SboxInst.T11 ;
    wire \SboxInst.T12 ;
    wire \SboxInst.T13 ;
    wire \SboxInst.T14 ;
    wire \SboxInst.T15 ;
    wire \SboxInst.T16 ;
    wire \SboxInst.T17 ;
    wire \SboxInst.T18 ;
    wire \SboxInst.T19 ;
    wire \SboxInst.T20 ;
    wire \SboxInst.T21 ;
    wire \SboxInst.T22 ;
    wire \SboxInst.T23 ;
    wire \SboxInst.T24 ;
    wire \SboxInst.T25 ;
    wire \SboxInst.T26 ;
    wire \SboxInst.T27 ;
    wire \SboxInst.M1 ;
    wire \SboxInst.M2 ;
    wire \SboxInst.M3 ;
    wire \SboxInst.M4 ;
    wire \SboxInst.M5 ;
    wire \SboxInst.M6 ;
    wire \SboxInst.M7 ;
    wire \SboxInst.M8 ;
    wire \SboxInst.M9 ;
    wire \SboxInst.M10 ;
    wire \SboxInst.M11 ;
    wire \SboxInst.M12 ;
    wire \SboxInst.M13 ;
    wire \SboxInst.M14 ;
    wire \SboxInst.M15 ;
    wire \SboxInst.M16 ;
    wire \SboxInst.M17 ;
    wire \SboxInst.M18 ;
    wire \SboxInst.M19 ;
    wire \SboxInst.M20 ;
    wire \SboxInst.M21 ;
    wire \SboxInst.M22 ;
    wire \SboxInst.M23 ;
    wire \SboxInst.M24 ;
    wire \SboxInst.M25 ;
    wire \SboxInst.M26 ;
    wire \SboxInst.M27 ;
    wire \SboxInst.M28 ;
    wire \SboxInst.M29 ;
    wire \SboxInst.M30 ;
    wire \SboxInst.M31 ;
    wire \SboxInst.M32 ;
    wire \SboxInst.M33 ;
    wire \SboxInst.M34 ;
    wire \SboxInst.M35 ;
    wire \SboxInst.M36 ;
    wire \SboxInst.M37 ;
    wire \SboxInst.M38 ;
    wire \SboxInst.M39 ;
    wire \SboxInst.M40 ;
    wire \SboxInst.M41 ;
    wire \SboxInst.M42 ;
    wire \SboxInst.M43 ;
    wire \SboxInst.M44 ;
    wire \SboxInst.M45 ;
    wire \SboxInst.M46 ;
    wire \SboxInst.M47 ;
    wire \SboxInst.M48 ;
    wire \SboxInst.M49 ;
    wire \SboxInst.M50 ;
    wire \SboxInst.M51 ;
    wire \SboxInst.M52 ;
    wire \SboxInst.M53 ;
    wire \SboxInst.M54 ;
    wire \SboxInst.M55 ;
    wire \SboxInst.M56 ;
    wire \SboxInst.M57 ;
    wire \SboxInst.M58 ;
    wire \SboxInst.M59 ;
    wire \SboxInst.M60 ;
    wire \SboxInst.M61 ;
    wire \SboxInst.M62 ;
    wire \SboxInst.M63 ;
    wire \SboxInst.L0 ;
    wire \SboxInst.L1 ;
    wire \SboxInst.L2 ;
    wire \SboxInst.L3 ;
    wire \SboxInst.L4 ;
    wire \SboxInst.L5 ;
    wire \SboxInst.L6 ;
    wire \SboxInst.L7 ;
    wire \SboxInst.L8 ;
    wire \SboxInst.L9 ;
    wire \SboxInst.L10 ;
    wire \SboxInst.L11 ;
    wire \SboxInst.L12 ;
    wire \SboxInst.L13 ;
    wire \SboxInst.L14 ;
    wire \SboxInst.L15 ;
    wire \SboxInst.L16 ;
    wire \SboxInst.L17 ;
    wire \SboxInst.L18 ;
    wire \SboxInst.L19 ;
    wire \SboxInst.L20 ;
    wire \SboxInst.L21 ;
    wire \SboxInst.L22 ;
    wire \SboxInst.L23 ;
    wire \SboxInst.L24 ;
    wire \SboxInst.L25 ;
    wire \SboxInst.L26 ;
    wire \SboxInst.L27 ;
    wire \SboxInst.L28 ;
    wire \SboxInst.L29 ;
    wire \M2.gen_loop_0__M.X ;
    wire \M2.gen_loop_0__M.Y ;
    wire \M2.gen_loop_1__M.X ;
    wire \M2.gen_loop_1__M.Y ;
    wire \M2.gen_loop_2__M.X ;
    wire \M2.gen_loop_2__M.Y ;
    wire \M2.gen_loop_3__M.X ;
    wire \M2.gen_loop_3__M.Y ;
    wire new_AGEMA_signal_864 ;
    wire new_AGEMA_signal_865 ;
    wire new_AGEMA_signal_866 ;
    wire new_AGEMA_signal_873 ;
    wire new_AGEMA_signal_874 ;
    wire new_AGEMA_signal_875 ;
    wire new_AGEMA_signal_882 ;
    wire new_AGEMA_signal_883 ;
    wire new_AGEMA_signal_884 ;
    wire new_AGEMA_signal_891 ;
    wire new_AGEMA_signal_892 ;
    wire new_AGEMA_signal_893 ;
    wire new_AGEMA_signal_900 ;
    wire new_AGEMA_signal_901 ;
    wire new_AGEMA_signal_902 ;
    wire new_AGEMA_signal_909 ;
    wire new_AGEMA_signal_910 ;
    wire new_AGEMA_signal_911 ;
    wire new_AGEMA_signal_918 ;
    wire new_AGEMA_signal_919 ;
    wire new_AGEMA_signal_920 ;
    wire new_AGEMA_signal_927 ;
    wire new_AGEMA_signal_928 ;
    wire new_AGEMA_signal_929 ;
    wire new_AGEMA_signal_930 ;
    wire new_AGEMA_signal_932 ;
    wire new_AGEMA_signal_933 ;
    wire new_AGEMA_signal_935 ;
    wire new_AGEMA_signal_936 ;
    wire new_AGEMA_signal_938 ;
    wire new_AGEMA_signal_939 ;
    wire new_AGEMA_signal_941 ;
    wire new_AGEMA_signal_943 ;
    wire new_AGEMA_signal_944 ;
    wire new_AGEMA_signal_945 ;
    wire new_AGEMA_signal_946 ;
    wire new_AGEMA_signal_947 ;
    wire new_AGEMA_signal_948 ;
    wire new_AGEMA_signal_949 ;
    wire new_AGEMA_signal_950 ;
    wire new_AGEMA_signal_951 ;
    wire new_AGEMA_signal_952 ;
    wire new_AGEMA_signal_953 ;
    wire new_AGEMA_signal_954 ;
    wire new_AGEMA_signal_955 ;
    wire new_AGEMA_signal_956 ;
    wire new_AGEMA_signal_957 ;
    wire new_AGEMA_signal_958 ;
    wire new_AGEMA_signal_959 ;
    wire new_AGEMA_signal_960 ;
    wire new_AGEMA_signal_961 ;
    wire new_AGEMA_signal_962 ;
    wire new_AGEMA_signal_963 ;
    wire new_AGEMA_signal_964 ;
    wire new_AGEMA_signal_965 ;
    wire new_AGEMA_signal_966 ;
    wire new_AGEMA_signal_967 ;
    wire new_AGEMA_signal_968 ;
    wire new_AGEMA_signal_969 ;
    wire new_AGEMA_signal_970 ;
    wire new_AGEMA_signal_971 ;
    wire new_AGEMA_signal_972 ;
    wire new_AGEMA_signal_973 ;
    wire new_AGEMA_signal_974 ;
    wire new_AGEMA_signal_975 ;
    wire new_AGEMA_signal_976 ;
    wire new_AGEMA_signal_977 ;
    wire new_AGEMA_signal_978 ;
    wire new_AGEMA_signal_979 ;
    wire new_AGEMA_signal_980 ;
    wire new_AGEMA_signal_981 ;
    wire new_AGEMA_signal_982 ;
    wire new_AGEMA_signal_983 ;
    wire new_AGEMA_signal_984 ;
    wire new_AGEMA_signal_985 ;
    wire new_AGEMA_signal_986 ;
    wire new_AGEMA_signal_987 ;
    wire new_AGEMA_signal_988 ;
    wire new_AGEMA_signal_989 ;
    wire new_AGEMA_signal_990 ;
    wire new_AGEMA_signal_991 ;
    wire new_AGEMA_signal_992 ;
    wire new_AGEMA_signal_993 ;
    wire new_AGEMA_signal_994 ;
    wire new_AGEMA_signal_995 ;
    wire new_AGEMA_signal_996 ;
    wire new_AGEMA_signal_997 ;
    wire new_AGEMA_signal_998 ;
    wire new_AGEMA_signal_999 ;
    wire new_AGEMA_signal_1000 ;
    wire new_AGEMA_signal_1001 ;
    wire new_AGEMA_signal_1002 ;
    wire new_AGEMA_signal_1003 ;
    wire new_AGEMA_signal_1004 ;
    wire new_AGEMA_signal_1005 ;
    wire new_AGEMA_signal_1006 ;
    wire new_AGEMA_signal_1007 ;
    wire new_AGEMA_signal_1008 ;
    wire new_AGEMA_signal_1009 ;
    wire new_AGEMA_signal_1010 ;
    wire new_AGEMA_signal_1011 ;
    wire new_AGEMA_signal_1012 ;
    wire new_AGEMA_signal_1013 ;
    wire new_AGEMA_signal_1014 ;
    wire new_AGEMA_signal_1015 ;
    wire new_AGEMA_signal_1016 ;
    wire new_AGEMA_signal_1017 ;
    wire new_AGEMA_signal_1018 ;
    wire new_AGEMA_signal_1019 ;
    wire new_AGEMA_signal_1020 ;
    wire new_AGEMA_signal_1021 ;
    wire new_AGEMA_signal_1022 ;
    wire new_AGEMA_signal_1023 ;
    wire new_AGEMA_signal_1024 ;
    wire new_AGEMA_signal_1025 ;
    wire new_AGEMA_signal_1026 ;
    wire new_AGEMA_signal_1027 ;
    wire new_AGEMA_signal_1028 ;
    wire new_AGEMA_signal_1029 ;
    wire new_AGEMA_signal_1030 ;
    wire new_AGEMA_signal_1031 ;
    wire new_AGEMA_signal_1032 ;
    wire new_AGEMA_signal_1033 ;
    wire new_AGEMA_signal_1034 ;
    wire new_AGEMA_signal_1035 ;
    wire new_AGEMA_signal_1036 ;
    wire new_AGEMA_signal_1037 ;
    wire new_AGEMA_signal_1038 ;
    wire new_AGEMA_signal_1039 ;
    wire new_AGEMA_signal_1040 ;
    wire new_AGEMA_signal_1041 ;
    wire new_AGEMA_signal_1042 ;
    wire new_AGEMA_signal_1043 ;
    wire new_AGEMA_signal_1044 ;
    wire new_AGEMA_signal_1045 ;
    wire new_AGEMA_signal_1046 ;
    wire new_AGEMA_signal_1047 ;
    wire new_AGEMA_signal_1048 ;
    wire new_AGEMA_signal_1049 ;
    wire new_AGEMA_signal_1050 ;
    wire new_AGEMA_signal_1051 ;
    wire new_AGEMA_signal_1052 ;
    wire new_AGEMA_signal_1053 ;
    wire new_AGEMA_signal_1054 ;
    wire new_AGEMA_signal_1055 ;
    wire new_AGEMA_signal_1056 ;
    wire new_AGEMA_signal_1057 ;
    wire new_AGEMA_signal_1058 ;
    wire new_AGEMA_signal_1059 ;
    wire new_AGEMA_signal_1060 ;
    wire new_AGEMA_signal_1061 ;
    wire new_AGEMA_signal_1062 ;
    wire new_AGEMA_signal_1063 ;
    wire new_AGEMA_signal_1064 ;
    wire new_AGEMA_signal_1065 ;
    wire new_AGEMA_signal_1066 ;
    wire new_AGEMA_signal_1067 ;
    wire new_AGEMA_signal_1068 ;
    wire new_AGEMA_signal_1069 ;
    wire new_AGEMA_signal_1070 ;
    wire new_AGEMA_signal_1071 ;
    wire new_AGEMA_signal_1072 ;
    wire new_AGEMA_signal_1073 ;
    wire new_AGEMA_signal_1074 ;
    wire new_AGEMA_signal_1075 ;
    wire new_AGEMA_signal_1076 ;
    wire new_AGEMA_signal_1077 ;
    wire new_AGEMA_signal_1078 ;
    wire new_AGEMA_signal_1079 ;
    wire new_AGEMA_signal_1080 ;
    wire new_AGEMA_signal_1081 ;
    wire new_AGEMA_signal_1082 ;
    wire new_AGEMA_signal_1083 ;
    wire new_AGEMA_signal_1084 ;
    wire new_AGEMA_signal_1085 ;
    wire new_AGEMA_signal_1086 ;
    wire new_AGEMA_signal_1087 ;
    wire new_AGEMA_signal_1088 ;
    wire new_AGEMA_signal_1089 ;
    wire new_AGEMA_signal_1090 ;
    wire new_AGEMA_signal_1091 ;
    wire new_AGEMA_signal_1092 ;
    wire new_AGEMA_signal_1093 ;
    wire new_AGEMA_signal_1094 ;
    wire new_AGEMA_signal_1095 ;
    wire new_AGEMA_signal_1096 ;
    wire new_AGEMA_signal_1097 ;
    wire new_AGEMA_signal_1098 ;
    wire new_AGEMA_signal_1099 ;
    wire new_AGEMA_signal_1100 ;
    wire new_AGEMA_signal_1101 ;
    wire new_AGEMA_signal_1102 ;
    wire new_AGEMA_signal_1103 ;
    wire new_AGEMA_signal_1104 ;
    wire new_AGEMA_signal_1105 ;
    wire new_AGEMA_signal_1106 ;
    wire new_AGEMA_signal_1107 ;
    wire new_AGEMA_signal_1108 ;
    wire new_AGEMA_signal_1109 ;
    wire new_AGEMA_signal_1110 ;
    wire new_AGEMA_signal_1111 ;
    wire new_AGEMA_signal_1112 ;
    wire new_AGEMA_signal_1113 ;
    wire new_AGEMA_signal_1114 ;
    wire new_AGEMA_signal_1115 ;
    wire new_AGEMA_signal_1116 ;
    wire new_AGEMA_signal_1117 ;
    wire new_AGEMA_signal_1118 ;
    wire new_AGEMA_signal_1119 ;
    wire new_AGEMA_signal_1120 ;
    wire new_AGEMA_signal_1121 ;
    wire new_AGEMA_signal_1122 ;
    wire new_AGEMA_signal_1123 ;
    wire new_AGEMA_signal_1124 ;
    wire new_AGEMA_signal_1125 ;
    wire new_AGEMA_signal_1126 ;
    wire new_AGEMA_signal_1127 ;
    wire new_AGEMA_signal_1128 ;
    wire new_AGEMA_signal_1129 ;
    wire new_AGEMA_signal_1130 ;
    wire new_AGEMA_signal_1131 ;
    wire new_AGEMA_signal_1132 ;
    wire new_AGEMA_signal_1133 ;
    wire new_AGEMA_signal_1134 ;
    wire new_AGEMA_signal_1135 ;
    wire new_AGEMA_signal_1136 ;
    wire new_AGEMA_signal_1137 ;
    wire new_AGEMA_signal_1138 ;
    wire new_AGEMA_signal_1139 ;
    wire new_AGEMA_signal_1140 ;
    wire new_AGEMA_signal_1141 ;
    wire new_AGEMA_signal_1142 ;
    wire new_AGEMA_signal_1143 ;
    wire new_AGEMA_signal_1144 ;
    wire new_AGEMA_signal_1145 ;
    wire new_AGEMA_signal_1146 ;
    wire new_AGEMA_signal_1147 ;
    wire new_AGEMA_signal_1148 ;
    wire new_AGEMA_signal_1149 ;
    wire new_AGEMA_signal_1150 ;
    wire new_AGEMA_signal_1151 ;
    wire new_AGEMA_signal_1152 ;
    wire new_AGEMA_signal_1153 ;
    wire new_AGEMA_signal_1154 ;
    wire new_AGEMA_signal_1155 ;
    wire new_AGEMA_signal_1156 ;
    wire new_AGEMA_signal_1157 ;
    wire new_AGEMA_signal_1158 ;
    wire new_AGEMA_signal_1159 ;
    wire new_AGEMA_signal_1160 ;
    wire new_AGEMA_signal_1161 ;
    wire new_AGEMA_signal_1162 ;
    wire new_AGEMA_signal_1163 ;
    wire new_AGEMA_signal_1164 ;
    wire new_AGEMA_signal_1165 ;
    wire new_AGEMA_signal_1166 ;
    wire new_AGEMA_signal_1167 ;
    wire new_AGEMA_signal_1168 ;
    wire new_AGEMA_signal_1169 ;
    wire new_AGEMA_signal_1170 ;
    wire new_AGEMA_signal_1171 ;
    wire new_AGEMA_signal_1172 ;
    wire new_AGEMA_signal_1173 ;
    wire new_AGEMA_signal_1174 ;
    wire new_AGEMA_signal_1175 ;
    wire new_AGEMA_signal_1176 ;
    wire new_AGEMA_signal_1177 ;
    wire new_AGEMA_signal_1178 ;
    wire new_AGEMA_signal_1179 ;
    wire new_AGEMA_signal_1180 ;
    wire new_AGEMA_signal_1181 ;
    wire new_AGEMA_signal_1182 ;
    wire new_AGEMA_signal_1183 ;
    wire new_AGEMA_signal_1184 ;
    wire new_AGEMA_signal_1185 ;
    wire new_AGEMA_signal_1186 ;
    wire new_AGEMA_signal_1187 ;
    wire new_AGEMA_signal_1188 ;
    wire new_AGEMA_signal_1189 ;
    wire new_AGEMA_signal_1190 ;
    wire new_AGEMA_signal_1191 ;
    wire new_AGEMA_signal_1192 ;
    wire new_AGEMA_signal_1193 ;
    wire new_AGEMA_signal_1194 ;
    wire new_AGEMA_signal_1195 ;
    wire new_AGEMA_signal_1196 ;
    wire new_AGEMA_signal_1197 ;
    wire new_AGEMA_signal_1198 ;
    wire new_AGEMA_signal_1199 ;
    wire new_AGEMA_signal_1200 ;
    wire new_AGEMA_signal_1201 ;
    wire new_AGEMA_signal_1202 ;
    wire new_AGEMA_signal_1203 ;
    wire new_AGEMA_signal_1204 ;
    wire new_AGEMA_signal_1205 ;
    wire new_AGEMA_signal_1206 ;
    wire new_AGEMA_signal_1207 ;
    wire new_AGEMA_signal_1208 ;
    wire new_AGEMA_signal_1209 ;
    wire new_AGEMA_signal_1210 ;
    wire new_AGEMA_signal_1211 ;
    wire new_AGEMA_signal_1212 ;
    wire new_AGEMA_signal_1213 ;
    wire new_AGEMA_signal_1214 ;
    wire new_AGEMA_signal_1215 ;
    wire new_AGEMA_signal_1216 ;
    wire new_AGEMA_signal_1217 ;
    wire new_AGEMA_signal_1218 ;
    wire new_AGEMA_signal_1219 ;
    wire new_AGEMA_signal_1220 ;
    wire new_AGEMA_signal_1221 ;
    wire new_AGEMA_signal_1222 ;
    wire new_AGEMA_signal_1223 ;
    wire new_AGEMA_signal_1224 ;
    wire new_AGEMA_signal_1225 ;
    wire new_AGEMA_signal_1226 ;
    wire new_AGEMA_signal_1227 ;
    wire new_AGEMA_signal_1228 ;
    wire new_AGEMA_signal_1229 ;
    wire new_AGEMA_signal_1230 ;
    wire new_AGEMA_signal_1231 ;
    wire new_AGEMA_signal_1232 ;
    wire new_AGEMA_signal_1233 ;
    wire new_AGEMA_signal_1234 ;
    wire new_AGEMA_signal_1235 ;
    wire new_AGEMA_signal_1236 ;
    wire new_AGEMA_signal_1237 ;
    wire new_AGEMA_signal_1238 ;
    wire new_AGEMA_signal_1239 ;
    wire new_AGEMA_signal_1240 ;
    wire new_AGEMA_signal_1241 ;
    wire new_AGEMA_signal_1242 ;
    wire new_AGEMA_signal_1243 ;
    wire new_AGEMA_signal_1244 ;
    wire new_AGEMA_signal_1245 ;
    wire new_AGEMA_signal_1246 ;
    wire new_AGEMA_signal_1247 ;
    wire new_AGEMA_signal_1248 ;
    wire new_AGEMA_signal_1249 ;
    wire new_AGEMA_signal_1250 ;
    wire new_AGEMA_signal_1251 ;
    wire new_AGEMA_signal_1252 ;
    wire new_AGEMA_signal_1253 ;
    wire new_AGEMA_signal_1254 ;
    wire new_AGEMA_signal_1255 ;
    wire new_AGEMA_signal_1256 ;
    wire new_AGEMA_signal_1257 ;
    wire new_AGEMA_signal_1258 ;
    wire new_AGEMA_signal_1259 ;
    wire new_AGEMA_signal_1260 ;
    wire new_AGEMA_signal_1261 ;
    wire new_AGEMA_signal_1262 ;
    wire new_AGEMA_signal_1263 ;
    wire new_AGEMA_signal_1264 ;
    wire new_AGEMA_signal_1265 ;
    wire new_AGEMA_signal_1266 ;
    wire new_AGEMA_signal_1267 ;
    wire new_AGEMA_signal_1268 ;
    wire new_AGEMA_signal_1269 ;
    wire new_AGEMA_signal_1270 ;
    wire new_AGEMA_signal_1271 ;
    wire new_AGEMA_signal_1272 ;
    wire new_AGEMA_signal_1273 ;
    wire new_AGEMA_signal_1274 ;
    wire new_AGEMA_signal_1275 ;
    wire new_AGEMA_signal_1276 ;
    wire new_AGEMA_signal_1277 ;
    wire new_AGEMA_signal_1278 ;
    wire new_AGEMA_signal_1279 ;
    wire new_AGEMA_signal_1280 ;
    wire new_AGEMA_signal_1281 ;
    wire new_AGEMA_signal_1282 ;
    wire new_AGEMA_signal_1283 ;
    wire new_AGEMA_signal_1284 ;
    wire new_AGEMA_signal_1285 ;
    wire new_AGEMA_signal_1286 ;
    wire new_AGEMA_signal_1287 ;
    wire new_AGEMA_signal_1288 ;
    wire new_AGEMA_signal_1289 ;
    wire new_AGEMA_signal_1290 ;
    wire new_AGEMA_signal_1291 ;
    wire new_AGEMA_signal_1292 ;
    wire new_AGEMA_signal_1293 ;
    wire new_AGEMA_signal_1294 ;
    wire new_AGEMA_signal_1295 ;
    wire new_AGEMA_signal_1296 ;
    wire new_AGEMA_signal_1297 ;
    wire new_AGEMA_signal_1298 ;
    wire new_AGEMA_signal_1299 ;
    wire new_AGEMA_signal_1300 ;
    wire new_AGEMA_signal_1301 ;
    wire new_AGEMA_signal_1302 ;
    wire new_AGEMA_signal_1303 ;
    wire new_AGEMA_signal_1304 ;
    wire new_AGEMA_signal_1305 ;
    wire new_AGEMA_signal_1306 ;
    wire new_AGEMA_signal_1307 ;
    wire new_AGEMA_signal_1308 ;
    wire new_AGEMA_signal_1309 ;
    wire new_AGEMA_signal_1310 ;
    wire new_AGEMA_signal_1311 ;
    wire new_AGEMA_signal_1312 ;
    wire new_AGEMA_signal_1313 ;
    wire new_AGEMA_signal_1314 ;
    wire new_AGEMA_signal_1315 ;
    wire new_AGEMA_signal_1316 ;
    wire new_AGEMA_signal_1317 ;
    wire new_AGEMA_signal_1318 ;
    wire new_AGEMA_signal_1319 ;
    wire new_AGEMA_signal_1320 ;
    wire new_AGEMA_signal_1321 ;
    wire new_AGEMA_signal_1322 ;
    wire new_AGEMA_signal_1323 ;
    wire new_AGEMA_signal_1324 ;
    wire new_AGEMA_signal_1325 ;
    wire new_AGEMA_signal_1326 ;
    wire new_AGEMA_signal_1327 ;
    wire new_AGEMA_signal_1328 ;
    wire new_AGEMA_signal_1329 ;
    wire new_AGEMA_signal_1330 ;
    wire new_AGEMA_signal_1331 ;
    wire new_AGEMA_signal_1332 ;
    wire new_AGEMA_signal_1333 ;
    wire new_AGEMA_signal_1334 ;
    wire new_AGEMA_signal_1335 ;
    wire new_AGEMA_signal_1336 ;
    wire new_AGEMA_signal_1337 ;
    wire new_AGEMA_signal_1338 ;
    wire new_AGEMA_signal_1339 ;
    wire new_AGEMA_signal_1340 ;
    wire new_AGEMA_signal_1341 ;
    wire new_AGEMA_signal_1342 ;
    wire new_AGEMA_signal_1343 ;
    wire new_AGEMA_signal_1344 ;
    wire new_AGEMA_signal_1345 ;
    wire new_AGEMA_signal_1346 ;
    wire new_AGEMA_signal_1347 ;
    wire new_AGEMA_signal_1348 ;
    wire new_AGEMA_signal_1349 ;
    wire new_AGEMA_signal_1350 ;
    wire new_AGEMA_signal_1351 ;
    wire new_AGEMA_signal_1352 ;
    wire new_AGEMA_signal_1353 ;
    wire new_AGEMA_signal_1354 ;
    wire new_AGEMA_signal_1355 ;
    wire new_AGEMA_signal_1356 ;
    wire new_AGEMA_signal_1357 ;
    wire new_AGEMA_signal_1358 ;
    wire new_AGEMA_signal_1359 ;
    wire new_AGEMA_signal_1360 ;
    wire new_AGEMA_signal_1361 ;

    /* cells in depth 0 */
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \M1.gen_loop_0__M.X1.U1 ( .A0_t (value_in_s0_t[0]), .A0_f (value_in_s0_f[0]), .A1_t (value_in_s1_t[0]), .A1_f (value_in_s1_f[0]), .B0_t (value_out_s0_t[0]), .B0_f (value_out_s0_f[0]), .B1_t (value_out_s1_t[0]), .B1_f (value_out_s1_f[0]), .Z0_t (\M1.gen_loop_0__M.X ), .Z0_f (new_AGEMA_signal_864), .Z1_t (new_AGEMA_signal_865), .Z1_f (new_AGEMA_signal_866) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \M1.gen_loop_0__M.A.U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (Inc_out[3]), .A1_f (new_AGEMA_signal_953), .B0_t (\M1.gen_loop_0__M.X ), .B0_f (new_AGEMA_signal_864), .B1_t (new_AGEMA_signal_865), .B1_f (new_AGEMA_signal_866), .Z0_t (\M1.gen_loop_0__M.Y ), .Z0_f (new_AGEMA_signal_954), .Z1_t (new_AGEMA_signal_955), .Z1_f (new_AGEMA_signal_956) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \M1.gen_loop_0__M.X2.U1 ( .A0_t (\M1.gen_loop_0__M.Y ), .A0_f (new_AGEMA_signal_954), .A1_t (new_AGEMA_signal_955), .A1_f (new_AGEMA_signal_956), .B0_t (value_in_s0_t[0]), .B0_f (value_in_s0_f[0]), .B1_t (value_in_s1_t[0]), .B1_f (value_in_s1_f[0]), .Z0_t (Sbox_in[0]), .Z0_f (new_AGEMA_signal_978), .Z1_t (new_AGEMA_signal_979), .Z1_f (new_AGEMA_signal_980) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \M1.gen_loop_1__M.X1.U1 ( .A0_t (value_in_s0_t[1]), .A0_f (value_in_s0_f[1]), .A1_t (value_in_s1_t[1]), .A1_f (value_in_s1_f[1]), .B0_t (value_out_s0_t[1]), .B0_f (value_out_s0_f[1]), .B1_t (value_out_s1_t[1]), .B1_f (value_out_s1_f[1]), .Z0_t (\M1.gen_loop_1__M.X ), .Z0_f (new_AGEMA_signal_873), .Z1_t (new_AGEMA_signal_874), .Z1_f (new_AGEMA_signal_875) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \M1.gen_loop_1__M.A.U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (Inc_out[3]), .A1_f (new_AGEMA_signal_953), .B0_t (\M1.gen_loop_1__M.X ), .B0_f (new_AGEMA_signal_873), .B1_t (new_AGEMA_signal_874), .B1_f (new_AGEMA_signal_875), .Z0_t (\M1.gen_loop_1__M.Y ), .Z0_f (new_AGEMA_signal_957), .Z1_t (new_AGEMA_signal_958), .Z1_f (new_AGEMA_signal_959) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \M1.gen_loop_1__M.X2.U1 ( .A0_t (\M1.gen_loop_1__M.Y ), .A0_f (new_AGEMA_signal_957), .A1_t (new_AGEMA_signal_958), .A1_f (new_AGEMA_signal_959), .B0_t (value_in_s0_t[1]), .B0_f (value_in_s0_f[1]), .B1_t (value_in_s1_t[1]), .B1_f (value_in_s1_f[1]), .Z0_t (Sbox_in[1]), .Z0_f (new_AGEMA_signal_981), .Z1_t (new_AGEMA_signal_982), .Z1_f (new_AGEMA_signal_983) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \M1.gen_loop_2__M.X1.U1 ( .A0_t (value_in_s0_t[2]), .A0_f (value_in_s0_f[2]), .A1_t (value_in_s1_t[2]), .A1_f (value_in_s1_f[2]), .B0_t (value_out_s0_t[2]), .B0_f (value_out_s0_f[2]), .B1_t (value_out_s1_t[2]), .B1_f (value_out_s1_f[2]), .Z0_t (\M1.gen_loop_2__M.X ), .Z0_f (new_AGEMA_signal_882), .Z1_t (new_AGEMA_signal_883), .Z1_f (new_AGEMA_signal_884) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \M1.gen_loop_2__M.A.U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (Inc_out[3]), .A1_f (new_AGEMA_signal_953), .B0_t (\M1.gen_loop_2__M.X ), .B0_f (new_AGEMA_signal_882), .B1_t (new_AGEMA_signal_883), .B1_f (new_AGEMA_signal_884), .Z0_t (\M1.gen_loop_2__M.Y ), .Z0_f (new_AGEMA_signal_960), .Z1_t (new_AGEMA_signal_961), .Z1_f (new_AGEMA_signal_962) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \M1.gen_loop_2__M.X2.U1 ( .A0_t (\M1.gen_loop_2__M.Y ), .A0_f (new_AGEMA_signal_960), .A1_t (new_AGEMA_signal_961), .A1_f (new_AGEMA_signal_962), .B0_t (value_in_s0_t[2]), .B0_f (value_in_s0_f[2]), .B1_t (value_in_s1_t[2]), .B1_f (value_in_s1_f[2]), .Z0_t (Sbox_in[2]), .Z0_f (new_AGEMA_signal_984), .Z1_t (new_AGEMA_signal_985), .Z1_f (new_AGEMA_signal_986) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \M1.gen_loop_3__M.X1.U1 ( .A0_t (value_in_s0_t[3]), .A0_f (value_in_s0_f[3]), .A1_t (value_in_s1_t[3]), .A1_f (value_in_s1_f[3]), .B0_t (value_out_s0_t[3]), .B0_f (value_out_s0_f[3]), .B1_t (value_out_s1_t[3]), .B1_f (value_out_s1_f[3]), .Z0_t (\M1.gen_loop_3__M.X ), .Z0_f (new_AGEMA_signal_891), .Z1_t (new_AGEMA_signal_892), .Z1_f (new_AGEMA_signal_893) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \M1.gen_loop_3__M.A.U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (Inc_out[3]), .A1_f (new_AGEMA_signal_953), .B0_t (\M1.gen_loop_3__M.X ), .B0_f (new_AGEMA_signal_891), .B1_t (new_AGEMA_signal_892), .B1_f (new_AGEMA_signal_893), .Z0_t (\M1.gen_loop_3__M.Y ), .Z0_f (new_AGEMA_signal_963), .Z1_t (new_AGEMA_signal_964), .Z1_f (new_AGEMA_signal_965) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \M1.gen_loop_3__M.X2.U1 ( .A0_t (\M1.gen_loop_3__M.Y ), .A0_f (new_AGEMA_signal_963), .A1_t (new_AGEMA_signal_964), .A1_f (new_AGEMA_signal_965), .B0_t (value_in_s0_t[3]), .B0_f (value_in_s0_f[3]), .B1_t (value_in_s1_t[3]), .B1_f (value_in_s1_f[3]), .Z0_t (Sbox_in[3]), .Z0_f (new_AGEMA_signal_987), .Z1_t (new_AGEMA_signal_988), .Z1_f (new_AGEMA_signal_989) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \M1.gen_loop_4__M.X1.U1 ( .A0_t (value_in_s0_t[4]), .A0_f (value_in_s0_f[4]), .A1_t (value_in_s1_t[4]), .A1_f (value_in_s1_f[4]), .B0_t (value_out_s0_t[4]), .B0_f (value_out_s0_f[4]), .B1_t (value_out_s1_t[4]), .B1_f (value_out_s1_f[4]), .Z0_t (\M1.gen_loop_4__M.X ), .Z0_f (new_AGEMA_signal_900), .Z1_t (new_AGEMA_signal_901), .Z1_f (new_AGEMA_signal_902) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \M1.gen_loop_4__M.A.U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (Inc_out[3]), .A1_f (new_AGEMA_signal_953), .B0_t (\M1.gen_loop_4__M.X ), .B0_f (new_AGEMA_signal_900), .B1_t (new_AGEMA_signal_901), .B1_f (new_AGEMA_signal_902), .Z0_t (\M1.gen_loop_4__M.Y ), .Z0_f (new_AGEMA_signal_966), .Z1_t (new_AGEMA_signal_967), .Z1_f (new_AGEMA_signal_968) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \M1.gen_loop_4__M.X2.U1 ( .A0_t (\M1.gen_loop_4__M.Y ), .A0_f (new_AGEMA_signal_966), .A1_t (new_AGEMA_signal_967), .A1_f (new_AGEMA_signal_968), .B0_t (value_in_s0_t[4]), .B0_f (value_in_s0_f[4]), .B1_t (value_in_s1_t[4]), .B1_f (value_in_s1_f[4]), .Z0_t (Sbox_in[4]), .Z0_f (new_AGEMA_signal_990), .Z1_t (new_AGEMA_signal_991), .Z1_f (new_AGEMA_signal_992) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \M1.gen_loop_5__M.X1.U1 ( .A0_t (value_in_s0_t[5]), .A0_f (value_in_s0_f[5]), .A1_t (value_in_s1_t[5]), .A1_f (value_in_s1_f[5]), .B0_t (value_out_s0_t[5]), .B0_f (value_out_s0_f[5]), .B1_t (value_out_s1_t[5]), .B1_f (value_out_s1_f[5]), .Z0_t (\M1.gen_loop_5__M.X ), .Z0_f (new_AGEMA_signal_909), .Z1_t (new_AGEMA_signal_910), .Z1_f (new_AGEMA_signal_911) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \M1.gen_loop_5__M.A.U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (Inc_out[3]), .A1_f (new_AGEMA_signal_953), .B0_t (\M1.gen_loop_5__M.X ), .B0_f (new_AGEMA_signal_909), .B1_t (new_AGEMA_signal_910), .B1_f (new_AGEMA_signal_911), .Z0_t (\M1.gen_loop_5__M.Y ), .Z0_f (new_AGEMA_signal_969), .Z1_t (new_AGEMA_signal_970), .Z1_f (new_AGEMA_signal_971) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \M1.gen_loop_5__M.X2.U1 ( .A0_t (\M1.gen_loop_5__M.Y ), .A0_f (new_AGEMA_signal_969), .A1_t (new_AGEMA_signal_970), .A1_f (new_AGEMA_signal_971), .B0_t (value_in_s0_t[5]), .B0_f (value_in_s0_f[5]), .B1_t (value_in_s1_t[5]), .B1_f (value_in_s1_f[5]), .Z0_t (Sbox_in[5]), .Z0_f (new_AGEMA_signal_993), .Z1_t (new_AGEMA_signal_994), .Z1_f (new_AGEMA_signal_995) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \M1.gen_loop_6__M.X1.U1 ( .A0_t (value_in_s0_t[6]), .A0_f (value_in_s0_f[6]), .A1_t (value_in_s1_t[6]), .A1_f (value_in_s1_f[6]), .B0_t (value_out_s0_t[6]), .B0_f (value_out_s0_f[6]), .B1_t (value_out_s1_t[6]), .B1_f (value_out_s1_f[6]), .Z0_t (\M1.gen_loop_6__M.X ), .Z0_f (new_AGEMA_signal_918), .Z1_t (new_AGEMA_signal_919), .Z1_f (new_AGEMA_signal_920) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \M1.gen_loop_6__M.A.U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (Inc_out[3]), .A1_f (new_AGEMA_signal_953), .B0_t (\M1.gen_loop_6__M.X ), .B0_f (new_AGEMA_signal_918), .B1_t (new_AGEMA_signal_919), .B1_f (new_AGEMA_signal_920), .Z0_t (\M1.gen_loop_6__M.Y ), .Z0_f (new_AGEMA_signal_972), .Z1_t (new_AGEMA_signal_973), .Z1_f (new_AGEMA_signal_974) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \M1.gen_loop_6__M.X2.U1 ( .A0_t (\M1.gen_loop_6__M.Y ), .A0_f (new_AGEMA_signal_972), .A1_t (new_AGEMA_signal_973), .A1_f (new_AGEMA_signal_974), .B0_t (value_in_s0_t[6]), .B0_f (value_in_s0_f[6]), .B1_t (value_in_s1_t[6]), .B1_f (value_in_s1_f[6]), .Z0_t (Sbox_in[6]), .Z0_f (new_AGEMA_signal_996), .Z1_t (new_AGEMA_signal_997), .Z1_f (new_AGEMA_signal_998) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \M1.gen_loop_7__M.X1.U1 ( .A0_t (value_in_s0_t[7]), .A0_f (value_in_s0_f[7]), .A1_t (value_in_s1_t[7]), .A1_f (value_in_s1_f[7]), .B0_t (value_out_s0_t[7]), .B0_f (value_out_s0_f[7]), .B1_t (value_out_s1_t[7]), .B1_f (value_out_s1_f[7]), .Z0_t (\M1.gen_loop_7__M.X ), .Z0_f (new_AGEMA_signal_927), .Z1_t (new_AGEMA_signal_928), .Z1_f (new_AGEMA_signal_929) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \M1.gen_loop_7__M.A.U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (Inc_out[3]), .A1_f (new_AGEMA_signal_953), .B0_t (\M1.gen_loop_7__M.X ), .B0_f (new_AGEMA_signal_927), .B1_t (new_AGEMA_signal_928), .B1_f (new_AGEMA_signal_929), .Z0_t (\M1.gen_loop_7__M.Y ), .Z0_f (new_AGEMA_signal_975), .Z1_t (new_AGEMA_signal_976), .Z1_f (new_AGEMA_signal_977) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \M1.gen_loop_7__M.X2.U1 ( .A0_t (\M1.gen_loop_7__M.Y ), .A0_f (new_AGEMA_signal_975), .A1_t (new_AGEMA_signal_976), .A1_f (new_AGEMA_signal_977), .B0_t (value_in_s0_t[7]), .B0_f (value_in_s0_f[7]), .B1_t (value_in_s1_t[7]), .B1_f (value_in_s1_f[7]), .Z0_t (Sbox_in[7]), .Z0_f (new_AGEMA_signal_999), .Z1_t (new_AGEMA_signal_1000), .Z1_f (new_AGEMA_signal_1001) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_T1.U1 ( .A0_t (Sbox_in[7]), .A0_f (new_AGEMA_signal_999), .A1_t (new_AGEMA_signal_1000), .A1_f (new_AGEMA_signal_1001), .B0_t (Sbox_in[4]), .B0_f (new_AGEMA_signal_990), .B1_t (new_AGEMA_signal_991), .B1_f (new_AGEMA_signal_992), .Z0_t (\SboxInst.T1 ), .Z0_f (new_AGEMA_signal_1002), .Z1_t (new_AGEMA_signal_1003), .Z1_f (new_AGEMA_signal_1004) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_T2.U1 ( .A0_t (Sbox_in[7]), .A0_f (new_AGEMA_signal_999), .A1_t (new_AGEMA_signal_1000), .A1_f (new_AGEMA_signal_1001), .B0_t (Sbox_in[2]), .B0_f (new_AGEMA_signal_984), .B1_t (new_AGEMA_signal_985), .B1_f (new_AGEMA_signal_986), .Z0_t (\SboxInst.T2 ), .Z0_f (new_AGEMA_signal_1005), .Z1_t (new_AGEMA_signal_1006), .Z1_f (new_AGEMA_signal_1007) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_T3.U1 ( .A0_t (Sbox_in[7]), .A0_f (new_AGEMA_signal_999), .A1_t (new_AGEMA_signal_1000), .A1_f (new_AGEMA_signal_1001), .B0_t (Sbox_in[1]), .B0_f (new_AGEMA_signal_981), .B1_t (new_AGEMA_signal_982), .B1_f (new_AGEMA_signal_983), .Z0_t (\SboxInst.T3 ), .Z0_f (new_AGEMA_signal_1008), .Z1_t (new_AGEMA_signal_1009), .Z1_f (new_AGEMA_signal_1010) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_T4.U1 ( .A0_t (Sbox_in[4]), .A0_f (new_AGEMA_signal_990), .A1_t (new_AGEMA_signal_991), .A1_f (new_AGEMA_signal_992), .B0_t (Sbox_in[2]), .B0_f (new_AGEMA_signal_984), .B1_t (new_AGEMA_signal_985), .B1_f (new_AGEMA_signal_986), .Z0_t (\SboxInst.T4 ), .Z0_f (new_AGEMA_signal_1011), .Z1_t (new_AGEMA_signal_1012), .Z1_f (new_AGEMA_signal_1013) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_T5.U1 ( .A0_t (Sbox_in[3]), .A0_f (new_AGEMA_signal_987), .A1_t (new_AGEMA_signal_988), .A1_f (new_AGEMA_signal_989), .B0_t (Sbox_in[1]), .B0_f (new_AGEMA_signal_981), .B1_t (new_AGEMA_signal_982), .B1_f (new_AGEMA_signal_983), .Z0_t (\SboxInst.T5 ), .Z0_f (new_AGEMA_signal_1014), .Z1_t (new_AGEMA_signal_1015), .Z1_f (new_AGEMA_signal_1016) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_T6.U1 ( .A0_t (\SboxInst.T1 ), .A0_f (new_AGEMA_signal_1002), .A1_t (new_AGEMA_signal_1003), .A1_f (new_AGEMA_signal_1004), .B0_t (\SboxInst.T5 ), .B0_f (new_AGEMA_signal_1014), .B1_t (new_AGEMA_signal_1015), .B1_f (new_AGEMA_signal_1016), .Z0_t (\SboxInst.T6 ), .Z0_f (new_AGEMA_signal_1032), .Z1_t (new_AGEMA_signal_1033), .Z1_f (new_AGEMA_signal_1034) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_T7.U1 ( .A0_t (Sbox_in[6]), .A0_f (new_AGEMA_signal_996), .A1_t (new_AGEMA_signal_997), .A1_f (new_AGEMA_signal_998), .B0_t (Sbox_in[5]), .B0_f (new_AGEMA_signal_993), .B1_t (new_AGEMA_signal_994), .B1_f (new_AGEMA_signal_995), .Z0_t (\SboxInst.T7 ), .Z0_f (new_AGEMA_signal_1017), .Z1_t (new_AGEMA_signal_1018), .Z1_f (new_AGEMA_signal_1019) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_T8.U1 ( .A0_t (Sbox_in[0]), .A0_f (new_AGEMA_signal_978), .A1_t (new_AGEMA_signal_979), .A1_f (new_AGEMA_signal_980), .B0_t (\SboxInst.T6 ), .B0_f (new_AGEMA_signal_1032), .B1_t (new_AGEMA_signal_1033), .B1_f (new_AGEMA_signal_1034), .Z0_t (\SboxInst.T8 ), .Z0_f (new_AGEMA_signal_1056), .Z1_t (new_AGEMA_signal_1057), .Z1_f (new_AGEMA_signal_1058) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_T9.U1 ( .A0_t (Sbox_in[0]), .A0_f (new_AGEMA_signal_978), .A1_t (new_AGEMA_signal_979), .A1_f (new_AGEMA_signal_980), .B0_t (\SboxInst.T7 ), .B0_f (new_AGEMA_signal_1017), .B1_t (new_AGEMA_signal_1018), .B1_f (new_AGEMA_signal_1019), .Z0_t (\SboxInst.T9 ), .Z0_f (new_AGEMA_signal_1035), .Z1_t (new_AGEMA_signal_1036), .Z1_f (new_AGEMA_signal_1037) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_T10.U1 ( .A0_t (\SboxInst.T6 ), .A0_f (new_AGEMA_signal_1032), .A1_t (new_AGEMA_signal_1033), .A1_f (new_AGEMA_signal_1034), .B0_t (\SboxInst.T7 ), .B0_f (new_AGEMA_signal_1017), .B1_t (new_AGEMA_signal_1018), .B1_f (new_AGEMA_signal_1019), .Z0_t (\SboxInst.T10 ), .Z0_f (new_AGEMA_signal_1059), .Z1_t (new_AGEMA_signal_1060), .Z1_f (new_AGEMA_signal_1061) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_T11.U1 ( .A0_t (Sbox_in[6]), .A0_f (new_AGEMA_signal_996), .A1_t (new_AGEMA_signal_997), .A1_f (new_AGEMA_signal_998), .B0_t (Sbox_in[2]), .B0_f (new_AGEMA_signal_984), .B1_t (new_AGEMA_signal_985), .B1_f (new_AGEMA_signal_986), .Z0_t (\SboxInst.T11 ), .Z0_f (new_AGEMA_signal_1020), .Z1_t (new_AGEMA_signal_1021), .Z1_f (new_AGEMA_signal_1022) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_T12.U1 ( .A0_t (Sbox_in[5]), .A0_f (new_AGEMA_signal_993), .A1_t (new_AGEMA_signal_994), .A1_f (new_AGEMA_signal_995), .B0_t (Sbox_in[2]), .B0_f (new_AGEMA_signal_984), .B1_t (new_AGEMA_signal_985), .B1_f (new_AGEMA_signal_986), .Z0_t (\SboxInst.T12 ), .Z0_f (new_AGEMA_signal_1023), .Z1_t (new_AGEMA_signal_1024), .Z1_f (new_AGEMA_signal_1025) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_T13.U1 ( .A0_t (\SboxInst.T3 ), .A0_f (new_AGEMA_signal_1008), .A1_t (new_AGEMA_signal_1009), .A1_f (new_AGEMA_signal_1010), .B0_t (\SboxInst.T4 ), .B0_f (new_AGEMA_signal_1011), .B1_t (new_AGEMA_signal_1012), .B1_f (new_AGEMA_signal_1013), .Z0_t (\SboxInst.T13 ), .Z0_f (new_AGEMA_signal_1038), .Z1_t (new_AGEMA_signal_1039), .Z1_f (new_AGEMA_signal_1040) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_T14.U1 ( .A0_t (\SboxInst.T6 ), .A0_f (new_AGEMA_signal_1032), .A1_t (new_AGEMA_signal_1033), .A1_f (new_AGEMA_signal_1034), .B0_t (\SboxInst.T11 ), .B0_f (new_AGEMA_signal_1020), .B1_t (new_AGEMA_signal_1021), .B1_f (new_AGEMA_signal_1022), .Z0_t (\SboxInst.T14 ), .Z0_f (new_AGEMA_signal_1062), .Z1_t (new_AGEMA_signal_1063), .Z1_f (new_AGEMA_signal_1064) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_T15.U1 ( .A0_t (\SboxInst.T5 ), .A0_f (new_AGEMA_signal_1014), .A1_t (new_AGEMA_signal_1015), .A1_f (new_AGEMA_signal_1016), .B0_t (\SboxInst.T11 ), .B0_f (new_AGEMA_signal_1020), .B1_t (new_AGEMA_signal_1021), .B1_f (new_AGEMA_signal_1022), .Z0_t (\SboxInst.T15 ), .Z0_f (new_AGEMA_signal_1041), .Z1_t (new_AGEMA_signal_1042), .Z1_f (new_AGEMA_signal_1043) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_T16.U1 ( .A0_t (\SboxInst.T5 ), .A0_f (new_AGEMA_signal_1014), .A1_t (new_AGEMA_signal_1015), .A1_f (new_AGEMA_signal_1016), .B0_t (\SboxInst.T12 ), .B0_f (new_AGEMA_signal_1023), .B1_t (new_AGEMA_signal_1024), .B1_f (new_AGEMA_signal_1025), .Z0_t (\SboxInst.T16 ), .Z0_f (new_AGEMA_signal_1044), .Z1_t (new_AGEMA_signal_1045), .Z1_f (new_AGEMA_signal_1046) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_T17.U1 ( .A0_t (\SboxInst.T9 ), .A0_f (new_AGEMA_signal_1035), .A1_t (new_AGEMA_signal_1036), .A1_f (new_AGEMA_signal_1037), .B0_t (\SboxInst.T16 ), .B0_f (new_AGEMA_signal_1044), .B1_t (new_AGEMA_signal_1045), .B1_f (new_AGEMA_signal_1046), .Z0_t (\SboxInst.T17 ), .Z0_f (new_AGEMA_signal_1065), .Z1_t (new_AGEMA_signal_1066), .Z1_f (new_AGEMA_signal_1067) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_T18.U1 ( .A0_t (Sbox_in[4]), .A0_f (new_AGEMA_signal_990), .A1_t (new_AGEMA_signal_991), .A1_f (new_AGEMA_signal_992), .B0_t (Sbox_in[0]), .B0_f (new_AGEMA_signal_978), .B1_t (new_AGEMA_signal_979), .B1_f (new_AGEMA_signal_980), .Z0_t (\SboxInst.T18 ), .Z0_f (new_AGEMA_signal_1026), .Z1_t (new_AGEMA_signal_1027), .Z1_f (new_AGEMA_signal_1028) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_T19.U1 ( .A0_t (\SboxInst.T7 ), .A0_f (new_AGEMA_signal_1017), .A1_t (new_AGEMA_signal_1018), .A1_f (new_AGEMA_signal_1019), .B0_t (\SboxInst.T18 ), .B0_f (new_AGEMA_signal_1026), .B1_t (new_AGEMA_signal_1027), .B1_f (new_AGEMA_signal_1028), .Z0_t (\SboxInst.T19 ), .Z0_f (new_AGEMA_signal_1047), .Z1_t (new_AGEMA_signal_1048), .Z1_f (new_AGEMA_signal_1049) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_T20.U1 ( .A0_t (\SboxInst.T1 ), .A0_f (new_AGEMA_signal_1002), .A1_t (new_AGEMA_signal_1003), .A1_f (new_AGEMA_signal_1004), .B0_t (\SboxInst.T19 ), .B0_f (new_AGEMA_signal_1047), .B1_t (new_AGEMA_signal_1048), .B1_f (new_AGEMA_signal_1049), .Z0_t (\SboxInst.T20 ), .Z0_f (new_AGEMA_signal_1068), .Z1_t (new_AGEMA_signal_1069), .Z1_f (new_AGEMA_signal_1070) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_T21.U1 ( .A0_t (Sbox_in[1]), .A0_f (new_AGEMA_signal_981), .A1_t (new_AGEMA_signal_982), .A1_f (new_AGEMA_signal_983), .B0_t (Sbox_in[0]), .B0_f (new_AGEMA_signal_978), .B1_t (new_AGEMA_signal_979), .B1_f (new_AGEMA_signal_980), .Z0_t (\SboxInst.T21 ), .Z0_f (new_AGEMA_signal_1029), .Z1_t (new_AGEMA_signal_1030), .Z1_f (new_AGEMA_signal_1031) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_T22.U1 ( .A0_t (\SboxInst.T7 ), .A0_f (new_AGEMA_signal_1017), .A1_t (new_AGEMA_signal_1018), .A1_f (new_AGEMA_signal_1019), .B0_t (\SboxInst.T21 ), .B0_f (new_AGEMA_signal_1029), .B1_t (new_AGEMA_signal_1030), .B1_f (new_AGEMA_signal_1031), .Z0_t (\SboxInst.T22 ), .Z0_f (new_AGEMA_signal_1050), .Z1_t (new_AGEMA_signal_1051), .Z1_f (new_AGEMA_signal_1052) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_T23.U1 ( .A0_t (\SboxInst.T2 ), .A0_f (new_AGEMA_signal_1005), .A1_t (new_AGEMA_signal_1006), .A1_f (new_AGEMA_signal_1007), .B0_t (\SboxInst.T22 ), .B0_f (new_AGEMA_signal_1050), .B1_t (new_AGEMA_signal_1051), .B1_f (new_AGEMA_signal_1052), .Z0_t (\SboxInst.T23 ), .Z0_f (new_AGEMA_signal_1071), .Z1_t (new_AGEMA_signal_1072), .Z1_f (new_AGEMA_signal_1073) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_T24.U1 ( .A0_t (\SboxInst.T2 ), .A0_f (new_AGEMA_signal_1005), .A1_t (new_AGEMA_signal_1006), .A1_f (new_AGEMA_signal_1007), .B0_t (\SboxInst.T10 ), .B0_f (new_AGEMA_signal_1059), .B1_t (new_AGEMA_signal_1060), .B1_f (new_AGEMA_signal_1061), .Z0_t (\SboxInst.T24 ), .Z0_f (new_AGEMA_signal_1095), .Z1_t (new_AGEMA_signal_1096), .Z1_f (new_AGEMA_signal_1097) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_T25.U1 ( .A0_t (\SboxInst.T20 ), .A0_f (new_AGEMA_signal_1068), .A1_t (new_AGEMA_signal_1069), .A1_f (new_AGEMA_signal_1070), .B0_t (\SboxInst.T17 ), .B0_f (new_AGEMA_signal_1065), .B1_t (new_AGEMA_signal_1066), .B1_f (new_AGEMA_signal_1067), .Z0_t (\SboxInst.T25 ), .Z0_f (new_AGEMA_signal_1098), .Z1_t (new_AGEMA_signal_1099), .Z1_f (new_AGEMA_signal_1100) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_T26.U1 ( .A0_t (\SboxInst.T3 ), .A0_f (new_AGEMA_signal_1008), .A1_t (new_AGEMA_signal_1009), .A1_f (new_AGEMA_signal_1010), .B0_t (\SboxInst.T16 ), .B0_f (new_AGEMA_signal_1044), .B1_t (new_AGEMA_signal_1045), .B1_f (new_AGEMA_signal_1046), .Z0_t (\SboxInst.T26 ), .Z0_f (new_AGEMA_signal_1074), .Z1_t (new_AGEMA_signal_1075), .Z1_f (new_AGEMA_signal_1076) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_T27.U1 ( .A0_t (\SboxInst.T1 ), .A0_f (new_AGEMA_signal_1002), .A1_t (new_AGEMA_signal_1003), .A1_f (new_AGEMA_signal_1004), .B0_t (\SboxInst.T12 ), .B0_f (new_AGEMA_signal_1023), .B1_t (new_AGEMA_signal_1024), .B1_f (new_AGEMA_signal_1025), .Z0_t (\SboxInst.T27 ), .Z0_f (new_AGEMA_signal_1053), .Z1_t (new_AGEMA_signal_1054), .Z1_f (new_AGEMA_signal_1055) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M1.U1 ( .A0_t (\SboxInst.T13 ), .A0_f (new_AGEMA_signal_1038), .A1_t (new_AGEMA_signal_1039), .A1_f (new_AGEMA_signal_1040), .B0_t (\SboxInst.T6 ), .B0_f (new_AGEMA_signal_1032), .B1_t (new_AGEMA_signal_1033), .B1_f (new_AGEMA_signal_1034), .Z0_t (\SboxInst.M1 ), .Z0_f (new_AGEMA_signal_1077), .Z1_t (new_AGEMA_signal_1078), .Z1_f (new_AGEMA_signal_1079) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M2.U1 ( .A0_t (\SboxInst.T23 ), .A0_f (new_AGEMA_signal_1071), .A1_t (new_AGEMA_signal_1072), .A1_f (new_AGEMA_signal_1073), .B0_t (\SboxInst.T8 ), .B0_f (new_AGEMA_signal_1056), .B1_t (new_AGEMA_signal_1057), .B1_f (new_AGEMA_signal_1058), .Z0_t (\SboxInst.M2 ), .Z0_f (new_AGEMA_signal_1101), .Z1_t (new_AGEMA_signal_1102), .Z1_f (new_AGEMA_signal_1103) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_M3.U1 ( .A0_t (\SboxInst.T14 ), .A0_f (new_AGEMA_signal_1062), .A1_t (new_AGEMA_signal_1063), .A1_f (new_AGEMA_signal_1064), .B0_t (\SboxInst.M1 ), .B0_f (new_AGEMA_signal_1077), .B1_t (new_AGEMA_signal_1078), .B1_f (new_AGEMA_signal_1079), .Z0_t (\SboxInst.M3 ), .Z0_f (new_AGEMA_signal_1104), .Z1_t (new_AGEMA_signal_1105), .Z1_f (new_AGEMA_signal_1106) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M4.U1 ( .A0_t (\SboxInst.T19 ), .A0_f (new_AGEMA_signal_1047), .A1_t (new_AGEMA_signal_1048), .A1_f (new_AGEMA_signal_1049), .B0_t (Sbox_in[0]), .B0_f (new_AGEMA_signal_978), .B1_t (new_AGEMA_signal_979), .B1_f (new_AGEMA_signal_980), .Z0_t (\SboxInst.M4 ), .Z0_f (new_AGEMA_signal_1080), .Z1_t (new_AGEMA_signal_1081), .Z1_f (new_AGEMA_signal_1082) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_M5.U1 ( .A0_t (\SboxInst.M4 ), .A0_f (new_AGEMA_signal_1080), .A1_t (new_AGEMA_signal_1081), .A1_f (new_AGEMA_signal_1082), .B0_t (\SboxInst.M1 ), .B0_f (new_AGEMA_signal_1077), .B1_t (new_AGEMA_signal_1078), .B1_f (new_AGEMA_signal_1079), .Z0_t (\SboxInst.M5 ), .Z0_f (new_AGEMA_signal_1107), .Z1_t (new_AGEMA_signal_1108), .Z1_f (new_AGEMA_signal_1109) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M6.U1 ( .A0_t (\SboxInst.T3 ), .A0_f (new_AGEMA_signal_1008), .A1_t (new_AGEMA_signal_1009), .A1_f (new_AGEMA_signal_1010), .B0_t (\SboxInst.T16 ), .B0_f (new_AGEMA_signal_1044), .B1_t (new_AGEMA_signal_1045), .B1_f (new_AGEMA_signal_1046), .Z0_t (\SboxInst.M6 ), .Z0_f (new_AGEMA_signal_1083), .Z1_t (new_AGEMA_signal_1084), .Z1_f (new_AGEMA_signal_1085) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M7.U1 ( .A0_t (\SboxInst.T22 ), .A0_f (new_AGEMA_signal_1050), .A1_t (new_AGEMA_signal_1051), .A1_f (new_AGEMA_signal_1052), .B0_t (\SboxInst.T9 ), .B0_f (new_AGEMA_signal_1035), .B1_t (new_AGEMA_signal_1036), .B1_f (new_AGEMA_signal_1037), .Z0_t (\SboxInst.M7 ), .Z0_f (new_AGEMA_signal_1086), .Z1_t (new_AGEMA_signal_1087), .Z1_f (new_AGEMA_signal_1088) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_M8.U1 ( .A0_t (\SboxInst.T26 ), .A0_f (new_AGEMA_signal_1074), .A1_t (new_AGEMA_signal_1075), .A1_f (new_AGEMA_signal_1076), .B0_t (\SboxInst.M6 ), .B0_f (new_AGEMA_signal_1083), .B1_t (new_AGEMA_signal_1084), .B1_f (new_AGEMA_signal_1085), .Z0_t (\SboxInst.M8 ), .Z0_f (new_AGEMA_signal_1110), .Z1_t (new_AGEMA_signal_1111), .Z1_f (new_AGEMA_signal_1112) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M9.U1 ( .A0_t (\SboxInst.T20 ), .A0_f (new_AGEMA_signal_1068), .A1_t (new_AGEMA_signal_1069), .A1_f (new_AGEMA_signal_1070), .B0_t (\SboxInst.T17 ), .B0_f (new_AGEMA_signal_1065), .B1_t (new_AGEMA_signal_1066), .B1_f (new_AGEMA_signal_1067), .Z0_t (\SboxInst.M9 ), .Z0_f (new_AGEMA_signal_1113), .Z1_t (new_AGEMA_signal_1114), .Z1_f (new_AGEMA_signal_1115) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_M10.U1 ( .A0_t (\SboxInst.M9 ), .A0_f (new_AGEMA_signal_1113), .A1_t (new_AGEMA_signal_1114), .A1_f (new_AGEMA_signal_1115), .B0_t (\SboxInst.M6 ), .B0_f (new_AGEMA_signal_1083), .B1_t (new_AGEMA_signal_1084), .B1_f (new_AGEMA_signal_1085), .Z0_t (\SboxInst.M10 ), .Z0_f (new_AGEMA_signal_1122), .Z1_t (new_AGEMA_signal_1123), .Z1_f (new_AGEMA_signal_1124) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M11.U1 ( .A0_t (\SboxInst.T1 ), .A0_f (new_AGEMA_signal_1002), .A1_t (new_AGEMA_signal_1003), .A1_f (new_AGEMA_signal_1004), .B0_t (\SboxInst.T15 ), .B0_f (new_AGEMA_signal_1041), .B1_t (new_AGEMA_signal_1042), .B1_f (new_AGEMA_signal_1043), .Z0_t (\SboxInst.M11 ), .Z0_f (new_AGEMA_signal_1089), .Z1_t (new_AGEMA_signal_1090), .Z1_f (new_AGEMA_signal_1091) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M12.U1 ( .A0_t (\SboxInst.T4 ), .A0_f (new_AGEMA_signal_1011), .A1_t (new_AGEMA_signal_1012), .A1_f (new_AGEMA_signal_1013), .B0_t (\SboxInst.T27 ), .B0_f (new_AGEMA_signal_1053), .B1_t (new_AGEMA_signal_1054), .B1_f (new_AGEMA_signal_1055), .Z0_t (\SboxInst.M12 ), .Z0_f (new_AGEMA_signal_1092), .Z1_t (new_AGEMA_signal_1093), .Z1_f (new_AGEMA_signal_1094) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_M13.U1 ( .A0_t (\SboxInst.M12 ), .A0_f (new_AGEMA_signal_1092), .A1_t (new_AGEMA_signal_1093), .A1_f (new_AGEMA_signal_1094), .B0_t (\SboxInst.M11 ), .B0_f (new_AGEMA_signal_1089), .B1_t (new_AGEMA_signal_1090), .B1_f (new_AGEMA_signal_1091), .Z0_t (\SboxInst.M13 ), .Z0_f (new_AGEMA_signal_1116), .Z1_t (new_AGEMA_signal_1117), .Z1_f (new_AGEMA_signal_1118) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M14.U1 ( .A0_t (\SboxInst.T2 ), .A0_f (new_AGEMA_signal_1005), .A1_t (new_AGEMA_signal_1006), .A1_f (new_AGEMA_signal_1007), .B0_t (\SboxInst.T10 ), .B0_f (new_AGEMA_signal_1059), .B1_t (new_AGEMA_signal_1060), .B1_f (new_AGEMA_signal_1061), .Z0_t (\SboxInst.M14 ), .Z0_f (new_AGEMA_signal_1119), .Z1_t (new_AGEMA_signal_1120), .Z1_f (new_AGEMA_signal_1121) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_M15.U1 ( .A0_t (\SboxInst.M14 ), .A0_f (new_AGEMA_signal_1119), .A1_t (new_AGEMA_signal_1120), .A1_f (new_AGEMA_signal_1121), .B0_t (\SboxInst.M11 ), .B0_f (new_AGEMA_signal_1089), .B1_t (new_AGEMA_signal_1090), .B1_f (new_AGEMA_signal_1091), .Z0_t (\SboxInst.M15 ), .Z0_f (new_AGEMA_signal_1125), .Z1_t (new_AGEMA_signal_1126), .Z1_f (new_AGEMA_signal_1127) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_M16.U1 ( .A0_t (\SboxInst.M3 ), .A0_f (new_AGEMA_signal_1104), .A1_t (new_AGEMA_signal_1105), .A1_f (new_AGEMA_signal_1106), .B0_t (\SboxInst.M2 ), .B0_f (new_AGEMA_signal_1101), .B1_t (new_AGEMA_signal_1102), .B1_f (new_AGEMA_signal_1103), .Z0_t (\SboxInst.M16 ), .Z0_f (new_AGEMA_signal_1128), .Z1_t (new_AGEMA_signal_1129), .Z1_f (new_AGEMA_signal_1130) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_M17.U1 ( .A0_t (\SboxInst.M5 ), .A0_f (new_AGEMA_signal_1107), .A1_t (new_AGEMA_signal_1108), .A1_f (new_AGEMA_signal_1109), .B0_t (\SboxInst.T24 ), .B0_f (new_AGEMA_signal_1095), .B1_t (new_AGEMA_signal_1096), .B1_f (new_AGEMA_signal_1097), .Z0_t (\SboxInst.M17 ), .Z0_f (new_AGEMA_signal_1131), .Z1_t (new_AGEMA_signal_1132), .Z1_f (new_AGEMA_signal_1133) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_M18.U1 ( .A0_t (\SboxInst.M8 ), .A0_f (new_AGEMA_signal_1110), .A1_t (new_AGEMA_signal_1111), .A1_f (new_AGEMA_signal_1112), .B0_t (\SboxInst.M7 ), .B0_f (new_AGEMA_signal_1086), .B1_t (new_AGEMA_signal_1087), .B1_f (new_AGEMA_signal_1088), .Z0_t (\SboxInst.M18 ), .Z0_f (new_AGEMA_signal_1134), .Z1_t (new_AGEMA_signal_1135), .Z1_f (new_AGEMA_signal_1136) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_M19.U1 ( .A0_t (\SboxInst.M10 ), .A0_f (new_AGEMA_signal_1122), .A1_t (new_AGEMA_signal_1123), .A1_f (new_AGEMA_signal_1124), .B0_t (\SboxInst.M15 ), .B0_f (new_AGEMA_signal_1125), .B1_t (new_AGEMA_signal_1126), .B1_f (new_AGEMA_signal_1127), .Z0_t (\SboxInst.M19 ), .Z0_f (new_AGEMA_signal_1137), .Z1_t (new_AGEMA_signal_1138), .Z1_f (new_AGEMA_signal_1139) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_M20.U1 ( .A0_t (\SboxInst.M16 ), .A0_f (new_AGEMA_signal_1128), .A1_t (new_AGEMA_signal_1129), .A1_f (new_AGEMA_signal_1130), .B0_t (\SboxInst.M13 ), .B0_f (new_AGEMA_signal_1116), .B1_t (new_AGEMA_signal_1117), .B1_f (new_AGEMA_signal_1118), .Z0_t (\SboxInst.M20 ), .Z0_f (new_AGEMA_signal_1140), .Z1_t (new_AGEMA_signal_1141), .Z1_f (new_AGEMA_signal_1142) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_M21.U1 ( .A0_t (\SboxInst.M17 ), .A0_f (new_AGEMA_signal_1131), .A1_t (new_AGEMA_signal_1132), .A1_f (new_AGEMA_signal_1133), .B0_t (\SboxInst.M15 ), .B0_f (new_AGEMA_signal_1125), .B1_t (new_AGEMA_signal_1126), .B1_f (new_AGEMA_signal_1127), .Z0_t (\SboxInst.M21 ), .Z0_f (new_AGEMA_signal_1143), .Z1_t (new_AGEMA_signal_1144), .Z1_f (new_AGEMA_signal_1145) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_M22.U1 ( .A0_t (\SboxInst.M18 ), .A0_f (new_AGEMA_signal_1134), .A1_t (new_AGEMA_signal_1135), .A1_f (new_AGEMA_signal_1136), .B0_t (\SboxInst.M13 ), .B0_f (new_AGEMA_signal_1116), .B1_t (new_AGEMA_signal_1117), .B1_f (new_AGEMA_signal_1118), .Z0_t (\SboxInst.M22 ), .Z0_f (new_AGEMA_signal_1146), .Z1_t (new_AGEMA_signal_1147), .Z1_f (new_AGEMA_signal_1148) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_M23.U1 ( .A0_t (\SboxInst.M19 ), .A0_f (new_AGEMA_signal_1137), .A1_t (new_AGEMA_signal_1138), .A1_f (new_AGEMA_signal_1139), .B0_t (\SboxInst.T25 ), .B0_f (new_AGEMA_signal_1098), .B1_t (new_AGEMA_signal_1099), .B1_f (new_AGEMA_signal_1100), .Z0_t (\SboxInst.M23 ), .Z0_f (new_AGEMA_signal_1149), .Z1_t (new_AGEMA_signal_1150), .Z1_f (new_AGEMA_signal_1151) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_M24.U1 ( .A0_t (\SboxInst.M22 ), .A0_f (new_AGEMA_signal_1146), .A1_t (new_AGEMA_signal_1147), .A1_f (new_AGEMA_signal_1148), .B0_t (\SboxInst.M23 ), .B0_f (new_AGEMA_signal_1149), .B1_t (new_AGEMA_signal_1150), .B1_f (new_AGEMA_signal_1151), .Z0_t (\SboxInst.M24 ), .Z0_f (new_AGEMA_signal_1161), .Z1_t (new_AGEMA_signal_1162), .Z1_f (new_AGEMA_signal_1163) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M25.U1 ( .A0_t (\SboxInst.M22 ), .A0_f (new_AGEMA_signal_1146), .A1_t (new_AGEMA_signal_1147), .A1_f (new_AGEMA_signal_1148), .B0_t (\SboxInst.M20 ), .B0_f (new_AGEMA_signal_1140), .B1_t (new_AGEMA_signal_1141), .B1_f (new_AGEMA_signal_1142), .Z0_t (\SboxInst.M25 ), .Z0_f (new_AGEMA_signal_1152), .Z1_t (new_AGEMA_signal_1153), .Z1_f (new_AGEMA_signal_1154) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_M26.U1 ( .A0_t (\SboxInst.M21 ), .A0_f (new_AGEMA_signal_1143), .A1_t (new_AGEMA_signal_1144), .A1_f (new_AGEMA_signal_1145), .B0_t (\SboxInst.M25 ), .B0_f (new_AGEMA_signal_1152), .B1_t (new_AGEMA_signal_1153), .B1_f (new_AGEMA_signal_1154), .Z0_t (\SboxInst.M26 ), .Z0_f (new_AGEMA_signal_1164), .Z1_t (new_AGEMA_signal_1165), .Z1_f (new_AGEMA_signal_1166) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_M27.U1 ( .A0_t (\SboxInst.M20 ), .A0_f (new_AGEMA_signal_1140), .A1_t (new_AGEMA_signal_1141), .A1_f (new_AGEMA_signal_1142), .B0_t (\SboxInst.M21 ), .B0_f (new_AGEMA_signal_1143), .B1_t (new_AGEMA_signal_1144), .B1_f (new_AGEMA_signal_1145), .Z0_t (\SboxInst.M27 ), .Z0_f (new_AGEMA_signal_1155), .Z1_t (new_AGEMA_signal_1156), .Z1_f (new_AGEMA_signal_1157) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_M28.U1 ( .A0_t (\SboxInst.M23 ), .A0_f (new_AGEMA_signal_1149), .A1_t (new_AGEMA_signal_1150), .A1_f (new_AGEMA_signal_1151), .B0_t (\SboxInst.M25 ), .B0_f (new_AGEMA_signal_1152), .B1_t (new_AGEMA_signal_1153), .B1_f (new_AGEMA_signal_1154), .Z0_t (\SboxInst.M28 ), .Z0_f (new_AGEMA_signal_1167), .Z1_t (new_AGEMA_signal_1168), .Z1_f (new_AGEMA_signal_1169) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M29.U1 ( .A0_t (\SboxInst.M28 ), .A0_f (new_AGEMA_signal_1167), .A1_t (new_AGEMA_signal_1168), .A1_f (new_AGEMA_signal_1169), .B0_t (\SboxInst.M27 ), .B0_f (new_AGEMA_signal_1155), .B1_t (new_AGEMA_signal_1156), .B1_f (new_AGEMA_signal_1157), .Z0_t (\SboxInst.M29 ), .Z0_f (new_AGEMA_signal_1176), .Z1_t (new_AGEMA_signal_1177), .Z1_f (new_AGEMA_signal_1178) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M30.U1 ( .A0_t (\SboxInst.M26 ), .A0_f (new_AGEMA_signal_1164), .A1_t (new_AGEMA_signal_1165), .A1_f (new_AGEMA_signal_1166), .B0_t (\SboxInst.M24 ), .B0_f (new_AGEMA_signal_1161), .B1_t (new_AGEMA_signal_1162), .B1_f (new_AGEMA_signal_1163), .Z0_t (\SboxInst.M30 ), .Z0_f (new_AGEMA_signal_1179), .Z1_t (new_AGEMA_signal_1180), .Z1_f (new_AGEMA_signal_1181) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M31.U1 ( .A0_t (\SboxInst.M20 ), .A0_f (new_AGEMA_signal_1140), .A1_t (new_AGEMA_signal_1141), .A1_f (new_AGEMA_signal_1142), .B0_t (\SboxInst.M23 ), .B0_f (new_AGEMA_signal_1149), .B1_t (new_AGEMA_signal_1150), .B1_f (new_AGEMA_signal_1151), .Z0_t (\SboxInst.M31 ), .Z0_f (new_AGEMA_signal_1170), .Z1_t (new_AGEMA_signal_1171), .Z1_f (new_AGEMA_signal_1172) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M32.U1 ( .A0_t (\SboxInst.M27 ), .A0_f (new_AGEMA_signal_1155), .A1_t (new_AGEMA_signal_1156), .A1_f (new_AGEMA_signal_1157), .B0_t (\SboxInst.M31 ), .B0_f (new_AGEMA_signal_1170), .B1_t (new_AGEMA_signal_1171), .B1_f (new_AGEMA_signal_1172), .Z0_t (\SboxInst.M32 ), .Z0_f (new_AGEMA_signal_1182), .Z1_t (new_AGEMA_signal_1183), .Z1_f (new_AGEMA_signal_1184) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_M33.U1 ( .A0_t (\SboxInst.M27 ), .A0_f (new_AGEMA_signal_1155), .A1_t (new_AGEMA_signal_1156), .A1_f (new_AGEMA_signal_1157), .B0_t (\SboxInst.M25 ), .B0_f (new_AGEMA_signal_1152), .B1_t (new_AGEMA_signal_1153), .B1_f (new_AGEMA_signal_1154), .Z0_t (\SboxInst.M33 ), .Z0_f (new_AGEMA_signal_1173), .Z1_t (new_AGEMA_signal_1174), .Z1_f (new_AGEMA_signal_1175) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M34.U1 ( .A0_t (\SboxInst.M21 ), .A0_f (new_AGEMA_signal_1143), .A1_t (new_AGEMA_signal_1144), .A1_f (new_AGEMA_signal_1145), .B0_t (\SboxInst.M22 ), .B0_f (new_AGEMA_signal_1146), .B1_t (new_AGEMA_signal_1147), .B1_f (new_AGEMA_signal_1148), .Z0_t (\SboxInst.M34 ), .Z0_f (new_AGEMA_signal_1158), .Z1_t (new_AGEMA_signal_1159), .Z1_f (new_AGEMA_signal_1160) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M35.U1 ( .A0_t (\SboxInst.M24 ), .A0_f (new_AGEMA_signal_1161), .A1_t (new_AGEMA_signal_1162), .A1_f (new_AGEMA_signal_1163), .B0_t (\SboxInst.M34 ), .B0_f (new_AGEMA_signal_1158), .B1_t (new_AGEMA_signal_1159), .B1_f (new_AGEMA_signal_1160), .Z0_t (\SboxInst.M35 ), .Z0_f (new_AGEMA_signal_1185), .Z1_t (new_AGEMA_signal_1186), .Z1_f (new_AGEMA_signal_1187) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_M36.U1 ( .A0_t (\SboxInst.M24 ), .A0_f (new_AGEMA_signal_1161), .A1_t (new_AGEMA_signal_1162), .A1_f (new_AGEMA_signal_1163), .B0_t (\SboxInst.M25 ), .B0_f (new_AGEMA_signal_1152), .B1_t (new_AGEMA_signal_1153), .B1_f (new_AGEMA_signal_1154), .Z0_t (\SboxInst.M36 ), .Z0_f (new_AGEMA_signal_1188), .Z1_t (new_AGEMA_signal_1189), .Z1_f (new_AGEMA_signal_1190) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_M37.U1 ( .A0_t (\SboxInst.M21 ), .A0_f (new_AGEMA_signal_1143), .A1_t (new_AGEMA_signal_1144), .A1_f (new_AGEMA_signal_1145), .B0_t (\SboxInst.M29 ), .B0_f (new_AGEMA_signal_1176), .B1_t (new_AGEMA_signal_1177), .B1_f (new_AGEMA_signal_1178), .Z0_t (\SboxInst.M37 ), .Z0_f (new_AGEMA_signal_1191), .Z1_t (new_AGEMA_signal_1192), .Z1_f (new_AGEMA_signal_1193) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_M38.U1 ( .A0_t (\SboxInst.M32 ), .A0_f (new_AGEMA_signal_1182), .A1_t (new_AGEMA_signal_1183), .A1_f (new_AGEMA_signal_1184), .B0_t (\SboxInst.M33 ), .B0_f (new_AGEMA_signal_1173), .B1_t (new_AGEMA_signal_1174), .B1_f (new_AGEMA_signal_1175), .Z0_t (\SboxInst.M38 ), .Z0_f (new_AGEMA_signal_1194), .Z1_t (new_AGEMA_signal_1195), .Z1_f (new_AGEMA_signal_1196) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_M39.U1 ( .A0_t (\SboxInst.M23 ), .A0_f (new_AGEMA_signal_1149), .A1_t (new_AGEMA_signal_1150), .A1_f (new_AGEMA_signal_1151), .B0_t (\SboxInst.M30 ), .B0_f (new_AGEMA_signal_1179), .B1_t (new_AGEMA_signal_1180), .B1_f (new_AGEMA_signal_1181), .Z0_t (\SboxInst.M39 ), .Z0_f (new_AGEMA_signal_1197), .Z1_t (new_AGEMA_signal_1198), .Z1_f (new_AGEMA_signal_1199) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_M40.U1 ( .A0_t (\SboxInst.M35 ), .A0_f (new_AGEMA_signal_1185), .A1_t (new_AGEMA_signal_1186), .A1_f (new_AGEMA_signal_1187), .B0_t (\SboxInst.M36 ), .B0_f (new_AGEMA_signal_1188), .B1_t (new_AGEMA_signal_1189), .B1_f (new_AGEMA_signal_1190), .Z0_t (\SboxInst.M40 ), .Z0_f (new_AGEMA_signal_1200), .Z1_t (new_AGEMA_signal_1201), .Z1_f (new_AGEMA_signal_1202) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_M41.U1 ( .A0_t (\SboxInst.M38 ), .A0_f (new_AGEMA_signal_1194), .A1_t (new_AGEMA_signal_1195), .A1_f (new_AGEMA_signal_1196), .B0_t (\SboxInst.M40 ), .B0_f (new_AGEMA_signal_1200), .B1_t (new_AGEMA_signal_1201), .B1_f (new_AGEMA_signal_1202), .Z0_t (\SboxInst.M41 ), .Z0_f (new_AGEMA_signal_1203), .Z1_t (new_AGEMA_signal_1204), .Z1_f (new_AGEMA_signal_1205) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_M42.U1 ( .A0_t (\SboxInst.M37 ), .A0_f (new_AGEMA_signal_1191), .A1_t (new_AGEMA_signal_1192), .A1_f (new_AGEMA_signal_1193), .B0_t (\SboxInst.M39 ), .B0_f (new_AGEMA_signal_1197), .B1_t (new_AGEMA_signal_1198), .B1_f (new_AGEMA_signal_1199), .Z0_t (\SboxInst.M42 ), .Z0_f (new_AGEMA_signal_1206), .Z1_t (new_AGEMA_signal_1207), .Z1_f (new_AGEMA_signal_1208) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_M43.U1 ( .A0_t (\SboxInst.M37 ), .A0_f (new_AGEMA_signal_1191), .A1_t (new_AGEMA_signal_1192), .A1_f (new_AGEMA_signal_1193), .B0_t (\SboxInst.M38 ), .B0_f (new_AGEMA_signal_1194), .B1_t (new_AGEMA_signal_1195), .B1_f (new_AGEMA_signal_1196), .Z0_t (\SboxInst.M43 ), .Z0_f (new_AGEMA_signal_1209), .Z1_t (new_AGEMA_signal_1210), .Z1_f (new_AGEMA_signal_1211) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_M44.U1 ( .A0_t (\SboxInst.M39 ), .A0_f (new_AGEMA_signal_1197), .A1_t (new_AGEMA_signal_1198), .A1_f (new_AGEMA_signal_1199), .B0_t (\SboxInst.M40 ), .B0_f (new_AGEMA_signal_1200), .B1_t (new_AGEMA_signal_1201), .B1_f (new_AGEMA_signal_1202), .Z0_t (\SboxInst.M44 ), .Z0_f (new_AGEMA_signal_1212), .Z1_t (new_AGEMA_signal_1213), .Z1_f (new_AGEMA_signal_1214) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_M45.U1 ( .A0_t (\SboxInst.M42 ), .A0_f (new_AGEMA_signal_1206), .A1_t (new_AGEMA_signal_1207), .A1_f (new_AGEMA_signal_1208), .B0_t (\SboxInst.M41 ), .B0_f (new_AGEMA_signal_1203), .B1_t (new_AGEMA_signal_1204), .B1_f (new_AGEMA_signal_1205), .Z0_t (\SboxInst.M45 ), .Z0_f (new_AGEMA_signal_1239), .Z1_t (new_AGEMA_signal_1240), .Z1_f (new_AGEMA_signal_1241) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M46.U1 ( .A0_t (\SboxInst.M44 ), .A0_f (new_AGEMA_signal_1212), .A1_t (new_AGEMA_signal_1213), .A1_f (new_AGEMA_signal_1214), .B0_t (\SboxInst.T6 ), .B0_f (new_AGEMA_signal_1032), .B1_t (new_AGEMA_signal_1033), .B1_f (new_AGEMA_signal_1034), .Z0_t (\SboxInst.M46 ), .Z0_f (new_AGEMA_signal_1242), .Z1_t (new_AGEMA_signal_1243), .Z1_f (new_AGEMA_signal_1244) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M47.U1 ( .A0_t (\SboxInst.M40 ), .A0_f (new_AGEMA_signal_1200), .A1_t (new_AGEMA_signal_1201), .A1_f (new_AGEMA_signal_1202), .B0_t (\SboxInst.T8 ), .B0_f (new_AGEMA_signal_1056), .B1_t (new_AGEMA_signal_1057), .B1_f (new_AGEMA_signal_1058), .Z0_t (\SboxInst.M47 ), .Z0_f (new_AGEMA_signal_1215), .Z1_t (new_AGEMA_signal_1216), .Z1_f (new_AGEMA_signal_1217) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M48.U1 ( .A0_t (\SboxInst.M39 ), .A0_f (new_AGEMA_signal_1197), .A1_t (new_AGEMA_signal_1198), .A1_f (new_AGEMA_signal_1199), .B0_t (Sbox_in[0]), .B0_f (new_AGEMA_signal_978), .B1_t (new_AGEMA_signal_979), .B1_f (new_AGEMA_signal_980), .Z0_t (\SboxInst.M48 ), .Z0_f (new_AGEMA_signal_1218), .Z1_t (new_AGEMA_signal_1219), .Z1_f (new_AGEMA_signal_1220) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M49.U1 ( .A0_t (\SboxInst.M43 ), .A0_f (new_AGEMA_signal_1209), .A1_t (new_AGEMA_signal_1210), .A1_f (new_AGEMA_signal_1211), .B0_t (\SboxInst.T16 ), .B0_f (new_AGEMA_signal_1044), .B1_t (new_AGEMA_signal_1045), .B1_f (new_AGEMA_signal_1046), .Z0_t (\SboxInst.M49 ), .Z0_f (new_AGEMA_signal_1245), .Z1_t (new_AGEMA_signal_1246), .Z1_f (new_AGEMA_signal_1247) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M50.U1 ( .A0_t (\SboxInst.M38 ), .A0_f (new_AGEMA_signal_1194), .A1_t (new_AGEMA_signal_1195), .A1_f (new_AGEMA_signal_1196), .B0_t (\SboxInst.T9 ), .B0_f (new_AGEMA_signal_1035), .B1_t (new_AGEMA_signal_1036), .B1_f (new_AGEMA_signal_1037), .Z0_t (\SboxInst.M50 ), .Z0_f (new_AGEMA_signal_1221), .Z1_t (new_AGEMA_signal_1222), .Z1_f (new_AGEMA_signal_1223) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M51.U1 ( .A0_t (\SboxInst.M37 ), .A0_f (new_AGEMA_signal_1191), .A1_t (new_AGEMA_signal_1192), .A1_f (new_AGEMA_signal_1193), .B0_t (\SboxInst.T17 ), .B0_f (new_AGEMA_signal_1065), .B1_t (new_AGEMA_signal_1066), .B1_f (new_AGEMA_signal_1067), .Z0_t (\SboxInst.M51 ), .Z0_f (new_AGEMA_signal_1224), .Z1_t (new_AGEMA_signal_1225), .Z1_f (new_AGEMA_signal_1226) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M52.U1 ( .A0_t (\SboxInst.M42 ), .A0_f (new_AGEMA_signal_1206), .A1_t (new_AGEMA_signal_1207), .A1_f (new_AGEMA_signal_1208), .B0_t (\SboxInst.T15 ), .B0_f (new_AGEMA_signal_1041), .B1_t (new_AGEMA_signal_1042), .B1_f (new_AGEMA_signal_1043), .Z0_t (\SboxInst.M52 ), .Z0_f (new_AGEMA_signal_1248), .Z1_t (new_AGEMA_signal_1249), .Z1_f (new_AGEMA_signal_1250) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M53.U1 ( .A0_t (\SboxInst.M45 ), .A0_f (new_AGEMA_signal_1239), .A1_t (new_AGEMA_signal_1240), .A1_f (new_AGEMA_signal_1241), .B0_t (\SboxInst.T27 ), .B0_f (new_AGEMA_signal_1053), .B1_t (new_AGEMA_signal_1054), .B1_f (new_AGEMA_signal_1055), .Z0_t (\SboxInst.M53 ), .Z0_f (new_AGEMA_signal_1275), .Z1_t (new_AGEMA_signal_1276), .Z1_f (new_AGEMA_signal_1277) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M54.U1 ( .A0_t (\SboxInst.M41 ), .A0_f (new_AGEMA_signal_1203), .A1_t (new_AGEMA_signal_1204), .A1_f (new_AGEMA_signal_1205), .B0_t (\SboxInst.T10 ), .B0_f (new_AGEMA_signal_1059), .B1_t (new_AGEMA_signal_1060), .B1_f (new_AGEMA_signal_1061), .Z0_t (\SboxInst.M54 ), .Z0_f (new_AGEMA_signal_1251), .Z1_t (new_AGEMA_signal_1252), .Z1_f (new_AGEMA_signal_1253) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M55.U1 ( .A0_t (\SboxInst.M44 ), .A0_f (new_AGEMA_signal_1212), .A1_t (new_AGEMA_signal_1213), .A1_f (new_AGEMA_signal_1214), .B0_t (\SboxInst.T13 ), .B0_f (new_AGEMA_signal_1038), .B1_t (new_AGEMA_signal_1039), .B1_f (new_AGEMA_signal_1040), .Z0_t (\SboxInst.M55 ), .Z0_f (new_AGEMA_signal_1254), .Z1_t (new_AGEMA_signal_1255), .Z1_f (new_AGEMA_signal_1256) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M56.U1 ( .A0_t (\SboxInst.M40 ), .A0_f (new_AGEMA_signal_1200), .A1_t (new_AGEMA_signal_1201), .A1_f (new_AGEMA_signal_1202), .B0_t (\SboxInst.T23 ), .B0_f (new_AGEMA_signal_1071), .B1_t (new_AGEMA_signal_1072), .B1_f (new_AGEMA_signal_1073), .Z0_t (\SboxInst.M56 ), .Z0_f (new_AGEMA_signal_1227), .Z1_t (new_AGEMA_signal_1228), .Z1_f (new_AGEMA_signal_1229) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M57.U1 ( .A0_t (\SboxInst.M39 ), .A0_f (new_AGEMA_signal_1197), .A1_t (new_AGEMA_signal_1198), .A1_f (new_AGEMA_signal_1199), .B0_t (\SboxInst.T19 ), .B0_f (new_AGEMA_signal_1047), .B1_t (new_AGEMA_signal_1048), .B1_f (new_AGEMA_signal_1049), .Z0_t (\SboxInst.M57 ), .Z0_f (new_AGEMA_signal_1230), .Z1_t (new_AGEMA_signal_1231), .Z1_f (new_AGEMA_signal_1232) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M58.U1 ( .A0_t (\SboxInst.M43 ), .A0_f (new_AGEMA_signal_1209), .A1_t (new_AGEMA_signal_1210), .A1_f (new_AGEMA_signal_1211), .B0_t (\SboxInst.T3 ), .B0_f (new_AGEMA_signal_1008), .B1_t (new_AGEMA_signal_1009), .B1_f (new_AGEMA_signal_1010), .Z0_t (\SboxInst.M58 ), .Z0_f (new_AGEMA_signal_1257), .Z1_t (new_AGEMA_signal_1258), .Z1_f (new_AGEMA_signal_1259) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M59.U1 ( .A0_t (\SboxInst.M38 ), .A0_f (new_AGEMA_signal_1194), .A1_t (new_AGEMA_signal_1195), .A1_f (new_AGEMA_signal_1196), .B0_t (\SboxInst.T22 ), .B0_f (new_AGEMA_signal_1050), .B1_t (new_AGEMA_signal_1051), .B1_f (new_AGEMA_signal_1052), .Z0_t (\SboxInst.M59 ), .Z0_f (new_AGEMA_signal_1233), .Z1_t (new_AGEMA_signal_1234), .Z1_f (new_AGEMA_signal_1235) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M60.U1 ( .A0_t (\SboxInst.M37 ), .A0_f (new_AGEMA_signal_1191), .A1_t (new_AGEMA_signal_1192), .A1_f (new_AGEMA_signal_1193), .B0_t (\SboxInst.T20 ), .B0_f (new_AGEMA_signal_1068), .B1_t (new_AGEMA_signal_1069), .B1_f (new_AGEMA_signal_1070), .Z0_t (\SboxInst.M60 ), .Z0_f (new_AGEMA_signal_1236), .Z1_t (new_AGEMA_signal_1237), .Z1_f (new_AGEMA_signal_1238) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M61.U1 ( .A0_t (\SboxInst.M42 ), .A0_f (new_AGEMA_signal_1206), .A1_t (new_AGEMA_signal_1207), .A1_f (new_AGEMA_signal_1208), .B0_t (\SboxInst.T1 ), .B0_f (new_AGEMA_signal_1002), .B1_t (new_AGEMA_signal_1003), .B1_f (new_AGEMA_signal_1004), .Z0_t (\SboxInst.M61 ), .Z0_f (new_AGEMA_signal_1260), .Z1_t (new_AGEMA_signal_1261), .Z1_f (new_AGEMA_signal_1262) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M62.U1 ( .A0_t (\SboxInst.M45 ), .A0_f (new_AGEMA_signal_1239), .A1_t (new_AGEMA_signal_1240), .A1_f (new_AGEMA_signal_1241), .B0_t (\SboxInst.T4 ), .B0_f (new_AGEMA_signal_1011), .B1_t (new_AGEMA_signal_1012), .B1_f (new_AGEMA_signal_1013), .Z0_t (\SboxInst.M62 ), .Z0_f (new_AGEMA_signal_1278), .Z1_t (new_AGEMA_signal_1279), .Z1_f (new_AGEMA_signal_1280) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M63.U1 ( .A0_t (\SboxInst.M41 ), .A0_f (new_AGEMA_signal_1203), .A1_t (new_AGEMA_signal_1204), .A1_f (new_AGEMA_signal_1205), .B0_t (\SboxInst.T2 ), .B0_f (new_AGEMA_signal_1005), .B1_t (new_AGEMA_signal_1006), .B1_f (new_AGEMA_signal_1007), .Z0_t (\SboxInst.M63 ), .Z0_f (new_AGEMA_signal_1263), .Z1_t (new_AGEMA_signal_1264), .Z1_f (new_AGEMA_signal_1265) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_L0.U1 ( .A0_t (\SboxInst.M61 ), .A0_f (new_AGEMA_signal_1260), .A1_t (new_AGEMA_signal_1261), .A1_f (new_AGEMA_signal_1262), .B0_t (\SboxInst.M62 ), .B0_f (new_AGEMA_signal_1278), .B1_t (new_AGEMA_signal_1279), .B1_f (new_AGEMA_signal_1280), .Z0_t (\SboxInst.L0 ), .Z0_f (new_AGEMA_signal_1305), .Z1_t (new_AGEMA_signal_1306), .Z1_f (new_AGEMA_signal_1307) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_L1.U1 ( .A0_t (\SboxInst.M50 ), .A0_f (new_AGEMA_signal_1221), .A1_t (new_AGEMA_signal_1222), .A1_f (new_AGEMA_signal_1223), .B0_t (\SboxInst.M56 ), .B0_f (new_AGEMA_signal_1227), .B1_t (new_AGEMA_signal_1228), .B1_f (new_AGEMA_signal_1229), .Z0_t (\SboxInst.L1 ), .Z0_f (new_AGEMA_signal_1266), .Z1_t (new_AGEMA_signal_1267), .Z1_f (new_AGEMA_signal_1268) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_L2.U1 ( .A0_t (\SboxInst.M46 ), .A0_f (new_AGEMA_signal_1242), .A1_t (new_AGEMA_signal_1243), .A1_f (new_AGEMA_signal_1244), .B0_t (\SboxInst.M48 ), .B0_f (new_AGEMA_signal_1218), .B1_t (new_AGEMA_signal_1219), .B1_f (new_AGEMA_signal_1220), .Z0_t (\SboxInst.L2 ), .Z0_f (new_AGEMA_signal_1281), .Z1_t (new_AGEMA_signal_1282), .Z1_f (new_AGEMA_signal_1283) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_L3.U1 ( .A0_t (\SboxInst.M47 ), .A0_f (new_AGEMA_signal_1215), .A1_t (new_AGEMA_signal_1216), .A1_f (new_AGEMA_signal_1217), .B0_t (\SboxInst.M55 ), .B0_f (new_AGEMA_signal_1254), .B1_t (new_AGEMA_signal_1255), .B1_f (new_AGEMA_signal_1256), .Z0_t (\SboxInst.L3 ), .Z0_f (new_AGEMA_signal_1284), .Z1_t (new_AGEMA_signal_1285), .Z1_f (new_AGEMA_signal_1286) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_L4.U1 ( .A0_t (\SboxInst.M54 ), .A0_f (new_AGEMA_signal_1251), .A1_t (new_AGEMA_signal_1252), .A1_f (new_AGEMA_signal_1253), .B0_t (\SboxInst.M58 ), .B0_f (new_AGEMA_signal_1257), .B1_t (new_AGEMA_signal_1258), .B1_f (new_AGEMA_signal_1259), .Z0_t (\SboxInst.L4 ), .Z0_f (new_AGEMA_signal_1287), .Z1_t (new_AGEMA_signal_1288), .Z1_f (new_AGEMA_signal_1289) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_L5.U1 ( .A0_t (\SboxInst.M49 ), .A0_f (new_AGEMA_signal_1245), .A1_t (new_AGEMA_signal_1246), .A1_f (new_AGEMA_signal_1247), .B0_t (\SboxInst.M61 ), .B0_f (new_AGEMA_signal_1260), .B1_t (new_AGEMA_signal_1261), .B1_f (new_AGEMA_signal_1262), .Z0_t (\SboxInst.L5 ), .Z0_f (new_AGEMA_signal_1290), .Z1_t (new_AGEMA_signal_1291), .Z1_f (new_AGEMA_signal_1292) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_L6.U1 ( .A0_t (\SboxInst.M62 ), .A0_f (new_AGEMA_signal_1278), .A1_t (new_AGEMA_signal_1279), .A1_f (new_AGEMA_signal_1280), .B0_t (\SboxInst.L5 ), .B0_f (new_AGEMA_signal_1290), .B1_t (new_AGEMA_signal_1291), .B1_f (new_AGEMA_signal_1292), .Z0_t (\SboxInst.L6 ), .Z0_f (new_AGEMA_signal_1308), .Z1_t (new_AGEMA_signal_1309), .Z1_f (new_AGEMA_signal_1310) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_L7.U1 ( .A0_t (\SboxInst.M46 ), .A0_f (new_AGEMA_signal_1242), .A1_t (new_AGEMA_signal_1243), .A1_f (new_AGEMA_signal_1244), .B0_t (\SboxInst.L3 ), .B0_f (new_AGEMA_signal_1284), .B1_t (new_AGEMA_signal_1285), .B1_f (new_AGEMA_signal_1286), .Z0_t (\SboxInst.L7 ), .Z0_f (new_AGEMA_signal_1311), .Z1_t (new_AGEMA_signal_1312), .Z1_f (new_AGEMA_signal_1313) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_L8.U1 ( .A0_t (\SboxInst.M51 ), .A0_f (new_AGEMA_signal_1224), .A1_t (new_AGEMA_signal_1225), .A1_f (new_AGEMA_signal_1226), .B0_t (\SboxInst.M59 ), .B0_f (new_AGEMA_signal_1233), .B1_t (new_AGEMA_signal_1234), .B1_f (new_AGEMA_signal_1235), .Z0_t (\SboxInst.L8 ), .Z0_f (new_AGEMA_signal_1269), .Z1_t (new_AGEMA_signal_1270), .Z1_f (new_AGEMA_signal_1271) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_L9.U1 ( .A0_t (\SboxInst.M52 ), .A0_f (new_AGEMA_signal_1248), .A1_t (new_AGEMA_signal_1249), .A1_f (new_AGEMA_signal_1250), .B0_t (\SboxInst.M53 ), .B0_f (new_AGEMA_signal_1275), .B1_t (new_AGEMA_signal_1276), .B1_f (new_AGEMA_signal_1277), .Z0_t (\SboxInst.L9 ), .Z0_f (new_AGEMA_signal_1314), .Z1_t (new_AGEMA_signal_1315), .Z1_f (new_AGEMA_signal_1316) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_L10.U1 ( .A0_t (\SboxInst.M53 ), .A0_f (new_AGEMA_signal_1275), .A1_t (new_AGEMA_signal_1276), .A1_f (new_AGEMA_signal_1277), .B0_t (\SboxInst.L4 ), .B0_f (new_AGEMA_signal_1287), .B1_t (new_AGEMA_signal_1288), .B1_f (new_AGEMA_signal_1289), .Z0_t (\SboxInst.L10 ), .Z0_f (new_AGEMA_signal_1317), .Z1_t (new_AGEMA_signal_1318), .Z1_f (new_AGEMA_signal_1319) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_L11.U1 ( .A0_t (\SboxInst.M60 ), .A0_f (new_AGEMA_signal_1236), .A1_t (new_AGEMA_signal_1237), .A1_f (new_AGEMA_signal_1238), .B0_t (\SboxInst.L2 ), .B0_f (new_AGEMA_signal_1281), .B1_t (new_AGEMA_signal_1282), .B1_f (new_AGEMA_signal_1283), .Z0_t (\SboxInst.L11 ), .Z0_f (new_AGEMA_signal_1320), .Z1_t (new_AGEMA_signal_1321), .Z1_f (new_AGEMA_signal_1322) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_L12.U1 ( .A0_t (\SboxInst.M48 ), .A0_f (new_AGEMA_signal_1218), .A1_t (new_AGEMA_signal_1219), .A1_f (new_AGEMA_signal_1220), .B0_t (\SboxInst.M51 ), .B0_f (new_AGEMA_signal_1224), .B1_t (new_AGEMA_signal_1225), .B1_f (new_AGEMA_signal_1226), .Z0_t (\SboxInst.L12 ), .Z0_f (new_AGEMA_signal_1272), .Z1_t (new_AGEMA_signal_1273), .Z1_f (new_AGEMA_signal_1274) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_L13.U1 ( .A0_t (\SboxInst.M50 ), .A0_f (new_AGEMA_signal_1221), .A1_t (new_AGEMA_signal_1222), .A1_f (new_AGEMA_signal_1223), .B0_t (\SboxInst.L0 ), .B0_f (new_AGEMA_signal_1305), .B1_t (new_AGEMA_signal_1306), .B1_f (new_AGEMA_signal_1307), .Z0_t (\SboxInst.L13 ), .Z0_f (new_AGEMA_signal_1332), .Z1_t (new_AGEMA_signal_1333), .Z1_f (new_AGEMA_signal_1334) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_L14.U1 ( .A0_t (\SboxInst.M52 ), .A0_f (new_AGEMA_signal_1248), .A1_t (new_AGEMA_signal_1249), .A1_f (new_AGEMA_signal_1250), .B0_t (\SboxInst.M61 ), .B0_f (new_AGEMA_signal_1260), .B1_t (new_AGEMA_signal_1261), .B1_f (new_AGEMA_signal_1262), .Z0_t (\SboxInst.L14 ), .Z0_f (new_AGEMA_signal_1293), .Z1_t (new_AGEMA_signal_1294), .Z1_f (new_AGEMA_signal_1295) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_L15.U1 ( .A0_t (\SboxInst.M55 ), .A0_f (new_AGEMA_signal_1254), .A1_t (new_AGEMA_signal_1255), .A1_f (new_AGEMA_signal_1256), .B0_t (\SboxInst.L1 ), .B0_f (new_AGEMA_signal_1266), .B1_t (new_AGEMA_signal_1267), .B1_f (new_AGEMA_signal_1268), .Z0_t (\SboxInst.L15 ), .Z0_f (new_AGEMA_signal_1296), .Z1_t (new_AGEMA_signal_1297), .Z1_f (new_AGEMA_signal_1298) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_L16.U1 ( .A0_t (\SboxInst.M56 ), .A0_f (new_AGEMA_signal_1227), .A1_t (new_AGEMA_signal_1228), .A1_f (new_AGEMA_signal_1229), .B0_t (\SboxInst.L0 ), .B0_f (new_AGEMA_signal_1305), .B1_t (new_AGEMA_signal_1306), .B1_f (new_AGEMA_signal_1307), .Z0_t (\SboxInst.L16 ), .Z0_f (new_AGEMA_signal_1335), .Z1_t (new_AGEMA_signal_1336), .Z1_f (new_AGEMA_signal_1337) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_L17.U1 ( .A0_t (\SboxInst.M57 ), .A0_f (new_AGEMA_signal_1230), .A1_t (new_AGEMA_signal_1231), .A1_f (new_AGEMA_signal_1232), .B0_t (\SboxInst.L1 ), .B0_f (new_AGEMA_signal_1266), .B1_t (new_AGEMA_signal_1267), .B1_f (new_AGEMA_signal_1268), .Z0_t (\SboxInst.L17 ), .Z0_f (new_AGEMA_signal_1299), .Z1_t (new_AGEMA_signal_1300), .Z1_f (new_AGEMA_signal_1301) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_L18.U1 ( .A0_t (\SboxInst.M58 ), .A0_f (new_AGEMA_signal_1257), .A1_t (new_AGEMA_signal_1258), .A1_f (new_AGEMA_signal_1259), .B0_t (\SboxInst.L8 ), .B0_f (new_AGEMA_signal_1269), .B1_t (new_AGEMA_signal_1270), .B1_f (new_AGEMA_signal_1271), .Z0_t (\SboxInst.L18 ), .Z0_f (new_AGEMA_signal_1302), .Z1_t (new_AGEMA_signal_1303), .Z1_f (new_AGEMA_signal_1304) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_L19.U1 ( .A0_t (\SboxInst.M63 ), .A0_f (new_AGEMA_signal_1263), .A1_t (new_AGEMA_signal_1264), .A1_f (new_AGEMA_signal_1265), .B0_t (\SboxInst.L4 ), .B0_f (new_AGEMA_signal_1287), .B1_t (new_AGEMA_signal_1288), .B1_f (new_AGEMA_signal_1289), .Z0_t (\SboxInst.L19 ), .Z0_f (new_AGEMA_signal_1323), .Z1_t (new_AGEMA_signal_1324), .Z1_f (new_AGEMA_signal_1325) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_L20.U1 ( .A0_t (\SboxInst.L0 ), .A0_f (new_AGEMA_signal_1305), .A1_t (new_AGEMA_signal_1306), .A1_f (new_AGEMA_signal_1307), .B0_t (\SboxInst.L1 ), .B0_f (new_AGEMA_signal_1266), .B1_t (new_AGEMA_signal_1267), .B1_f (new_AGEMA_signal_1268), .Z0_t (\SboxInst.L20 ), .Z0_f (new_AGEMA_signal_1338), .Z1_t (new_AGEMA_signal_1339), .Z1_f (new_AGEMA_signal_1340) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_L21.U1 ( .A0_t (\SboxInst.L1 ), .A0_f (new_AGEMA_signal_1266), .A1_t (new_AGEMA_signal_1267), .A1_f (new_AGEMA_signal_1268), .B0_t (\SboxInst.L7 ), .B0_f (new_AGEMA_signal_1311), .B1_t (new_AGEMA_signal_1312), .B1_f (new_AGEMA_signal_1313), .Z0_t (\SboxInst.L21 ), .Z0_f (new_AGEMA_signal_1341), .Z1_t (new_AGEMA_signal_1342), .Z1_f (new_AGEMA_signal_1343) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_L22.U1 ( .A0_t (\SboxInst.L3 ), .A0_f (new_AGEMA_signal_1284), .A1_t (new_AGEMA_signal_1285), .A1_f (new_AGEMA_signal_1286), .B0_t (\SboxInst.L12 ), .B0_f (new_AGEMA_signal_1272), .B1_t (new_AGEMA_signal_1273), .B1_f (new_AGEMA_signal_1274), .Z0_t (\SboxInst.L22 ), .Z0_f (new_AGEMA_signal_1326), .Z1_t (new_AGEMA_signal_1327), .Z1_f (new_AGEMA_signal_1328) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_L23.U1 ( .A0_t (\SboxInst.L18 ), .A0_f (new_AGEMA_signal_1302), .A1_t (new_AGEMA_signal_1303), .A1_f (new_AGEMA_signal_1304), .B0_t (\SboxInst.L2 ), .B0_f (new_AGEMA_signal_1281), .B1_t (new_AGEMA_signal_1282), .B1_f (new_AGEMA_signal_1283), .Z0_t (\SboxInst.L23 ), .Z0_f (new_AGEMA_signal_1329), .Z1_t (new_AGEMA_signal_1330), .Z1_f (new_AGEMA_signal_1331) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_L24.U1 ( .A0_t (\SboxInst.L15 ), .A0_f (new_AGEMA_signal_1296), .A1_t (new_AGEMA_signal_1297), .A1_f (new_AGEMA_signal_1298), .B0_t (\SboxInst.L9 ), .B0_f (new_AGEMA_signal_1314), .B1_t (new_AGEMA_signal_1315), .B1_f (new_AGEMA_signal_1316), .Z0_t (\SboxInst.L24 ), .Z0_f (new_AGEMA_signal_1344), .Z1_t (new_AGEMA_signal_1345), .Z1_f (new_AGEMA_signal_1346) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_L25.U1 ( .A0_t (\SboxInst.L6 ), .A0_f (new_AGEMA_signal_1308), .A1_t (new_AGEMA_signal_1309), .A1_f (new_AGEMA_signal_1310), .B0_t (\SboxInst.L10 ), .B0_f (new_AGEMA_signal_1317), .B1_t (new_AGEMA_signal_1318), .B1_f (new_AGEMA_signal_1319), .Z0_t (\SboxInst.L25 ), .Z0_f (new_AGEMA_signal_1347), .Z1_t (new_AGEMA_signal_1348), .Z1_f (new_AGEMA_signal_1349) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_L26.U1 ( .A0_t (\SboxInst.L7 ), .A0_f (new_AGEMA_signal_1311), .A1_t (new_AGEMA_signal_1312), .A1_f (new_AGEMA_signal_1313), .B0_t (\SboxInst.L9 ), .B0_f (new_AGEMA_signal_1314), .B1_t (new_AGEMA_signal_1315), .B1_f (new_AGEMA_signal_1316), .Z0_t (\SboxInst.L26 ), .Z0_f (new_AGEMA_signal_1350), .Z1_t (new_AGEMA_signal_1351), .Z1_f (new_AGEMA_signal_1352) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_L27.U1 ( .A0_t (\SboxInst.L8 ), .A0_f (new_AGEMA_signal_1269), .A1_t (new_AGEMA_signal_1270), .A1_f (new_AGEMA_signal_1271), .B0_t (\SboxInst.L10 ), .B0_f (new_AGEMA_signal_1317), .B1_t (new_AGEMA_signal_1318), .B1_f (new_AGEMA_signal_1319), .Z0_t (\SboxInst.L27 ), .Z0_f (new_AGEMA_signal_1353), .Z1_t (new_AGEMA_signal_1354), .Z1_f (new_AGEMA_signal_1355) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_L28.U1 ( .A0_t (\SboxInst.L11 ), .A0_f (new_AGEMA_signal_1320), .A1_t (new_AGEMA_signal_1321), .A1_f (new_AGEMA_signal_1322), .B0_t (\SboxInst.L14 ), .B0_f (new_AGEMA_signal_1293), .B1_t (new_AGEMA_signal_1294), .B1_f (new_AGEMA_signal_1295), .Z0_t (\SboxInst.L28 ), .Z0_f (new_AGEMA_signal_1356), .Z1_t (new_AGEMA_signal_1357), .Z1_f (new_AGEMA_signal_1358) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_L29.U1 ( .A0_t (\SboxInst.L11 ), .A0_f (new_AGEMA_signal_1320), .A1_t (new_AGEMA_signal_1321), .A1_f (new_AGEMA_signal_1322), .B0_t (\SboxInst.L17 ), .B0_f (new_AGEMA_signal_1299), .B1_t (new_AGEMA_signal_1300), .B1_f (new_AGEMA_signal_1301), .Z0_t (\SboxInst.L29 ), .Z0_f (new_AGEMA_signal_1359), .Z1_t (new_AGEMA_signal_1360), .Z1_f (new_AGEMA_signal_1361) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) \SboxInst.XOR_S0.U1 ( .A0_t (\SboxInst.L6 ), .A0_f (new_AGEMA_signal_1308), .A1_t (new_AGEMA_signal_1309), .A1_f (new_AGEMA_signal_1310), .B0_t (\SboxInst.L24 ), .B0_f (new_AGEMA_signal_1344), .B1_t (new_AGEMA_signal_1345), .B1_f (new_AGEMA_signal_1346), .Z0_t (value_out_s0_t[7]), .Z0_f (value_out_s0_f[7]), .Z1_t (value_out_s1_t[7]), .Z1_f (value_out_s1_f[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) \SboxInst.XOR_S1.U1 ( .A0_t (\SboxInst.L16 ), .A0_f (new_AGEMA_signal_1335), .A1_t (new_AGEMA_signal_1336), .A1_f (new_AGEMA_signal_1337), .B0_t (\SboxInst.L26 ), .B0_f (new_AGEMA_signal_1350), .B1_t (new_AGEMA_signal_1351), .B1_f (new_AGEMA_signal_1352), .Z0_t (value_out_s0_t[6]), .Z0_f (value_out_s0_f[6]), .Z1_t (value_out_s1_t[6]), .Z1_f (value_out_s1_f[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) \SboxInst.XOR_S2.U1 ( .A0_t (\SboxInst.L19 ), .A0_f (new_AGEMA_signal_1323), .A1_t (new_AGEMA_signal_1324), .A1_f (new_AGEMA_signal_1325), .B0_t (\SboxInst.L28 ), .B0_f (new_AGEMA_signal_1356), .B1_t (new_AGEMA_signal_1357), .B1_f (new_AGEMA_signal_1358), .Z0_t (value_out_s0_t[5]), .Z0_f (value_out_s0_f[5]), .Z1_t (value_out_s1_t[5]), .Z1_f (value_out_s1_f[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) \SboxInst.XOR_S3.U1 ( .A0_t (\SboxInst.L6 ), .A0_f (new_AGEMA_signal_1308), .A1_t (new_AGEMA_signal_1309), .A1_f (new_AGEMA_signal_1310), .B0_t (\SboxInst.L21 ), .B0_f (new_AGEMA_signal_1341), .B1_t (new_AGEMA_signal_1342), .B1_f (new_AGEMA_signal_1343), .Z0_t (value_out_s0_t[4]), .Z0_f (value_out_s0_f[4]), .Z1_t (value_out_s1_t[4]), .Z1_f (value_out_s1_f[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) \SboxInst.XOR_S4.U1 ( .A0_t (\SboxInst.L20 ), .A0_f (new_AGEMA_signal_1338), .A1_t (new_AGEMA_signal_1339), .A1_f (new_AGEMA_signal_1340), .B0_t (\SboxInst.L22 ), .B0_f (new_AGEMA_signal_1326), .B1_t (new_AGEMA_signal_1327), .B1_f (new_AGEMA_signal_1328), .Z0_t (value_out_s0_t[3]), .Z0_f (value_out_s0_f[3]), .Z1_t (value_out_s1_t[3]), .Z1_f (value_out_s1_f[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) \SboxInst.XOR_S5.U1 ( .A0_t (\SboxInst.L25 ), .A0_f (new_AGEMA_signal_1347), .A1_t (new_AGEMA_signal_1348), .A1_f (new_AGEMA_signal_1349), .B0_t (\SboxInst.L29 ), .B0_f (new_AGEMA_signal_1359), .B1_t (new_AGEMA_signal_1360), .B1_f (new_AGEMA_signal_1361), .Z0_t (value_out_s0_t[2]), .Z0_f (value_out_s0_f[2]), .Z1_t (value_out_s1_t[2]), .Z1_f (value_out_s1_f[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) \SboxInst.XOR_S6.U1 ( .A0_t (\SboxInst.L13 ), .A0_f (new_AGEMA_signal_1332), .A1_t (new_AGEMA_signal_1333), .A1_f (new_AGEMA_signal_1334), .B0_t (\SboxInst.L27 ), .B0_f (new_AGEMA_signal_1353), .B1_t (new_AGEMA_signal_1354), .B1_f (new_AGEMA_signal_1355), .Z0_t (value_out_s0_t[1]), .Z0_f (value_out_s0_f[1]), .Z1_t (value_out_s1_t[1]), .Z1_f (value_out_s1_f[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) \SboxInst.XOR_S7.U1 ( .A0_t (\SboxInst.L6 ), .A0_f (new_AGEMA_signal_1308), .A1_t (new_AGEMA_signal_1309), .A1_f (new_AGEMA_signal_1310), .B0_t (\SboxInst.L23 ), .B0_f (new_AGEMA_signal_1329), .B1_t (new_AGEMA_signal_1330), .B1_f (new_AGEMA_signal_1331), .Z0_t (value_out_s0_t[0]), .Z0_f (value_out_s0_f[0]), .Z1_t (value_out_s1_t[0]), .Z1_f (value_out_s1_f[0]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) \M2.gen_loop_0__M.X1.U1 ( .A0_t (Inc_Reg[0]), .A0_f (new_AGEMA_signal_930), .B0_t (start_t[0]), .B0_f (start_f[0]), .Z0_t (\M2.gen_loop_0__M.X ), .Z0_f (new_AGEMA_signal_932) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) \M2.gen_loop_0__M.A.U1 ( .A0_t (rst_t), .A0_f (rst_f), .B0_t (\M2.gen_loop_0__M.X ), .B0_f (new_AGEMA_signal_932), .Z0_t (\M2.gen_loop_0__M.Y ), .Z0_f (new_AGEMA_signal_943) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) \M2.gen_loop_0__M.X2.U1 ( .A0_t (\M2.gen_loop_0__M.Y ), .A0_f (new_AGEMA_signal_943), .B0_t (Inc_Reg[0]), .B0_f (new_AGEMA_signal_930), .Z0_t (Inc_in[0]), .Z0_f (new_AGEMA_signal_947) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) \M2.gen_loop_1__M.X1.U1 ( .A0_t (Inc_Reg[1]), .A0_f (new_AGEMA_signal_933), .B0_t (start_t[1]), .B0_f (start_f[1]), .Z0_t (\M2.gen_loop_1__M.X ), .Z0_f (new_AGEMA_signal_935) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) \M2.gen_loop_1__M.A.U1 ( .A0_t (rst_t), .A0_f (rst_f), .B0_t (\M2.gen_loop_1__M.X ), .B0_f (new_AGEMA_signal_935), .Z0_t (\M2.gen_loop_1__M.Y ), .Z0_f (new_AGEMA_signal_944) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) \M2.gen_loop_1__M.X2.U1 ( .A0_t (\M2.gen_loop_1__M.Y ), .A0_f (new_AGEMA_signal_944), .B0_t (Inc_Reg[1]), .B0_f (new_AGEMA_signal_933), .Z0_t (Inc_in[1]), .Z0_f (new_AGEMA_signal_948) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) \M2.gen_loop_2__M.X1.U1 ( .A0_t (Inc_Reg[2]), .A0_f (new_AGEMA_signal_936), .B0_t (start_t[2]), .B0_f (start_f[2]), .Z0_t (\M2.gen_loop_2__M.X ), .Z0_f (new_AGEMA_signal_938) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) \M2.gen_loop_2__M.A.U1 ( .A0_t (rst_t), .A0_f (rst_f), .B0_t (\M2.gen_loop_2__M.X ), .B0_f (new_AGEMA_signal_938), .Z0_t (\M2.gen_loop_2__M.Y ), .Z0_f (new_AGEMA_signal_945) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) \M2.gen_loop_2__M.X2.U1 ( .A0_t (\M2.gen_loop_2__M.Y ), .A0_f (new_AGEMA_signal_945), .B0_t (Inc_Reg[2]), .B0_f (new_AGEMA_signal_936), .Z0_t (Inc_in[2]), .Z0_f (new_AGEMA_signal_949) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) \M2.gen_loop_3__M.X1.U1 ( .A0_t (Inc_Reg[3]), .A0_f (new_AGEMA_signal_939), .B0_t (start_t[3]), .B0_f (start_f[3]), .Z0_t (\M2.gen_loop_3__M.X ), .Z0_f (new_AGEMA_signal_941) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) \M2.gen_loop_3__M.A.U1 ( .A0_t (rst_t), .A0_f (rst_f), .B0_t (\M2.gen_loop_3__M.X ), .B0_f (new_AGEMA_signal_941), .Z0_t (\M2.gen_loop_3__M.Y ), .Z0_f (new_AGEMA_signal_946) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) \M2.gen_loop_3__M.X2.U1 ( .A0_t (\M2.gen_loop_3__M.Y ), .A0_f (new_AGEMA_signal_946), .B0_t (Inc_Reg[3]), .B0_f (new_AGEMA_signal_939), .Z0_t (Inc_in[3]), .Z0_f (new_AGEMA_signal_950) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) U10 ( .A0_t (Inc_in[0]), .A0_f (new_AGEMA_signal_947), .B0_t (Inc_in[1]), .B0_f (new_AGEMA_signal_948), .Z0_t (n9), .Z0_f (new_AGEMA_signal_951) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b1), .NL(1'b0)) U12 ( .A0_t (Inc_in[1]), .A0_f (new_AGEMA_signal_948), .B0_t (Inc_in[0]), .B0_f (new_AGEMA_signal_947), .Z0_t (Inc_Reg[1]), .Z0_f (new_AGEMA_signal_933) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1), .NL(1'b0)) U13 ( .A0_t (n9), .A0_f (new_AGEMA_signal_951), .B0_t (Inc_in[2]), .B0_f (new_AGEMA_signal_949), .Z0_t (Inc_Reg[2]), .Z0_f (new_AGEMA_signal_936) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) U14 ( .A0_t (n9), .A0_f (new_AGEMA_signal_951), .B0_t (Inc_in[2]), .B0_f (new_AGEMA_signal_949), .Z0_t (n10), .Z0_f (new_AGEMA_signal_952) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b0)) U15 ( .A0_t (Inc_in[3]), .A0_f (new_AGEMA_signal_950), .B0_t (n10), .B0_f (new_AGEMA_signal_952), .Z0_t (Inc_out[3]), .Z0_f (new_AGEMA_signal_953) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1), .NL(1'b0)) new_AGEMA_gate_182 ( .A0_t (Inc_in[0]), .A0_f (new_AGEMA_signal_947), .B0_t (1'b0), .B0_f (1'b1), .Z0_t (Inc_Reg[0]), .Z0_f (new_AGEMA_signal_930) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1), .NL(1'b0)) new_AGEMA_gate_183 ( .A0_t (Inc_out[3]), .A0_f (new_AGEMA_signal_953), .B0_t (1'b0), .B0_f (1'b1), .Z0_t (Inc_Reg[3]), .Z0_f (new_AGEMA_signal_939) ) ;

    /* register cells */
endmodule
