module eFPGA_top
    #(
        parameter include_eFPGA=1,
        parameter NumberOfRows=60,
        parameter NumberOfCols=39,
        parameter FrameBitsPerRow=32,
        parameter MaxFramesPerCol=20,
        parameter desync_flag=20,
        parameter FrameSelectWidth=7,
        parameter RowSelectWidth=7
    )
    (
        //External IO port
        output [240-1:0] A_config_C,
        output [240-1:0] B_config_C,
        output [60-1:0] I_top_0_t,
        output [60-1:0] I_top_0_f,
        output [60-1:0] I_top_1_t,
        output [60-1:0] I_top_1_f,
        output [60-1:0] T_top,
        input [60-1:0] O_top_0_t,
        input [60-1:0] O_top_0_f,
        input [60-1:0] O_top_1_t,
        input [60-1:0] O_top_1_f,
        output [60-1:0] ctrl_I_top_0_t,
        output [60-1:0] ctrl_I_top_0_f,
        output [60-1:0] ctrl_T_top,
        input [60-1:0] ctrl_O_top_0_t,
        input [60-1:0] ctrl_O_top_0_f,

        //Custom ports (*SAUBER*)
        input rst,
        output f_detected,
        output prech1,
        output prech2,
        input prng_rst,
        input [79:0] key_t,
        input [79:0] key_f,
        input [79:0] iv_t,
        input [79:0] iv_f,

        //Config related ports
        input CLK,
        input resetn,
        input SelfWriteStrobe,
        input [31:0] SelfWriteData,
        input Rx,
        output ComActive,
        output ReceiveLED,
        input s_clk,
        input s_data
);

 //Custom signal declarations for SAUBER
wire[59:0] F_masked1_top;
wire[59:0] F_masked2_top;
wire[59:0] F_ctrl_top;
wire[1499:0] R_t_top;
wire[1499:0] R_f_top;


 //Signal declarations
wire[(NumberOfRows*FrameBitsPerRow)-1:0] FrameRegister;
wire[(MaxFramesPerCol*NumberOfCols)-1:0] FrameSelect;
wire[(FrameBitsPerRow*(NumberOfRows+2))-1:0] FrameData;
wire[FrameBitsPerRow-1:0] FrameAddressRegister;
wire LongFrameStrobe;
wire[31:0] LocalWriteData;
wire LocalWriteStrobe;
wire[RowSelectWidth-1:0] RowSelect;
wire resten;
`ifndef EMULATION

eFPGA_Config
    #(
    .RowSelectWidth(RowSelectWidth),
    .NumberOfRows(NumberOfRows),
    .desync_flag(desync_flag),
    .FrameBitsPerRow(FrameBitsPerRow)
    )
    eFPGA_Config_inst
    (
    .CLK(CLK),
    .resetn(resetn),
    .Rx(Rx),
    .ComActive(ComActive),
    .ReceiveLED(ReceiveLED),
    .s_clk(s_clk),
    .s_data(s_data),
    .SelfWriteData(SelfWriteData),
    .SelfWriteStrobe(SelfWriteStrobe),
    .ConfigWriteData(LocalWriteData),
    .ConfigWriteStrobe(LocalWriteStrobe),
    .FrameAddressRegister(FrameAddressRegister),
    .LongFrameStrobe(LongFrameStrobe),
    .RowSelect(RowSelect)
);


Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(1)
    )
    inst_Frame_Data_Reg_0
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[0*FrameBitsPerRow+FrameBitsPerRow-1:0*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(2)
    )
    inst_Frame_Data_Reg_1
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[1*FrameBitsPerRow+FrameBitsPerRow-1:1*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(3)
    )
    inst_Frame_Data_Reg_2
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[2*FrameBitsPerRow+FrameBitsPerRow-1:2*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(4)
    )
    inst_Frame_Data_Reg_3
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[3*FrameBitsPerRow+FrameBitsPerRow-1:3*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(5)
    )
    inst_Frame_Data_Reg_4
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[4*FrameBitsPerRow+FrameBitsPerRow-1:4*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(6)
    )
    inst_Frame_Data_Reg_5
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[5*FrameBitsPerRow+FrameBitsPerRow-1:5*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(7)
    )
    inst_Frame_Data_Reg_6
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[6*FrameBitsPerRow+FrameBitsPerRow-1:6*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(8)
    )
    inst_Frame_Data_Reg_7
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[7*FrameBitsPerRow+FrameBitsPerRow-1:7*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(9)
    )
    inst_Frame_Data_Reg_8
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[8*FrameBitsPerRow+FrameBitsPerRow-1:8*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(10)
    )
    inst_Frame_Data_Reg_9
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[9*FrameBitsPerRow+FrameBitsPerRow-1:9*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(11)
    )
    inst_Frame_Data_Reg_10
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[10*FrameBitsPerRow+FrameBitsPerRow-1:10*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(12)
    )
    inst_Frame_Data_Reg_11
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[11*FrameBitsPerRow+FrameBitsPerRow-1:11*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(13)
    )
    inst_Frame_Data_Reg_12
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[12*FrameBitsPerRow+FrameBitsPerRow-1:12*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(14)
    )
    inst_Frame_Data_Reg_13
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[13*FrameBitsPerRow+FrameBitsPerRow-1:13*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(15)
    )
    inst_Frame_Data_Reg_14
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[14*FrameBitsPerRow+FrameBitsPerRow-1:14*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(16)
    )
    inst_Frame_Data_Reg_15
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[15*FrameBitsPerRow+FrameBitsPerRow-1:15*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(17)
    )
    inst_Frame_Data_Reg_16
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[16*FrameBitsPerRow+FrameBitsPerRow-1:16*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(18)
    )
    inst_Frame_Data_Reg_17
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[17*FrameBitsPerRow+FrameBitsPerRow-1:17*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(19)
    )
    inst_Frame_Data_Reg_18
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[18*FrameBitsPerRow+FrameBitsPerRow-1:18*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(20)
    )
    inst_Frame_Data_Reg_19
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[19*FrameBitsPerRow+FrameBitsPerRow-1:19*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(21)
    )
    inst_Frame_Data_Reg_20
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[20*FrameBitsPerRow+FrameBitsPerRow-1:20*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(22)
    )
    inst_Frame_Data_Reg_21
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[21*FrameBitsPerRow+FrameBitsPerRow-1:21*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(23)
    )
    inst_Frame_Data_Reg_22
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[22*FrameBitsPerRow+FrameBitsPerRow-1:22*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(24)
    )
    inst_Frame_Data_Reg_23
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[23*FrameBitsPerRow+FrameBitsPerRow-1:23*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(25)
    )
    inst_Frame_Data_Reg_24
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[24*FrameBitsPerRow+FrameBitsPerRow-1:24*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(26)
    )
    inst_Frame_Data_Reg_25
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[25*FrameBitsPerRow+FrameBitsPerRow-1:25*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(27)
    )
    inst_Frame_Data_Reg_26
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[26*FrameBitsPerRow+FrameBitsPerRow-1:26*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(28)
    )
    inst_Frame_Data_Reg_27
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[27*FrameBitsPerRow+FrameBitsPerRow-1:27*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(29)
    )
    inst_Frame_Data_Reg_28
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[28*FrameBitsPerRow+FrameBitsPerRow-1:28*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(30)
    )
    inst_Frame_Data_Reg_29
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[29*FrameBitsPerRow+FrameBitsPerRow-1:29*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(31)
    )
    inst_Frame_Data_Reg_30
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[30*FrameBitsPerRow+FrameBitsPerRow-1:30*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(32)
    )
    inst_Frame_Data_Reg_31
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[31*FrameBitsPerRow+FrameBitsPerRow-1:31*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(33)
    )
    inst_Frame_Data_Reg_32
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[32*FrameBitsPerRow+FrameBitsPerRow-1:32*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(34)
    )
    inst_Frame_Data_Reg_33
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[33*FrameBitsPerRow+FrameBitsPerRow-1:33*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(35)
    )
    inst_Frame_Data_Reg_34
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[34*FrameBitsPerRow+FrameBitsPerRow-1:34*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(36)
    )
    inst_Frame_Data_Reg_35
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[35*FrameBitsPerRow+FrameBitsPerRow-1:35*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(37)
    )
    inst_Frame_Data_Reg_36
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[36*FrameBitsPerRow+FrameBitsPerRow-1:36*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(38)
    )
    inst_Frame_Data_Reg_37
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[37*FrameBitsPerRow+FrameBitsPerRow-1:37*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(39)
    )
    inst_Frame_Data_Reg_38
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[38*FrameBitsPerRow+FrameBitsPerRow-1:38*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(40)
    )
    inst_Frame_Data_Reg_39
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[39*FrameBitsPerRow+FrameBitsPerRow-1:39*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(41)
    )
    inst_Frame_Data_Reg_40
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[40*FrameBitsPerRow+FrameBitsPerRow-1:40*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(42)
    )
    inst_Frame_Data_Reg_41
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[41*FrameBitsPerRow+FrameBitsPerRow-1:41*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(43)
    )
    inst_Frame_Data_Reg_42
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[42*FrameBitsPerRow+FrameBitsPerRow-1:42*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(44)
    )
    inst_Frame_Data_Reg_43
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[43*FrameBitsPerRow+FrameBitsPerRow-1:43*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(45)
    )
    inst_Frame_Data_Reg_44
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[44*FrameBitsPerRow+FrameBitsPerRow-1:44*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(46)
    )
    inst_Frame_Data_Reg_45
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[45*FrameBitsPerRow+FrameBitsPerRow-1:45*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(47)
    )
    inst_Frame_Data_Reg_46
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[46*FrameBitsPerRow+FrameBitsPerRow-1:46*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(48)
    )
    inst_Frame_Data_Reg_47
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[47*FrameBitsPerRow+FrameBitsPerRow-1:47*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(49)
    )
    inst_Frame_Data_Reg_48
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[48*FrameBitsPerRow+FrameBitsPerRow-1:48*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(50)
    )
    inst_Frame_Data_Reg_49
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[49*FrameBitsPerRow+FrameBitsPerRow-1:49*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(51)
    )
    inst_Frame_Data_Reg_50
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[50*FrameBitsPerRow+FrameBitsPerRow-1:50*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(52)
    )
    inst_Frame_Data_Reg_51
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[51*FrameBitsPerRow+FrameBitsPerRow-1:51*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(53)
    )
    inst_Frame_Data_Reg_52
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[52*FrameBitsPerRow+FrameBitsPerRow-1:52*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(54)
    )
    inst_Frame_Data_Reg_53
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[53*FrameBitsPerRow+FrameBitsPerRow-1:53*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(55)
    )
    inst_Frame_Data_Reg_54
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[54*FrameBitsPerRow+FrameBitsPerRow-1:54*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(56)
    )
    inst_Frame_Data_Reg_55
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[55*FrameBitsPerRow+FrameBitsPerRow-1:55*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(57)
    )
    inst_Frame_Data_Reg_56
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[56*FrameBitsPerRow+FrameBitsPerRow-1:56*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(58)
    )
    inst_Frame_Data_Reg_57
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[57*FrameBitsPerRow+FrameBitsPerRow-1:57*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(59)
    )
    inst_Frame_Data_Reg_58
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[58*FrameBitsPerRow+FrameBitsPerRow-1:58*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);

Frame_Data_Reg
    #(
    .FrameBitsPerRow(FrameBitsPerRow),
    .RowSelectWidth(RowSelectWidth),
    .Row(60)
    )
    inst_Frame_Data_Reg_59
    (
    .FrameData_I(LocalWriteData),
    .FrameData_O(FrameRegister[59*FrameBitsPerRow+FrameBitsPerRow-1:59*FrameBitsPerRow]),
    .RowSelect(RowSelect),
    .CLK(CLK)
);


Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(0)
    )
    inst_Frame_Select_0
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[0*MaxFramesPerCol+MaxFramesPerCol-1:0*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(1)
    )
    inst_Frame_Select_1
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[1*MaxFramesPerCol+MaxFramesPerCol-1:1*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(2)
    )
    inst_Frame_Select_2
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[2*MaxFramesPerCol+MaxFramesPerCol-1:2*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(3)
    )
    inst_Frame_Select_3
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[3*MaxFramesPerCol+MaxFramesPerCol-1:3*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(4)
    )
    inst_Frame_Select_4
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[4*MaxFramesPerCol+MaxFramesPerCol-1:4*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(5)
    )
    inst_Frame_Select_5
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[5*MaxFramesPerCol+MaxFramesPerCol-1:5*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(6)
    )
    inst_Frame_Select_6
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[6*MaxFramesPerCol+MaxFramesPerCol-1:6*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(7)
    )
    inst_Frame_Select_7
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[7*MaxFramesPerCol+MaxFramesPerCol-1:7*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(8)
    )
    inst_Frame_Select_8
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[8*MaxFramesPerCol+MaxFramesPerCol-1:8*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(9)
    )
    inst_Frame_Select_9
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[9*MaxFramesPerCol+MaxFramesPerCol-1:9*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(10)
    )
    inst_Frame_Select_10
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[10*MaxFramesPerCol+MaxFramesPerCol-1:10*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(11)
    )
    inst_Frame_Select_11
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[11*MaxFramesPerCol+MaxFramesPerCol-1:11*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(12)
    )
    inst_Frame_Select_12
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[12*MaxFramesPerCol+MaxFramesPerCol-1:12*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(13)
    )
    inst_Frame_Select_13
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[13*MaxFramesPerCol+MaxFramesPerCol-1:13*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(14)
    )
    inst_Frame_Select_14
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[14*MaxFramesPerCol+MaxFramesPerCol-1:14*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(15)
    )
    inst_Frame_Select_15
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[15*MaxFramesPerCol+MaxFramesPerCol-1:15*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(16)
    )
    inst_Frame_Select_16
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[16*MaxFramesPerCol+MaxFramesPerCol-1:16*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(17)
    )
    inst_Frame_Select_17
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[17*MaxFramesPerCol+MaxFramesPerCol-1:17*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(18)
    )
    inst_Frame_Select_18
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[18*MaxFramesPerCol+MaxFramesPerCol-1:18*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(19)
    )
    inst_Frame_Select_19
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[19*MaxFramesPerCol+MaxFramesPerCol-1:19*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(20)
    )
    inst_Frame_Select_20
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[20*MaxFramesPerCol+MaxFramesPerCol-1:20*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(21)
    )
    inst_Frame_Select_21
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[21*MaxFramesPerCol+MaxFramesPerCol-1:21*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(22)
    )
    inst_Frame_Select_22
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[22*MaxFramesPerCol+MaxFramesPerCol-1:22*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(23)
    )
    inst_Frame_Select_23
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[23*MaxFramesPerCol+MaxFramesPerCol-1:23*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(24)
    )
    inst_Frame_Select_24
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[24*MaxFramesPerCol+MaxFramesPerCol-1:24*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(25)
    )
    inst_Frame_Select_25
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[25*MaxFramesPerCol+MaxFramesPerCol-1:25*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(26)
    )
    inst_Frame_Select_26
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[26*MaxFramesPerCol+MaxFramesPerCol-1:26*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(27)
    )
    inst_Frame_Select_27
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[27*MaxFramesPerCol+MaxFramesPerCol-1:27*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(28)
    )
    inst_Frame_Select_28
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[28*MaxFramesPerCol+MaxFramesPerCol-1:28*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(29)
    )
    inst_Frame_Select_29
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[29*MaxFramesPerCol+MaxFramesPerCol-1:29*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(30)
    )
    inst_Frame_Select_30
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[30*MaxFramesPerCol+MaxFramesPerCol-1:30*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(31)
    )
    inst_Frame_Select_31
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[31*MaxFramesPerCol+MaxFramesPerCol-1:31*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(32)
    )
    inst_Frame_Select_32
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[32*MaxFramesPerCol+MaxFramesPerCol-1:32*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(33)
    )
    inst_Frame_Select_33
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[33*MaxFramesPerCol+MaxFramesPerCol-1:33*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(34)
    )
    inst_Frame_Select_34
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[34*MaxFramesPerCol+MaxFramesPerCol-1:34*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(35)
    )
    inst_Frame_Select_35
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[35*MaxFramesPerCol+MaxFramesPerCol-1:35*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(36)
    )
    inst_Frame_Select_36
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[36*MaxFramesPerCol+MaxFramesPerCol-1:36*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(37)
    )
    inst_Frame_Select_37
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[37*MaxFramesPerCol+MaxFramesPerCol-1:37*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);

Frame_Select
    #(
    .MaxFramesPerCol(MaxFramesPerCol),
    .FrameSelectWidth(FrameSelectWidth),
    .Col(38)
    )
    inst_Frame_Select_38
    (
    .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
    .FrameStrobe_O(FrameSelect[38*MaxFramesPerCol+MaxFramesPerCol-1:38*MaxFramesPerCol]),
    .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
    .FrameStrobe(LongFrameStrobe)
);


`endif
eFPGA eFPGA_inst (
    .Tile_X3Y1_R_t(R_t_top[0]),
    .Tile_X3Y1_R_f(R_f_top[0]),
    .Tile_X6Y1_R_t(R_t_top[1]),
    .Tile_X6Y1_R_f(R_f_top[1]),
    .Tile_X9Y1_R_t(R_t_top[2]),
    .Tile_X9Y1_R_f(R_f_top[2]),
    .Tile_X12Y1_R_t(R_t_top[3]),
    .Tile_X12Y1_R_f(R_f_top[3]),
    .Tile_X15Y1_R_t(R_t_top[4]),
    .Tile_X15Y1_R_f(R_f_top[4]),
    .Tile_X18Y1_R_t(R_t_top[5]),
    .Tile_X18Y1_R_f(R_f_top[5]),
    .Tile_X21Y1_R_t(R_t_top[6]),
    .Tile_X21Y1_R_f(R_f_top[6]),
    .Tile_X24Y1_R_t(R_t_top[7]),
    .Tile_X24Y1_R_f(R_f_top[7]),
    .Tile_X27Y1_R_t(R_t_top[8]),
    .Tile_X27Y1_R_f(R_f_top[8]),
    .Tile_X30Y1_R_t(R_t_top[9]),
    .Tile_X30Y1_R_f(R_f_top[9]),
    .Tile_X33Y1_R_t(R_t_top[10]),
    .Tile_X33Y1_R_f(R_f_top[10]),
    .Tile_X36Y1_R_t(R_t_top[11]),
    .Tile_X36Y1_R_f(R_f_top[11]),
    .Tile_X39Y1_R_t(R_t_top[12]),
    .Tile_X39Y1_R_f(R_f_top[12]),
    .Tile_X42Y1_R_t(R_t_top[13]),
    .Tile_X42Y1_R_f(R_f_top[13]),
    .Tile_X45Y1_R_t(R_t_top[14]),
    .Tile_X45Y1_R_f(R_f_top[14]),
    .Tile_X48Y1_R_t(R_t_top[15]),
    .Tile_X48Y1_R_f(R_f_top[15]),
    .Tile_X51Y1_R_t(R_t_top[16]),
    .Tile_X51Y1_R_f(R_f_top[16]),
    .Tile_X54Y1_R_t(R_t_top[17]),
    .Tile_X54Y1_R_f(R_f_top[17]),
    .Tile_X57Y1_R_t(R_t_top[18]),
    .Tile_X57Y1_R_f(R_f_top[18]),
    .Tile_X60Y1_R_t(R_t_top[19]),
    .Tile_X60Y1_R_f(R_f_top[19]),
    .Tile_X63Y1_R_t(R_t_top[20]),
    .Tile_X63Y1_R_f(R_f_top[20]),
    .Tile_X66Y1_R_t(R_t_top[21]),
    .Tile_X66Y1_R_f(R_f_top[21]),
    .Tile_X69Y1_R_t(R_t_top[22]),
    .Tile_X69Y1_R_f(R_f_top[22]),
    .Tile_X72Y1_R_t(R_t_top[23]),
    .Tile_X72Y1_R_f(R_f_top[23]),
    .Tile_X75Y1_R_t(R_t_top[24]),
    .Tile_X75Y1_R_f(R_f_top[24]),
    .Tile_X3Y2_R_t(R_t_top[25]),
    .Tile_X3Y2_R_f(R_f_top[25]),
    .Tile_X6Y2_R_t(R_t_top[26]),
    .Tile_X6Y2_R_f(R_f_top[26]),
    .Tile_X9Y2_R_t(R_t_top[27]),
    .Tile_X9Y2_R_f(R_f_top[27]),
    .Tile_X12Y2_R_t(R_t_top[28]),
    .Tile_X12Y2_R_f(R_f_top[28]),
    .Tile_X15Y2_R_t(R_t_top[29]),
    .Tile_X15Y2_R_f(R_f_top[29]),
    .Tile_X18Y2_R_t(R_t_top[30]),
    .Tile_X18Y2_R_f(R_f_top[30]),
    .Tile_X21Y2_R_t(R_t_top[31]),
    .Tile_X21Y2_R_f(R_f_top[31]),
    .Tile_X24Y2_R_t(R_t_top[32]),
    .Tile_X24Y2_R_f(R_f_top[32]),
    .Tile_X27Y2_R_t(R_t_top[33]),
    .Tile_X27Y2_R_f(R_f_top[33]),
    .Tile_X30Y2_R_t(R_t_top[34]),
    .Tile_X30Y2_R_f(R_f_top[34]),
    .Tile_X33Y2_R_t(R_t_top[35]),
    .Tile_X33Y2_R_f(R_f_top[35]),
    .Tile_X36Y2_R_t(R_t_top[36]),
    .Tile_X36Y2_R_f(R_f_top[36]),
    .Tile_X39Y2_R_t(R_t_top[37]),
    .Tile_X39Y2_R_f(R_f_top[37]),
    .Tile_X42Y2_R_t(R_t_top[38]),
    .Tile_X42Y2_R_f(R_f_top[38]),
    .Tile_X45Y2_R_t(R_t_top[39]),
    .Tile_X45Y2_R_f(R_f_top[39]),
    .Tile_X48Y2_R_t(R_t_top[40]),
    .Tile_X48Y2_R_f(R_f_top[40]),
    .Tile_X51Y2_R_t(R_t_top[41]),
    .Tile_X51Y2_R_f(R_f_top[41]),
    .Tile_X54Y2_R_t(R_t_top[42]),
    .Tile_X54Y2_R_f(R_f_top[42]),
    .Tile_X57Y2_R_t(R_t_top[43]),
    .Tile_X57Y2_R_f(R_f_top[43]),
    .Tile_X60Y2_R_t(R_t_top[44]),
    .Tile_X60Y2_R_f(R_f_top[44]),
    .Tile_X63Y2_R_t(R_t_top[45]),
    .Tile_X63Y2_R_f(R_f_top[45]),
    .Tile_X66Y2_R_t(R_t_top[46]),
    .Tile_X66Y2_R_f(R_f_top[46]),
    .Tile_X69Y2_R_t(R_t_top[47]),
    .Tile_X69Y2_R_f(R_f_top[47]),
    .Tile_X72Y2_R_t(R_t_top[48]),
    .Tile_X72Y2_R_f(R_f_top[48]),
    .Tile_X75Y2_R_t(R_t_top[49]),
    .Tile_X75Y2_R_f(R_f_top[49]),
    .Tile_X3Y3_R_t(R_t_top[50]),
    .Tile_X3Y3_R_f(R_f_top[50]),
    .Tile_X6Y3_R_t(R_t_top[51]),
    .Tile_X6Y3_R_f(R_f_top[51]),
    .Tile_X9Y3_R_t(R_t_top[52]),
    .Tile_X9Y3_R_f(R_f_top[52]),
    .Tile_X12Y3_R_t(R_t_top[53]),
    .Tile_X12Y3_R_f(R_f_top[53]),
    .Tile_X15Y3_R_t(R_t_top[54]),
    .Tile_X15Y3_R_f(R_f_top[54]),
    .Tile_X18Y3_R_t(R_t_top[55]),
    .Tile_X18Y3_R_f(R_f_top[55]),
    .Tile_X21Y3_R_t(R_t_top[56]),
    .Tile_X21Y3_R_f(R_f_top[56]),
    .Tile_X24Y3_R_t(R_t_top[57]),
    .Tile_X24Y3_R_f(R_f_top[57]),
    .Tile_X27Y3_R_t(R_t_top[58]),
    .Tile_X27Y3_R_f(R_f_top[58]),
    .Tile_X30Y3_R_t(R_t_top[59]),
    .Tile_X30Y3_R_f(R_f_top[59]),
    .Tile_X33Y3_R_t(R_t_top[60]),
    .Tile_X33Y3_R_f(R_f_top[60]),
    .Tile_X36Y3_R_t(R_t_top[61]),
    .Tile_X36Y3_R_f(R_f_top[61]),
    .Tile_X39Y3_R_t(R_t_top[62]),
    .Tile_X39Y3_R_f(R_f_top[62]),
    .Tile_X42Y3_R_t(R_t_top[63]),
    .Tile_X42Y3_R_f(R_f_top[63]),
    .Tile_X45Y3_R_t(R_t_top[64]),
    .Tile_X45Y3_R_f(R_f_top[64]),
    .Tile_X48Y3_R_t(R_t_top[65]),
    .Tile_X48Y3_R_f(R_f_top[65]),
    .Tile_X51Y3_R_t(R_t_top[66]),
    .Tile_X51Y3_R_f(R_f_top[66]),
    .Tile_X54Y3_R_t(R_t_top[67]),
    .Tile_X54Y3_R_f(R_f_top[67]),
    .Tile_X57Y3_R_t(R_t_top[68]),
    .Tile_X57Y3_R_f(R_f_top[68]),
    .Tile_X60Y3_R_t(R_t_top[69]),
    .Tile_X60Y3_R_f(R_f_top[69]),
    .Tile_X63Y3_R_t(R_t_top[70]),
    .Tile_X63Y3_R_f(R_f_top[70]),
    .Tile_X66Y3_R_t(R_t_top[71]),
    .Tile_X66Y3_R_f(R_f_top[71]),
    .Tile_X69Y3_R_t(R_t_top[72]),
    .Tile_X69Y3_R_f(R_f_top[72]),
    .Tile_X72Y3_R_t(R_t_top[73]),
    .Tile_X72Y3_R_f(R_f_top[73]),
    .Tile_X75Y3_R_t(R_t_top[74]),
    .Tile_X75Y3_R_f(R_f_top[74]),
    .Tile_X3Y4_R_t(R_t_top[75]),
    .Tile_X3Y4_R_f(R_f_top[75]),
    .Tile_X6Y4_R_t(R_t_top[76]),
    .Tile_X6Y4_R_f(R_f_top[76]),
    .Tile_X9Y4_R_t(R_t_top[77]),
    .Tile_X9Y4_R_f(R_f_top[77]),
    .Tile_X12Y4_R_t(R_t_top[78]),
    .Tile_X12Y4_R_f(R_f_top[78]),
    .Tile_X15Y4_R_t(R_t_top[79]),
    .Tile_X15Y4_R_f(R_f_top[79]),
    .Tile_X18Y4_R_t(R_t_top[80]),
    .Tile_X18Y4_R_f(R_f_top[80]),
    .Tile_X21Y4_R_t(R_t_top[81]),
    .Tile_X21Y4_R_f(R_f_top[81]),
    .Tile_X24Y4_R_t(R_t_top[82]),
    .Tile_X24Y4_R_f(R_f_top[82]),
    .Tile_X27Y4_R_t(R_t_top[83]),
    .Tile_X27Y4_R_f(R_f_top[83]),
    .Tile_X30Y4_R_t(R_t_top[84]),
    .Tile_X30Y4_R_f(R_f_top[84]),
    .Tile_X33Y4_R_t(R_t_top[85]),
    .Tile_X33Y4_R_f(R_f_top[85]),
    .Tile_X36Y4_R_t(R_t_top[86]),
    .Tile_X36Y4_R_f(R_f_top[86]),
    .Tile_X39Y4_R_t(R_t_top[87]),
    .Tile_X39Y4_R_f(R_f_top[87]),
    .Tile_X42Y4_R_t(R_t_top[88]),
    .Tile_X42Y4_R_f(R_f_top[88]),
    .Tile_X45Y4_R_t(R_t_top[89]),
    .Tile_X45Y4_R_f(R_f_top[89]),
    .Tile_X48Y4_R_t(R_t_top[90]),
    .Tile_X48Y4_R_f(R_f_top[90]),
    .Tile_X51Y4_R_t(R_t_top[91]),
    .Tile_X51Y4_R_f(R_f_top[91]),
    .Tile_X54Y4_R_t(R_t_top[92]),
    .Tile_X54Y4_R_f(R_f_top[92]),
    .Tile_X57Y4_R_t(R_t_top[93]),
    .Tile_X57Y4_R_f(R_f_top[93]),
    .Tile_X60Y4_R_t(R_t_top[94]),
    .Tile_X60Y4_R_f(R_f_top[94]),
    .Tile_X63Y4_R_t(R_t_top[95]),
    .Tile_X63Y4_R_f(R_f_top[95]),
    .Tile_X66Y4_R_t(R_t_top[96]),
    .Tile_X66Y4_R_f(R_f_top[96]),
    .Tile_X69Y4_R_t(R_t_top[97]),
    .Tile_X69Y4_R_f(R_f_top[97]),
    .Tile_X72Y4_R_t(R_t_top[98]),
    .Tile_X72Y4_R_f(R_f_top[98]),
    .Tile_X75Y4_R_t(R_t_top[99]),
    .Tile_X75Y4_R_f(R_f_top[99]),
    .Tile_X3Y5_R_t(R_t_top[100]),
    .Tile_X3Y5_R_f(R_f_top[100]),
    .Tile_X6Y5_R_t(R_t_top[101]),
    .Tile_X6Y5_R_f(R_f_top[101]),
    .Tile_X9Y5_R_t(R_t_top[102]),
    .Tile_X9Y5_R_f(R_f_top[102]),
    .Tile_X12Y5_R_t(R_t_top[103]),
    .Tile_X12Y5_R_f(R_f_top[103]),
    .Tile_X15Y5_R_t(R_t_top[104]),
    .Tile_X15Y5_R_f(R_f_top[104]),
    .Tile_X18Y5_R_t(R_t_top[105]),
    .Tile_X18Y5_R_f(R_f_top[105]),
    .Tile_X21Y5_R_t(R_t_top[106]),
    .Tile_X21Y5_R_f(R_f_top[106]),
    .Tile_X24Y5_R_t(R_t_top[107]),
    .Tile_X24Y5_R_f(R_f_top[107]),
    .Tile_X27Y5_R_t(R_t_top[108]),
    .Tile_X27Y5_R_f(R_f_top[108]),
    .Tile_X30Y5_R_t(R_t_top[109]),
    .Tile_X30Y5_R_f(R_f_top[109]),
    .Tile_X33Y5_R_t(R_t_top[110]),
    .Tile_X33Y5_R_f(R_f_top[110]),
    .Tile_X36Y5_R_t(R_t_top[111]),
    .Tile_X36Y5_R_f(R_f_top[111]),
    .Tile_X39Y5_R_t(R_t_top[112]),
    .Tile_X39Y5_R_f(R_f_top[112]),
    .Tile_X42Y5_R_t(R_t_top[113]),
    .Tile_X42Y5_R_f(R_f_top[113]),
    .Tile_X45Y5_R_t(R_t_top[114]),
    .Tile_X45Y5_R_f(R_f_top[114]),
    .Tile_X48Y5_R_t(R_t_top[115]),
    .Tile_X48Y5_R_f(R_f_top[115]),
    .Tile_X51Y5_R_t(R_t_top[116]),
    .Tile_X51Y5_R_f(R_f_top[116]),
    .Tile_X54Y5_R_t(R_t_top[117]),
    .Tile_X54Y5_R_f(R_f_top[117]),
    .Tile_X57Y5_R_t(R_t_top[118]),
    .Tile_X57Y5_R_f(R_f_top[118]),
    .Tile_X60Y5_R_t(R_t_top[119]),
    .Tile_X60Y5_R_f(R_f_top[119]),
    .Tile_X63Y5_R_t(R_t_top[120]),
    .Tile_X63Y5_R_f(R_f_top[120]),
    .Tile_X66Y5_R_t(R_t_top[121]),
    .Tile_X66Y5_R_f(R_f_top[121]),
    .Tile_X69Y5_R_t(R_t_top[122]),
    .Tile_X69Y5_R_f(R_f_top[122]),
    .Tile_X72Y5_R_t(R_t_top[123]),
    .Tile_X72Y5_R_f(R_f_top[123]),
    .Tile_X75Y5_R_t(R_t_top[124]),
    .Tile_X75Y5_R_f(R_f_top[124]),
    .Tile_X3Y6_R_t(R_t_top[125]),
    .Tile_X3Y6_R_f(R_f_top[125]),
    .Tile_X6Y6_R_t(R_t_top[126]),
    .Tile_X6Y6_R_f(R_f_top[126]),
    .Tile_X9Y6_R_t(R_t_top[127]),
    .Tile_X9Y6_R_f(R_f_top[127]),
    .Tile_X12Y6_R_t(R_t_top[128]),
    .Tile_X12Y6_R_f(R_f_top[128]),
    .Tile_X15Y6_R_t(R_t_top[129]),
    .Tile_X15Y6_R_f(R_f_top[129]),
    .Tile_X18Y6_R_t(R_t_top[130]),
    .Tile_X18Y6_R_f(R_f_top[130]),
    .Tile_X21Y6_R_t(R_t_top[131]),
    .Tile_X21Y6_R_f(R_f_top[131]),
    .Tile_X24Y6_R_t(R_t_top[132]),
    .Tile_X24Y6_R_f(R_f_top[132]),
    .Tile_X27Y6_R_t(R_t_top[133]),
    .Tile_X27Y6_R_f(R_f_top[133]),
    .Tile_X30Y6_R_t(R_t_top[134]),
    .Tile_X30Y6_R_f(R_f_top[134]),
    .Tile_X33Y6_R_t(R_t_top[135]),
    .Tile_X33Y6_R_f(R_f_top[135]),
    .Tile_X36Y6_R_t(R_t_top[136]),
    .Tile_X36Y6_R_f(R_f_top[136]),
    .Tile_X39Y6_R_t(R_t_top[137]),
    .Tile_X39Y6_R_f(R_f_top[137]),
    .Tile_X42Y6_R_t(R_t_top[138]),
    .Tile_X42Y6_R_f(R_f_top[138]),
    .Tile_X45Y6_R_t(R_t_top[139]),
    .Tile_X45Y6_R_f(R_f_top[139]),
    .Tile_X48Y6_R_t(R_t_top[140]),
    .Tile_X48Y6_R_f(R_f_top[140]),
    .Tile_X51Y6_R_t(R_t_top[141]),
    .Tile_X51Y6_R_f(R_f_top[141]),
    .Tile_X54Y6_R_t(R_t_top[142]),
    .Tile_X54Y6_R_f(R_f_top[142]),
    .Tile_X57Y6_R_t(R_t_top[143]),
    .Tile_X57Y6_R_f(R_f_top[143]),
    .Tile_X60Y6_R_t(R_t_top[144]),
    .Tile_X60Y6_R_f(R_f_top[144]),
    .Tile_X63Y6_R_t(R_t_top[145]),
    .Tile_X63Y6_R_f(R_f_top[145]),
    .Tile_X66Y6_R_t(R_t_top[146]),
    .Tile_X66Y6_R_f(R_f_top[146]),
    .Tile_X69Y6_R_t(R_t_top[147]),
    .Tile_X69Y6_R_f(R_f_top[147]),
    .Tile_X72Y6_R_t(R_t_top[148]),
    .Tile_X72Y6_R_f(R_f_top[148]),
    .Tile_X75Y6_R_t(R_t_top[149]),
    .Tile_X75Y6_R_f(R_f_top[149]),
    .Tile_X3Y7_R_t(R_t_top[150]),
    .Tile_X3Y7_R_f(R_f_top[150]),
    .Tile_X6Y7_R_t(R_t_top[151]),
    .Tile_X6Y7_R_f(R_f_top[151]),
    .Tile_X9Y7_R_t(R_t_top[152]),
    .Tile_X9Y7_R_f(R_f_top[152]),
    .Tile_X12Y7_R_t(R_t_top[153]),
    .Tile_X12Y7_R_f(R_f_top[153]),
    .Tile_X15Y7_R_t(R_t_top[154]),
    .Tile_X15Y7_R_f(R_f_top[154]),
    .Tile_X18Y7_R_t(R_t_top[155]),
    .Tile_X18Y7_R_f(R_f_top[155]),
    .Tile_X21Y7_R_t(R_t_top[156]),
    .Tile_X21Y7_R_f(R_f_top[156]),
    .Tile_X24Y7_R_t(R_t_top[157]),
    .Tile_X24Y7_R_f(R_f_top[157]),
    .Tile_X27Y7_R_t(R_t_top[158]),
    .Tile_X27Y7_R_f(R_f_top[158]),
    .Tile_X30Y7_R_t(R_t_top[159]),
    .Tile_X30Y7_R_f(R_f_top[159]),
    .Tile_X33Y7_R_t(R_t_top[160]),
    .Tile_X33Y7_R_f(R_f_top[160]),
    .Tile_X36Y7_R_t(R_t_top[161]),
    .Tile_X36Y7_R_f(R_f_top[161]),
    .Tile_X39Y7_R_t(R_t_top[162]),
    .Tile_X39Y7_R_f(R_f_top[162]),
    .Tile_X42Y7_R_t(R_t_top[163]),
    .Tile_X42Y7_R_f(R_f_top[163]),
    .Tile_X45Y7_R_t(R_t_top[164]),
    .Tile_X45Y7_R_f(R_f_top[164]),
    .Tile_X48Y7_R_t(R_t_top[165]),
    .Tile_X48Y7_R_f(R_f_top[165]),
    .Tile_X51Y7_R_t(R_t_top[166]),
    .Tile_X51Y7_R_f(R_f_top[166]),
    .Tile_X54Y7_R_t(R_t_top[167]),
    .Tile_X54Y7_R_f(R_f_top[167]),
    .Tile_X57Y7_R_t(R_t_top[168]),
    .Tile_X57Y7_R_f(R_f_top[168]),
    .Tile_X60Y7_R_t(R_t_top[169]),
    .Tile_X60Y7_R_f(R_f_top[169]),
    .Tile_X63Y7_R_t(R_t_top[170]),
    .Tile_X63Y7_R_f(R_f_top[170]),
    .Tile_X66Y7_R_t(R_t_top[171]),
    .Tile_X66Y7_R_f(R_f_top[171]),
    .Tile_X69Y7_R_t(R_t_top[172]),
    .Tile_X69Y7_R_f(R_f_top[172]),
    .Tile_X72Y7_R_t(R_t_top[173]),
    .Tile_X72Y7_R_f(R_f_top[173]),
    .Tile_X75Y7_R_t(R_t_top[174]),
    .Tile_X75Y7_R_f(R_f_top[174]),
    .Tile_X3Y8_R_t(R_t_top[175]),
    .Tile_X3Y8_R_f(R_f_top[175]),
    .Tile_X6Y8_R_t(R_t_top[176]),
    .Tile_X6Y8_R_f(R_f_top[176]),
    .Tile_X9Y8_R_t(R_t_top[177]),
    .Tile_X9Y8_R_f(R_f_top[177]),
    .Tile_X12Y8_R_t(R_t_top[178]),
    .Tile_X12Y8_R_f(R_f_top[178]),
    .Tile_X15Y8_R_t(R_t_top[179]),
    .Tile_X15Y8_R_f(R_f_top[179]),
    .Tile_X18Y8_R_t(R_t_top[180]),
    .Tile_X18Y8_R_f(R_f_top[180]),
    .Tile_X21Y8_R_t(R_t_top[181]),
    .Tile_X21Y8_R_f(R_f_top[181]),
    .Tile_X24Y8_R_t(R_t_top[182]),
    .Tile_X24Y8_R_f(R_f_top[182]),
    .Tile_X27Y8_R_t(R_t_top[183]),
    .Tile_X27Y8_R_f(R_f_top[183]),
    .Tile_X30Y8_R_t(R_t_top[184]),
    .Tile_X30Y8_R_f(R_f_top[184]),
    .Tile_X33Y8_R_t(R_t_top[185]),
    .Tile_X33Y8_R_f(R_f_top[185]),
    .Tile_X36Y8_R_t(R_t_top[186]),
    .Tile_X36Y8_R_f(R_f_top[186]),
    .Tile_X39Y8_R_t(R_t_top[187]),
    .Tile_X39Y8_R_f(R_f_top[187]),
    .Tile_X42Y8_R_t(R_t_top[188]),
    .Tile_X42Y8_R_f(R_f_top[188]),
    .Tile_X45Y8_R_t(R_t_top[189]),
    .Tile_X45Y8_R_f(R_f_top[189]),
    .Tile_X48Y8_R_t(R_t_top[190]),
    .Tile_X48Y8_R_f(R_f_top[190]),
    .Tile_X51Y8_R_t(R_t_top[191]),
    .Tile_X51Y8_R_f(R_f_top[191]),
    .Tile_X54Y8_R_t(R_t_top[192]),
    .Tile_X54Y8_R_f(R_f_top[192]),
    .Tile_X57Y8_R_t(R_t_top[193]),
    .Tile_X57Y8_R_f(R_f_top[193]),
    .Tile_X60Y8_R_t(R_t_top[194]),
    .Tile_X60Y8_R_f(R_f_top[194]),
    .Tile_X63Y8_R_t(R_t_top[195]),
    .Tile_X63Y8_R_f(R_f_top[195]),
    .Tile_X66Y8_R_t(R_t_top[196]),
    .Tile_X66Y8_R_f(R_f_top[196]),
    .Tile_X69Y8_R_t(R_t_top[197]),
    .Tile_X69Y8_R_f(R_f_top[197]),
    .Tile_X72Y8_R_t(R_t_top[198]),
    .Tile_X72Y8_R_f(R_f_top[198]),
    .Tile_X75Y8_R_t(R_t_top[199]),
    .Tile_X75Y8_R_f(R_f_top[199]),
    .Tile_X3Y9_R_t(R_t_top[200]),
    .Tile_X3Y9_R_f(R_f_top[200]),
    .Tile_X6Y9_R_t(R_t_top[201]),
    .Tile_X6Y9_R_f(R_f_top[201]),
    .Tile_X9Y9_R_t(R_t_top[202]),
    .Tile_X9Y9_R_f(R_f_top[202]),
    .Tile_X12Y9_R_t(R_t_top[203]),
    .Tile_X12Y9_R_f(R_f_top[203]),
    .Tile_X15Y9_R_t(R_t_top[204]),
    .Tile_X15Y9_R_f(R_f_top[204]),
    .Tile_X18Y9_R_t(R_t_top[205]),
    .Tile_X18Y9_R_f(R_f_top[205]),
    .Tile_X21Y9_R_t(R_t_top[206]),
    .Tile_X21Y9_R_f(R_f_top[206]),
    .Tile_X24Y9_R_t(R_t_top[207]),
    .Tile_X24Y9_R_f(R_f_top[207]),
    .Tile_X27Y9_R_t(R_t_top[208]),
    .Tile_X27Y9_R_f(R_f_top[208]),
    .Tile_X30Y9_R_t(R_t_top[209]),
    .Tile_X30Y9_R_f(R_f_top[209]),
    .Tile_X33Y9_R_t(R_t_top[210]),
    .Tile_X33Y9_R_f(R_f_top[210]),
    .Tile_X36Y9_R_t(R_t_top[211]),
    .Tile_X36Y9_R_f(R_f_top[211]),
    .Tile_X39Y9_R_t(R_t_top[212]),
    .Tile_X39Y9_R_f(R_f_top[212]),
    .Tile_X42Y9_R_t(R_t_top[213]),
    .Tile_X42Y9_R_f(R_f_top[213]),
    .Tile_X45Y9_R_t(R_t_top[214]),
    .Tile_X45Y9_R_f(R_f_top[214]),
    .Tile_X48Y9_R_t(R_t_top[215]),
    .Tile_X48Y9_R_f(R_f_top[215]),
    .Tile_X51Y9_R_t(R_t_top[216]),
    .Tile_X51Y9_R_f(R_f_top[216]),
    .Tile_X54Y9_R_t(R_t_top[217]),
    .Tile_X54Y9_R_f(R_f_top[217]),
    .Tile_X57Y9_R_t(R_t_top[218]),
    .Tile_X57Y9_R_f(R_f_top[218]),
    .Tile_X60Y9_R_t(R_t_top[219]),
    .Tile_X60Y9_R_f(R_f_top[219]),
    .Tile_X63Y9_R_t(R_t_top[220]),
    .Tile_X63Y9_R_f(R_f_top[220]),
    .Tile_X66Y9_R_t(R_t_top[221]),
    .Tile_X66Y9_R_f(R_f_top[221]),
    .Tile_X69Y9_R_t(R_t_top[222]),
    .Tile_X69Y9_R_f(R_f_top[222]),
    .Tile_X72Y9_R_t(R_t_top[223]),
    .Tile_X72Y9_R_f(R_f_top[223]),
    .Tile_X75Y9_R_t(R_t_top[224]),
    .Tile_X75Y9_R_f(R_f_top[224]),
    .Tile_X3Y10_R_t(R_t_top[225]),
    .Tile_X3Y10_R_f(R_f_top[225]),
    .Tile_X6Y10_R_t(R_t_top[226]),
    .Tile_X6Y10_R_f(R_f_top[226]),
    .Tile_X9Y10_R_t(R_t_top[227]),
    .Tile_X9Y10_R_f(R_f_top[227]),
    .Tile_X12Y10_R_t(R_t_top[228]),
    .Tile_X12Y10_R_f(R_f_top[228]),
    .Tile_X15Y10_R_t(R_t_top[229]),
    .Tile_X15Y10_R_f(R_f_top[229]),
    .Tile_X18Y10_R_t(R_t_top[230]),
    .Tile_X18Y10_R_f(R_f_top[230]),
    .Tile_X21Y10_R_t(R_t_top[231]),
    .Tile_X21Y10_R_f(R_f_top[231]),
    .Tile_X24Y10_R_t(R_t_top[232]),
    .Tile_X24Y10_R_f(R_f_top[232]),
    .Tile_X27Y10_R_t(R_t_top[233]),
    .Tile_X27Y10_R_f(R_f_top[233]),
    .Tile_X30Y10_R_t(R_t_top[234]),
    .Tile_X30Y10_R_f(R_f_top[234]),
    .Tile_X33Y10_R_t(R_t_top[235]),
    .Tile_X33Y10_R_f(R_f_top[235]),
    .Tile_X36Y10_R_t(R_t_top[236]),
    .Tile_X36Y10_R_f(R_f_top[236]),
    .Tile_X39Y10_R_t(R_t_top[237]),
    .Tile_X39Y10_R_f(R_f_top[237]),
    .Tile_X42Y10_R_t(R_t_top[238]),
    .Tile_X42Y10_R_f(R_f_top[238]),
    .Tile_X45Y10_R_t(R_t_top[239]),
    .Tile_X45Y10_R_f(R_f_top[239]),
    .Tile_X48Y10_R_t(R_t_top[240]),
    .Tile_X48Y10_R_f(R_f_top[240]),
    .Tile_X51Y10_R_t(R_t_top[241]),
    .Tile_X51Y10_R_f(R_f_top[241]),
    .Tile_X54Y10_R_t(R_t_top[242]),
    .Tile_X54Y10_R_f(R_f_top[242]),
    .Tile_X57Y10_R_t(R_t_top[243]),
    .Tile_X57Y10_R_f(R_f_top[243]),
    .Tile_X60Y10_R_t(R_t_top[244]),
    .Tile_X60Y10_R_f(R_f_top[244]),
    .Tile_X63Y10_R_t(R_t_top[245]),
    .Tile_X63Y10_R_f(R_f_top[245]),
    .Tile_X66Y10_R_t(R_t_top[246]),
    .Tile_X66Y10_R_f(R_f_top[246]),
    .Tile_X69Y10_R_t(R_t_top[247]),
    .Tile_X69Y10_R_f(R_f_top[247]),
    .Tile_X72Y10_R_t(R_t_top[248]),
    .Tile_X72Y10_R_f(R_f_top[248]),
    .Tile_X75Y10_R_t(R_t_top[249]),
    .Tile_X75Y10_R_f(R_f_top[249]),
    .Tile_X3Y11_R_t(R_t_top[250]),
    .Tile_X3Y11_R_f(R_f_top[250]),
    .Tile_X6Y11_R_t(R_t_top[251]),
    .Tile_X6Y11_R_f(R_f_top[251]),
    .Tile_X9Y11_R_t(R_t_top[252]),
    .Tile_X9Y11_R_f(R_f_top[252]),
    .Tile_X12Y11_R_t(R_t_top[253]),
    .Tile_X12Y11_R_f(R_f_top[253]),
    .Tile_X15Y11_R_t(R_t_top[254]),
    .Tile_X15Y11_R_f(R_f_top[254]),
    .Tile_X18Y11_R_t(R_t_top[255]),
    .Tile_X18Y11_R_f(R_f_top[255]),
    .Tile_X21Y11_R_t(R_t_top[256]),
    .Tile_X21Y11_R_f(R_f_top[256]),
    .Tile_X24Y11_R_t(R_t_top[257]),
    .Tile_X24Y11_R_f(R_f_top[257]),
    .Tile_X27Y11_R_t(R_t_top[258]),
    .Tile_X27Y11_R_f(R_f_top[258]),
    .Tile_X30Y11_R_t(R_t_top[259]),
    .Tile_X30Y11_R_f(R_f_top[259]),
    .Tile_X33Y11_R_t(R_t_top[260]),
    .Tile_X33Y11_R_f(R_f_top[260]),
    .Tile_X36Y11_R_t(R_t_top[261]),
    .Tile_X36Y11_R_f(R_f_top[261]),
    .Tile_X39Y11_R_t(R_t_top[262]),
    .Tile_X39Y11_R_f(R_f_top[262]),
    .Tile_X42Y11_R_t(R_t_top[263]),
    .Tile_X42Y11_R_f(R_f_top[263]),
    .Tile_X45Y11_R_t(R_t_top[264]),
    .Tile_X45Y11_R_f(R_f_top[264]),
    .Tile_X48Y11_R_t(R_t_top[265]),
    .Tile_X48Y11_R_f(R_f_top[265]),
    .Tile_X51Y11_R_t(R_t_top[266]),
    .Tile_X51Y11_R_f(R_f_top[266]),
    .Tile_X54Y11_R_t(R_t_top[267]),
    .Tile_X54Y11_R_f(R_f_top[267]),
    .Tile_X57Y11_R_t(R_t_top[268]),
    .Tile_X57Y11_R_f(R_f_top[268]),
    .Tile_X60Y11_R_t(R_t_top[269]),
    .Tile_X60Y11_R_f(R_f_top[269]),
    .Tile_X63Y11_R_t(R_t_top[270]),
    .Tile_X63Y11_R_f(R_f_top[270]),
    .Tile_X66Y11_R_t(R_t_top[271]),
    .Tile_X66Y11_R_f(R_f_top[271]),
    .Tile_X69Y11_R_t(R_t_top[272]),
    .Tile_X69Y11_R_f(R_f_top[272]),
    .Tile_X72Y11_R_t(R_t_top[273]),
    .Tile_X72Y11_R_f(R_f_top[273]),
    .Tile_X75Y11_R_t(R_t_top[274]),
    .Tile_X75Y11_R_f(R_f_top[274]),
    .Tile_X3Y12_R_t(R_t_top[275]),
    .Tile_X3Y12_R_f(R_f_top[275]),
    .Tile_X6Y12_R_t(R_t_top[276]),
    .Tile_X6Y12_R_f(R_f_top[276]),
    .Tile_X9Y12_R_t(R_t_top[277]),
    .Tile_X9Y12_R_f(R_f_top[277]),
    .Tile_X12Y12_R_t(R_t_top[278]),
    .Tile_X12Y12_R_f(R_f_top[278]),
    .Tile_X15Y12_R_t(R_t_top[279]),
    .Tile_X15Y12_R_f(R_f_top[279]),
    .Tile_X18Y12_R_t(R_t_top[280]),
    .Tile_X18Y12_R_f(R_f_top[280]),
    .Tile_X21Y12_R_t(R_t_top[281]),
    .Tile_X21Y12_R_f(R_f_top[281]),
    .Tile_X24Y12_R_t(R_t_top[282]),
    .Tile_X24Y12_R_f(R_f_top[282]),
    .Tile_X27Y12_R_t(R_t_top[283]),
    .Tile_X27Y12_R_f(R_f_top[283]),
    .Tile_X30Y12_R_t(R_t_top[284]),
    .Tile_X30Y12_R_f(R_f_top[284]),
    .Tile_X33Y12_R_t(R_t_top[285]),
    .Tile_X33Y12_R_f(R_f_top[285]),
    .Tile_X36Y12_R_t(R_t_top[286]),
    .Tile_X36Y12_R_f(R_f_top[286]),
    .Tile_X39Y12_R_t(R_t_top[287]),
    .Tile_X39Y12_R_f(R_f_top[287]),
    .Tile_X42Y12_R_t(R_t_top[288]),
    .Tile_X42Y12_R_f(R_f_top[288]),
    .Tile_X45Y12_R_t(R_t_top[289]),
    .Tile_X45Y12_R_f(R_f_top[289]),
    .Tile_X48Y12_R_t(R_t_top[290]),
    .Tile_X48Y12_R_f(R_f_top[290]),
    .Tile_X51Y12_R_t(R_t_top[291]),
    .Tile_X51Y12_R_f(R_f_top[291]),
    .Tile_X54Y12_R_t(R_t_top[292]),
    .Tile_X54Y12_R_f(R_f_top[292]),
    .Tile_X57Y12_R_t(R_t_top[293]),
    .Tile_X57Y12_R_f(R_f_top[293]),
    .Tile_X60Y12_R_t(R_t_top[294]),
    .Tile_X60Y12_R_f(R_f_top[294]),
    .Tile_X63Y12_R_t(R_t_top[295]),
    .Tile_X63Y12_R_f(R_f_top[295]),
    .Tile_X66Y12_R_t(R_t_top[296]),
    .Tile_X66Y12_R_f(R_f_top[296]),
    .Tile_X69Y12_R_t(R_t_top[297]),
    .Tile_X69Y12_R_f(R_f_top[297]),
    .Tile_X72Y12_R_t(R_t_top[298]),
    .Tile_X72Y12_R_f(R_f_top[298]),
    .Tile_X75Y12_R_t(R_t_top[299]),
    .Tile_X75Y12_R_f(R_f_top[299]),
    .Tile_X3Y13_R_t(R_t_top[300]),
    .Tile_X3Y13_R_f(R_f_top[300]),
    .Tile_X6Y13_R_t(R_t_top[301]),
    .Tile_X6Y13_R_f(R_f_top[301]),
    .Tile_X9Y13_R_t(R_t_top[302]),
    .Tile_X9Y13_R_f(R_f_top[302]),
    .Tile_X12Y13_R_t(R_t_top[303]),
    .Tile_X12Y13_R_f(R_f_top[303]),
    .Tile_X15Y13_R_t(R_t_top[304]),
    .Tile_X15Y13_R_f(R_f_top[304]),
    .Tile_X18Y13_R_t(R_t_top[305]),
    .Tile_X18Y13_R_f(R_f_top[305]),
    .Tile_X21Y13_R_t(R_t_top[306]),
    .Tile_X21Y13_R_f(R_f_top[306]),
    .Tile_X24Y13_R_t(R_t_top[307]),
    .Tile_X24Y13_R_f(R_f_top[307]),
    .Tile_X27Y13_R_t(R_t_top[308]),
    .Tile_X27Y13_R_f(R_f_top[308]),
    .Tile_X30Y13_R_t(R_t_top[309]),
    .Tile_X30Y13_R_f(R_f_top[309]),
    .Tile_X33Y13_R_t(R_t_top[310]),
    .Tile_X33Y13_R_f(R_f_top[310]),
    .Tile_X36Y13_R_t(R_t_top[311]),
    .Tile_X36Y13_R_f(R_f_top[311]),
    .Tile_X39Y13_R_t(R_t_top[312]),
    .Tile_X39Y13_R_f(R_f_top[312]),
    .Tile_X42Y13_R_t(R_t_top[313]),
    .Tile_X42Y13_R_f(R_f_top[313]),
    .Tile_X45Y13_R_t(R_t_top[314]),
    .Tile_X45Y13_R_f(R_f_top[314]),
    .Tile_X48Y13_R_t(R_t_top[315]),
    .Tile_X48Y13_R_f(R_f_top[315]),
    .Tile_X51Y13_R_t(R_t_top[316]),
    .Tile_X51Y13_R_f(R_f_top[316]),
    .Tile_X54Y13_R_t(R_t_top[317]),
    .Tile_X54Y13_R_f(R_f_top[317]),
    .Tile_X57Y13_R_t(R_t_top[318]),
    .Tile_X57Y13_R_f(R_f_top[318]),
    .Tile_X60Y13_R_t(R_t_top[319]),
    .Tile_X60Y13_R_f(R_f_top[319]),
    .Tile_X63Y13_R_t(R_t_top[320]),
    .Tile_X63Y13_R_f(R_f_top[320]),
    .Tile_X66Y13_R_t(R_t_top[321]),
    .Tile_X66Y13_R_f(R_f_top[321]),
    .Tile_X69Y13_R_t(R_t_top[322]),
    .Tile_X69Y13_R_f(R_f_top[322]),
    .Tile_X72Y13_R_t(R_t_top[323]),
    .Tile_X72Y13_R_f(R_f_top[323]),
    .Tile_X75Y13_R_t(R_t_top[324]),
    .Tile_X75Y13_R_f(R_f_top[324]),
    .Tile_X3Y14_R_t(R_t_top[325]),
    .Tile_X3Y14_R_f(R_f_top[325]),
    .Tile_X6Y14_R_t(R_t_top[326]),
    .Tile_X6Y14_R_f(R_f_top[326]),
    .Tile_X9Y14_R_t(R_t_top[327]),
    .Tile_X9Y14_R_f(R_f_top[327]),
    .Tile_X12Y14_R_t(R_t_top[328]),
    .Tile_X12Y14_R_f(R_f_top[328]),
    .Tile_X15Y14_R_t(R_t_top[329]),
    .Tile_X15Y14_R_f(R_f_top[329]),
    .Tile_X18Y14_R_t(R_t_top[330]),
    .Tile_X18Y14_R_f(R_f_top[330]),
    .Tile_X21Y14_R_t(R_t_top[331]),
    .Tile_X21Y14_R_f(R_f_top[331]),
    .Tile_X24Y14_R_t(R_t_top[332]),
    .Tile_X24Y14_R_f(R_f_top[332]),
    .Tile_X27Y14_R_t(R_t_top[333]),
    .Tile_X27Y14_R_f(R_f_top[333]),
    .Tile_X30Y14_R_t(R_t_top[334]),
    .Tile_X30Y14_R_f(R_f_top[334]),
    .Tile_X33Y14_R_t(R_t_top[335]),
    .Tile_X33Y14_R_f(R_f_top[335]),
    .Tile_X36Y14_R_t(R_t_top[336]),
    .Tile_X36Y14_R_f(R_f_top[336]),
    .Tile_X39Y14_R_t(R_t_top[337]),
    .Tile_X39Y14_R_f(R_f_top[337]),
    .Tile_X42Y14_R_t(R_t_top[338]),
    .Tile_X42Y14_R_f(R_f_top[338]),
    .Tile_X45Y14_R_t(R_t_top[339]),
    .Tile_X45Y14_R_f(R_f_top[339]),
    .Tile_X48Y14_R_t(R_t_top[340]),
    .Tile_X48Y14_R_f(R_f_top[340]),
    .Tile_X51Y14_R_t(R_t_top[341]),
    .Tile_X51Y14_R_f(R_f_top[341]),
    .Tile_X54Y14_R_t(R_t_top[342]),
    .Tile_X54Y14_R_f(R_f_top[342]),
    .Tile_X57Y14_R_t(R_t_top[343]),
    .Tile_X57Y14_R_f(R_f_top[343]),
    .Tile_X60Y14_R_t(R_t_top[344]),
    .Tile_X60Y14_R_f(R_f_top[344]),
    .Tile_X63Y14_R_t(R_t_top[345]),
    .Tile_X63Y14_R_f(R_f_top[345]),
    .Tile_X66Y14_R_t(R_t_top[346]),
    .Tile_X66Y14_R_f(R_f_top[346]),
    .Tile_X69Y14_R_t(R_t_top[347]),
    .Tile_X69Y14_R_f(R_f_top[347]),
    .Tile_X72Y14_R_t(R_t_top[348]),
    .Tile_X72Y14_R_f(R_f_top[348]),
    .Tile_X75Y14_R_t(R_t_top[349]),
    .Tile_X75Y14_R_f(R_f_top[349]),
    .Tile_X3Y15_R_t(R_t_top[350]),
    .Tile_X3Y15_R_f(R_f_top[350]),
    .Tile_X6Y15_R_t(R_t_top[351]),
    .Tile_X6Y15_R_f(R_f_top[351]),
    .Tile_X9Y15_R_t(R_t_top[352]),
    .Tile_X9Y15_R_f(R_f_top[352]),
    .Tile_X12Y15_R_t(R_t_top[353]),
    .Tile_X12Y15_R_f(R_f_top[353]),
    .Tile_X15Y15_R_t(R_t_top[354]),
    .Tile_X15Y15_R_f(R_f_top[354]),
    .Tile_X18Y15_R_t(R_t_top[355]),
    .Tile_X18Y15_R_f(R_f_top[355]),
    .Tile_X21Y15_R_t(R_t_top[356]),
    .Tile_X21Y15_R_f(R_f_top[356]),
    .Tile_X24Y15_R_t(R_t_top[357]),
    .Tile_X24Y15_R_f(R_f_top[357]),
    .Tile_X27Y15_R_t(R_t_top[358]),
    .Tile_X27Y15_R_f(R_f_top[358]),
    .Tile_X30Y15_R_t(R_t_top[359]),
    .Tile_X30Y15_R_f(R_f_top[359]),
    .Tile_X33Y15_R_t(R_t_top[360]),
    .Tile_X33Y15_R_f(R_f_top[360]),
    .Tile_X36Y15_R_t(R_t_top[361]),
    .Tile_X36Y15_R_f(R_f_top[361]),
    .Tile_X39Y15_R_t(R_t_top[362]),
    .Tile_X39Y15_R_f(R_f_top[362]),
    .Tile_X42Y15_R_t(R_t_top[363]),
    .Tile_X42Y15_R_f(R_f_top[363]),
    .Tile_X45Y15_R_t(R_t_top[364]),
    .Tile_X45Y15_R_f(R_f_top[364]),
    .Tile_X48Y15_R_t(R_t_top[365]),
    .Tile_X48Y15_R_f(R_f_top[365]),
    .Tile_X51Y15_R_t(R_t_top[366]),
    .Tile_X51Y15_R_f(R_f_top[366]),
    .Tile_X54Y15_R_t(R_t_top[367]),
    .Tile_X54Y15_R_f(R_f_top[367]),
    .Tile_X57Y15_R_t(R_t_top[368]),
    .Tile_X57Y15_R_f(R_f_top[368]),
    .Tile_X60Y15_R_t(R_t_top[369]),
    .Tile_X60Y15_R_f(R_f_top[369]),
    .Tile_X63Y15_R_t(R_t_top[370]),
    .Tile_X63Y15_R_f(R_f_top[370]),
    .Tile_X66Y15_R_t(R_t_top[371]),
    .Tile_X66Y15_R_f(R_f_top[371]),
    .Tile_X69Y15_R_t(R_t_top[372]),
    .Tile_X69Y15_R_f(R_f_top[372]),
    .Tile_X72Y15_R_t(R_t_top[373]),
    .Tile_X72Y15_R_f(R_f_top[373]),
    .Tile_X75Y15_R_t(R_t_top[374]),
    .Tile_X75Y15_R_f(R_f_top[374]),
    .Tile_X3Y16_R_t(R_t_top[375]),
    .Tile_X3Y16_R_f(R_f_top[375]),
    .Tile_X6Y16_R_t(R_t_top[376]),
    .Tile_X6Y16_R_f(R_f_top[376]),
    .Tile_X9Y16_R_t(R_t_top[377]),
    .Tile_X9Y16_R_f(R_f_top[377]),
    .Tile_X12Y16_R_t(R_t_top[378]),
    .Tile_X12Y16_R_f(R_f_top[378]),
    .Tile_X15Y16_R_t(R_t_top[379]),
    .Tile_X15Y16_R_f(R_f_top[379]),
    .Tile_X18Y16_R_t(R_t_top[380]),
    .Tile_X18Y16_R_f(R_f_top[380]),
    .Tile_X21Y16_R_t(R_t_top[381]),
    .Tile_X21Y16_R_f(R_f_top[381]),
    .Tile_X24Y16_R_t(R_t_top[382]),
    .Tile_X24Y16_R_f(R_f_top[382]),
    .Tile_X27Y16_R_t(R_t_top[383]),
    .Tile_X27Y16_R_f(R_f_top[383]),
    .Tile_X30Y16_R_t(R_t_top[384]),
    .Tile_X30Y16_R_f(R_f_top[384]),
    .Tile_X33Y16_R_t(R_t_top[385]),
    .Tile_X33Y16_R_f(R_f_top[385]),
    .Tile_X36Y16_R_t(R_t_top[386]),
    .Tile_X36Y16_R_f(R_f_top[386]),
    .Tile_X39Y16_R_t(R_t_top[387]),
    .Tile_X39Y16_R_f(R_f_top[387]),
    .Tile_X42Y16_R_t(R_t_top[388]),
    .Tile_X42Y16_R_f(R_f_top[388]),
    .Tile_X45Y16_R_t(R_t_top[389]),
    .Tile_X45Y16_R_f(R_f_top[389]),
    .Tile_X48Y16_R_t(R_t_top[390]),
    .Tile_X48Y16_R_f(R_f_top[390]),
    .Tile_X51Y16_R_t(R_t_top[391]),
    .Tile_X51Y16_R_f(R_f_top[391]),
    .Tile_X54Y16_R_t(R_t_top[392]),
    .Tile_X54Y16_R_f(R_f_top[392]),
    .Tile_X57Y16_R_t(R_t_top[393]),
    .Tile_X57Y16_R_f(R_f_top[393]),
    .Tile_X60Y16_R_t(R_t_top[394]),
    .Tile_X60Y16_R_f(R_f_top[394]),
    .Tile_X63Y16_R_t(R_t_top[395]),
    .Tile_X63Y16_R_f(R_f_top[395]),
    .Tile_X66Y16_R_t(R_t_top[396]),
    .Tile_X66Y16_R_f(R_f_top[396]),
    .Tile_X69Y16_R_t(R_t_top[397]),
    .Tile_X69Y16_R_f(R_f_top[397]),
    .Tile_X72Y16_R_t(R_t_top[398]),
    .Tile_X72Y16_R_f(R_f_top[398]),
    .Tile_X75Y16_R_t(R_t_top[399]),
    .Tile_X75Y16_R_f(R_f_top[399]),
    .Tile_X3Y17_R_t(R_t_top[400]),
    .Tile_X3Y17_R_f(R_f_top[400]),
    .Tile_X6Y17_R_t(R_t_top[401]),
    .Tile_X6Y17_R_f(R_f_top[401]),
    .Tile_X9Y17_R_t(R_t_top[402]),
    .Tile_X9Y17_R_f(R_f_top[402]),
    .Tile_X12Y17_R_t(R_t_top[403]),
    .Tile_X12Y17_R_f(R_f_top[403]),
    .Tile_X15Y17_R_t(R_t_top[404]),
    .Tile_X15Y17_R_f(R_f_top[404]),
    .Tile_X18Y17_R_t(R_t_top[405]),
    .Tile_X18Y17_R_f(R_f_top[405]),
    .Tile_X21Y17_R_t(R_t_top[406]),
    .Tile_X21Y17_R_f(R_f_top[406]),
    .Tile_X24Y17_R_t(R_t_top[407]),
    .Tile_X24Y17_R_f(R_f_top[407]),
    .Tile_X27Y17_R_t(R_t_top[408]),
    .Tile_X27Y17_R_f(R_f_top[408]),
    .Tile_X30Y17_R_t(R_t_top[409]),
    .Tile_X30Y17_R_f(R_f_top[409]),
    .Tile_X33Y17_R_t(R_t_top[410]),
    .Tile_X33Y17_R_f(R_f_top[410]),
    .Tile_X36Y17_R_t(R_t_top[411]),
    .Tile_X36Y17_R_f(R_f_top[411]),
    .Tile_X39Y17_R_t(R_t_top[412]),
    .Tile_X39Y17_R_f(R_f_top[412]),
    .Tile_X42Y17_R_t(R_t_top[413]),
    .Tile_X42Y17_R_f(R_f_top[413]),
    .Tile_X45Y17_R_t(R_t_top[414]),
    .Tile_X45Y17_R_f(R_f_top[414]),
    .Tile_X48Y17_R_t(R_t_top[415]),
    .Tile_X48Y17_R_f(R_f_top[415]),
    .Tile_X51Y17_R_t(R_t_top[416]),
    .Tile_X51Y17_R_f(R_f_top[416]),
    .Tile_X54Y17_R_t(R_t_top[417]),
    .Tile_X54Y17_R_f(R_f_top[417]),
    .Tile_X57Y17_R_t(R_t_top[418]),
    .Tile_X57Y17_R_f(R_f_top[418]),
    .Tile_X60Y17_R_t(R_t_top[419]),
    .Tile_X60Y17_R_f(R_f_top[419]),
    .Tile_X63Y17_R_t(R_t_top[420]),
    .Tile_X63Y17_R_f(R_f_top[420]),
    .Tile_X66Y17_R_t(R_t_top[421]),
    .Tile_X66Y17_R_f(R_f_top[421]),
    .Tile_X69Y17_R_t(R_t_top[422]),
    .Tile_X69Y17_R_f(R_f_top[422]),
    .Tile_X72Y17_R_t(R_t_top[423]),
    .Tile_X72Y17_R_f(R_f_top[423]),
    .Tile_X75Y17_R_t(R_t_top[424]),
    .Tile_X75Y17_R_f(R_f_top[424]),
    .Tile_X3Y18_R_t(R_t_top[425]),
    .Tile_X3Y18_R_f(R_f_top[425]),
    .Tile_X6Y18_R_t(R_t_top[426]),
    .Tile_X6Y18_R_f(R_f_top[426]),
    .Tile_X9Y18_R_t(R_t_top[427]),
    .Tile_X9Y18_R_f(R_f_top[427]),
    .Tile_X12Y18_R_t(R_t_top[428]),
    .Tile_X12Y18_R_f(R_f_top[428]),
    .Tile_X15Y18_R_t(R_t_top[429]),
    .Tile_X15Y18_R_f(R_f_top[429]),
    .Tile_X18Y18_R_t(R_t_top[430]),
    .Tile_X18Y18_R_f(R_f_top[430]),
    .Tile_X21Y18_R_t(R_t_top[431]),
    .Tile_X21Y18_R_f(R_f_top[431]),
    .Tile_X24Y18_R_t(R_t_top[432]),
    .Tile_X24Y18_R_f(R_f_top[432]),
    .Tile_X27Y18_R_t(R_t_top[433]),
    .Tile_X27Y18_R_f(R_f_top[433]),
    .Tile_X30Y18_R_t(R_t_top[434]),
    .Tile_X30Y18_R_f(R_f_top[434]),
    .Tile_X33Y18_R_t(R_t_top[435]),
    .Tile_X33Y18_R_f(R_f_top[435]),
    .Tile_X36Y18_R_t(R_t_top[436]),
    .Tile_X36Y18_R_f(R_f_top[436]),
    .Tile_X39Y18_R_t(R_t_top[437]),
    .Tile_X39Y18_R_f(R_f_top[437]),
    .Tile_X42Y18_R_t(R_t_top[438]),
    .Tile_X42Y18_R_f(R_f_top[438]),
    .Tile_X45Y18_R_t(R_t_top[439]),
    .Tile_X45Y18_R_f(R_f_top[439]),
    .Tile_X48Y18_R_t(R_t_top[440]),
    .Tile_X48Y18_R_f(R_f_top[440]),
    .Tile_X51Y18_R_t(R_t_top[441]),
    .Tile_X51Y18_R_f(R_f_top[441]),
    .Tile_X54Y18_R_t(R_t_top[442]),
    .Tile_X54Y18_R_f(R_f_top[442]),
    .Tile_X57Y18_R_t(R_t_top[443]),
    .Tile_X57Y18_R_f(R_f_top[443]),
    .Tile_X60Y18_R_t(R_t_top[444]),
    .Tile_X60Y18_R_f(R_f_top[444]),
    .Tile_X63Y18_R_t(R_t_top[445]),
    .Tile_X63Y18_R_f(R_f_top[445]),
    .Tile_X66Y18_R_t(R_t_top[446]),
    .Tile_X66Y18_R_f(R_f_top[446]),
    .Tile_X69Y18_R_t(R_t_top[447]),
    .Tile_X69Y18_R_f(R_f_top[447]),
    .Tile_X72Y18_R_t(R_t_top[448]),
    .Tile_X72Y18_R_f(R_f_top[448]),
    .Tile_X75Y18_R_t(R_t_top[449]),
    .Tile_X75Y18_R_f(R_f_top[449]),
    .Tile_X3Y19_R_t(R_t_top[450]),
    .Tile_X3Y19_R_f(R_f_top[450]),
    .Tile_X6Y19_R_t(R_t_top[451]),
    .Tile_X6Y19_R_f(R_f_top[451]),
    .Tile_X9Y19_R_t(R_t_top[452]),
    .Tile_X9Y19_R_f(R_f_top[452]),
    .Tile_X12Y19_R_t(R_t_top[453]),
    .Tile_X12Y19_R_f(R_f_top[453]),
    .Tile_X15Y19_R_t(R_t_top[454]),
    .Tile_X15Y19_R_f(R_f_top[454]),
    .Tile_X18Y19_R_t(R_t_top[455]),
    .Tile_X18Y19_R_f(R_f_top[455]),
    .Tile_X21Y19_R_t(R_t_top[456]),
    .Tile_X21Y19_R_f(R_f_top[456]),
    .Tile_X24Y19_R_t(R_t_top[457]),
    .Tile_X24Y19_R_f(R_f_top[457]),
    .Tile_X27Y19_R_t(R_t_top[458]),
    .Tile_X27Y19_R_f(R_f_top[458]),
    .Tile_X30Y19_R_t(R_t_top[459]),
    .Tile_X30Y19_R_f(R_f_top[459]),
    .Tile_X33Y19_R_t(R_t_top[460]),
    .Tile_X33Y19_R_f(R_f_top[460]),
    .Tile_X36Y19_R_t(R_t_top[461]),
    .Tile_X36Y19_R_f(R_f_top[461]),
    .Tile_X39Y19_R_t(R_t_top[462]),
    .Tile_X39Y19_R_f(R_f_top[462]),
    .Tile_X42Y19_R_t(R_t_top[463]),
    .Tile_X42Y19_R_f(R_f_top[463]),
    .Tile_X45Y19_R_t(R_t_top[464]),
    .Tile_X45Y19_R_f(R_f_top[464]),
    .Tile_X48Y19_R_t(R_t_top[465]),
    .Tile_X48Y19_R_f(R_f_top[465]),
    .Tile_X51Y19_R_t(R_t_top[466]),
    .Tile_X51Y19_R_f(R_f_top[466]),
    .Tile_X54Y19_R_t(R_t_top[467]),
    .Tile_X54Y19_R_f(R_f_top[467]),
    .Tile_X57Y19_R_t(R_t_top[468]),
    .Tile_X57Y19_R_f(R_f_top[468]),
    .Tile_X60Y19_R_t(R_t_top[469]),
    .Tile_X60Y19_R_f(R_f_top[469]),
    .Tile_X63Y19_R_t(R_t_top[470]),
    .Tile_X63Y19_R_f(R_f_top[470]),
    .Tile_X66Y19_R_t(R_t_top[471]),
    .Tile_X66Y19_R_f(R_f_top[471]),
    .Tile_X69Y19_R_t(R_t_top[472]),
    .Tile_X69Y19_R_f(R_f_top[472]),
    .Tile_X72Y19_R_t(R_t_top[473]),
    .Tile_X72Y19_R_f(R_f_top[473]),
    .Tile_X75Y19_R_t(R_t_top[474]),
    .Tile_X75Y19_R_f(R_f_top[474]),
    .Tile_X3Y20_R_t(R_t_top[475]),
    .Tile_X3Y20_R_f(R_f_top[475]),
    .Tile_X6Y20_R_t(R_t_top[476]),
    .Tile_X6Y20_R_f(R_f_top[476]),
    .Tile_X9Y20_R_t(R_t_top[477]),
    .Tile_X9Y20_R_f(R_f_top[477]),
    .Tile_X12Y20_R_t(R_t_top[478]),
    .Tile_X12Y20_R_f(R_f_top[478]),
    .Tile_X15Y20_R_t(R_t_top[479]),
    .Tile_X15Y20_R_f(R_f_top[479]),
    .Tile_X18Y20_R_t(R_t_top[480]),
    .Tile_X18Y20_R_f(R_f_top[480]),
    .Tile_X21Y20_R_t(R_t_top[481]),
    .Tile_X21Y20_R_f(R_f_top[481]),
    .Tile_X24Y20_R_t(R_t_top[482]),
    .Tile_X24Y20_R_f(R_f_top[482]),
    .Tile_X27Y20_R_t(R_t_top[483]),
    .Tile_X27Y20_R_f(R_f_top[483]),
    .Tile_X30Y20_R_t(R_t_top[484]),
    .Tile_X30Y20_R_f(R_f_top[484]),
    .Tile_X33Y20_R_t(R_t_top[485]),
    .Tile_X33Y20_R_f(R_f_top[485]),
    .Tile_X36Y20_R_t(R_t_top[486]),
    .Tile_X36Y20_R_f(R_f_top[486]),
    .Tile_X39Y20_R_t(R_t_top[487]),
    .Tile_X39Y20_R_f(R_f_top[487]),
    .Tile_X42Y20_R_t(R_t_top[488]),
    .Tile_X42Y20_R_f(R_f_top[488]),
    .Tile_X45Y20_R_t(R_t_top[489]),
    .Tile_X45Y20_R_f(R_f_top[489]),
    .Tile_X48Y20_R_t(R_t_top[490]),
    .Tile_X48Y20_R_f(R_f_top[490]),
    .Tile_X51Y20_R_t(R_t_top[491]),
    .Tile_X51Y20_R_f(R_f_top[491]),
    .Tile_X54Y20_R_t(R_t_top[492]),
    .Tile_X54Y20_R_f(R_f_top[492]),
    .Tile_X57Y20_R_t(R_t_top[493]),
    .Tile_X57Y20_R_f(R_f_top[493]),
    .Tile_X60Y20_R_t(R_t_top[494]),
    .Tile_X60Y20_R_f(R_f_top[494]),
    .Tile_X63Y20_R_t(R_t_top[495]),
    .Tile_X63Y20_R_f(R_f_top[495]),
    .Tile_X66Y20_R_t(R_t_top[496]),
    .Tile_X66Y20_R_f(R_f_top[496]),
    .Tile_X69Y20_R_t(R_t_top[497]),
    .Tile_X69Y20_R_f(R_f_top[497]),
    .Tile_X72Y20_R_t(R_t_top[498]),
    .Tile_X72Y20_R_f(R_f_top[498]),
    .Tile_X75Y20_R_t(R_t_top[499]),
    .Tile_X75Y20_R_f(R_f_top[499]),
    .Tile_X3Y21_R_t(R_t_top[500]),
    .Tile_X3Y21_R_f(R_f_top[500]),
    .Tile_X6Y21_R_t(R_t_top[501]),
    .Tile_X6Y21_R_f(R_f_top[501]),
    .Tile_X9Y21_R_t(R_t_top[502]),
    .Tile_X9Y21_R_f(R_f_top[502]),
    .Tile_X12Y21_R_t(R_t_top[503]),
    .Tile_X12Y21_R_f(R_f_top[503]),
    .Tile_X15Y21_R_t(R_t_top[504]),
    .Tile_X15Y21_R_f(R_f_top[504]),
    .Tile_X18Y21_R_t(R_t_top[505]),
    .Tile_X18Y21_R_f(R_f_top[505]),
    .Tile_X21Y21_R_t(R_t_top[506]),
    .Tile_X21Y21_R_f(R_f_top[506]),
    .Tile_X24Y21_R_t(R_t_top[507]),
    .Tile_X24Y21_R_f(R_f_top[507]),
    .Tile_X27Y21_R_t(R_t_top[508]),
    .Tile_X27Y21_R_f(R_f_top[508]),
    .Tile_X30Y21_R_t(R_t_top[509]),
    .Tile_X30Y21_R_f(R_f_top[509]),
    .Tile_X33Y21_R_t(R_t_top[510]),
    .Tile_X33Y21_R_f(R_f_top[510]),
    .Tile_X36Y21_R_t(R_t_top[511]),
    .Tile_X36Y21_R_f(R_f_top[511]),
    .Tile_X39Y21_R_t(R_t_top[512]),
    .Tile_X39Y21_R_f(R_f_top[512]),
    .Tile_X42Y21_R_t(R_t_top[513]),
    .Tile_X42Y21_R_f(R_f_top[513]),
    .Tile_X45Y21_R_t(R_t_top[514]),
    .Tile_X45Y21_R_f(R_f_top[514]),
    .Tile_X48Y21_R_t(R_t_top[515]),
    .Tile_X48Y21_R_f(R_f_top[515]),
    .Tile_X51Y21_R_t(R_t_top[516]),
    .Tile_X51Y21_R_f(R_f_top[516]),
    .Tile_X54Y21_R_t(R_t_top[517]),
    .Tile_X54Y21_R_f(R_f_top[517]),
    .Tile_X57Y21_R_t(R_t_top[518]),
    .Tile_X57Y21_R_f(R_f_top[518]),
    .Tile_X60Y21_R_t(R_t_top[519]),
    .Tile_X60Y21_R_f(R_f_top[519]),
    .Tile_X63Y21_R_t(R_t_top[520]),
    .Tile_X63Y21_R_f(R_f_top[520]),
    .Tile_X66Y21_R_t(R_t_top[521]),
    .Tile_X66Y21_R_f(R_f_top[521]),
    .Tile_X69Y21_R_t(R_t_top[522]),
    .Tile_X69Y21_R_f(R_f_top[522]),
    .Tile_X72Y21_R_t(R_t_top[523]),
    .Tile_X72Y21_R_f(R_f_top[523]),
    .Tile_X75Y21_R_t(R_t_top[524]),
    .Tile_X75Y21_R_f(R_f_top[524]),
    .Tile_X3Y22_R_t(R_t_top[525]),
    .Tile_X3Y22_R_f(R_f_top[525]),
    .Tile_X6Y22_R_t(R_t_top[526]),
    .Tile_X6Y22_R_f(R_f_top[526]),
    .Tile_X9Y22_R_t(R_t_top[527]),
    .Tile_X9Y22_R_f(R_f_top[527]),
    .Tile_X12Y22_R_t(R_t_top[528]),
    .Tile_X12Y22_R_f(R_f_top[528]),
    .Tile_X15Y22_R_t(R_t_top[529]),
    .Tile_X15Y22_R_f(R_f_top[529]),
    .Tile_X18Y22_R_t(R_t_top[530]),
    .Tile_X18Y22_R_f(R_f_top[530]),
    .Tile_X21Y22_R_t(R_t_top[531]),
    .Tile_X21Y22_R_f(R_f_top[531]),
    .Tile_X24Y22_R_t(R_t_top[532]),
    .Tile_X24Y22_R_f(R_f_top[532]),
    .Tile_X27Y22_R_t(R_t_top[533]),
    .Tile_X27Y22_R_f(R_f_top[533]),
    .Tile_X30Y22_R_t(R_t_top[534]),
    .Tile_X30Y22_R_f(R_f_top[534]),
    .Tile_X33Y22_R_t(R_t_top[535]),
    .Tile_X33Y22_R_f(R_f_top[535]),
    .Tile_X36Y22_R_t(R_t_top[536]),
    .Tile_X36Y22_R_f(R_f_top[536]),
    .Tile_X39Y22_R_t(R_t_top[537]),
    .Tile_X39Y22_R_f(R_f_top[537]),
    .Tile_X42Y22_R_t(R_t_top[538]),
    .Tile_X42Y22_R_f(R_f_top[538]),
    .Tile_X45Y22_R_t(R_t_top[539]),
    .Tile_X45Y22_R_f(R_f_top[539]),
    .Tile_X48Y22_R_t(R_t_top[540]),
    .Tile_X48Y22_R_f(R_f_top[540]),
    .Tile_X51Y22_R_t(R_t_top[541]),
    .Tile_X51Y22_R_f(R_f_top[541]),
    .Tile_X54Y22_R_t(R_t_top[542]),
    .Tile_X54Y22_R_f(R_f_top[542]),
    .Tile_X57Y22_R_t(R_t_top[543]),
    .Tile_X57Y22_R_f(R_f_top[543]),
    .Tile_X60Y22_R_t(R_t_top[544]),
    .Tile_X60Y22_R_f(R_f_top[544]),
    .Tile_X63Y22_R_t(R_t_top[545]),
    .Tile_X63Y22_R_f(R_f_top[545]),
    .Tile_X66Y22_R_t(R_t_top[546]),
    .Tile_X66Y22_R_f(R_f_top[546]),
    .Tile_X69Y22_R_t(R_t_top[547]),
    .Tile_X69Y22_R_f(R_f_top[547]),
    .Tile_X72Y22_R_t(R_t_top[548]),
    .Tile_X72Y22_R_f(R_f_top[548]),
    .Tile_X75Y22_R_t(R_t_top[549]),
    .Tile_X75Y22_R_f(R_f_top[549]),
    .Tile_X3Y23_R_t(R_t_top[550]),
    .Tile_X3Y23_R_f(R_f_top[550]),
    .Tile_X6Y23_R_t(R_t_top[551]),
    .Tile_X6Y23_R_f(R_f_top[551]),
    .Tile_X9Y23_R_t(R_t_top[552]),
    .Tile_X9Y23_R_f(R_f_top[552]),
    .Tile_X12Y23_R_t(R_t_top[553]),
    .Tile_X12Y23_R_f(R_f_top[553]),
    .Tile_X15Y23_R_t(R_t_top[554]),
    .Tile_X15Y23_R_f(R_f_top[554]),
    .Tile_X18Y23_R_t(R_t_top[555]),
    .Tile_X18Y23_R_f(R_f_top[555]),
    .Tile_X21Y23_R_t(R_t_top[556]),
    .Tile_X21Y23_R_f(R_f_top[556]),
    .Tile_X24Y23_R_t(R_t_top[557]),
    .Tile_X24Y23_R_f(R_f_top[557]),
    .Tile_X27Y23_R_t(R_t_top[558]),
    .Tile_X27Y23_R_f(R_f_top[558]),
    .Tile_X30Y23_R_t(R_t_top[559]),
    .Tile_X30Y23_R_f(R_f_top[559]),
    .Tile_X33Y23_R_t(R_t_top[560]),
    .Tile_X33Y23_R_f(R_f_top[560]),
    .Tile_X36Y23_R_t(R_t_top[561]),
    .Tile_X36Y23_R_f(R_f_top[561]),
    .Tile_X39Y23_R_t(R_t_top[562]),
    .Tile_X39Y23_R_f(R_f_top[562]),
    .Tile_X42Y23_R_t(R_t_top[563]),
    .Tile_X42Y23_R_f(R_f_top[563]),
    .Tile_X45Y23_R_t(R_t_top[564]),
    .Tile_X45Y23_R_f(R_f_top[564]),
    .Tile_X48Y23_R_t(R_t_top[565]),
    .Tile_X48Y23_R_f(R_f_top[565]),
    .Tile_X51Y23_R_t(R_t_top[566]),
    .Tile_X51Y23_R_f(R_f_top[566]),
    .Tile_X54Y23_R_t(R_t_top[567]),
    .Tile_X54Y23_R_f(R_f_top[567]),
    .Tile_X57Y23_R_t(R_t_top[568]),
    .Tile_X57Y23_R_f(R_f_top[568]),
    .Tile_X60Y23_R_t(R_t_top[569]),
    .Tile_X60Y23_R_f(R_f_top[569]),
    .Tile_X63Y23_R_t(R_t_top[570]),
    .Tile_X63Y23_R_f(R_f_top[570]),
    .Tile_X66Y23_R_t(R_t_top[571]),
    .Tile_X66Y23_R_f(R_f_top[571]),
    .Tile_X69Y23_R_t(R_t_top[572]),
    .Tile_X69Y23_R_f(R_f_top[572]),
    .Tile_X72Y23_R_t(R_t_top[573]),
    .Tile_X72Y23_R_f(R_f_top[573]),
    .Tile_X75Y23_R_t(R_t_top[574]),
    .Tile_X75Y23_R_f(R_f_top[574]),
    .Tile_X3Y24_R_t(R_t_top[575]),
    .Tile_X3Y24_R_f(R_f_top[575]),
    .Tile_X6Y24_R_t(R_t_top[576]),
    .Tile_X6Y24_R_f(R_f_top[576]),
    .Tile_X9Y24_R_t(R_t_top[577]),
    .Tile_X9Y24_R_f(R_f_top[577]),
    .Tile_X12Y24_R_t(R_t_top[578]),
    .Tile_X12Y24_R_f(R_f_top[578]),
    .Tile_X15Y24_R_t(R_t_top[579]),
    .Tile_X15Y24_R_f(R_f_top[579]),
    .Tile_X18Y24_R_t(R_t_top[580]),
    .Tile_X18Y24_R_f(R_f_top[580]),
    .Tile_X21Y24_R_t(R_t_top[581]),
    .Tile_X21Y24_R_f(R_f_top[581]),
    .Tile_X24Y24_R_t(R_t_top[582]),
    .Tile_X24Y24_R_f(R_f_top[582]),
    .Tile_X27Y24_R_t(R_t_top[583]),
    .Tile_X27Y24_R_f(R_f_top[583]),
    .Tile_X30Y24_R_t(R_t_top[584]),
    .Tile_X30Y24_R_f(R_f_top[584]),
    .Tile_X33Y24_R_t(R_t_top[585]),
    .Tile_X33Y24_R_f(R_f_top[585]),
    .Tile_X36Y24_R_t(R_t_top[586]),
    .Tile_X36Y24_R_f(R_f_top[586]),
    .Tile_X39Y24_R_t(R_t_top[587]),
    .Tile_X39Y24_R_f(R_f_top[587]),
    .Tile_X42Y24_R_t(R_t_top[588]),
    .Tile_X42Y24_R_f(R_f_top[588]),
    .Tile_X45Y24_R_t(R_t_top[589]),
    .Tile_X45Y24_R_f(R_f_top[589]),
    .Tile_X48Y24_R_t(R_t_top[590]),
    .Tile_X48Y24_R_f(R_f_top[590]),
    .Tile_X51Y24_R_t(R_t_top[591]),
    .Tile_X51Y24_R_f(R_f_top[591]),
    .Tile_X54Y24_R_t(R_t_top[592]),
    .Tile_X54Y24_R_f(R_f_top[592]),
    .Tile_X57Y24_R_t(R_t_top[593]),
    .Tile_X57Y24_R_f(R_f_top[593]),
    .Tile_X60Y24_R_t(R_t_top[594]),
    .Tile_X60Y24_R_f(R_f_top[594]),
    .Tile_X63Y24_R_t(R_t_top[595]),
    .Tile_X63Y24_R_f(R_f_top[595]),
    .Tile_X66Y24_R_t(R_t_top[596]),
    .Tile_X66Y24_R_f(R_f_top[596]),
    .Tile_X69Y24_R_t(R_t_top[597]),
    .Tile_X69Y24_R_f(R_f_top[597]),
    .Tile_X72Y24_R_t(R_t_top[598]),
    .Tile_X72Y24_R_f(R_f_top[598]),
    .Tile_X75Y24_R_t(R_t_top[599]),
    .Tile_X75Y24_R_f(R_f_top[599]),
    .Tile_X3Y25_R_t(R_t_top[600]),
    .Tile_X3Y25_R_f(R_f_top[600]),
    .Tile_X6Y25_R_t(R_t_top[601]),
    .Tile_X6Y25_R_f(R_f_top[601]),
    .Tile_X9Y25_R_t(R_t_top[602]),
    .Tile_X9Y25_R_f(R_f_top[602]),
    .Tile_X12Y25_R_t(R_t_top[603]),
    .Tile_X12Y25_R_f(R_f_top[603]),
    .Tile_X15Y25_R_t(R_t_top[604]),
    .Tile_X15Y25_R_f(R_f_top[604]),
    .Tile_X18Y25_R_t(R_t_top[605]),
    .Tile_X18Y25_R_f(R_f_top[605]),
    .Tile_X21Y25_R_t(R_t_top[606]),
    .Tile_X21Y25_R_f(R_f_top[606]),
    .Tile_X24Y25_R_t(R_t_top[607]),
    .Tile_X24Y25_R_f(R_f_top[607]),
    .Tile_X27Y25_R_t(R_t_top[608]),
    .Tile_X27Y25_R_f(R_f_top[608]),
    .Tile_X30Y25_R_t(R_t_top[609]),
    .Tile_X30Y25_R_f(R_f_top[609]),
    .Tile_X33Y25_R_t(R_t_top[610]),
    .Tile_X33Y25_R_f(R_f_top[610]),
    .Tile_X36Y25_R_t(R_t_top[611]),
    .Tile_X36Y25_R_f(R_f_top[611]),
    .Tile_X39Y25_R_t(R_t_top[612]),
    .Tile_X39Y25_R_f(R_f_top[612]),
    .Tile_X42Y25_R_t(R_t_top[613]),
    .Tile_X42Y25_R_f(R_f_top[613]),
    .Tile_X45Y25_R_t(R_t_top[614]),
    .Tile_X45Y25_R_f(R_f_top[614]),
    .Tile_X48Y25_R_t(R_t_top[615]),
    .Tile_X48Y25_R_f(R_f_top[615]),
    .Tile_X51Y25_R_t(R_t_top[616]),
    .Tile_X51Y25_R_f(R_f_top[616]),
    .Tile_X54Y25_R_t(R_t_top[617]),
    .Tile_X54Y25_R_f(R_f_top[617]),
    .Tile_X57Y25_R_t(R_t_top[618]),
    .Tile_X57Y25_R_f(R_f_top[618]),
    .Tile_X60Y25_R_t(R_t_top[619]),
    .Tile_X60Y25_R_f(R_f_top[619]),
    .Tile_X63Y25_R_t(R_t_top[620]),
    .Tile_X63Y25_R_f(R_f_top[620]),
    .Tile_X66Y25_R_t(R_t_top[621]),
    .Tile_X66Y25_R_f(R_f_top[621]),
    .Tile_X69Y25_R_t(R_t_top[622]),
    .Tile_X69Y25_R_f(R_f_top[622]),
    .Tile_X72Y25_R_t(R_t_top[623]),
    .Tile_X72Y25_R_f(R_f_top[623]),
    .Tile_X75Y25_R_t(R_t_top[624]),
    .Tile_X75Y25_R_f(R_f_top[624]),
    .Tile_X3Y26_R_t(R_t_top[625]),
    .Tile_X3Y26_R_f(R_f_top[625]),
    .Tile_X6Y26_R_t(R_t_top[626]),
    .Tile_X6Y26_R_f(R_f_top[626]),
    .Tile_X9Y26_R_t(R_t_top[627]),
    .Tile_X9Y26_R_f(R_f_top[627]),
    .Tile_X12Y26_R_t(R_t_top[628]),
    .Tile_X12Y26_R_f(R_f_top[628]),
    .Tile_X15Y26_R_t(R_t_top[629]),
    .Tile_X15Y26_R_f(R_f_top[629]),
    .Tile_X18Y26_R_t(R_t_top[630]),
    .Tile_X18Y26_R_f(R_f_top[630]),
    .Tile_X21Y26_R_t(R_t_top[631]),
    .Tile_X21Y26_R_f(R_f_top[631]),
    .Tile_X24Y26_R_t(R_t_top[632]),
    .Tile_X24Y26_R_f(R_f_top[632]),
    .Tile_X27Y26_R_t(R_t_top[633]),
    .Tile_X27Y26_R_f(R_f_top[633]),
    .Tile_X30Y26_R_t(R_t_top[634]),
    .Tile_X30Y26_R_f(R_f_top[634]),
    .Tile_X33Y26_R_t(R_t_top[635]),
    .Tile_X33Y26_R_f(R_f_top[635]),
    .Tile_X36Y26_R_t(R_t_top[636]),
    .Tile_X36Y26_R_f(R_f_top[636]),
    .Tile_X39Y26_R_t(R_t_top[637]),
    .Tile_X39Y26_R_f(R_f_top[637]),
    .Tile_X42Y26_R_t(R_t_top[638]),
    .Tile_X42Y26_R_f(R_f_top[638]),
    .Tile_X45Y26_R_t(R_t_top[639]),
    .Tile_X45Y26_R_f(R_f_top[639]),
    .Tile_X48Y26_R_t(R_t_top[640]),
    .Tile_X48Y26_R_f(R_f_top[640]),
    .Tile_X51Y26_R_t(R_t_top[641]),
    .Tile_X51Y26_R_f(R_f_top[641]),
    .Tile_X54Y26_R_t(R_t_top[642]),
    .Tile_X54Y26_R_f(R_f_top[642]),
    .Tile_X57Y26_R_t(R_t_top[643]),
    .Tile_X57Y26_R_f(R_f_top[643]),
    .Tile_X60Y26_R_t(R_t_top[644]),
    .Tile_X60Y26_R_f(R_f_top[644]),
    .Tile_X63Y26_R_t(R_t_top[645]),
    .Tile_X63Y26_R_f(R_f_top[645]),
    .Tile_X66Y26_R_t(R_t_top[646]),
    .Tile_X66Y26_R_f(R_f_top[646]),
    .Tile_X69Y26_R_t(R_t_top[647]),
    .Tile_X69Y26_R_f(R_f_top[647]),
    .Tile_X72Y26_R_t(R_t_top[648]),
    .Tile_X72Y26_R_f(R_f_top[648]),
    .Tile_X75Y26_R_t(R_t_top[649]),
    .Tile_X75Y26_R_f(R_f_top[649]),
    .Tile_X3Y27_R_t(R_t_top[650]),
    .Tile_X3Y27_R_f(R_f_top[650]),
    .Tile_X6Y27_R_t(R_t_top[651]),
    .Tile_X6Y27_R_f(R_f_top[651]),
    .Tile_X9Y27_R_t(R_t_top[652]),
    .Tile_X9Y27_R_f(R_f_top[652]),
    .Tile_X12Y27_R_t(R_t_top[653]),
    .Tile_X12Y27_R_f(R_f_top[653]),
    .Tile_X15Y27_R_t(R_t_top[654]),
    .Tile_X15Y27_R_f(R_f_top[654]),
    .Tile_X18Y27_R_t(R_t_top[655]),
    .Tile_X18Y27_R_f(R_f_top[655]),
    .Tile_X21Y27_R_t(R_t_top[656]),
    .Tile_X21Y27_R_f(R_f_top[656]),
    .Tile_X24Y27_R_t(R_t_top[657]),
    .Tile_X24Y27_R_f(R_f_top[657]),
    .Tile_X27Y27_R_t(R_t_top[658]),
    .Tile_X27Y27_R_f(R_f_top[658]),
    .Tile_X30Y27_R_t(R_t_top[659]),
    .Tile_X30Y27_R_f(R_f_top[659]),
    .Tile_X33Y27_R_t(R_t_top[660]),
    .Tile_X33Y27_R_f(R_f_top[660]),
    .Tile_X36Y27_R_t(R_t_top[661]),
    .Tile_X36Y27_R_f(R_f_top[661]),
    .Tile_X39Y27_R_t(R_t_top[662]),
    .Tile_X39Y27_R_f(R_f_top[662]),
    .Tile_X42Y27_R_t(R_t_top[663]),
    .Tile_X42Y27_R_f(R_f_top[663]),
    .Tile_X45Y27_R_t(R_t_top[664]),
    .Tile_X45Y27_R_f(R_f_top[664]),
    .Tile_X48Y27_R_t(R_t_top[665]),
    .Tile_X48Y27_R_f(R_f_top[665]),
    .Tile_X51Y27_R_t(R_t_top[666]),
    .Tile_X51Y27_R_f(R_f_top[666]),
    .Tile_X54Y27_R_t(R_t_top[667]),
    .Tile_X54Y27_R_f(R_f_top[667]),
    .Tile_X57Y27_R_t(R_t_top[668]),
    .Tile_X57Y27_R_f(R_f_top[668]),
    .Tile_X60Y27_R_t(R_t_top[669]),
    .Tile_X60Y27_R_f(R_f_top[669]),
    .Tile_X63Y27_R_t(R_t_top[670]),
    .Tile_X63Y27_R_f(R_f_top[670]),
    .Tile_X66Y27_R_t(R_t_top[671]),
    .Tile_X66Y27_R_f(R_f_top[671]),
    .Tile_X69Y27_R_t(R_t_top[672]),
    .Tile_X69Y27_R_f(R_f_top[672]),
    .Tile_X72Y27_R_t(R_t_top[673]),
    .Tile_X72Y27_R_f(R_f_top[673]),
    .Tile_X75Y27_R_t(R_t_top[674]),
    .Tile_X75Y27_R_f(R_f_top[674]),
    .Tile_X3Y28_R_t(R_t_top[675]),
    .Tile_X3Y28_R_f(R_f_top[675]),
    .Tile_X6Y28_R_t(R_t_top[676]),
    .Tile_X6Y28_R_f(R_f_top[676]),
    .Tile_X9Y28_R_t(R_t_top[677]),
    .Tile_X9Y28_R_f(R_f_top[677]),
    .Tile_X12Y28_R_t(R_t_top[678]),
    .Tile_X12Y28_R_f(R_f_top[678]),
    .Tile_X15Y28_R_t(R_t_top[679]),
    .Tile_X15Y28_R_f(R_f_top[679]),
    .Tile_X18Y28_R_t(R_t_top[680]),
    .Tile_X18Y28_R_f(R_f_top[680]),
    .Tile_X21Y28_R_t(R_t_top[681]),
    .Tile_X21Y28_R_f(R_f_top[681]),
    .Tile_X24Y28_R_t(R_t_top[682]),
    .Tile_X24Y28_R_f(R_f_top[682]),
    .Tile_X27Y28_R_t(R_t_top[683]),
    .Tile_X27Y28_R_f(R_f_top[683]),
    .Tile_X30Y28_R_t(R_t_top[684]),
    .Tile_X30Y28_R_f(R_f_top[684]),
    .Tile_X33Y28_R_t(R_t_top[685]),
    .Tile_X33Y28_R_f(R_f_top[685]),
    .Tile_X36Y28_R_t(R_t_top[686]),
    .Tile_X36Y28_R_f(R_f_top[686]),
    .Tile_X39Y28_R_t(R_t_top[687]),
    .Tile_X39Y28_R_f(R_f_top[687]),
    .Tile_X42Y28_R_t(R_t_top[688]),
    .Tile_X42Y28_R_f(R_f_top[688]),
    .Tile_X45Y28_R_t(R_t_top[689]),
    .Tile_X45Y28_R_f(R_f_top[689]),
    .Tile_X48Y28_R_t(R_t_top[690]),
    .Tile_X48Y28_R_f(R_f_top[690]),
    .Tile_X51Y28_R_t(R_t_top[691]),
    .Tile_X51Y28_R_f(R_f_top[691]),
    .Tile_X54Y28_R_t(R_t_top[692]),
    .Tile_X54Y28_R_f(R_f_top[692]),
    .Tile_X57Y28_R_t(R_t_top[693]),
    .Tile_X57Y28_R_f(R_f_top[693]),
    .Tile_X60Y28_R_t(R_t_top[694]),
    .Tile_X60Y28_R_f(R_f_top[694]),
    .Tile_X63Y28_R_t(R_t_top[695]),
    .Tile_X63Y28_R_f(R_f_top[695]),
    .Tile_X66Y28_R_t(R_t_top[696]),
    .Tile_X66Y28_R_f(R_f_top[696]),
    .Tile_X69Y28_R_t(R_t_top[697]),
    .Tile_X69Y28_R_f(R_f_top[697]),
    .Tile_X72Y28_R_t(R_t_top[698]),
    .Tile_X72Y28_R_f(R_f_top[698]),
    .Tile_X75Y28_R_t(R_t_top[699]),
    .Tile_X75Y28_R_f(R_f_top[699]),
    .Tile_X3Y29_R_t(R_t_top[700]),
    .Tile_X3Y29_R_f(R_f_top[700]),
    .Tile_X6Y29_R_t(R_t_top[701]),
    .Tile_X6Y29_R_f(R_f_top[701]),
    .Tile_X9Y29_R_t(R_t_top[702]),
    .Tile_X9Y29_R_f(R_f_top[702]),
    .Tile_X12Y29_R_t(R_t_top[703]),
    .Tile_X12Y29_R_f(R_f_top[703]),
    .Tile_X15Y29_R_t(R_t_top[704]),
    .Tile_X15Y29_R_f(R_f_top[704]),
    .Tile_X18Y29_R_t(R_t_top[705]),
    .Tile_X18Y29_R_f(R_f_top[705]),
    .Tile_X21Y29_R_t(R_t_top[706]),
    .Tile_X21Y29_R_f(R_f_top[706]),
    .Tile_X24Y29_R_t(R_t_top[707]),
    .Tile_X24Y29_R_f(R_f_top[707]),
    .Tile_X27Y29_R_t(R_t_top[708]),
    .Tile_X27Y29_R_f(R_f_top[708]),
    .Tile_X30Y29_R_t(R_t_top[709]),
    .Tile_X30Y29_R_f(R_f_top[709]),
    .Tile_X33Y29_R_t(R_t_top[710]),
    .Tile_X33Y29_R_f(R_f_top[710]),
    .Tile_X36Y29_R_t(R_t_top[711]),
    .Tile_X36Y29_R_f(R_f_top[711]),
    .Tile_X39Y29_R_t(R_t_top[712]),
    .Tile_X39Y29_R_f(R_f_top[712]),
    .Tile_X42Y29_R_t(R_t_top[713]),
    .Tile_X42Y29_R_f(R_f_top[713]),
    .Tile_X45Y29_R_t(R_t_top[714]),
    .Tile_X45Y29_R_f(R_f_top[714]),
    .Tile_X48Y29_R_t(R_t_top[715]),
    .Tile_X48Y29_R_f(R_f_top[715]),
    .Tile_X51Y29_R_t(R_t_top[716]),
    .Tile_X51Y29_R_f(R_f_top[716]),
    .Tile_X54Y29_R_t(R_t_top[717]),
    .Tile_X54Y29_R_f(R_f_top[717]),
    .Tile_X57Y29_R_t(R_t_top[718]),
    .Tile_X57Y29_R_f(R_f_top[718]),
    .Tile_X60Y29_R_t(R_t_top[719]),
    .Tile_X60Y29_R_f(R_f_top[719]),
    .Tile_X63Y29_R_t(R_t_top[720]),
    .Tile_X63Y29_R_f(R_f_top[720]),
    .Tile_X66Y29_R_t(R_t_top[721]),
    .Tile_X66Y29_R_f(R_f_top[721]),
    .Tile_X69Y29_R_t(R_t_top[722]),
    .Tile_X69Y29_R_f(R_f_top[722]),
    .Tile_X72Y29_R_t(R_t_top[723]),
    .Tile_X72Y29_R_f(R_f_top[723]),
    .Tile_X75Y29_R_t(R_t_top[724]),
    .Tile_X75Y29_R_f(R_f_top[724]),
    .Tile_X3Y30_R_t(R_t_top[725]),
    .Tile_X3Y30_R_f(R_f_top[725]),
    .Tile_X6Y30_R_t(R_t_top[726]),
    .Tile_X6Y30_R_f(R_f_top[726]),
    .Tile_X9Y30_R_t(R_t_top[727]),
    .Tile_X9Y30_R_f(R_f_top[727]),
    .Tile_X12Y30_R_t(R_t_top[728]),
    .Tile_X12Y30_R_f(R_f_top[728]),
    .Tile_X15Y30_R_t(R_t_top[729]),
    .Tile_X15Y30_R_f(R_f_top[729]),
    .Tile_X18Y30_R_t(R_t_top[730]),
    .Tile_X18Y30_R_f(R_f_top[730]),
    .Tile_X21Y30_R_t(R_t_top[731]),
    .Tile_X21Y30_R_f(R_f_top[731]),
    .Tile_X24Y30_R_t(R_t_top[732]),
    .Tile_X24Y30_R_f(R_f_top[732]),
    .Tile_X27Y30_R_t(R_t_top[733]),
    .Tile_X27Y30_R_f(R_f_top[733]),
    .Tile_X30Y30_R_t(R_t_top[734]),
    .Tile_X30Y30_R_f(R_f_top[734]),
    .Tile_X33Y30_R_t(R_t_top[735]),
    .Tile_X33Y30_R_f(R_f_top[735]),
    .Tile_X36Y30_R_t(R_t_top[736]),
    .Tile_X36Y30_R_f(R_f_top[736]),
    .Tile_X39Y30_R_t(R_t_top[737]),
    .Tile_X39Y30_R_f(R_f_top[737]),
    .Tile_X42Y30_R_t(R_t_top[738]),
    .Tile_X42Y30_R_f(R_f_top[738]),
    .Tile_X45Y30_R_t(R_t_top[739]),
    .Tile_X45Y30_R_f(R_f_top[739]),
    .Tile_X48Y30_R_t(R_t_top[740]),
    .Tile_X48Y30_R_f(R_f_top[740]),
    .Tile_X51Y30_R_t(R_t_top[741]),
    .Tile_X51Y30_R_f(R_f_top[741]),
    .Tile_X54Y30_R_t(R_t_top[742]),
    .Tile_X54Y30_R_f(R_f_top[742]),
    .Tile_X57Y30_R_t(R_t_top[743]),
    .Tile_X57Y30_R_f(R_f_top[743]),
    .Tile_X60Y30_R_t(R_t_top[744]),
    .Tile_X60Y30_R_f(R_f_top[744]),
    .Tile_X63Y30_R_t(R_t_top[745]),
    .Tile_X63Y30_R_f(R_f_top[745]),
    .Tile_X66Y30_R_t(R_t_top[746]),
    .Tile_X66Y30_R_f(R_f_top[746]),
    .Tile_X69Y30_R_t(R_t_top[747]),
    .Tile_X69Y30_R_f(R_f_top[747]),
    .Tile_X72Y30_R_t(R_t_top[748]),
    .Tile_X72Y30_R_f(R_f_top[748]),
    .Tile_X75Y30_R_t(R_t_top[749]),
    .Tile_X75Y30_R_f(R_f_top[749]),
    .Tile_X3Y31_R_t(R_t_top[750]),
    .Tile_X3Y31_R_f(R_f_top[750]),
    .Tile_X6Y31_R_t(R_t_top[751]),
    .Tile_X6Y31_R_f(R_f_top[751]),
    .Tile_X9Y31_R_t(R_t_top[752]),
    .Tile_X9Y31_R_f(R_f_top[752]),
    .Tile_X12Y31_R_t(R_t_top[753]),
    .Tile_X12Y31_R_f(R_f_top[753]),
    .Tile_X15Y31_R_t(R_t_top[754]),
    .Tile_X15Y31_R_f(R_f_top[754]),
    .Tile_X18Y31_R_t(R_t_top[755]),
    .Tile_X18Y31_R_f(R_f_top[755]),
    .Tile_X21Y31_R_t(R_t_top[756]),
    .Tile_X21Y31_R_f(R_f_top[756]),
    .Tile_X24Y31_R_t(R_t_top[757]),
    .Tile_X24Y31_R_f(R_f_top[757]),
    .Tile_X27Y31_R_t(R_t_top[758]),
    .Tile_X27Y31_R_f(R_f_top[758]),
    .Tile_X30Y31_R_t(R_t_top[759]),
    .Tile_X30Y31_R_f(R_f_top[759]),
    .Tile_X33Y31_R_t(R_t_top[760]),
    .Tile_X33Y31_R_f(R_f_top[760]),
    .Tile_X36Y31_R_t(R_t_top[761]),
    .Tile_X36Y31_R_f(R_f_top[761]),
    .Tile_X39Y31_R_t(R_t_top[762]),
    .Tile_X39Y31_R_f(R_f_top[762]),
    .Tile_X42Y31_R_t(R_t_top[763]),
    .Tile_X42Y31_R_f(R_f_top[763]),
    .Tile_X45Y31_R_t(R_t_top[764]),
    .Tile_X45Y31_R_f(R_f_top[764]),
    .Tile_X48Y31_R_t(R_t_top[765]),
    .Tile_X48Y31_R_f(R_f_top[765]),
    .Tile_X51Y31_R_t(R_t_top[766]),
    .Tile_X51Y31_R_f(R_f_top[766]),
    .Tile_X54Y31_R_t(R_t_top[767]),
    .Tile_X54Y31_R_f(R_f_top[767]),
    .Tile_X57Y31_R_t(R_t_top[768]),
    .Tile_X57Y31_R_f(R_f_top[768]),
    .Tile_X60Y31_R_t(R_t_top[769]),
    .Tile_X60Y31_R_f(R_f_top[769]),
    .Tile_X63Y31_R_t(R_t_top[770]),
    .Tile_X63Y31_R_f(R_f_top[770]),
    .Tile_X66Y31_R_t(R_t_top[771]),
    .Tile_X66Y31_R_f(R_f_top[771]),
    .Tile_X69Y31_R_t(R_t_top[772]),
    .Tile_X69Y31_R_f(R_f_top[772]),
    .Tile_X72Y31_R_t(R_t_top[773]),
    .Tile_X72Y31_R_f(R_f_top[773]),
    .Tile_X75Y31_R_t(R_t_top[774]),
    .Tile_X75Y31_R_f(R_f_top[774]),
    .Tile_X3Y32_R_t(R_t_top[775]),
    .Tile_X3Y32_R_f(R_f_top[775]),
    .Tile_X6Y32_R_t(R_t_top[776]),
    .Tile_X6Y32_R_f(R_f_top[776]),
    .Tile_X9Y32_R_t(R_t_top[777]),
    .Tile_X9Y32_R_f(R_f_top[777]),
    .Tile_X12Y32_R_t(R_t_top[778]),
    .Tile_X12Y32_R_f(R_f_top[778]),
    .Tile_X15Y32_R_t(R_t_top[779]),
    .Tile_X15Y32_R_f(R_f_top[779]),
    .Tile_X18Y32_R_t(R_t_top[780]),
    .Tile_X18Y32_R_f(R_f_top[780]),
    .Tile_X21Y32_R_t(R_t_top[781]),
    .Tile_X21Y32_R_f(R_f_top[781]),
    .Tile_X24Y32_R_t(R_t_top[782]),
    .Tile_X24Y32_R_f(R_f_top[782]),
    .Tile_X27Y32_R_t(R_t_top[783]),
    .Tile_X27Y32_R_f(R_f_top[783]),
    .Tile_X30Y32_R_t(R_t_top[784]),
    .Tile_X30Y32_R_f(R_f_top[784]),
    .Tile_X33Y32_R_t(R_t_top[785]),
    .Tile_X33Y32_R_f(R_f_top[785]),
    .Tile_X36Y32_R_t(R_t_top[786]),
    .Tile_X36Y32_R_f(R_f_top[786]),
    .Tile_X39Y32_R_t(R_t_top[787]),
    .Tile_X39Y32_R_f(R_f_top[787]),
    .Tile_X42Y32_R_t(R_t_top[788]),
    .Tile_X42Y32_R_f(R_f_top[788]),
    .Tile_X45Y32_R_t(R_t_top[789]),
    .Tile_X45Y32_R_f(R_f_top[789]),
    .Tile_X48Y32_R_t(R_t_top[790]),
    .Tile_X48Y32_R_f(R_f_top[790]),
    .Tile_X51Y32_R_t(R_t_top[791]),
    .Tile_X51Y32_R_f(R_f_top[791]),
    .Tile_X54Y32_R_t(R_t_top[792]),
    .Tile_X54Y32_R_f(R_f_top[792]),
    .Tile_X57Y32_R_t(R_t_top[793]),
    .Tile_X57Y32_R_f(R_f_top[793]),
    .Tile_X60Y32_R_t(R_t_top[794]),
    .Tile_X60Y32_R_f(R_f_top[794]),
    .Tile_X63Y32_R_t(R_t_top[795]),
    .Tile_X63Y32_R_f(R_f_top[795]),
    .Tile_X66Y32_R_t(R_t_top[796]),
    .Tile_X66Y32_R_f(R_f_top[796]),
    .Tile_X69Y32_R_t(R_t_top[797]),
    .Tile_X69Y32_R_f(R_f_top[797]),
    .Tile_X72Y32_R_t(R_t_top[798]),
    .Tile_X72Y32_R_f(R_f_top[798]),
    .Tile_X75Y32_R_t(R_t_top[799]),
    .Tile_X75Y32_R_f(R_f_top[799]),
    .Tile_X3Y33_R_t(R_t_top[800]),
    .Tile_X3Y33_R_f(R_f_top[800]),
    .Tile_X6Y33_R_t(R_t_top[801]),
    .Tile_X6Y33_R_f(R_f_top[801]),
    .Tile_X9Y33_R_t(R_t_top[802]),
    .Tile_X9Y33_R_f(R_f_top[802]),
    .Tile_X12Y33_R_t(R_t_top[803]),
    .Tile_X12Y33_R_f(R_f_top[803]),
    .Tile_X15Y33_R_t(R_t_top[804]),
    .Tile_X15Y33_R_f(R_f_top[804]),
    .Tile_X18Y33_R_t(R_t_top[805]),
    .Tile_X18Y33_R_f(R_f_top[805]),
    .Tile_X21Y33_R_t(R_t_top[806]),
    .Tile_X21Y33_R_f(R_f_top[806]),
    .Tile_X24Y33_R_t(R_t_top[807]),
    .Tile_X24Y33_R_f(R_f_top[807]),
    .Tile_X27Y33_R_t(R_t_top[808]),
    .Tile_X27Y33_R_f(R_f_top[808]),
    .Tile_X30Y33_R_t(R_t_top[809]),
    .Tile_X30Y33_R_f(R_f_top[809]),
    .Tile_X33Y33_R_t(R_t_top[810]),
    .Tile_X33Y33_R_f(R_f_top[810]),
    .Tile_X36Y33_R_t(R_t_top[811]),
    .Tile_X36Y33_R_f(R_f_top[811]),
    .Tile_X39Y33_R_t(R_t_top[812]),
    .Tile_X39Y33_R_f(R_f_top[812]),
    .Tile_X42Y33_R_t(R_t_top[813]),
    .Tile_X42Y33_R_f(R_f_top[813]),
    .Tile_X45Y33_R_t(R_t_top[814]),
    .Tile_X45Y33_R_f(R_f_top[814]),
    .Tile_X48Y33_R_t(R_t_top[815]),
    .Tile_X48Y33_R_f(R_f_top[815]),
    .Tile_X51Y33_R_t(R_t_top[816]),
    .Tile_X51Y33_R_f(R_f_top[816]),
    .Tile_X54Y33_R_t(R_t_top[817]),
    .Tile_X54Y33_R_f(R_f_top[817]),
    .Tile_X57Y33_R_t(R_t_top[818]),
    .Tile_X57Y33_R_f(R_f_top[818]),
    .Tile_X60Y33_R_t(R_t_top[819]),
    .Tile_X60Y33_R_f(R_f_top[819]),
    .Tile_X63Y33_R_t(R_t_top[820]),
    .Tile_X63Y33_R_f(R_f_top[820]),
    .Tile_X66Y33_R_t(R_t_top[821]),
    .Tile_X66Y33_R_f(R_f_top[821]),
    .Tile_X69Y33_R_t(R_t_top[822]),
    .Tile_X69Y33_R_f(R_f_top[822]),
    .Tile_X72Y33_R_t(R_t_top[823]),
    .Tile_X72Y33_R_f(R_f_top[823]),
    .Tile_X75Y33_R_t(R_t_top[824]),
    .Tile_X75Y33_R_f(R_f_top[824]),
    .Tile_X3Y34_R_t(R_t_top[825]),
    .Tile_X3Y34_R_f(R_f_top[825]),
    .Tile_X6Y34_R_t(R_t_top[826]),
    .Tile_X6Y34_R_f(R_f_top[826]),
    .Tile_X9Y34_R_t(R_t_top[827]),
    .Tile_X9Y34_R_f(R_f_top[827]),
    .Tile_X12Y34_R_t(R_t_top[828]),
    .Tile_X12Y34_R_f(R_f_top[828]),
    .Tile_X15Y34_R_t(R_t_top[829]),
    .Tile_X15Y34_R_f(R_f_top[829]),
    .Tile_X18Y34_R_t(R_t_top[830]),
    .Tile_X18Y34_R_f(R_f_top[830]),
    .Tile_X21Y34_R_t(R_t_top[831]),
    .Tile_X21Y34_R_f(R_f_top[831]),
    .Tile_X24Y34_R_t(R_t_top[832]),
    .Tile_X24Y34_R_f(R_f_top[832]),
    .Tile_X27Y34_R_t(R_t_top[833]),
    .Tile_X27Y34_R_f(R_f_top[833]),
    .Tile_X30Y34_R_t(R_t_top[834]),
    .Tile_X30Y34_R_f(R_f_top[834]),
    .Tile_X33Y34_R_t(R_t_top[835]),
    .Tile_X33Y34_R_f(R_f_top[835]),
    .Tile_X36Y34_R_t(R_t_top[836]),
    .Tile_X36Y34_R_f(R_f_top[836]),
    .Tile_X39Y34_R_t(R_t_top[837]),
    .Tile_X39Y34_R_f(R_f_top[837]),
    .Tile_X42Y34_R_t(R_t_top[838]),
    .Tile_X42Y34_R_f(R_f_top[838]),
    .Tile_X45Y34_R_t(R_t_top[839]),
    .Tile_X45Y34_R_f(R_f_top[839]),
    .Tile_X48Y34_R_t(R_t_top[840]),
    .Tile_X48Y34_R_f(R_f_top[840]),
    .Tile_X51Y34_R_t(R_t_top[841]),
    .Tile_X51Y34_R_f(R_f_top[841]),
    .Tile_X54Y34_R_t(R_t_top[842]),
    .Tile_X54Y34_R_f(R_f_top[842]),
    .Tile_X57Y34_R_t(R_t_top[843]),
    .Tile_X57Y34_R_f(R_f_top[843]),
    .Tile_X60Y34_R_t(R_t_top[844]),
    .Tile_X60Y34_R_f(R_f_top[844]),
    .Tile_X63Y34_R_t(R_t_top[845]),
    .Tile_X63Y34_R_f(R_f_top[845]),
    .Tile_X66Y34_R_t(R_t_top[846]),
    .Tile_X66Y34_R_f(R_f_top[846]),
    .Tile_X69Y34_R_t(R_t_top[847]),
    .Tile_X69Y34_R_f(R_f_top[847]),
    .Tile_X72Y34_R_t(R_t_top[848]),
    .Tile_X72Y34_R_f(R_f_top[848]),
    .Tile_X75Y34_R_t(R_t_top[849]),
    .Tile_X75Y34_R_f(R_f_top[849]),
    .Tile_X3Y35_R_t(R_t_top[850]),
    .Tile_X3Y35_R_f(R_f_top[850]),
    .Tile_X6Y35_R_t(R_t_top[851]),
    .Tile_X6Y35_R_f(R_f_top[851]),
    .Tile_X9Y35_R_t(R_t_top[852]),
    .Tile_X9Y35_R_f(R_f_top[852]),
    .Tile_X12Y35_R_t(R_t_top[853]),
    .Tile_X12Y35_R_f(R_f_top[853]),
    .Tile_X15Y35_R_t(R_t_top[854]),
    .Tile_X15Y35_R_f(R_f_top[854]),
    .Tile_X18Y35_R_t(R_t_top[855]),
    .Tile_X18Y35_R_f(R_f_top[855]),
    .Tile_X21Y35_R_t(R_t_top[856]),
    .Tile_X21Y35_R_f(R_f_top[856]),
    .Tile_X24Y35_R_t(R_t_top[857]),
    .Tile_X24Y35_R_f(R_f_top[857]),
    .Tile_X27Y35_R_t(R_t_top[858]),
    .Tile_X27Y35_R_f(R_f_top[858]),
    .Tile_X30Y35_R_t(R_t_top[859]),
    .Tile_X30Y35_R_f(R_f_top[859]),
    .Tile_X33Y35_R_t(R_t_top[860]),
    .Tile_X33Y35_R_f(R_f_top[860]),
    .Tile_X36Y35_R_t(R_t_top[861]),
    .Tile_X36Y35_R_f(R_f_top[861]),
    .Tile_X39Y35_R_t(R_t_top[862]),
    .Tile_X39Y35_R_f(R_f_top[862]),
    .Tile_X42Y35_R_t(R_t_top[863]),
    .Tile_X42Y35_R_f(R_f_top[863]),
    .Tile_X45Y35_R_t(R_t_top[864]),
    .Tile_X45Y35_R_f(R_f_top[864]),
    .Tile_X48Y35_R_t(R_t_top[865]),
    .Tile_X48Y35_R_f(R_f_top[865]),
    .Tile_X51Y35_R_t(R_t_top[866]),
    .Tile_X51Y35_R_f(R_f_top[866]),
    .Tile_X54Y35_R_t(R_t_top[867]),
    .Tile_X54Y35_R_f(R_f_top[867]),
    .Tile_X57Y35_R_t(R_t_top[868]),
    .Tile_X57Y35_R_f(R_f_top[868]),
    .Tile_X60Y35_R_t(R_t_top[869]),
    .Tile_X60Y35_R_f(R_f_top[869]),
    .Tile_X63Y35_R_t(R_t_top[870]),
    .Tile_X63Y35_R_f(R_f_top[870]),
    .Tile_X66Y35_R_t(R_t_top[871]),
    .Tile_X66Y35_R_f(R_f_top[871]),
    .Tile_X69Y35_R_t(R_t_top[872]),
    .Tile_X69Y35_R_f(R_f_top[872]),
    .Tile_X72Y35_R_t(R_t_top[873]),
    .Tile_X72Y35_R_f(R_f_top[873]),
    .Tile_X75Y35_R_t(R_t_top[874]),
    .Tile_X75Y35_R_f(R_f_top[874]),
    .Tile_X3Y36_R_t(R_t_top[875]),
    .Tile_X3Y36_R_f(R_f_top[875]),
    .Tile_X6Y36_R_t(R_t_top[876]),
    .Tile_X6Y36_R_f(R_f_top[876]),
    .Tile_X9Y36_R_t(R_t_top[877]),
    .Tile_X9Y36_R_f(R_f_top[877]),
    .Tile_X12Y36_R_t(R_t_top[878]),
    .Tile_X12Y36_R_f(R_f_top[878]),
    .Tile_X15Y36_R_t(R_t_top[879]),
    .Tile_X15Y36_R_f(R_f_top[879]),
    .Tile_X18Y36_R_t(R_t_top[880]),
    .Tile_X18Y36_R_f(R_f_top[880]),
    .Tile_X21Y36_R_t(R_t_top[881]),
    .Tile_X21Y36_R_f(R_f_top[881]),
    .Tile_X24Y36_R_t(R_t_top[882]),
    .Tile_X24Y36_R_f(R_f_top[882]),
    .Tile_X27Y36_R_t(R_t_top[883]),
    .Tile_X27Y36_R_f(R_f_top[883]),
    .Tile_X30Y36_R_t(R_t_top[884]),
    .Tile_X30Y36_R_f(R_f_top[884]),
    .Tile_X33Y36_R_t(R_t_top[885]),
    .Tile_X33Y36_R_f(R_f_top[885]),
    .Tile_X36Y36_R_t(R_t_top[886]),
    .Tile_X36Y36_R_f(R_f_top[886]),
    .Tile_X39Y36_R_t(R_t_top[887]),
    .Tile_X39Y36_R_f(R_f_top[887]),
    .Tile_X42Y36_R_t(R_t_top[888]),
    .Tile_X42Y36_R_f(R_f_top[888]),
    .Tile_X45Y36_R_t(R_t_top[889]),
    .Tile_X45Y36_R_f(R_f_top[889]),
    .Tile_X48Y36_R_t(R_t_top[890]),
    .Tile_X48Y36_R_f(R_f_top[890]),
    .Tile_X51Y36_R_t(R_t_top[891]),
    .Tile_X51Y36_R_f(R_f_top[891]),
    .Tile_X54Y36_R_t(R_t_top[892]),
    .Tile_X54Y36_R_f(R_f_top[892]),
    .Tile_X57Y36_R_t(R_t_top[893]),
    .Tile_X57Y36_R_f(R_f_top[893]),
    .Tile_X60Y36_R_t(R_t_top[894]),
    .Tile_X60Y36_R_f(R_f_top[894]),
    .Tile_X63Y36_R_t(R_t_top[895]),
    .Tile_X63Y36_R_f(R_f_top[895]),
    .Tile_X66Y36_R_t(R_t_top[896]),
    .Tile_X66Y36_R_f(R_f_top[896]),
    .Tile_X69Y36_R_t(R_t_top[897]),
    .Tile_X69Y36_R_f(R_f_top[897]),
    .Tile_X72Y36_R_t(R_t_top[898]),
    .Tile_X72Y36_R_f(R_f_top[898]),
    .Tile_X75Y36_R_t(R_t_top[899]),
    .Tile_X75Y36_R_f(R_f_top[899]),
    .Tile_X3Y37_R_t(R_t_top[900]),
    .Tile_X3Y37_R_f(R_f_top[900]),
    .Tile_X6Y37_R_t(R_t_top[901]),
    .Tile_X6Y37_R_f(R_f_top[901]),
    .Tile_X9Y37_R_t(R_t_top[902]),
    .Tile_X9Y37_R_f(R_f_top[902]),
    .Tile_X12Y37_R_t(R_t_top[903]),
    .Tile_X12Y37_R_f(R_f_top[903]),
    .Tile_X15Y37_R_t(R_t_top[904]),
    .Tile_X15Y37_R_f(R_f_top[904]),
    .Tile_X18Y37_R_t(R_t_top[905]),
    .Tile_X18Y37_R_f(R_f_top[905]),
    .Tile_X21Y37_R_t(R_t_top[906]),
    .Tile_X21Y37_R_f(R_f_top[906]),
    .Tile_X24Y37_R_t(R_t_top[907]),
    .Tile_X24Y37_R_f(R_f_top[907]),
    .Tile_X27Y37_R_t(R_t_top[908]),
    .Tile_X27Y37_R_f(R_f_top[908]),
    .Tile_X30Y37_R_t(R_t_top[909]),
    .Tile_X30Y37_R_f(R_f_top[909]),
    .Tile_X33Y37_R_t(R_t_top[910]),
    .Tile_X33Y37_R_f(R_f_top[910]),
    .Tile_X36Y37_R_t(R_t_top[911]),
    .Tile_X36Y37_R_f(R_f_top[911]),
    .Tile_X39Y37_R_t(R_t_top[912]),
    .Tile_X39Y37_R_f(R_f_top[912]),
    .Tile_X42Y37_R_t(R_t_top[913]),
    .Tile_X42Y37_R_f(R_f_top[913]),
    .Tile_X45Y37_R_t(R_t_top[914]),
    .Tile_X45Y37_R_f(R_f_top[914]),
    .Tile_X48Y37_R_t(R_t_top[915]),
    .Tile_X48Y37_R_f(R_f_top[915]),
    .Tile_X51Y37_R_t(R_t_top[916]),
    .Tile_X51Y37_R_f(R_f_top[916]),
    .Tile_X54Y37_R_t(R_t_top[917]),
    .Tile_X54Y37_R_f(R_f_top[917]),
    .Tile_X57Y37_R_t(R_t_top[918]),
    .Tile_X57Y37_R_f(R_f_top[918]),
    .Tile_X60Y37_R_t(R_t_top[919]),
    .Tile_X60Y37_R_f(R_f_top[919]),
    .Tile_X63Y37_R_t(R_t_top[920]),
    .Tile_X63Y37_R_f(R_f_top[920]),
    .Tile_X66Y37_R_t(R_t_top[921]),
    .Tile_X66Y37_R_f(R_f_top[921]),
    .Tile_X69Y37_R_t(R_t_top[922]),
    .Tile_X69Y37_R_f(R_f_top[922]),
    .Tile_X72Y37_R_t(R_t_top[923]),
    .Tile_X72Y37_R_f(R_f_top[923]),
    .Tile_X75Y37_R_t(R_t_top[924]),
    .Tile_X75Y37_R_f(R_f_top[924]),
    .Tile_X3Y38_R_t(R_t_top[925]),
    .Tile_X3Y38_R_f(R_f_top[925]),
    .Tile_X6Y38_R_t(R_t_top[926]),
    .Tile_X6Y38_R_f(R_f_top[926]),
    .Tile_X9Y38_R_t(R_t_top[927]),
    .Tile_X9Y38_R_f(R_f_top[927]),
    .Tile_X12Y38_R_t(R_t_top[928]),
    .Tile_X12Y38_R_f(R_f_top[928]),
    .Tile_X15Y38_R_t(R_t_top[929]),
    .Tile_X15Y38_R_f(R_f_top[929]),
    .Tile_X18Y38_R_t(R_t_top[930]),
    .Tile_X18Y38_R_f(R_f_top[930]),
    .Tile_X21Y38_R_t(R_t_top[931]),
    .Tile_X21Y38_R_f(R_f_top[931]),
    .Tile_X24Y38_R_t(R_t_top[932]),
    .Tile_X24Y38_R_f(R_f_top[932]),
    .Tile_X27Y38_R_t(R_t_top[933]),
    .Tile_X27Y38_R_f(R_f_top[933]),
    .Tile_X30Y38_R_t(R_t_top[934]),
    .Tile_X30Y38_R_f(R_f_top[934]),
    .Tile_X33Y38_R_t(R_t_top[935]),
    .Tile_X33Y38_R_f(R_f_top[935]),
    .Tile_X36Y38_R_t(R_t_top[936]),
    .Tile_X36Y38_R_f(R_f_top[936]),
    .Tile_X39Y38_R_t(R_t_top[937]),
    .Tile_X39Y38_R_f(R_f_top[937]),
    .Tile_X42Y38_R_t(R_t_top[938]),
    .Tile_X42Y38_R_f(R_f_top[938]),
    .Tile_X45Y38_R_t(R_t_top[939]),
    .Tile_X45Y38_R_f(R_f_top[939]),
    .Tile_X48Y38_R_t(R_t_top[940]),
    .Tile_X48Y38_R_f(R_f_top[940]),
    .Tile_X51Y38_R_t(R_t_top[941]),
    .Tile_X51Y38_R_f(R_f_top[941]),
    .Tile_X54Y38_R_t(R_t_top[942]),
    .Tile_X54Y38_R_f(R_f_top[942]),
    .Tile_X57Y38_R_t(R_t_top[943]),
    .Tile_X57Y38_R_f(R_f_top[943]),
    .Tile_X60Y38_R_t(R_t_top[944]),
    .Tile_X60Y38_R_f(R_f_top[944]),
    .Tile_X63Y38_R_t(R_t_top[945]),
    .Tile_X63Y38_R_f(R_f_top[945]),
    .Tile_X66Y38_R_t(R_t_top[946]),
    .Tile_X66Y38_R_f(R_f_top[946]),
    .Tile_X69Y38_R_t(R_t_top[947]),
    .Tile_X69Y38_R_f(R_f_top[947]),
    .Tile_X72Y38_R_t(R_t_top[948]),
    .Tile_X72Y38_R_f(R_f_top[948]),
    .Tile_X75Y38_R_t(R_t_top[949]),
    .Tile_X75Y38_R_f(R_f_top[949]),
    .Tile_X3Y39_R_t(R_t_top[950]),
    .Tile_X3Y39_R_f(R_f_top[950]),
    .Tile_X6Y39_R_t(R_t_top[951]),
    .Tile_X6Y39_R_f(R_f_top[951]),
    .Tile_X9Y39_R_t(R_t_top[952]),
    .Tile_X9Y39_R_f(R_f_top[952]),
    .Tile_X12Y39_R_t(R_t_top[953]),
    .Tile_X12Y39_R_f(R_f_top[953]),
    .Tile_X15Y39_R_t(R_t_top[954]),
    .Tile_X15Y39_R_f(R_f_top[954]),
    .Tile_X18Y39_R_t(R_t_top[955]),
    .Tile_X18Y39_R_f(R_f_top[955]),
    .Tile_X21Y39_R_t(R_t_top[956]),
    .Tile_X21Y39_R_f(R_f_top[956]),
    .Tile_X24Y39_R_t(R_t_top[957]),
    .Tile_X24Y39_R_f(R_f_top[957]),
    .Tile_X27Y39_R_t(R_t_top[958]),
    .Tile_X27Y39_R_f(R_f_top[958]),
    .Tile_X30Y39_R_t(R_t_top[959]),
    .Tile_X30Y39_R_f(R_f_top[959]),
    .Tile_X33Y39_R_t(R_t_top[960]),
    .Tile_X33Y39_R_f(R_f_top[960]),
    .Tile_X36Y39_R_t(R_t_top[961]),
    .Tile_X36Y39_R_f(R_f_top[961]),
    .Tile_X39Y39_R_t(R_t_top[962]),
    .Tile_X39Y39_R_f(R_f_top[962]),
    .Tile_X42Y39_R_t(R_t_top[963]),
    .Tile_X42Y39_R_f(R_f_top[963]),
    .Tile_X45Y39_R_t(R_t_top[964]),
    .Tile_X45Y39_R_f(R_f_top[964]),
    .Tile_X48Y39_R_t(R_t_top[965]),
    .Tile_X48Y39_R_f(R_f_top[965]),
    .Tile_X51Y39_R_t(R_t_top[966]),
    .Tile_X51Y39_R_f(R_f_top[966]),
    .Tile_X54Y39_R_t(R_t_top[967]),
    .Tile_X54Y39_R_f(R_f_top[967]),
    .Tile_X57Y39_R_t(R_t_top[968]),
    .Tile_X57Y39_R_f(R_f_top[968]),
    .Tile_X60Y39_R_t(R_t_top[969]),
    .Tile_X60Y39_R_f(R_f_top[969]),
    .Tile_X63Y39_R_t(R_t_top[970]),
    .Tile_X63Y39_R_f(R_f_top[970]),
    .Tile_X66Y39_R_t(R_t_top[971]),
    .Tile_X66Y39_R_f(R_f_top[971]),
    .Tile_X69Y39_R_t(R_t_top[972]),
    .Tile_X69Y39_R_f(R_f_top[972]),
    .Tile_X72Y39_R_t(R_t_top[973]),
    .Tile_X72Y39_R_f(R_f_top[973]),
    .Tile_X75Y39_R_t(R_t_top[974]),
    .Tile_X75Y39_R_f(R_f_top[974]),
    .Tile_X3Y40_R_t(R_t_top[975]),
    .Tile_X3Y40_R_f(R_f_top[975]),
    .Tile_X6Y40_R_t(R_t_top[976]),
    .Tile_X6Y40_R_f(R_f_top[976]),
    .Tile_X9Y40_R_t(R_t_top[977]),
    .Tile_X9Y40_R_f(R_f_top[977]),
    .Tile_X12Y40_R_t(R_t_top[978]),
    .Tile_X12Y40_R_f(R_f_top[978]),
    .Tile_X15Y40_R_t(R_t_top[979]),
    .Tile_X15Y40_R_f(R_f_top[979]),
    .Tile_X18Y40_R_t(R_t_top[980]),
    .Tile_X18Y40_R_f(R_f_top[980]),
    .Tile_X21Y40_R_t(R_t_top[981]),
    .Tile_X21Y40_R_f(R_f_top[981]),
    .Tile_X24Y40_R_t(R_t_top[982]),
    .Tile_X24Y40_R_f(R_f_top[982]),
    .Tile_X27Y40_R_t(R_t_top[983]),
    .Tile_X27Y40_R_f(R_f_top[983]),
    .Tile_X30Y40_R_t(R_t_top[984]),
    .Tile_X30Y40_R_f(R_f_top[984]),
    .Tile_X33Y40_R_t(R_t_top[985]),
    .Tile_X33Y40_R_f(R_f_top[985]),
    .Tile_X36Y40_R_t(R_t_top[986]),
    .Tile_X36Y40_R_f(R_f_top[986]),
    .Tile_X39Y40_R_t(R_t_top[987]),
    .Tile_X39Y40_R_f(R_f_top[987]),
    .Tile_X42Y40_R_t(R_t_top[988]),
    .Tile_X42Y40_R_f(R_f_top[988]),
    .Tile_X45Y40_R_t(R_t_top[989]),
    .Tile_X45Y40_R_f(R_f_top[989]),
    .Tile_X48Y40_R_t(R_t_top[990]),
    .Tile_X48Y40_R_f(R_f_top[990]),
    .Tile_X51Y40_R_t(R_t_top[991]),
    .Tile_X51Y40_R_f(R_f_top[991]),
    .Tile_X54Y40_R_t(R_t_top[992]),
    .Tile_X54Y40_R_f(R_f_top[992]),
    .Tile_X57Y40_R_t(R_t_top[993]),
    .Tile_X57Y40_R_f(R_f_top[993]),
    .Tile_X60Y40_R_t(R_t_top[994]),
    .Tile_X60Y40_R_f(R_f_top[994]),
    .Tile_X63Y40_R_t(R_t_top[995]),
    .Tile_X63Y40_R_f(R_f_top[995]),
    .Tile_X66Y40_R_t(R_t_top[996]),
    .Tile_X66Y40_R_f(R_f_top[996]),
    .Tile_X69Y40_R_t(R_t_top[997]),
    .Tile_X69Y40_R_f(R_f_top[997]),
    .Tile_X72Y40_R_t(R_t_top[998]),
    .Tile_X72Y40_R_f(R_f_top[998]),
    .Tile_X75Y40_R_t(R_t_top[999]),
    .Tile_X75Y40_R_f(R_f_top[999]),
    .Tile_X3Y41_R_t(R_t_top[1000]),
    .Tile_X3Y41_R_f(R_f_top[1000]),
    .Tile_X6Y41_R_t(R_t_top[1001]),
    .Tile_X6Y41_R_f(R_f_top[1001]),
    .Tile_X9Y41_R_t(R_t_top[1002]),
    .Tile_X9Y41_R_f(R_f_top[1002]),
    .Tile_X12Y41_R_t(R_t_top[1003]),
    .Tile_X12Y41_R_f(R_f_top[1003]),
    .Tile_X15Y41_R_t(R_t_top[1004]),
    .Tile_X15Y41_R_f(R_f_top[1004]),
    .Tile_X18Y41_R_t(R_t_top[1005]),
    .Tile_X18Y41_R_f(R_f_top[1005]),
    .Tile_X21Y41_R_t(R_t_top[1006]),
    .Tile_X21Y41_R_f(R_f_top[1006]),
    .Tile_X24Y41_R_t(R_t_top[1007]),
    .Tile_X24Y41_R_f(R_f_top[1007]),
    .Tile_X27Y41_R_t(R_t_top[1008]),
    .Tile_X27Y41_R_f(R_f_top[1008]),
    .Tile_X30Y41_R_t(R_t_top[1009]),
    .Tile_X30Y41_R_f(R_f_top[1009]),
    .Tile_X33Y41_R_t(R_t_top[1010]),
    .Tile_X33Y41_R_f(R_f_top[1010]),
    .Tile_X36Y41_R_t(R_t_top[1011]),
    .Tile_X36Y41_R_f(R_f_top[1011]),
    .Tile_X39Y41_R_t(R_t_top[1012]),
    .Tile_X39Y41_R_f(R_f_top[1012]),
    .Tile_X42Y41_R_t(R_t_top[1013]),
    .Tile_X42Y41_R_f(R_f_top[1013]),
    .Tile_X45Y41_R_t(R_t_top[1014]),
    .Tile_X45Y41_R_f(R_f_top[1014]),
    .Tile_X48Y41_R_t(R_t_top[1015]),
    .Tile_X48Y41_R_f(R_f_top[1015]),
    .Tile_X51Y41_R_t(R_t_top[1016]),
    .Tile_X51Y41_R_f(R_f_top[1016]),
    .Tile_X54Y41_R_t(R_t_top[1017]),
    .Tile_X54Y41_R_f(R_f_top[1017]),
    .Tile_X57Y41_R_t(R_t_top[1018]),
    .Tile_X57Y41_R_f(R_f_top[1018]),
    .Tile_X60Y41_R_t(R_t_top[1019]),
    .Tile_X60Y41_R_f(R_f_top[1019]),
    .Tile_X63Y41_R_t(R_t_top[1020]),
    .Tile_X63Y41_R_f(R_f_top[1020]),
    .Tile_X66Y41_R_t(R_t_top[1021]),
    .Tile_X66Y41_R_f(R_f_top[1021]),
    .Tile_X69Y41_R_t(R_t_top[1022]),
    .Tile_X69Y41_R_f(R_f_top[1022]),
    .Tile_X72Y41_R_t(R_t_top[1023]),
    .Tile_X72Y41_R_f(R_f_top[1023]),
    .Tile_X75Y41_R_t(R_t_top[1024]),
    .Tile_X75Y41_R_f(R_f_top[1024]),
    .Tile_X3Y42_R_t(R_t_top[1025]),
    .Tile_X3Y42_R_f(R_f_top[1025]),
    .Tile_X6Y42_R_t(R_t_top[1026]),
    .Tile_X6Y42_R_f(R_f_top[1026]),
    .Tile_X9Y42_R_t(R_t_top[1027]),
    .Tile_X9Y42_R_f(R_f_top[1027]),
    .Tile_X12Y42_R_t(R_t_top[1028]),
    .Tile_X12Y42_R_f(R_f_top[1028]),
    .Tile_X15Y42_R_t(R_t_top[1029]),
    .Tile_X15Y42_R_f(R_f_top[1029]),
    .Tile_X18Y42_R_t(R_t_top[1030]),
    .Tile_X18Y42_R_f(R_f_top[1030]),
    .Tile_X21Y42_R_t(R_t_top[1031]),
    .Tile_X21Y42_R_f(R_f_top[1031]),
    .Tile_X24Y42_R_t(R_t_top[1032]),
    .Tile_X24Y42_R_f(R_f_top[1032]),
    .Tile_X27Y42_R_t(R_t_top[1033]),
    .Tile_X27Y42_R_f(R_f_top[1033]),
    .Tile_X30Y42_R_t(R_t_top[1034]),
    .Tile_X30Y42_R_f(R_f_top[1034]),
    .Tile_X33Y42_R_t(R_t_top[1035]),
    .Tile_X33Y42_R_f(R_f_top[1035]),
    .Tile_X36Y42_R_t(R_t_top[1036]),
    .Tile_X36Y42_R_f(R_f_top[1036]),
    .Tile_X39Y42_R_t(R_t_top[1037]),
    .Tile_X39Y42_R_f(R_f_top[1037]),
    .Tile_X42Y42_R_t(R_t_top[1038]),
    .Tile_X42Y42_R_f(R_f_top[1038]),
    .Tile_X45Y42_R_t(R_t_top[1039]),
    .Tile_X45Y42_R_f(R_f_top[1039]),
    .Tile_X48Y42_R_t(R_t_top[1040]),
    .Tile_X48Y42_R_f(R_f_top[1040]),
    .Tile_X51Y42_R_t(R_t_top[1041]),
    .Tile_X51Y42_R_f(R_f_top[1041]),
    .Tile_X54Y42_R_t(R_t_top[1042]),
    .Tile_X54Y42_R_f(R_f_top[1042]),
    .Tile_X57Y42_R_t(R_t_top[1043]),
    .Tile_X57Y42_R_f(R_f_top[1043]),
    .Tile_X60Y42_R_t(R_t_top[1044]),
    .Tile_X60Y42_R_f(R_f_top[1044]),
    .Tile_X63Y42_R_t(R_t_top[1045]),
    .Tile_X63Y42_R_f(R_f_top[1045]),
    .Tile_X66Y42_R_t(R_t_top[1046]),
    .Tile_X66Y42_R_f(R_f_top[1046]),
    .Tile_X69Y42_R_t(R_t_top[1047]),
    .Tile_X69Y42_R_f(R_f_top[1047]),
    .Tile_X72Y42_R_t(R_t_top[1048]),
    .Tile_X72Y42_R_f(R_f_top[1048]),
    .Tile_X75Y42_R_t(R_t_top[1049]),
    .Tile_X75Y42_R_f(R_f_top[1049]),
    .Tile_X3Y43_R_t(R_t_top[1050]),
    .Tile_X3Y43_R_f(R_f_top[1050]),
    .Tile_X6Y43_R_t(R_t_top[1051]),
    .Tile_X6Y43_R_f(R_f_top[1051]),
    .Tile_X9Y43_R_t(R_t_top[1052]),
    .Tile_X9Y43_R_f(R_f_top[1052]),
    .Tile_X12Y43_R_t(R_t_top[1053]),
    .Tile_X12Y43_R_f(R_f_top[1053]),
    .Tile_X15Y43_R_t(R_t_top[1054]),
    .Tile_X15Y43_R_f(R_f_top[1054]),
    .Tile_X18Y43_R_t(R_t_top[1055]),
    .Tile_X18Y43_R_f(R_f_top[1055]),
    .Tile_X21Y43_R_t(R_t_top[1056]),
    .Tile_X21Y43_R_f(R_f_top[1056]),
    .Tile_X24Y43_R_t(R_t_top[1057]),
    .Tile_X24Y43_R_f(R_f_top[1057]),
    .Tile_X27Y43_R_t(R_t_top[1058]),
    .Tile_X27Y43_R_f(R_f_top[1058]),
    .Tile_X30Y43_R_t(R_t_top[1059]),
    .Tile_X30Y43_R_f(R_f_top[1059]),
    .Tile_X33Y43_R_t(R_t_top[1060]),
    .Tile_X33Y43_R_f(R_f_top[1060]),
    .Tile_X36Y43_R_t(R_t_top[1061]),
    .Tile_X36Y43_R_f(R_f_top[1061]),
    .Tile_X39Y43_R_t(R_t_top[1062]),
    .Tile_X39Y43_R_f(R_f_top[1062]),
    .Tile_X42Y43_R_t(R_t_top[1063]),
    .Tile_X42Y43_R_f(R_f_top[1063]),
    .Tile_X45Y43_R_t(R_t_top[1064]),
    .Tile_X45Y43_R_f(R_f_top[1064]),
    .Tile_X48Y43_R_t(R_t_top[1065]),
    .Tile_X48Y43_R_f(R_f_top[1065]),
    .Tile_X51Y43_R_t(R_t_top[1066]),
    .Tile_X51Y43_R_f(R_f_top[1066]),
    .Tile_X54Y43_R_t(R_t_top[1067]),
    .Tile_X54Y43_R_f(R_f_top[1067]),
    .Tile_X57Y43_R_t(R_t_top[1068]),
    .Tile_X57Y43_R_f(R_f_top[1068]),
    .Tile_X60Y43_R_t(R_t_top[1069]),
    .Tile_X60Y43_R_f(R_f_top[1069]),
    .Tile_X63Y43_R_t(R_t_top[1070]),
    .Tile_X63Y43_R_f(R_f_top[1070]),
    .Tile_X66Y43_R_t(R_t_top[1071]),
    .Tile_X66Y43_R_f(R_f_top[1071]),
    .Tile_X69Y43_R_t(R_t_top[1072]),
    .Tile_X69Y43_R_f(R_f_top[1072]),
    .Tile_X72Y43_R_t(R_t_top[1073]),
    .Tile_X72Y43_R_f(R_f_top[1073]),
    .Tile_X75Y43_R_t(R_t_top[1074]),
    .Tile_X75Y43_R_f(R_f_top[1074]),
    .Tile_X3Y44_R_t(R_t_top[1075]),
    .Tile_X3Y44_R_f(R_f_top[1075]),
    .Tile_X6Y44_R_t(R_t_top[1076]),
    .Tile_X6Y44_R_f(R_f_top[1076]),
    .Tile_X9Y44_R_t(R_t_top[1077]),
    .Tile_X9Y44_R_f(R_f_top[1077]),
    .Tile_X12Y44_R_t(R_t_top[1078]),
    .Tile_X12Y44_R_f(R_f_top[1078]),
    .Tile_X15Y44_R_t(R_t_top[1079]),
    .Tile_X15Y44_R_f(R_f_top[1079]),
    .Tile_X18Y44_R_t(R_t_top[1080]),
    .Tile_X18Y44_R_f(R_f_top[1080]),
    .Tile_X21Y44_R_t(R_t_top[1081]),
    .Tile_X21Y44_R_f(R_f_top[1081]),
    .Tile_X24Y44_R_t(R_t_top[1082]),
    .Tile_X24Y44_R_f(R_f_top[1082]),
    .Tile_X27Y44_R_t(R_t_top[1083]),
    .Tile_X27Y44_R_f(R_f_top[1083]),
    .Tile_X30Y44_R_t(R_t_top[1084]),
    .Tile_X30Y44_R_f(R_f_top[1084]),
    .Tile_X33Y44_R_t(R_t_top[1085]),
    .Tile_X33Y44_R_f(R_f_top[1085]),
    .Tile_X36Y44_R_t(R_t_top[1086]),
    .Tile_X36Y44_R_f(R_f_top[1086]),
    .Tile_X39Y44_R_t(R_t_top[1087]),
    .Tile_X39Y44_R_f(R_f_top[1087]),
    .Tile_X42Y44_R_t(R_t_top[1088]),
    .Tile_X42Y44_R_f(R_f_top[1088]),
    .Tile_X45Y44_R_t(R_t_top[1089]),
    .Tile_X45Y44_R_f(R_f_top[1089]),
    .Tile_X48Y44_R_t(R_t_top[1090]),
    .Tile_X48Y44_R_f(R_f_top[1090]),
    .Tile_X51Y44_R_t(R_t_top[1091]),
    .Tile_X51Y44_R_f(R_f_top[1091]),
    .Tile_X54Y44_R_t(R_t_top[1092]),
    .Tile_X54Y44_R_f(R_f_top[1092]),
    .Tile_X57Y44_R_t(R_t_top[1093]),
    .Tile_X57Y44_R_f(R_f_top[1093]),
    .Tile_X60Y44_R_t(R_t_top[1094]),
    .Tile_X60Y44_R_f(R_f_top[1094]),
    .Tile_X63Y44_R_t(R_t_top[1095]),
    .Tile_X63Y44_R_f(R_f_top[1095]),
    .Tile_X66Y44_R_t(R_t_top[1096]),
    .Tile_X66Y44_R_f(R_f_top[1096]),
    .Tile_X69Y44_R_t(R_t_top[1097]),
    .Tile_X69Y44_R_f(R_f_top[1097]),
    .Tile_X72Y44_R_t(R_t_top[1098]),
    .Tile_X72Y44_R_f(R_f_top[1098]),
    .Tile_X75Y44_R_t(R_t_top[1099]),
    .Tile_X75Y44_R_f(R_f_top[1099]),
    .Tile_X3Y45_R_t(R_t_top[1100]),
    .Tile_X3Y45_R_f(R_f_top[1100]),
    .Tile_X6Y45_R_t(R_t_top[1101]),
    .Tile_X6Y45_R_f(R_f_top[1101]),
    .Tile_X9Y45_R_t(R_t_top[1102]),
    .Tile_X9Y45_R_f(R_f_top[1102]),
    .Tile_X12Y45_R_t(R_t_top[1103]),
    .Tile_X12Y45_R_f(R_f_top[1103]),
    .Tile_X15Y45_R_t(R_t_top[1104]),
    .Tile_X15Y45_R_f(R_f_top[1104]),
    .Tile_X18Y45_R_t(R_t_top[1105]),
    .Tile_X18Y45_R_f(R_f_top[1105]),
    .Tile_X21Y45_R_t(R_t_top[1106]),
    .Tile_X21Y45_R_f(R_f_top[1106]),
    .Tile_X24Y45_R_t(R_t_top[1107]),
    .Tile_X24Y45_R_f(R_f_top[1107]),
    .Tile_X27Y45_R_t(R_t_top[1108]),
    .Tile_X27Y45_R_f(R_f_top[1108]),
    .Tile_X30Y45_R_t(R_t_top[1109]),
    .Tile_X30Y45_R_f(R_f_top[1109]),
    .Tile_X33Y45_R_t(R_t_top[1110]),
    .Tile_X33Y45_R_f(R_f_top[1110]),
    .Tile_X36Y45_R_t(R_t_top[1111]),
    .Tile_X36Y45_R_f(R_f_top[1111]),
    .Tile_X39Y45_R_t(R_t_top[1112]),
    .Tile_X39Y45_R_f(R_f_top[1112]),
    .Tile_X42Y45_R_t(R_t_top[1113]),
    .Tile_X42Y45_R_f(R_f_top[1113]),
    .Tile_X45Y45_R_t(R_t_top[1114]),
    .Tile_X45Y45_R_f(R_f_top[1114]),
    .Tile_X48Y45_R_t(R_t_top[1115]),
    .Tile_X48Y45_R_f(R_f_top[1115]),
    .Tile_X51Y45_R_t(R_t_top[1116]),
    .Tile_X51Y45_R_f(R_f_top[1116]),
    .Tile_X54Y45_R_t(R_t_top[1117]),
    .Tile_X54Y45_R_f(R_f_top[1117]),
    .Tile_X57Y45_R_t(R_t_top[1118]),
    .Tile_X57Y45_R_f(R_f_top[1118]),
    .Tile_X60Y45_R_t(R_t_top[1119]),
    .Tile_X60Y45_R_f(R_f_top[1119]),
    .Tile_X63Y45_R_t(R_t_top[1120]),
    .Tile_X63Y45_R_f(R_f_top[1120]),
    .Tile_X66Y45_R_t(R_t_top[1121]),
    .Tile_X66Y45_R_f(R_f_top[1121]),
    .Tile_X69Y45_R_t(R_t_top[1122]),
    .Tile_X69Y45_R_f(R_f_top[1122]),
    .Tile_X72Y45_R_t(R_t_top[1123]),
    .Tile_X72Y45_R_f(R_f_top[1123]),
    .Tile_X75Y45_R_t(R_t_top[1124]),
    .Tile_X75Y45_R_f(R_f_top[1124]),
    .Tile_X3Y46_R_t(R_t_top[1125]),
    .Tile_X3Y46_R_f(R_f_top[1125]),
    .Tile_X6Y46_R_t(R_t_top[1126]),
    .Tile_X6Y46_R_f(R_f_top[1126]),
    .Tile_X9Y46_R_t(R_t_top[1127]),
    .Tile_X9Y46_R_f(R_f_top[1127]),
    .Tile_X12Y46_R_t(R_t_top[1128]),
    .Tile_X12Y46_R_f(R_f_top[1128]),
    .Tile_X15Y46_R_t(R_t_top[1129]),
    .Tile_X15Y46_R_f(R_f_top[1129]),
    .Tile_X18Y46_R_t(R_t_top[1130]),
    .Tile_X18Y46_R_f(R_f_top[1130]),
    .Tile_X21Y46_R_t(R_t_top[1131]),
    .Tile_X21Y46_R_f(R_f_top[1131]),
    .Tile_X24Y46_R_t(R_t_top[1132]),
    .Tile_X24Y46_R_f(R_f_top[1132]),
    .Tile_X27Y46_R_t(R_t_top[1133]),
    .Tile_X27Y46_R_f(R_f_top[1133]),
    .Tile_X30Y46_R_t(R_t_top[1134]),
    .Tile_X30Y46_R_f(R_f_top[1134]),
    .Tile_X33Y46_R_t(R_t_top[1135]),
    .Tile_X33Y46_R_f(R_f_top[1135]),
    .Tile_X36Y46_R_t(R_t_top[1136]),
    .Tile_X36Y46_R_f(R_f_top[1136]),
    .Tile_X39Y46_R_t(R_t_top[1137]),
    .Tile_X39Y46_R_f(R_f_top[1137]),
    .Tile_X42Y46_R_t(R_t_top[1138]),
    .Tile_X42Y46_R_f(R_f_top[1138]),
    .Tile_X45Y46_R_t(R_t_top[1139]),
    .Tile_X45Y46_R_f(R_f_top[1139]),
    .Tile_X48Y46_R_t(R_t_top[1140]),
    .Tile_X48Y46_R_f(R_f_top[1140]),
    .Tile_X51Y46_R_t(R_t_top[1141]),
    .Tile_X51Y46_R_f(R_f_top[1141]),
    .Tile_X54Y46_R_t(R_t_top[1142]),
    .Tile_X54Y46_R_f(R_f_top[1142]),
    .Tile_X57Y46_R_t(R_t_top[1143]),
    .Tile_X57Y46_R_f(R_f_top[1143]),
    .Tile_X60Y46_R_t(R_t_top[1144]),
    .Tile_X60Y46_R_f(R_f_top[1144]),
    .Tile_X63Y46_R_t(R_t_top[1145]),
    .Tile_X63Y46_R_f(R_f_top[1145]),
    .Tile_X66Y46_R_t(R_t_top[1146]),
    .Tile_X66Y46_R_f(R_f_top[1146]),
    .Tile_X69Y46_R_t(R_t_top[1147]),
    .Tile_X69Y46_R_f(R_f_top[1147]),
    .Tile_X72Y46_R_t(R_t_top[1148]),
    .Tile_X72Y46_R_f(R_f_top[1148]),
    .Tile_X75Y46_R_t(R_t_top[1149]),
    .Tile_X75Y46_R_f(R_f_top[1149]),
    .Tile_X3Y47_R_t(R_t_top[1150]),
    .Tile_X3Y47_R_f(R_f_top[1150]),
    .Tile_X6Y47_R_t(R_t_top[1151]),
    .Tile_X6Y47_R_f(R_f_top[1151]),
    .Tile_X9Y47_R_t(R_t_top[1152]),
    .Tile_X9Y47_R_f(R_f_top[1152]),
    .Tile_X12Y47_R_t(R_t_top[1153]),
    .Tile_X12Y47_R_f(R_f_top[1153]),
    .Tile_X15Y47_R_t(R_t_top[1154]),
    .Tile_X15Y47_R_f(R_f_top[1154]),
    .Tile_X18Y47_R_t(R_t_top[1155]),
    .Tile_X18Y47_R_f(R_f_top[1155]),
    .Tile_X21Y47_R_t(R_t_top[1156]),
    .Tile_X21Y47_R_f(R_f_top[1156]),
    .Tile_X24Y47_R_t(R_t_top[1157]),
    .Tile_X24Y47_R_f(R_f_top[1157]),
    .Tile_X27Y47_R_t(R_t_top[1158]),
    .Tile_X27Y47_R_f(R_f_top[1158]),
    .Tile_X30Y47_R_t(R_t_top[1159]),
    .Tile_X30Y47_R_f(R_f_top[1159]),
    .Tile_X33Y47_R_t(R_t_top[1160]),
    .Tile_X33Y47_R_f(R_f_top[1160]),
    .Tile_X36Y47_R_t(R_t_top[1161]),
    .Tile_X36Y47_R_f(R_f_top[1161]),
    .Tile_X39Y47_R_t(R_t_top[1162]),
    .Tile_X39Y47_R_f(R_f_top[1162]),
    .Tile_X42Y47_R_t(R_t_top[1163]),
    .Tile_X42Y47_R_f(R_f_top[1163]),
    .Tile_X45Y47_R_t(R_t_top[1164]),
    .Tile_X45Y47_R_f(R_f_top[1164]),
    .Tile_X48Y47_R_t(R_t_top[1165]),
    .Tile_X48Y47_R_f(R_f_top[1165]),
    .Tile_X51Y47_R_t(R_t_top[1166]),
    .Tile_X51Y47_R_f(R_f_top[1166]),
    .Tile_X54Y47_R_t(R_t_top[1167]),
    .Tile_X54Y47_R_f(R_f_top[1167]),
    .Tile_X57Y47_R_t(R_t_top[1168]),
    .Tile_X57Y47_R_f(R_f_top[1168]),
    .Tile_X60Y47_R_t(R_t_top[1169]),
    .Tile_X60Y47_R_f(R_f_top[1169]),
    .Tile_X63Y47_R_t(R_t_top[1170]),
    .Tile_X63Y47_R_f(R_f_top[1170]),
    .Tile_X66Y47_R_t(R_t_top[1171]),
    .Tile_X66Y47_R_f(R_f_top[1171]),
    .Tile_X69Y47_R_t(R_t_top[1172]),
    .Tile_X69Y47_R_f(R_f_top[1172]),
    .Tile_X72Y47_R_t(R_t_top[1173]),
    .Tile_X72Y47_R_f(R_f_top[1173]),
    .Tile_X75Y47_R_t(R_t_top[1174]),
    .Tile_X75Y47_R_f(R_f_top[1174]),
    .Tile_X3Y48_R_t(R_t_top[1175]),
    .Tile_X3Y48_R_f(R_f_top[1175]),
    .Tile_X6Y48_R_t(R_t_top[1176]),
    .Tile_X6Y48_R_f(R_f_top[1176]),
    .Tile_X9Y48_R_t(R_t_top[1177]),
    .Tile_X9Y48_R_f(R_f_top[1177]),
    .Tile_X12Y48_R_t(R_t_top[1178]),
    .Tile_X12Y48_R_f(R_f_top[1178]),
    .Tile_X15Y48_R_t(R_t_top[1179]),
    .Tile_X15Y48_R_f(R_f_top[1179]),
    .Tile_X18Y48_R_t(R_t_top[1180]),
    .Tile_X18Y48_R_f(R_f_top[1180]),
    .Tile_X21Y48_R_t(R_t_top[1181]),
    .Tile_X21Y48_R_f(R_f_top[1181]),
    .Tile_X24Y48_R_t(R_t_top[1182]),
    .Tile_X24Y48_R_f(R_f_top[1182]),
    .Tile_X27Y48_R_t(R_t_top[1183]),
    .Tile_X27Y48_R_f(R_f_top[1183]),
    .Tile_X30Y48_R_t(R_t_top[1184]),
    .Tile_X30Y48_R_f(R_f_top[1184]),
    .Tile_X33Y48_R_t(R_t_top[1185]),
    .Tile_X33Y48_R_f(R_f_top[1185]),
    .Tile_X36Y48_R_t(R_t_top[1186]),
    .Tile_X36Y48_R_f(R_f_top[1186]),
    .Tile_X39Y48_R_t(R_t_top[1187]),
    .Tile_X39Y48_R_f(R_f_top[1187]),
    .Tile_X42Y48_R_t(R_t_top[1188]),
    .Tile_X42Y48_R_f(R_f_top[1188]),
    .Tile_X45Y48_R_t(R_t_top[1189]),
    .Tile_X45Y48_R_f(R_f_top[1189]),
    .Tile_X48Y48_R_t(R_t_top[1190]),
    .Tile_X48Y48_R_f(R_f_top[1190]),
    .Tile_X51Y48_R_t(R_t_top[1191]),
    .Tile_X51Y48_R_f(R_f_top[1191]),
    .Tile_X54Y48_R_t(R_t_top[1192]),
    .Tile_X54Y48_R_f(R_f_top[1192]),
    .Tile_X57Y48_R_t(R_t_top[1193]),
    .Tile_X57Y48_R_f(R_f_top[1193]),
    .Tile_X60Y48_R_t(R_t_top[1194]),
    .Tile_X60Y48_R_f(R_f_top[1194]),
    .Tile_X63Y48_R_t(R_t_top[1195]),
    .Tile_X63Y48_R_f(R_f_top[1195]),
    .Tile_X66Y48_R_t(R_t_top[1196]),
    .Tile_X66Y48_R_f(R_f_top[1196]),
    .Tile_X69Y48_R_t(R_t_top[1197]),
    .Tile_X69Y48_R_f(R_f_top[1197]),
    .Tile_X72Y48_R_t(R_t_top[1198]),
    .Tile_X72Y48_R_f(R_f_top[1198]),
    .Tile_X75Y48_R_t(R_t_top[1199]),
    .Tile_X75Y48_R_f(R_f_top[1199]),
    .Tile_X3Y49_R_t(R_t_top[1200]),
    .Tile_X3Y49_R_f(R_f_top[1200]),
    .Tile_X6Y49_R_t(R_t_top[1201]),
    .Tile_X6Y49_R_f(R_f_top[1201]),
    .Tile_X9Y49_R_t(R_t_top[1202]),
    .Tile_X9Y49_R_f(R_f_top[1202]),
    .Tile_X12Y49_R_t(R_t_top[1203]),
    .Tile_X12Y49_R_f(R_f_top[1203]),
    .Tile_X15Y49_R_t(R_t_top[1204]),
    .Tile_X15Y49_R_f(R_f_top[1204]),
    .Tile_X18Y49_R_t(R_t_top[1205]),
    .Tile_X18Y49_R_f(R_f_top[1205]),
    .Tile_X21Y49_R_t(R_t_top[1206]),
    .Tile_X21Y49_R_f(R_f_top[1206]),
    .Tile_X24Y49_R_t(R_t_top[1207]),
    .Tile_X24Y49_R_f(R_f_top[1207]),
    .Tile_X27Y49_R_t(R_t_top[1208]),
    .Tile_X27Y49_R_f(R_f_top[1208]),
    .Tile_X30Y49_R_t(R_t_top[1209]),
    .Tile_X30Y49_R_f(R_f_top[1209]),
    .Tile_X33Y49_R_t(R_t_top[1210]),
    .Tile_X33Y49_R_f(R_f_top[1210]),
    .Tile_X36Y49_R_t(R_t_top[1211]),
    .Tile_X36Y49_R_f(R_f_top[1211]),
    .Tile_X39Y49_R_t(R_t_top[1212]),
    .Tile_X39Y49_R_f(R_f_top[1212]),
    .Tile_X42Y49_R_t(R_t_top[1213]),
    .Tile_X42Y49_R_f(R_f_top[1213]),
    .Tile_X45Y49_R_t(R_t_top[1214]),
    .Tile_X45Y49_R_f(R_f_top[1214]),
    .Tile_X48Y49_R_t(R_t_top[1215]),
    .Tile_X48Y49_R_f(R_f_top[1215]),
    .Tile_X51Y49_R_t(R_t_top[1216]),
    .Tile_X51Y49_R_f(R_f_top[1216]),
    .Tile_X54Y49_R_t(R_t_top[1217]),
    .Tile_X54Y49_R_f(R_f_top[1217]),
    .Tile_X57Y49_R_t(R_t_top[1218]),
    .Tile_X57Y49_R_f(R_f_top[1218]),
    .Tile_X60Y49_R_t(R_t_top[1219]),
    .Tile_X60Y49_R_f(R_f_top[1219]),
    .Tile_X63Y49_R_t(R_t_top[1220]),
    .Tile_X63Y49_R_f(R_f_top[1220]),
    .Tile_X66Y49_R_t(R_t_top[1221]),
    .Tile_X66Y49_R_f(R_f_top[1221]),
    .Tile_X69Y49_R_t(R_t_top[1222]),
    .Tile_X69Y49_R_f(R_f_top[1222]),
    .Tile_X72Y49_R_t(R_t_top[1223]),
    .Tile_X72Y49_R_f(R_f_top[1223]),
    .Tile_X75Y49_R_t(R_t_top[1224]),
    .Tile_X75Y49_R_f(R_f_top[1224]),
    .Tile_X3Y50_R_t(R_t_top[1225]),
    .Tile_X3Y50_R_f(R_f_top[1225]),
    .Tile_X6Y50_R_t(R_t_top[1226]),
    .Tile_X6Y50_R_f(R_f_top[1226]),
    .Tile_X9Y50_R_t(R_t_top[1227]),
    .Tile_X9Y50_R_f(R_f_top[1227]),
    .Tile_X12Y50_R_t(R_t_top[1228]),
    .Tile_X12Y50_R_f(R_f_top[1228]),
    .Tile_X15Y50_R_t(R_t_top[1229]),
    .Tile_X15Y50_R_f(R_f_top[1229]),
    .Tile_X18Y50_R_t(R_t_top[1230]),
    .Tile_X18Y50_R_f(R_f_top[1230]),
    .Tile_X21Y50_R_t(R_t_top[1231]),
    .Tile_X21Y50_R_f(R_f_top[1231]),
    .Tile_X24Y50_R_t(R_t_top[1232]),
    .Tile_X24Y50_R_f(R_f_top[1232]),
    .Tile_X27Y50_R_t(R_t_top[1233]),
    .Tile_X27Y50_R_f(R_f_top[1233]),
    .Tile_X30Y50_R_t(R_t_top[1234]),
    .Tile_X30Y50_R_f(R_f_top[1234]),
    .Tile_X33Y50_R_t(R_t_top[1235]),
    .Tile_X33Y50_R_f(R_f_top[1235]),
    .Tile_X36Y50_R_t(R_t_top[1236]),
    .Tile_X36Y50_R_f(R_f_top[1236]),
    .Tile_X39Y50_R_t(R_t_top[1237]),
    .Tile_X39Y50_R_f(R_f_top[1237]),
    .Tile_X42Y50_R_t(R_t_top[1238]),
    .Tile_X42Y50_R_f(R_f_top[1238]),
    .Tile_X45Y50_R_t(R_t_top[1239]),
    .Tile_X45Y50_R_f(R_f_top[1239]),
    .Tile_X48Y50_R_t(R_t_top[1240]),
    .Tile_X48Y50_R_f(R_f_top[1240]),
    .Tile_X51Y50_R_t(R_t_top[1241]),
    .Tile_X51Y50_R_f(R_f_top[1241]),
    .Tile_X54Y50_R_t(R_t_top[1242]),
    .Tile_X54Y50_R_f(R_f_top[1242]),
    .Tile_X57Y50_R_t(R_t_top[1243]),
    .Tile_X57Y50_R_f(R_f_top[1243]),
    .Tile_X60Y50_R_t(R_t_top[1244]),
    .Tile_X60Y50_R_f(R_f_top[1244]),
    .Tile_X63Y50_R_t(R_t_top[1245]),
    .Tile_X63Y50_R_f(R_f_top[1245]),
    .Tile_X66Y50_R_t(R_t_top[1246]),
    .Tile_X66Y50_R_f(R_f_top[1246]),
    .Tile_X69Y50_R_t(R_t_top[1247]),
    .Tile_X69Y50_R_f(R_f_top[1247]),
    .Tile_X72Y50_R_t(R_t_top[1248]),
    .Tile_X72Y50_R_f(R_f_top[1248]),
    .Tile_X75Y50_R_t(R_t_top[1249]),
    .Tile_X75Y50_R_f(R_f_top[1249]),
    .Tile_X3Y51_R_t(R_t_top[1250]),
    .Tile_X3Y51_R_f(R_f_top[1250]),
    .Tile_X6Y51_R_t(R_t_top[1251]),
    .Tile_X6Y51_R_f(R_f_top[1251]),
    .Tile_X9Y51_R_t(R_t_top[1252]),
    .Tile_X9Y51_R_f(R_f_top[1252]),
    .Tile_X12Y51_R_t(R_t_top[1253]),
    .Tile_X12Y51_R_f(R_f_top[1253]),
    .Tile_X15Y51_R_t(R_t_top[1254]),
    .Tile_X15Y51_R_f(R_f_top[1254]),
    .Tile_X18Y51_R_t(R_t_top[1255]),
    .Tile_X18Y51_R_f(R_f_top[1255]),
    .Tile_X21Y51_R_t(R_t_top[1256]),
    .Tile_X21Y51_R_f(R_f_top[1256]),
    .Tile_X24Y51_R_t(R_t_top[1257]),
    .Tile_X24Y51_R_f(R_f_top[1257]),
    .Tile_X27Y51_R_t(R_t_top[1258]),
    .Tile_X27Y51_R_f(R_f_top[1258]),
    .Tile_X30Y51_R_t(R_t_top[1259]),
    .Tile_X30Y51_R_f(R_f_top[1259]),
    .Tile_X33Y51_R_t(R_t_top[1260]),
    .Tile_X33Y51_R_f(R_f_top[1260]),
    .Tile_X36Y51_R_t(R_t_top[1261]),
    .Tile_X36Y51_R_f(R_f_top[1261]),
    .Tile_X39Y51_R_t(R_t_top[1262]),
    .Tile_X39Y51_R_f(R_f_top[1262]),
    .Tile_X42Y51_R_t(R_t_top[1263]),
    .Tile_X42Y51_R_f(R_f_top[1263]),
    .Tile_X45Y51_R_t(R_t_top[1264]),
    .Tile_X45Y51_R_f(R_f_top[1264]),
    .Tile_X48Y51_R_t(R_t_top[1265]),
    .Tile_X48Y51_R_f(R_f_top[1265]),
    .Tile_X51Y51_R_t(R_t_top[1266]),
    .Tile_X51Y51_R_f(R_f_top[1266]),
    .Tile_X54Y51_R_t(R_t_top[1267]),
    .Tile_X54Y51_R_f(R_f_top[1267]),
    .Tile_X57Y51_R_t(R_t_top[1268]),
    .Tile_X57Y51_R_f(R_f_top[1268]),
    .Tile_X60Y51_R_t(R_t_top[1269]),
    .Tile_X60Y51_R_f(R_f_top[1269]),
    .Tile_X63Y51_R_t(R_t_top[1270]),
    .Tile_X63Y51_R_f(R_f_top[1270]),
    .Tile_X66Y51_R_t(R_t_top[1271]),
    .Tile_X66Y51_R_f(R_f_top[1271]),
    .Tile_X69Y51_R_t(R_t_top[1272]),
    .Tile_X69Y51_R_f(R_f_top[1272]),
    .Tile_X72Y51_R_t(R_t_top[1273]),
    .Tile_X72Y51_R_f(R_f_top[1273]),
    .Tile_X75Y51_R_t(R_t_top[1274]),
    .Tile_X75Y51_R_f(R_f_top[1274]),
    .Tile_X3Y52_R_t(R_t_top[1275]),
    .Tile_X3Y52_R_f(R_f_top[1275]),
    .Tile_X6Y52_R_t(R_t_top[1276]),
    .Tile_X6Y52_R_f(R_f_top[1276]),
    .Tile_X9Y52_R_t(R_t_top[1277]),
    .Tile_X9Y52_R_f(R_f_top[1277]),
    .Tile_X12Y52_R_t(R_t_top[1278]),
    .Tile_X12Y52_R_f(R_f_top[1278]),
    .Tile_X15Y52_R_t(R_t_top[1279]),
    .Tile_X15Y52_R_f(R_f_top[1279]),
    .Tile_X18Y52_R_t(R_t_top[1280]),
    .Tile_X18Y52_R_f(R_f_top[1280]),
    .Tile_X21Y52_R_t(R_t_top[1281]),
    .Tile_X21Y52_R_f(R_f_top[1281]),
    .Tile_X24Y52_R_t(R_t_top[1282]),
    .Tile_X24Y52_R_f(R_f_top[1282]),
    .Tile_X27Y52_R_t(R_t_top[1283]),
    .Tile_X27Y52_R_f(R_f_top[1283]),
    .Tile_X30Y52_R_t(R_t_top[1284]),
    .Tile_X30Y52_R_f(R_f_top[1284]),
    .Tile_X33Y52_R_t(R_t_top[1285]),
    .Tile_X33Y52_R_f(R_f_top[1285]),
    .Tile_X36Y52_R_t(R_t_top[1286]),
    .Tile_X36Y52_R_f(R_f_top[1286]),
    .Tile_X39Y52_R_t(R_t_top[1287]),
    .Tile_X39Y52_R_f(R_f_top[1287]),
    .Tile_X42Y52_R_t(R_t_top[1288]),
    .Tile_X42Y52_R_f(R_f_top[1288]),
    .Tile_X45Y52_R_t(R_t_top[1289]),
    .Tile_X45Y52_R_f(R_f_top[1289]),
    .Tile_X48Y52_R_t(R_t_top[1290]),
    .Tile_X48Y52_R_f(R_f_top[1290]),
    .Tile_X51Y52_R_t(R_t_top[1291]),
    .Tile_X51Y52_R_f(R_f_top[1291]),
    .Tile_X54Y52_R_t(R_t_top[1292]),
    .Tile_X54Y52_R_f(R_f_top[1292]),
    .Tile_X57Y52_R_t(R_t_top[1293]),
    .Tile_X57Y52_R_f(R_f_top[1293]),
    .Tile_X60Y52_R_t(R_t_top[1294]),
    .Tile_X60Y52_R_f(R_f_top[1294]),
    .Tile_X63Y52_R_t(R_t_top[1295]),
    .Tile_X63Y52_R_f(R_f_top[1295]),
    .Tile_X66Y52_R_t(R_t_top[1296]),
    .Tile_X66Y52_R_f(R_f_top[1296]),
    .Tile_X69Y52_R_t(R_t_top[1297]),
    .Tile_X69Y52_R_f(R_f_top[1297]),
    .Tile_X72Y52_R_t(R_t_top[1298]),
    .Tile_X72Y52_R_f(R_f_top[1298]),
    .Tile_X75Y52_R_t(R_t_top[1299]),
    .Tile_X75Y52_R_f(R_f_top[1299]),
    .Tile_X3Y53_R_t(R_t_top[1300]),
    .Tile_X3Y53_R_f(R_f_top[1300]),
    .Tile_X6Y53_R_t(R_t_top[1301]),
    .Tile_X6Y53_R_f(R_f_top[1301]),
    .Tile_X9Y53_R_t(R_t_top[1302]),
    .Tile_X9Y53_R_f(R_f_top[1302]),
    .Tile_X12Y53_R_t(R_t_top[1303]),
    .Tile_X12Y53_R_f(R_f_top[1303]),
    .Tile_X15Y53_R_t(R_t_top[1304]),
    .Tile_X15Y53_R_f(R_f_top[1304]),
    .Tile_X18Y53_R_t(R_t_top[1305]),
    .Tile_X18Y53_R_f(R_f_top[1305]),
    .Tile_X21Y53_R_t(R_t_top[1306]),
    .Tile_X21Y53_R_f(R_f_top[1306]),
    .Tile_X24Y53_R_t(R_t_top[1307]),
    .Tile_X24Y53_R_f(R_f_top[1307]),
    .Tile_X27Y53_R_t(R_t_top[1308]),
    .Tile_X27Y53_R_f(R_f_top[1308]),
    .Tile_X30Y53_R_t(R_t_top[1309]),
    .Tile_X30Y53_R_f(R_f_top[1309]),
    .Tile_X33Y53_R_t(R_t_top[1310]),
    .Tile_X33Y53_R_f(R_f_top[1310]),
    .Tile_X36Y53_R_t(R_t_top[1311]),
    .Tile_X36Y53_R_f(R_f_top[1311]),
    .Tile_X39Y53_R_t(R_t_top[1312]),
    .Tile_X39Y53_R_f(R_f_top[1312]),
    .Tile_X42Y53_R_t(R_t_top[1313]),
    .Tile_X42Y53_R_f(R_f_top[1313]),
    .Tile_X45Y53_R_t(R_t_top[1314]),
    .Tile_X45Y53_R_f(R_f_top[1314]),
    .Tile_X48Y53_R_t(R_t_top[1315]),
    .Tile_X48Y53_R_f(R_f_top[1315]),
    .Tile_X51Y53_R_t(R_t_top[1316]),
    .Tile_X51Y53_R_f(R_f_top[1316]),
    .Tile_X54Y53_R_t(R_t_top[1317]),
    .Tile_X54Y53_R_f(R_f_top[1317]),
    .Tile_X57Y53_R_t(R_t_top[1318]),
    .Tile_X57Y53_R_f(R_f_top[1318]),
    .Tile_X60Y53_R_t(R_t_top[1319]),
    .Tile_X60Y53_R_f(R_f_top[1319]),
    .Tile_X63Y53_R_t(R_t_top[1320]),
    .Tile_X63Y53_R_f(R_f_top[1320]),
    .Tile_X66Y53_R_t(R_t_top[1321]),
    .Tile_X66Y53_R_f(R_f_top[1321]),
    .Tile_X69Y53_R_t(R_t_top[1322]),
    .Tile_X69Y53_R_f(R_f_top[1322]),
    .Tile_X72Y53_R_t(R_t_top[1323]),
    .Tile_X72Y53_R_f(R_f_top[1323]),
    .Tile_X75Y53_R_t(R_t_top[1324]),
    .Tile_X75Y53_R_f(R_f_top[1324]),
    .Tile_X3Y54_R_t(R_t_top[1325]),
    .Tile_X3Y54_R_f(R_f_top[1325]),
    .Tile_X6Y54_R_t(R_t_top[1326]),
    .Tile_X6Y54_R_f(R_f_top[1326]),
    .Tile_X9Y54_R_t(R_t_top[1327]),
    .Tile_X9Y54_R_f(R_f_top[1327]),
    .Tile_X12Y54_R_t(R_t_top[1328]),
    .Tile_X12Y54_R_f(R_f_top[1328]),
    .Tile_X15Y54_R_t(R_t_top[1329]),
    .Tile_X15Y54_R_f(R_f_top[1329]),
    .Tile_X18Y54_R_t(R_t_top[1330]),
    .Tile_X18Y54_R_f(R_f_top[1330]),
    .Tile_X21Y54_R_t(R_t_top[1331]),
    .Tile_X21Y54_R_f(R_f_top[1331]),
    .Tile_X24Y54_R_t(R_t_top[1332]),
    .Tile_X24Y54_R_f(R_f_top[1332]),
    .Tile_X27Y54_R_t(R_t_top[1333]),
    .Tile_X27Y54_R_f(R_f_top[1333]),
    .Tile_X30Y54_R_t(R_t_top[1334]),
    .Tile_X30Y54_R_f(R_f_top[1334]),
    .Tile_X33Y54_R_t(R_t_top[1335]),
    .Tile_X33Y54_R_f(R_f_top[1335]),
    .Tile_X36Y54_R_t(R_t_top[1336]),
    .Tile_X36Y54_R_f(R_f_top[1336]),
    .Tile_X39Y54_R_t(R_t_top[1337]),
    .Tile_X39Y54_R_f(R_f_top[1337]),
    .Tile_X42Y54_R_t(R_t_top[1338]),
    .Tile_X42Y54_R_f(R_f_top[1338]),
    .Tile_X45Y54_R_t(R_t_top[1339]),
    .Tile_X45Y54_R_f(R_f_top[1339]),
    .Tile_X48Y54_R_t(R_t_top[1340]),
    .Tile_X48Y54_R_f(R_f_top[1340]),
    .Tile_X51Y54_R_t(R_t_top[1341]),
    .Tile_X51Y54_R_f(R_f_top[1341]),
    .Tile_X54Y54_R_t(R_t_top[1342]),
    .Tile_X54Y54_R_f(R_f_top[1342]),
    .Tile_X57Y54_R_t(R_t_top[1343]),
    .Tile_X57Y54_R_f(R_f_top[1343]),
    .Tile_X60Y54_R_t(R_t_top[1344]),
    .Tile_X60Y54_R_f(R_f_top[1344]),
    .Tile_X63Y54_R_t(R_t_top[1345]),
    .Tile_X63Y54_R_f(R_f_top[1345]),
    .Tile_X66Y54_R_t(R_t_top[1346]),
    .Tile_X66Y54_R_f(R_f_top[1346]),
    .Tile_X69Y54_R_t(R_t_top[1347]),
    .Tile_X69Y54_R_f(R_f_top[1347]),
    .Tile_X72Y54_R_t(R_t_top[1348]),
    .Tile_X72Y54_R_f(R_f_top[1348]),
    .Tile_X75Y54_R_t(R_t_top[1349]),
    .Tile_X75Y54_R_f(R_f_top[1349]),
    .Tile_X3Y55_R_t(R_t_top[1350]),
    .Tile_X3Y55_R_f(R_f_top[1350]),
    .Tile_X6Y55_R_t(R_t_top[1351]),
    .Tile_X6Y55_R_f(R_f_top[1351]),
    .Tile_X9Y55_R_t(R_t_top[1352]),
    .Tile_X9Y55_R_f(R_f_top[1352]),
    .Tile_X12Y55_R_t(R_t_top[1353]),
    .Tile_X12Y55_R_f(R_f_top[1353]),
    .Tile_X15Y55_R_t(R_t_top[1354]),
    .Tile_X15Y55_R_f(R_f_top[1354]),
    .Tile_X18Y55_R_t(R_t_top[1355]),
    .Tile_X18Y55_R_f(R_f_top[1355]),
    .Tile_X21Y55_R_t(R_t_top[1356]),
    .Tile_X21Y55_R_f(R_f_top[1356]),
    .Tile_X24Y55_R_t(R_t_top[1357]),
    .Tile_X24Y55_R_f(R_f_top[1357]),
    .Tile_X27Y55_R_t(R_t_top[1358]),
    .Tile_X27Y55_R_f(R_f_top[1358]),
    .Tile_X30Y55_R_t(R_t_top[1359]),
    .Tile_X30Y55_R_f(R_f_top[1359]),
    .Tile_X33Y55_R_t(R_t_top[1360]),
    .Tile_X33Y55_R_f(R_f_top[1360]),
    .Tile_X36Y55_R_t(R_t_top[1361]),
    .Tile_X36Y55_R_f(R_f_top[1361]),
    .Tile_X39Y55_R_t(R_t_top[1362]),
    .Tile_X39Y55_R_f(R_f_top[1362]),
    .Tile_X42Y55_R_t(R_t_top[1363]),
    .Tile_X42Y55_R_f(R_f_top[1363]),
    .Tile_X45Y55_R_t(R_t_top[1364]),
    .Tile_X45Y55_R_f(R_f_top[1364]),
    .Tile_X48Y55_R_t(R_t_top[1365]),
    .Tile_X48Y55_R_f(R_f_top[1365]),
    .Tile_X51Y55_R_t(R_t_top[1366]),
    .Tile_X51Y55_R_f(R_f_top[1366]),
    .Tile_X54Y55_R_t(R_t_top[1367]),
    .Tile_X54Y55_R_f(R_f_top[1367]),
    .Tile_X57Y55_R_t(R_t_top[1368]),
    .Tile_X57Y55_R_f(R_f_top[1368]),
    .Tile_X60Y55_R_t(R_t_top[1369]),
    .Tile_X60Y55_R_f(R_f_top[1369]),
    .Tile_X63Y55_R_t(R_t_top[1370]),
    .Tile_X63Y55_R_f(R_f_top[1370]),
    .Tile_X66Y55_R_t(R_t_top[1371]),
    .Tile_X66Y55_R_f(R_f_top[1371]),
    .Tile_X69Y55_R_t(R_t_top[1372]),
    .Tile_X69Y55_R_f(R_f_top[1372]),
    .Tile_X72Y55_R_t(R_t_top[1373]),
    .Tile_X72Y55_R_f(R_f_top[1373]),
    .Tile_X75Y55_R_t(R_t_top[1374]),
    .Tile_X75Y55_R_f(R_f_top[1374]),
    .Tile_X3Y56_R_t(R_t_top[1375]),
    .Tile_X3Y56_R_f(R_f_top[1375]),
    .Tile_X6Y56_R_t(R_t_top[1376]),
    .Tile_X6Y56_R_f(R_f_top[1376]),
    .Tile_X9Y56_R_t(R_t_top[1377]),
    .Tile_X9Y56_R_f(R_f_top[1377]),
    .Tile_X12Y56_R_t(R_t_top[1378]),
    .Tile_X12Y56_R_f(R_f_top[1378]),
    .Tile_X15Y56_R_t(R_t_top[1379]),
    .Tile_X15Y56_R_f(R_f_top[1379]),
    .Tile_X18Y56_R_t(R_t_top[1380]),
    .Tile_X18Y56_R_f(R_f_top[1380]),
    .Tile_X21Y56_R_t(R_t_top[1381]),
    .Tile_X21Y56_R_f(R_f_top[1381]),
    .Tile_X24Y56_R_t(R_t_top[1382]),
    .Tile_X24Y56_R_f(R_f_top[1382]),
    .Tile_X27Y56_R_t(R_t_top[1383]),
    .Tile_X27Y56_R_f(R_f_top[1383]),
    .Tile_X30Y56_R_t(R_t_top[1384]),
    .Tile_X30Y56_R_f(R_f_top[1384]),
    .Tile_X33Y56_R_t(R_t_top[1385]),
    .Tile_X33Y56_R_f(R_f_top[1385]),
    .Tile_X36Y56_R_t(R_t_top[1386]),
    .Tile_X36Y56_R_f(R_f_top[1386]),
    .Tile_X39Y56_R_t(R_t_top[1387]),
    .Tile_X39Y56_R_f(R_f_top[1387]),
    .Tile_X42Y56_R_t(R_t_top[1388]),
    .Tile_X42Y56_R_f(R_f_top[1388]),
    .Tile_X45Y56_R_t(R_t_top[1389]),
    .Tile_X45Y56_R_f(R_f_top[1389]),
    .Tile_X48Y56_R_t(R_t_top[1390]),
    .Tile_X48Y56_R_f(R_f_top[1390]),
    .Tile_X51Y56_R_t(R_t_top[1391]),
    .Tile_X51Y56_R_f(R_f_top[1391]),
    .Tile_X54Y56_R_t(R_t_top[1392]),
    .Tile_X54Y56_R_f(R_f_top[1392]),
    .Tile_X57Y56_R_t(R_t_top[1393]),
    .Tile_X57Y56_R_f(R_f_top[1393]),
    .Tile_X60Y56_R_t(R_t_top[1394]),
    .Tile_X60Y56_R_f(R_f_top[1394]),
    .Tile_X63Y56_R_t(R_t_top[1395]),
    .Tile_X63Y56_R_f(R_f_top[1395]),
    .Tile_X66Y56_R_t(R_t_top[1396]),
    .Tile_X66Y56_R_f(R_f_top[1396]),
    .Tile_X69Y56_R_t(R_t_top[1397]),
    .Tile_X69Y56_R_f(R_f_top[1397]),
    .Tile_X72Y56_R_t(R_t_top[1398]),
    .Tile_X72Y56_R_f(R_f_top[1398]),
    .Tile_X75Y56_R_t(R_t_top[1399]),
    .Tile_X75Y56_R_f(R_f_top[1399]),
    .Tile_X3Y57_R_t(R_t_top[1400]),
    .Tile_X3Y57_R_f(R_f_top[1400]),
    .Tile_X6Y57_R_t(R_t_top[1401]),
    .Tile_X6Y57_R_f(R_f_top[1401]),
    .Tile_X9Y57_R_t(R_t_top[1402]),
    .Tile_X9Y57_R_f(R_f_top[1402]),
    .Tile_X12Y57_R_t(R_t_top[1403]),
    .Tile_X12Y57_R_f(R_f_top[1403]),
    .Tile_X15Y57_R_t(R_t_top[1404]),
    .Tile_X15Y57_R_f(R_f_top[1404]),
    .Tile_X18Y57_R_t(R_t_top[1405]),
    .Tile_X18Y57_R_f(R_f_top[1405]),
    .Tile_X21Y57_R_t(R_t_top[1406]),
    .Tile_X21Y57_R_f(R_f_top[1406]),
    .Tile_X24Y57_R_t(R_t_top[1407]),
    .Tile_X24Y57_R_f(R_f_top[1407]),
    .Tile_X27Y57_R_t(R_t_top[1408]),
    .Tile_X27Y57_R_f(R_f_top[1408]),
    .Tile_X30Y57_R_t(R_t_top[1409]),
    .Tile_X30Y57_R_f(R_f_top[1409]),
    .Tile_X33Y57_R_t(R_t_top[1410]),
    .Tile_X33Y57_R_f(R_f_top[1410]),
    .Tile_X36Y57_R_t(R_t_top[1411]),
    .Tile_X36Y57_R_f(R_f_top[1411]),
    .Tile_X39Y57_R_t(R_t_top[1412]),
    .Tile_X39Y57_R_f(R_f_top[1412]),
    .Tile_X42Y57_R_t(R_t_top[1413]),
    .Tile_X42Y57_R_f(R_f_top[1413]),
    .Tile_X45Y57_R_t(R_t_top[1414]),
    .Tile_X45Y57_R_f(R_f_top[1414]),
    .Tile_X48Y57_R_t(R_t_top[1415]),
    .Tile_X48Y57_R_f(R_f_top[1415]),
    .Tile_X51Y57_R_t(R_t_top[1416]),
    .Tile_X51Y57_R_f(R_f_top[1416]),
    .Tile_X54Y57_R_t(R_t_top[1417]),
    .Tile_X54Y57_R_f(R_f_top[1417]),
    .Tile_X57Y57_R_t(R_t_top[1418]),
    .Tile_X57Y57_R_f(R_f_top[1418]),
    .Tile_X60Y57_R_t(R_t_top[1419]),
    .Tile_X60Y57_R_f(R_f_top[1419]),
    .Tile_X63Y57_R_t(R_t_top[1420]),
    .Tile_X63Y57_R_f(R_f_top[1420]),
    .Tile_X66Y57_R_t(R_t_top[1421]),
    .Tile_X66Y57_R_f(R_f_top[1421]),
    .Tile_X69Y57_R_t(R_t_top[1422]),
    .Tile_X69Y57_R_f(R_f_top[1422]),
    .Tile_X72Y57_R_t(R_t_top[1423]),
    .Tile_X72Y57_R_f(R_f_top[1423]),
    .Tile_X75Y57_R_t(R_t_top[1424]),
    .Tile_X75Y57_R_f(R_f_top[1424]),
    .Tile_X3Y58_R_t(R_t_top[1425]),
    .Tile_X3Y58_R_f(R_f_top[1425]),
    .Tile_X6Y58_R_t(R_t_top[1426]),
    .Tile_X6Y58_R_f(R_f_top[1426]),
    .Tile_X9Y58_R_t(R_t_top[1427]),
    .Tile_X9Y58_R_f(R_f_top[1427]),
    .Tile_X12Y58_R_t(R_t_top[1428]),
    .Tile_X12Y58_R_f(R_f_top[1428]),
    .Tile_X15Y58_R_t(R_t_top[1429]),
    .Tile_X15Y58_R_f(R_f_top[1429]),
    .Tile_X18Y58_R_t(R_t_top[1430]),
    .Tile_X18Y58_R_f(R_f_top[1430]),
    .Tile_X21Y58_R_t(R_t_top[1431]),
    .Tile_X21Y58_R_f(R_f_top[1431]),
    .Tile_X24Y58_R_t(R_t_top[1432]),
    .Tile_X24Y58_R_f(R_f_top[1432]),
    .Tile_X27Y58_R_t(R_t_top[1433]),
    .Tile_X27Y58_R_f(R_f_top[1433]),
    .Tile_X30Y58_R_t(R_t_top[1434]),
    .Tile_X30Y58_R_f(R_f_top[1434]),
    .Tile_X33Y58_R_t(R_t_top[1435]),
    .Tile_X33Y58_R_f(R_f_top[1435]),
    .Tile_X36Y58_R_t(R_t_top[1436]),
    .Tile_X36Y58_R_f(R_f_top[1436]),
    .Tile_X39Y58_R_t(R_t_top[1437]),
    .Tile_X39Y58_R_f(R_f_top[1437]),
    .Tile_X42Y58_R_t(R_t_top[1438]),
    .Tile_X42Y58_R_f(R_f_top[1438]),
    .Tile_X45Y58_R_t(R_t_top[1439]),
    .Tile_X45Y58_R_f(R_f_top[1439]),
    .Tile_X48Y58_R_t(R_t_top[1440]),
    .Tile_X48Y58_R_f(R_f_top[1440]),
    .Tile_X51Y58_R_t(R_t_top[1441]),
    .Tile_X51Y58_R_f(R_f_top[1441]),
    .Tile_X54Y58_R_t(R_t_top[1442]),
    .Tile_X54Y58_R_f(R_f_top[1442]),
    .Tile_X57Y58_R_t(R_t_top[1443]),
    .Tile_X57Y58_R_f(R_f_top[1443]),
    .Tile_X60Y58_R_t(R_t_top[1444]),
    .Tile_X60Y58_R_f(R_f_top[1444]),
    .Tile_X63Y58_R_t(R_t_top[1445]),
    .Tile_X63Y58_R_f(R_f_top[1445]),
    .Tile_X66Y58_R_t(R_t_top[1446]),
    .Tile_X66Y58_R_f(R_f_top[1446]),
    .Tile_X69Y58_R_t(R_t_top[1447]),
    .Tile_X69Y58_R_f(R_f_top[1447]),
    .Tile_X72Y58_R_t(R_t_top[1448]),
    .Tile_X72Y58_R_f(R_f_top[1448]),
    .Tile_X75Y58_R_t(R_t_top[1449]),
    .Tile_X75Y58_R_f(R_f_top[1449]),
    .Tile_X3Y59_R_t(R_t_top[1450]),
    .Tile_X3Y59_R_f(R_f_top[1450]),
    .Tile_X6Y59_R_t(R_t_top[1451]),
    .Tile_X6Y59_R_f(R_f_top[1451]),
    .Tile_X9Y59_R_t(R_t_top[1452]),
    .Tile_X9Y59_R_f(R_f_top[1452]),
    .Tile_X12Y59_R_t(R_t_top[1453]),
    .Tile_X12Y59_R_f(R_f_top[1453]),
    .Tile_X15Y59_R_t(R_t_top[1454]),
    .Tile_X15Y59_R_f(R_f_top[1454]),
    .Tile_X18Y59_R_t(R_t_top[1455]),
    .Tile_X18Y59_R_f(R_f_top[1455]),
    .Tile_X21Y59_R_t(R_t_top[1456]),
    .Tile_X21Y59_R_f(R_f_top[1456]),
    .Tile_X24Y59_R_t(R_t_top[1457]),
    .Tile_X24Y59_R_f(R_f_top[1457]),
    .Tile_X27Y59_R_t(R_t_top[1458]),
    .Tile_X27Y59_R_f(R_f_top[1458]),
    .Tile_X30Y59_R_t(R_t_top[1459]),
    .Tile_X30Y59_R_f(R_f_top[1459]),
    .Tile_X33Y59_R_t(R_t_top[1460]),
    .Tile_X33Y59_R_f(R_f_top[1460]),
    .Tile_X36Y59_R_t(R_t_top[1461]),
    .Tile_X36Y59_R_f(R_f_top[1461]),
    .Tile_X39Y59_R_t(R_t_top[1462]),
    .Tile_X39Y59_R_f(R_f_top[1462]),
    .Tile_X42Y59_R_t(R_t_top[1463]),
    .Tile_X42Y59_R_f(R_f_top[1463]),
    .Tile_X45Y59_R_t(R_t_top[1464]),
    .Tile_X45Y59_R_f(R_f_top[1464]),
    .Tile_X48Y59_R_t(R_t_top[1465]),
    .Tile_X48Y59_R_f(R_f_top[1465]),
    .Tile_X51Y59_R_t(R_t_top[1466]),
    .Tile_X51Y59_R_f(R_f_top[1466]),
    .Tile_X54Y59_R_t(R_t_top[1467]),
    .Tile_X54Y59_R_f(R_f_top[1467]),
    .Tile_X57Y59_R_t(R_t_top[1468]),
    .Tile_X57Y59_R_f(R_f_top[1468]),
    .Tile_X60Y59_R_t(R_t_top[1469]),
    .Tile_X60Y59_R_f(R_f_top[1469]),
    .Tile_X63Y59_R_t(R_t_top[1470]),
    .Tile_X63Y59_R_f(R_f_top[1470]),
    .Tile_X66Y59_R_t(R_t_top[1471]),
    .Tile_X66Y59_R_f(R_f_top[1471]),
    .Tile_X69Y59_R_t(R_t_top[1472]),
    .Tile_X69Y59_R_f(R_f_top[1472]),
    .Tile_X72Y59_R_t(R_t_top[1473]),
    .Tile_X72Y59_R_f(R_f_top[1473]),
    .Tile_X75Y59_R_t(R_t_top[1474]),
    .Tile_X75Y59_R_f(R_f_top[1474]),
    .Tile_X3Y60_R_t(R_t_top[1475]),
    .Tile_X3Y60_R_f(R_f_top[1475]),
    .Tile_X6Y60_R_t(R_t_top[1476]),
    .Tile_X6Y60_R_f(R_f_top[1476]),
    .Tile_X9Y60_R_t(R_t_top[1477]),
    .Tile_X9Y60_R_f(R_f_top[1477]),
    .Tile_X12Y60_R_t(R_t_top[1478]),
    .Tile_X12Y60_R_f(R_f_top[1478]),
    .Tile_X15Y60_R_t(R_t_top[1479]),
    .Tile_X15Y60_R_f(R_f_top[1479]),
    .Tile_X18Y60_R_t(R_t_top[1480]),
    .Tile_X18Y60_R_f(R_f_top[1480]),
    .Tile_X21Y60_R_t(R_t_top[1481]),
    .Tile_X21Y60_R_f(R_f_top[1481]),
    .Tile_X24Y60_R_t(R_t_top[1482]),
    .Tile_X24Y60_R_f(R_f_top[1482]),
    .Tile_X27Y60_R_t(R_t_top[1483]),
    .Tile_X27Y60_R_f(R_f_top[1483]),
    .Tile_X30Y60_R_t(R_t_top[1484]),
    .Tile_X30Y60_R_f(R_f_top[1484]),
    .Tile_X33Y60_R_t(R_t_top[1485]),
    .Tile_X33Y60_R_f(R_f_top[1485]),
    .Tile_X36Y60_R_t(R_t_top[1486]),
    .Tile_X36Y60_R_f(R_f_top[1486]),
    .Tile_X39Y60_R_t(R_t_top[1487]),
    .Tile_X39Y60_R_f(R_f_top[1487]),
    .Tile_X42Y60_R_t(R_t_top[1488]),
    .Tile_X42Y60_R_f(R_f_top[1488]),
    .Tile_X45Y60_R_t(R_t_top[1489]),
    .Tile_X45Y60_R_f(R_f_top[1489]),
    .Tile_X48Y60_R_t(R_t_top[1490]),
    .Tile_X48Y60_R_f(R_f_top[1490]),
    .Tile_X51Y60_R_t(R_t_top[1491]),
    .Tile_X51Y60_R_f(R_f_top[1491]),
    .Tile_X54Y60_R_t(R_t_top[1492]),
    .Tile_X54Y60_R_f(R_f_top[1492]),
    .Tile_X57Y60_R_t(R_t_top[1493]),
    .Tile_X57Y60_R_f(R_f_top[1493]),
    .Tile_X60Y60_R_t(R_t_top[1494]),
    .Tile_X60Y60_R_f(R_f_top[1494]),
    .Tile_X63Y60_R_t(R_t_top[1495]),
    .Tile_X63Y60_R_f(R_f_top[1495]),
    .Tile_X66Y60_R_t(R_t_top[1496]),
    .Tile_X66Y60_R_f(R_f_top[1496]),
    .Tile_X69Y60_R_t(R_t_top[1497]),
    .Tile_X69Y60_R_f(R_f_top[1497]),
    .Tile_X72Y60_R_t(R_t_top[1498]),
    .Tile_X72Y60_R_f(R_f_top[1498]),
    .Tile_X75Y60_R_t(R_t_top[1499]),
    .Tile_X75Y60_R_f(R_f_top[1499]),
    .Tile_X0Y1_A_F_masked1(F_masked1_top[0]),
    .Tile_X0Y1_A_F_masked2(F_masked2_top[0]),
    .Tile_X0Y2_A_F_masked1(F_masked1_top[1]),
    .Tile_X0Y2_A_F_masked2(F_masked2_top[1]),
    .Tile_X0Y3_A_F_masked1(F_masked1_top[2]),
    .Tile_X0Y3_A_F_masked2(F_masked2_top[2]),
    .Tile_X0Y4_A_F_masked1(F_masked1_top[3]),
    .Tile_X0Y4_A_F_masked2(F_masked2_top[3]),
    .Tile_X0Y5_A_F_masked1(F_masked1_top[4]),
    .Tile_X0Y5_A_F_masked2(F_masked2_top[4]),
    .Tile_X0Y6_A_F_masked1(F_masked1_top[5]),
    .Tile_X0Y6_A_F_masked2(F_masked2_top[5]),
    .Tile_X0Y7_A_F_masked1(F_masked1_top[6]),
    .Tile_X0Y7_A_F_masked2(F_masked2_top[6]),
    .Tile_X0Y8_A_F_masked1(F_masked1_top[7]),
    .Tile_X0Y8_A_F_masked2(F_masked2_top[7]),
    .Tile_X0Y9_A_F_masked1(F_masked1_top[8]),
    .Tile_X0Y9_A_F_masked2(F_masked2_top[8]),
    .Tile_X0Y10_A_F_masked1(F_masked1_top[9]),
    .Tile_X0Y10_A_F_masked2(F_masked2_top[9]),
    .Tile_X0Y11_A_F_masked1(F_masked1_top[10]),
    .Tile_X0Y11_A_F_masked2(F_masked2_top[10]),
    .Tile_X0Y12_A_F_masked1(F_masked1_top[11]),
    .Tile_X0Y12_A_F_masked2(F_masked2_top[11]),
    .Tile_X0Y13_A_F_masked1(F_masked1_top[12]),
    .Tile_X0Y13_A_F_masked2(F_masked2_top[12]),
    .Tile_X0Y14_A_F_masked1(F_masked1_top[13]),
    .Tile_X0Y14_A_F_masked2(F_masked2_top[13]),
    .Tile_X0Y15_A_F_masked1(F_masked1_top[14]),
    .Tile_X0Y15_A_F_masked2(F_masked2_top[14]),
    .Tile_X0Y16_A_F_masked1(F_masked1_top[15]),
    .Tile_X0Y16_A_F_masked2(F_masked2_top[15]),
    .Tile_X0Y17_A_F_masked1(F_masked1_top[16]),
    .Tile_X0Y17_A_F_masked2(F_masked2_top[16]),
    .Tile_X0Y18_A_F_masked1(F_masked1_top[17]),
    .Tile_X0Y18_A_F_masked2(F_masked2_top[17]),
    .Tile_X0Y19_A_F_masked1(F_masked1_top[18]),
    .Tile_X0Y19_A_F_masked2(F_masked2_top[18]),
    .Tile_X0Y20_A_F_masked1(F_masked1_top[19]),
    .Tile_X0Y20_A_F_masked2(F_masked2_top[19]),
    .Tile_X0Y21_A_F_masked1(F_masked1_top[20]),
    .Tile_X0Y21_A_F_masked2(F_masked2_top[20]),
    .Tile_X0Y22_A_F_masked1(F_masked1_top[21]),
    .Tile_X0Y22_A_F_masked2(F_masked2_top[21]),
    .Tile_X0Y23_A_F_masked1(F_masked1_top[22]),
    .Tile_X0Y23_A_F_masked2(F_masked2_top[22]),
    .Tile_X0Y24_A_F_masked1(F_masked1_top[23]),
    .Tile_X0Y24_A_F_masked2(F_masked2_top[23]),
    .Tile_X0Y25_A_F_masked1(F_masked1_top[24]),
    .Tile_X0Y25_A_F_masked2(F_masked2_top[24]),
    .Tile_X0Y26_A_F_masked1(F_masked1_top[25]),
    .Tile_X0Y26_A_F_masked2(F_masked2_top[25]),
    .Tile_X0Y27_A_F_masked1(F_masked1_top[26]),
    .Tile_X0Y27_A_F_masked2(F_masked2_top[26]),
    .Tile_X0Y28_A_F_masked1(F_masked1_top[27]),
    .Tile_X0Y28_A_F_masked2(F_masked2_top[27]),
    .Tile_X0Y29_A_F_masked1(F_masked1_top[28]),
    .Tile_X0Y29_A_F_masked2(F_masked2_top[28]),
    .Tile_X0Y30_A_F_masked1(F_masked1_top[29]),
    .Tile_X0Y30_A_F_masked2(F_masked2_top[29]),
    .Tile_X0Y31_A_F_masked1(F_masked1_top[30]),
    .Tile_X0Y31_A_F_masked2(F_masked2_top[30]),
    .Tile_X0Y32_A_F_masked1(F_masked1_top[31]),
    .Tile_X0Y32_A_F_masked2(F_masked2_top[31]),
    .Tile_X0Y33_A_F_masked1(F_masked1_top[32]),
    .Tile_X0Y33_A_F_masked2(F_masked2_top[32]),
    .Tile_X0Y34_A_F_masked1(F_masked1_top[33]),
    .Tile_X0Y34_A_F_masked2(F_masked2_top[33]),
    .Tile_X0Y35_A_F_masked1(F_masked1_top[34]),
    .Tile_X0Y35_A_F_masked2(F_masked2_top[34]),
    .Tile_X0Y36_A_F_masked1(F_masked1_top[35]),
    .Tile_X0Y36_A_F_masked2(F_masked2_top[35]),
    .Tile_X0Y37_A_F_masked1(F_masked1_top[36]),
    .Tile_X0Y37_A_F_masked2(F_masked2_top[36]),
    .Tile_X0Y38_A_F_masked1(F_masked1_top[37]),
    .Tile_X0Y38_A_F_masked2(F_masked2_top[37]),
    .Tile_X0Y39_A_F_masked1(F_masked1_top[38]),
    .Tile_X0Y39_A_F_masked2(F_masked2_top[38]),
    .Tile_X0Y40_A_F_masked1(F_masked1_top[39]),
    .Tile_X0Y40_A_F_masked2(F_masked2_top[39]),
    .Tile_X0Y41_A_F_masked1(F_masked1_top[40]),
    .Tile_X0Y41_A_F_masked2(F_masked2_top[40]),
    .Tile_X0Y42_A_F_masked1(F_masked1_top[41]),
    .Tile_X0Y42_A_F_masked2(F_masked2_top[41]),
    .Tile_X0Y43_A_F_masked1(F_masked1_top[42]),
    .Tile_X0Y43_A_F_masked2(F_masked2_top[42]),
    .Tile_X0Y44_A_F_masked1(F_masked1_top[43]),
    .Tile_X0Y44_A_F_masked2(F_masked2_top[43]),
    .Tile_X0Y45_A_F_masked1(F_masked1_top[44]),
    .Tile_X0Y45_A_F_masked2(F_masked2_top[44]),
    .Tile_X0Y46_A_F_masked1(F_masked1_top[45]),
    .Tile_X0Y46_A_F_masked2(F_masked2_top[45]),
    .Tile_X0Y47_A_F_masked1(F_masked1_top[46]),
    .Tile_X0Y47_A_F_masked2(F_masked2_top[46]),
    .Tile_X0Y48_A_F_masked1(F_masked1_top[47]),
    .Tile_X0Y48_A_F_masked2(F_masked2_top[47]),
    .Tile_X0Y49_A_F_masked1(F_masked1_top[48]),
    .Tile_X0Y49_A_F_masked2(F_masked2_top[48]),
    .Tile_X0Y50_A_F_masked1(F_masked1_top[49]),
    .Tile_X0Y50_A_F_masked2(F_masked2_top[49]),
    .Tile_X0Y51_A_F_masked1(F_masked1_top[50]),
    .Tile_X0Y51_A_F_masked2(F_masked2_top[50]),
    .Tile_X0Y52_A_F_masked1(F_masked1_top[51]),
    .Tile_X0Y52_A_F_masked2(F_masked2_top[51]),
    .Tile_X0Y53_A_F_masked1(F_masked1_top[52]),
    .Tile_X0Y53_A_F_masked2(F_masked2_top[52]),
    .Tile_X0Y54_A_F_masked1(F_masked1_top[53]),
    .Tile_X0Y54_A_F_masked2(F_masked2_top[53]),
    .Tile_X0Y55_A_F_masked1(F_masked1_top[54]),
    .Tile_X0Y55_A_F_masked2(F_masked2_top[54]),
    .Tile_X0Y56_A_F_masked1(F_masked1_top[55]),
    .Tile_X0Y56_A_F_masked2(F_masked2_top[55]),
    .Tile_X0Y57_A_F_masked1(F_masked1_top[56]),
    .Tile_X0Y57_A_F_masked2(F_masked2_top[56]),
    .Tile_X0Y58_A_F_masked1(F_masked1_top[57]),
    .Tile_X0Y58_A_F_masked2(F_masked2_top[57]),
    .Tile_X0Y59_A_F_masked1(F_masked1_top[58]),
    .Tile_X0Y59_A_F_masked2(F_masked2_top[58]),
    .Tile_X0Y60_A_F_masked1(F_masked1_top[59]),
    .Tile_X0Y60_A_F_masked2(F_masked2_top[59]),
    .Tile_X38Y1_A_F_ctrl(F_ctrl_top[0]),
    .Tile_X38Y2_A_F_ctrl(F_ctrl_top[1]),
    .Tile_X38Y3_A_F_ctrl(F_ctrl_top[2]),
    .Tile_X38Y4_A_F_ctrl(F_ctrl_top[3]),
    .Tile_X38Y5_A_F_ctrl(F_ctrl_top[4]),
    .Tile_X38Y6_A_F_ctrl(F_ctrl_top[5]),
    .Tile_X38Y7_A_F_ctrl(F_ctrl_top[6]),
    .Tile_X38Y8_A_F_ctrl(F_ctrl_top[7]),
    .Tile_X38Y9_A_F_ctrl(F_ctrl_top[8]),
    .Tile_X38Y10_A_F_ctrl(F_ctrl_top[9]),
    .Tile_X38Y11_A_F_ctrl(F_ctrl_top[10]),
    .Tile_X38Y12_A_F_ctrl(F_ctrl_top[11]),
    .Tile_X38Y13_A_F_ctrl(F_ctrl_top[12]),
    .Tile_X38Y14_A_F_ctrl(F_ctrl_top[13]),
    .Tile_X38Y15_A_F_ctrl(F_ctrl_top[14]),
    .Tile_X38Y16_A_F_ctrl(F_ctrl_top[15]),
    .Tile_X38Y17_A_F_ctrl(F_ctrl_top[16]),
    .Tile_X38Y18_A_F_ctrl(F_ctrl_top[17]),
    .Tile_X38Y19_A_F_ctrl(F_ctrl_top[18]),
    .Tile_X38Y20_A_F_ctrl(F_ctrl_top[19]),
    .Tile_X38Y21_A_F_ctrl(F_ctrl_top[20]),
    .Tile_X38Y22_A_F_ctrl(F_ctrl_top[21]),
    .Tile_X38Y23_A_F_ctrl(F_ctrl_top[22]),
    .Tile_X38Y24_A_F_ctrl(F_ctrl_top[23]),
    .Tile_X38Y25_A_F_ctrl(F_ctrl_top[24]),
    .Tile_X38Y26_A_F_ctrl(F_ctrl_top[25]),
    .Tile_X38Y27_A_F_ctrl(F_ctrl_top[26]),
    .Tile_X38Y28_A_F_ctrl(F_ctrl_top[27]),
    .Tile_X38Y29_A_F_ctrl(F_ctrl_top[28]),
    .Tile_X38Y30_A_F_ctrl(F_ctrl_top[29]),
    .Tile_X38Y31_A_F_ctrl(F_ctrl_top[30]),
    .Tile_X38Y32_A_F_ctrl(F_ctrl_top[31]),
    .Tile_X38Y33_A_F_ctrl(F_ctrl_top[32]),
    .Tile_X38Y34_A_F_ctrl(F_ctrl_top[33]),
    .Tile_X38Y35_A_F_ctrl(F_ctrl_top[34]),
    .Tile_X38Y36_A_F_ctrl(F_ctrl_top[35]),
    .Tile_X38Y37_A_F_ctrl(F_ctrl_top[36]),
    .Tile_X38Y38_A_F_ctrl(F_ctrl_top[37]),
    .Tile_X38Y39_A_F_ctrl(F_ctrl_top[38]),
    .Tile_X38Y40_A_F_ctrl(F_ctrl_top[39]),
    .Tile_X38Y41_A_F_ctrl(F_ctrl_top[40]),
    .Tile_X38Y42_A_F_ctrl(F_ctrl_top[41]),
    .Tile_X38Y43_A_F_ctrl(F_ctrl_top[42]),
    .Tile_X38Y44_A_F_ctrl(F_ctrl_top[43]),
    .Tile_X38Y45_A_F_ctrl(F_ctrl_top[44]),
    .Tile_X38Y46_A_F_ctrl(F_ctrl_top[45]),
    .Tile_X38Y47_A_F_ctrl(F_ctrl_top[46]),
    .Tile_X38Y48_A_F_ctrl(F_ctrl_top[47]),
    .Tile_X38Y49_A_F_ctrl(F_ctrl_top[48]),
    .Tile_X38Y50_A_F_ctrl(F_ctrl_top[49]),
    .Tile_X38Y51_A_F_ctrl(F_ctrl_top[50]),
    .Tile_X38Y52_A_F_ctrl(F_ctrl_top[51]),
    .Tile_X38Y53_A_F_ctrl(F_ctrl_top[52]),
    .Tile_X38Y54_A_F_ctrl(F_ctrl_top[53]),
    .Tile_X38Y55_A_F_ctrl(F_ctrl_top[54]),
    .Tile_X38Y56_A_F_ctrl(F_ctrl_top[55]),
    .Tile_X38Y57_A_F_ctrl(F_ctrl_top[56]),
    .Tile_X38Y58_A_F_ctrl(F_ctrl_top[57]),
    .Tile_X38Y59_A_F_ctrl(F_ctrl_top[58]),
    .Tile_X38Y60_A_F_ctrl(F_ctrl_top[59]),
    .Tile_X0Y1_A_prech1(prech1),
    .Tile_X0Y1_A_prech2(prech2),
    .Tile_X38Y1_A_prech2(prech2),
    .Tile_X0Y2_A_prech1(prech1),
    .Tile_X0Y2_A_prech2(prech2),
    .Tile_X38Y2_A_prech2(prech2),
    .Tile_X0Y3_A_prech1(prech1),
    .Tile_X0Y3_A_prech2(prech2),
    .Tile_X38Y3_A_prech2(prech2),
    .Tile_X0Y4_A_prech1(prech1),
    .Tile_X0Y4_A_prech2(prech2),
    .Tile_X38Y4_A_prech2(prech2),
    .Tile_X0Y5_A_prech1(prech1),
    .Tile_X0Y5_A_prech2(prech2),
    .Tile_X38Y5_A_prech2(prech2),
    .Tile_X0Y6_A_prech1(prech1),
    .Tile_X0Y6_A_prech2(prech2),
    .Tile_X38Y6_A_prech2(prech2),
    .Tile_X0Y7_A_prech1(prech1),
    .Tile_X0Y7_A_prech2(prech2),
    .Tile_X38Y7_A_prech2(prech2),
    .Tile_X0Y8_A_prech1(prech1),
    .Tile_X0Y8_A_prech2(prech2),
    .Tile_X38Y8_A_prech2(prech2),
    .Tile_X0Y9_A_prech1(prech1),
    .Tile_X0Y9_A_prech2(prech2),
    .Tile_X38Y9_A_prech2(prech2),
    .Tile_X0Y10_A_prech1(prech1),
    .Tile_X0Y10_A_prech2(prech2),
    .Tile_X38Y10_A_prech2(prech2),
    .Tile_X0Y11_A_prech1(prech1),
    .Tile_X0Y11_A_prech2(prech2),
    .Tile_X38Y11_A_prech2(prech2),
    .Tile_X0Y12_A_prech1(prech1),
    .Tile_X0Y12_A_prech2(prech2),
    .Tile_X38Y12_A_prech2(prech2),
    .Tile_X0Y13_A_prech1(prech1),
    .Tile_X0Y13_A_prech2(prech2),
    .Tile_X38Y13_A_prech2(prech2),
    .Tile_X0Y14_A_prech1(prech1),
    .Tile_X0Y14_A_prech2(prech2),
    .Tile_X38Y14_A_prech2(prech2),
    .Tile_X0Y15_A_prech1(prech1),
    .Tile_X0Y15_A_prech2(prech2),
    .Tile_X38Y15_A_prech2(prech2),
    .Tile_X0Y16_A_prech1(prech1),
    .Tile_X0Y16_A_prech2(prech2),
    .Tile_X38Y16_A_prech2(prech2),
    .Tile_X0Y17_A_prech1(prech1),
    .Tile_X0Y17_A_prech2(prech2),
    .Tile_X38Y17_A_prech2(prech2),
    .Tile_X0Y18_A_prech1(prech1),
    .Tile_X0Y18_A_prech2(prech2),
    .Tile_X38Y18_A_prech2(prech2),
    .Tile_X0Y19_A_prech1(prech1),
    .Tile_X0Y19_A_prech2(prech2),
    .Tile_X38Y19_A_prech2(prech2),
    .Tile_X0Y20_A_prech1(prech1),
    .Tile_X0Y20_A_prech2(prech2),
    .Tile_X38Y20_A_prech2(prech2),
    .Tile_X0Y21_A_prech1(prech1),
    .Tile_X0Y21_A_prech2(prech2),
    .Tile_X38Y21_A_prech2(prech2),
    .Tile_X0Y22_A_prech1(prech1),
    .Tile_X0Y22_A_prech2(prech2),
    .Tile_X38Y22_A_prech2(prech2),
    .Tile_X0Y23_A_prech1(prech1),
    .Tile_X0Y23_A_prech2(prech2),
    .Tile_X38Y23_A_prech2(prech2),
    .Tile_X0Y24_A_prech1(prech1),
    .Tile_X0Y24_A_prech2(prech2),
    .Tile_X38Y24_A_prech2(prech2),
    .Tile_X0Y25_A_prech1(prech1),
    .Tile_X0Y25_A_prech2(prech2),
    .Tile_X38Y25_A_prech2(prech2),
    .Tile_X0Y26_A_prech1(prech1),
    .Tile_X0Y26_A_prech2(prech2),
    .Tile_X38Y26_A_prech2(prech2),
    .Tile_X0Y27_A_prech1(prech1),
    .Tile_X0Y27_A_prech2(prech2),
    .Tile_X38Y27_A_prech2(prech2),
    .Tile_X0Y28_A_prech1(prech1),
    .Tile_X0Y28_A_prech2(prech2),
    .Tile_X38Y28_A_prech2(prech2),
    .Tile_X0Y29_A_prech1(prech1),
    .Tile_X0Y29_A_prech2(prech2),
    .Tile_X38Y29_A_prech2(prech2),
    .Tile_X0Y30_A_prech1(prech1),
    .Tile_X0Y30_A_prech2(prech2),
    .Tile_X38Y30_A_prech2(prech2),
    .Tile_X0Y31_A_prech1(prech1),
    .Tile_X0Y31_A_prech2(prech2),
    .Tile_X38Y31_A_prech2(prech2),
    .Tile_X0Y32_A_prech1(prech1),
    .Tile_X0Y32_A_prech2(prech2),
    .Tile_X38Y32_A_prech2(prech2),
    .Tile_X0Y33_A_prech1(prech1),
    .Tile_X0Y33_A_prech2(prech2),
    .Tile_X38Y33_A_prech2(prech2),
    .Tile_X0Y34_A_prech1(prech1),
    .Tile_X0Y34_A_prech2(prech2),
    .Tile_X38Y34_A_prech2(prech2),
    .Tile_X0Y35_A_prech1(prech1),
    .Tile_X0Y35_A_prech2(prech2),
    .Tile_X38Y35_A_prech2(prech2),
    .Tile_X0Y36_A_prech1(prech1),
    .Tile_X0Y36_A_prech2(prech2),
    .Tile_X38Y36_A_prech2(prech2),
    .Tile_X0Y37_A_prech1(prech1),
    .Tile_X0Y37_A_prech2(prech2),
    .Tile_X38Y37_A_prech2(prech2),
    .Tile_X0Y38_A_prech1(prech1),
    .Tile_X0Y38_A_prech2(prech2),
    .Tile_X38Y38_A_prech2(prech2),
    .Tile_X0Y39_A_prech1(prech1),
    .Tile_X0Y39_A_prech2(prech2),
    .Tile_X38Y39_A_prech2(prech2),
    .Tile_X0Y40_A_prech1(prech1),
    .Tile_X0Y40_A_prech2(prech2),
    .Tile_X38Y40_A_prech2(prech2),
    .Tile_X0Y41_A_prech1(prech1),
    .Tile_X0Y41_A_prech2(prech2),
    .Tile_X38Y41_A_prech2(prech2),
    .Tile_X0Y42_A_prech1(prech1),
    .Tile_X0Y42_A_prech2(prech2),
    .Tile_X38Y42_A_prech2(prech2),
    .Tile_X0Y43_A_prech1(prech1),
    .Tile_X0Y43_A_prech2(prech2),
    .Tile_X38Y43_A_prech2(prech2),
    .Tile_X0Y44_A_prech1(prech1),
    .Tile_X0Y44_A_prech2(prech2),
    .Tile_X38Y44_A_prech2(prech2),
    .Tile_X0Y45_A_prech1(prech1),
    .Tile_X0Y45_A_prech2(prech2),
    .Tile_X38Y45_A_prech2(prech2),
    .Tile_X0Y46_A_prech1(prech1),
    .Tile_X0Y46_A_prech2(prech2),
    .Tile_X38Y46_A_prech2(prech2),
    .Tile_X0Y47_A_prech1(prech1),
    .Tile_X0Y47_A_prech2(prech2),
    .Tile_X38Y47_A_prech2(prech2),
    .Tile_X0Y48_A_prech1(prech1),
    .Tile_X0Y48_A_prech2(prech2),
    .Tile_X38Y48_A_prech2(prech2),
    .Tile_X0Y49_A_prech1(prech1),
    .Tile_X0Y49_A_prech2(prech2),
    .Tile_X38Y49_A_prech2(prech2),
    .Tile_X0Y50_A_prech1(prech1),
    .Tile_X0Y50_A_prech2(prech2),
    .Tile_X38Y50_A_prech2(prech2),
    .Tile_X0Y51_A_prech1(prech1),
    .Tile_X0Y51_A_prech2(prech2),
    .Tile_X38Y51_A_prech2(prech2),
    .Tile_X0Y52_A_prech1(prech1),
    .Tile_X0Y52_A_prech2(prech2),
    .Tile_X38Y52_A_prech2(prech2),
    .Tile_X0Y53_A_prech1(prech1),
    .Tile_X0Y53_A_prech2(prech2),
    .Tile_X38Y53_A_prech2(prech2),
    .Tile_X0Y54_A_prech1(prech1),
    .Tile_X0Y54_A_prech2(prech2),
    .Tile_X38Y54_A_prech2(prech2),
    .Tile_X0Y55_A_prech1(prech1),
    .Tile_X0Y55_A_prech2(prech2),
    .Tile_X38Y55_A_prech2(prech2),
    .Tile_X0Y56_A_prech1(prech1),
    .Tile_X0Y56_A_prech2(prech2),
    .Tile_X38Y56_A_prech2(prech2),
    .Tile_X0Y57_A_prech1(prech1),
    .Tile_X0Y57_A_prech2(prech2),
    .Tile_X38Y57_A_prech2(prech2),
    .Tile_X0Y58_A_prech1(prech1),
    .Tile_X0Y58_A_prech2(prech2),
    .Tile_X38Y58_A_prech2(prech2),
    .Tile_X0Y59_A_prech1(prech1),
    .Tile_X0Y59_A_prech2(prech2),
    .Tile_X38Y59_A_prech2(prech2),
    .Tile_X0Y60_A_prech1(prech1),
    .Tile_X0Y60_A_prech2(prech2),
    .Tile_X38Y60_A_prech2(prech2),
    .Tile_X0Y1_A_I_top_0_t(I_top_0_t[0]),
    .Tile_X0Y1_A_I_top_0_f(I_top_0_f[0]),
    .Tile_X0Y1_A_I_top_1_t(I_top_1_t[0]),
    .Tile_X0Y1_A_I_top_1_f(I_top_1_f[0]),
    .Tile_X0Y2_A_I_top_0_t(I_top_0_t[1]),
    .Tile_X0Y2_A_I_top_0_f(I_top_0_f[1]),
    .Tile_X0Y2_A_I_top_1_t(I_top_1_t[1]),
    .Tile_X0Y2_A_I_top_1_f(I_top_1_f[1]),
    .Tile_X0Y3_A_I_top_0_t(I_top_0_t[2]),
    .Tile_X0Y3_A_I_top_0_f(I_top_0_f[2]),
    .Tile_X0Y3_A_I_top_1_t(I_top_1_t[2]),
    .Tile_X0Y3_A_I_top_1_f(I_top_1_f[2]),
    .Tile_X0Y4_A_I_top_0_t(I_top_0_t[3]),
    .Tile_X0Y4_A_I_top_0_f(I_top_0_f[3]),
    .Tile_X0Y4_A_I_top_1_t(I_top_1_t[3]),
    .Tile_X0Y4_A_I_top_1_f(I_top_1_f[3]),
    .Tile_X0Y5_A_I_top_0_t(I_top_0_t[4]),
    .Tile_X0Y5_A_I_top_0_f(I_top_0_f[4]),
    .Tile_X0Y5_A_I_top_1_t(I_top_1_t[4]),
    .Tile_X0Y5_A_I_top_1_f(I_top_1_f[4]),
    .Tile_X0Y6_A_I_top_0_t(I_top_0_t[5]),
    .Tile_X0Y6_A_I_top_0_f(I_top_0_f[5]),
    .Tile_X0Y6_A_I_top_1_t(I_top_1_t[5]),
    .Tile_X0Y6_A_I_top_1_f(I_top_1_f[5]),
    .Tile_X0Y7_A_I_top_0_t(I_top_0_t[6]),
    .Tile_X0Y7_A_I_top_0_f(I_top_0_f[6]),
    .Tile_X0Y7_A_I_top_1_t(I_top_1_t[6]),
    .Tile_X0Y7_A_I_top_1_f(I_top_1_f[6]),
    .Tile_X0Y8_A_I_top_0_t(I_top_0_t[7]),
    .Tile_X0Y8_A_I_top_0_f(I_top_0_f[7]),
    .Tile_X0Y8_A_I_top_1_t(I_top_1_t[7]),
    .Tile_X0Y8_A_I_top_1_f(I_top_1_f[7]),
    .Tile_X0Y9_A_I_top_0_t(I_top_0_t[8]),
    .Tile_X0Y9_A_I_top_0_f(I_top_0_f[8]),
    .Tile_X0Y9_A_I_top_1_t(I_top_1_t[8]),
    .Tile_X0Y9_A_I_top_1_f(I_top_1_f[8]),
    .Tile_X0Y10_A_I_top_0_t(I_top_0_t[9]),
    .Tile_X0Y10_A_I_top_0_f(I_top_0_f[9]),
    .Tile_X0Y10_A_I_top_1_t(I_top_1_t[9]),
    .Tile_X0Y10_A_I_top_1_f(I_top_1_f[9]),
    .Tile_X0Y11_A_I_top_0_t(I_top_0_t[10]),
    .Tile_X0Y11_A_I_top_0_f(I_top_0_f[10]),
    .Tile_X0Y11_A_I_top_1_t(I_top_1_t[10]),
    .Tile_X0Y11_A_I_top_1_f(I_top_1_f[10]),
    .Tile_X0Y12_A_I_top_0_t(I_top_0_t[11]),
    .Tile_X0Y12_A_I_top_0_f(I_top_0_f[11]),
    .Tile_X0Y12_A_I_top_1_t(I_top_1_t[11]),
    .Tile_X0Y12_A_I_top_1_f(I_top_1_f[11]),
    .Tile_X0Y13_A_I_top_0_t(I_top_0_t[12]),
    .Tile_X0Y13_A_I_top_0_f(I_top_0_f[12]),
    .Tile_X0Y13_A_I_top_1_t(I_top_1_t[12]),
    .Tile_X0Y13_A_I_top_1_f(I_top_1_f[12]),
    .Tile_X0Y14_A_I_top_0_t(I_top_0_t[13]),
    .Tile_X0Y14_A_I_top_0_f(I_top_0_f[13]),
    .Tile_X0Y14_A_I_top_1_t(I_top_1_t[13]),
    .Tile_X0Y14_A_I_top_1_f(I_top_1_f[13]),
    .Tile_X0Y15_A_I_top_0_t(I_top_0_t[14]),
    .Tile_X0Y15_A_I_top_0_f(I_top_0_f[14]),
    .Tile_X0Y15_A_I_top_1_t(I_top_1_t[14]),
    .Tile_X0Y15_A_I_top_1_f(I_top_1_f[14]),
    .Tile_X0Y16_A_I_top_0_t(I_top_0_t[15]),
    .Tile_X0Y16_A_I_top_0_f(I_top_0_f[15]),
    .Tile_X0Y16_A_I_top_1_t(I_top_1_t[15]),
    .Tile_X0Y16_A_I_top_1_f(I_top_1_f[15]),
    .Tile_X0Y17_A_I_top_0_t(I_top_0_t[16]),
    .Tile_X0Y17_A_I_top_0_f(I_top_0_f[16]),
    .Tile_X0Y17_A_I_top_1_t(I_top_1_t[16]),
    .Tile_X0Y17_A_I_top_1_f(I_top_1_f[16]),
    .Tile_X0Y18_A_I_top_0_t(I_top_0_t[17]),
    .Tile_X0Y18_A_I_top_0_f(I_top_0_f[17]),
    .Tile_X0Y18_A_I_top_1_t(I_top_1_t[17]),
    .Tile_X0Y18_A_I_top_1_f(I_top_1_f[17]),
    .Tile_X0Y19_A_I_top_0_t(I_top_0_t[18]),
    .Tile_X0Y19_A_I_top_0_f(I_top_0_f[18]),
    .Tile_X0Y19_A_I_top_1_t(I_top_1_t[18]),
    .Tile_X0Y19_A_I_top_1_f(I_top_1_f[18]),
    .Tile_X0Y20_A_I_top_0_t(I_top_0_t[19]),
    .Tile_X0Y20_A_I_top_0_f(I_top_0_f[19]),
    .Tile_X0Y20_A_I_top_1_t(I_top_1_t[19]),
    .Tile_X0Y20_A_I_top_1_f(I_top_1_f[19]),
    .Tile_X0Y21_A_I_top_0_t(I_top_0_t[20]),
    .Tile_X0Y21_A_I_top_0_f(I_top_0_f[20]),
    .Tile_X0Y21_A_I_top_1_t(I_top_1_t[20]),
    .Tile_X0Y21_A_I_top_1_f(I_top_1_f[20]),
    .Tile_X0Y22_A_I_top_0_t(I_top_0_t[21]),
    .Tile_X0Y22_A_I_top_0_f(I_top_0_f[21]),
    .Tile_X0Y22_A_I_top_1_t(I_top_1_t[21]),
    .Tile_X0Y22_A_I_top_1_f(I_top_1_f[21]),
    .Tile_X0Y23_A_I_top_0_t(I_top_0_t[22]),
    .Tile_X0Y23_A_I_top_0_f(I_top_0_f[22]),
    .Tile_X0Y23_A_I_top_1_t(I_top_1_t[22]),
    .Tile_X0Y23_A_I_top_1_f(I_top_1_f[22]),
    .Tile_X0Y24_A_I_top_0_t(I_top_0_t[23]),
    .Tile_X0Y24_A_I_top_0_f(I_top_0_f[23]),
    .Tile_X0Y24_A_I_top_1_t(I_top_1_t[23]),
    .Tile_X0Y24_A_I_top_1_f(I_top_1_f[23]),
    .Tile_X0Y25_A_I_top_0_t(I_top_0_t[24]),
    .Tile_X0Y25_A_I_top_0_f(I_top_0_f[24]),
    .Tile_X0Y25_A_I_top_1_t(I_top_1_t[24]),
    .Tile_X0Y25_A_I_top_1_f(I_top_1_f[24]),
    .Tile_X0Y26_A_I_top_0_t(I_top_0_t[25]),
    .Tile_X0Y26_A_I_top_0_f(I_top_0_f[25]),
    .Tile_X0Y26_A_I_top_1_t(I_top_1_t[25]),
    .Tile_X0Y26_A_I_top_1_f(I_top_1_f[25]),
    .Tile_X0Y27_A_I_top_0_t(I_top_0_t[26]),
    .Tile_X0Y27_A_I_top_0_f(I_top_0_f[26]),
    .Tile_X0Y27_A_I_top_1_t(I_top_1_t[26]),
    .Tile_X0Y27_A_I_top_1_f(I_top_1_f[26]),
    .Tile_X0Y28_A_I_top_0_t(I_top_0_t[27]),
    .Tile_X0Y28_A_I_top_0_f(I_top_0_f[27]),
    .Tile_X0Y28_A_I_top_1_t(I_top_1_t[27]),
    .Tile_X0Y28_A_I_top_1_f(I_top_1_f[27]),
    .Tile_X0Y29_A_I_top_0_t(I_top_0_t[28]),
    .Tile_X0Y29_A_I_top_0_f(I_top_0_f[28]),
    .Tile_X0Y29_A_I_top_1_t(I_top_1_t[28]),
    .Tile_X0Y29_A_I_top_1_f(I_top_1_f[28]),
    .Tile_X0Y30_A_I_top_0_t(I_top_0_t[29]),
    .Tile_X0Y30_A_I_top_0_f(I_top_0_f[29]),
    .Tile_X0Y30_A_I_top_1_t(I_top_1_t[29]),
    .Tile_X0Y30_A_I_top_1_f(I_top_1_f[29]),
    .Tile_X0Y31_A_I_top_0_t(I_top_0_t[30]),
    .Tile_X0Y31_A_I_top_0_f(I_top_0_f[30]),
    .Tile_X0Y31_A_I_top_1_t(I_top_1_t[30]),
    .Tile_X0Y31_A_I_top_1_f(I_top_1_f[30]),
    .Tile_X0Y32_A_I_top_0_t(I_top_0_t[31]),
    .Tile_X0Y32_A_I_top_0_f(I_top_0_f[31]),
    .Tile_X0Y32_A_I_top_1_t(I_top_1_t[31]),
    .Tile_X0Y32_A_I_top_1_f(I_top_1_f[31]),
    .Tile_X0Y33_A_I_top_0_t(I_top_0_t[32]),
    .Tile_X0Y33_A_I_top_0_f(I_top_0_f[32]),
    .Tile_X0Y33_A_I_top_1_t(I_top_1_t[32]),
    .Tile_X0Y33_A_I_top_1_f(I_top_1_f[32]),
    .Tile_X0Y34_A_I_top_0_t(I_top_0_t[33]),
    .Tile_X0Y34_A_I_top_0_f(I_top_0_f[33]),
    .Tile_X0Y34_A_I_top_1_t(I_top_1_t[33]),
    .Tile_X0Y34_A_I_top_1_f(I_top_1_f[33]),
    .Tile_X0Y35_A_I_top_0_t(I_top_0_t[34]),
    .Tile_X0Y35_A_I_top_0_f(I_top_0_f[34]),
    .Tile_X0Y35_A_I_top_1_t(I_top_1_t[34]),
    .Tile_X0Y35_A_I_top_1_f(I_top_1_f[34]),
    .Tile_X0Y36_A_I_top_0_t(I_top_0_t[35]),
    .Tile_X0Y36_A_I_top_0_f(I_top_0_f[35]),
    .Tile_X0Y36_A_I_top_1_t(I_top_1_t[35]),
    .Tile_X0Y36_A_I_top_1_f(I_top_1_f[35]),
    .Tile_X0Y37_A_I_top_0_t(I_top_0_t[36]),
    .Tile_X0Y37_A_I_top_0_f(I_top_0_f[36]),
    .Tile_X0Y37_A_I_top_1_t(I_top_1_t[36]),
    .Tile_X0Y37_A_I_top_1_f(I_top_1_f[36]),
    .Tile_X0Y38_A_I_top_0_t(I_top_0_t[37]),
    .Tile_X0Y38_A_I_top_0_f(I_top_0_f[37]),
    .Tile_X0Y38_A_I_top_1_t(I_top_1_t[37]),
    .Tile_X0Y38_A_I_top_1_f(I_top_1_f[37]),
    .Tile_X0Y39_A_I_top_0_t(I_top_0_t[38]),
    .Tile_X0Y39_A_I_top_0_f(I_top_0_f[38]),
    .Tile_X0Y39_A_I_top_1_t(I_top_1_t[38]),
    .Tile_X0Y39_A_I_top_1_f(I_top_1_f[38]),
    .Tile_X0Y40_A_I_top_0_t(I_top_0_t[39]),
    .Tile_X0Y40_A_I_top_0_f(I_top_0_f[39]),
    .Tile_X0Y40_A_I_top_1_t(I_top_1_t[39]),
    .Tile_X0Y40_A_I_top_1_f(I_top_1_f[39]),
    .Tile_X0Y41_A_I_top_0_t(I_top_0_t[40]),
    .Tile_X0Y41_A_I_top_0_f(I_top_0_f[40]),
    .Tile_X0Y41_A_I_top_1_t(I_top_1_t[40]),
    .Tile_X0Y41_A_I_top_1_f(I_top_1_f[40]),
    .Tile_X0Y42_A_I_top_0_t(I_top_0_t[41]),
    .Tile_X0Y42_A_I_top_0_f(I_top_0_f[41]),
    .Tile_X0Y42_A_I_top_1_t(I_top_1_t[41]),
    .Tile_X0Y42_A_I_top_1_f(I_top_1_f[41]),
    .Tile_X0Y43_A_I_top_0_t(I_top_0_t[42]),
    .Tile_X0Y43_A_I_top_0_f(I_top_0_f[42]),
    .Tile_X0Y43_A_I_top_1_t(I_top_1_t[42]),
    .Tile_X0Y43_A_I_top_1_f(I_top_1_f[42]),
    .Tile_X0Y44_A_I_top_0_t(I_top_0_t[43]),
    .Tile_X0Y44_A_I_top_0_f(I_top_0_f[43]),
    .Tile_X0Y44_A_I_top_1_t(I_top_1_t[43]),
    .Tile_X0Y44_A_I_top_1_f(I_top_1_f[43]),
    .Tile_X0Y45_A_I_top_0_t(I_top_0_t[44]),
    .Tile_X0Y45_A_I_top_0_f(I_top_0_f[44]),
    .Tile_X0Y45_A_I_top_1_t(I_top_1_t[44]),
    .Tile_X0Y45_A_I_top_1_f(I_top_1_f[44]),
    .Tile_X0Y46_A_I_top_0_t(I_top_0_t[45]),
    .Tile_X0Y46_A_I_top_0_f(I_top_0_f[45]),
    .Tile_X0Y46_A_I_top_1_t(I_top_1_t[45]),
    .Tile_X0Y46_A_I_top_1_f(I_top_1_f[45]),
    .Tile_X0Y47_A_I_top_0_t(I_top_0_t[46]),
    .Tile_X0Y47_A_I_top_0_f(I_top_0_f[46]),
    .Tile_X0Y47_A_I_top_1_t(I_top_1_t[46]),
    .Tile_X0Y47_A_I_top_1_f(I_top_1_f[46]),
    .Tile_X0Y48_A_I_top_0_t(I_top_0_t[47]),
    .Tile_X0Y48_A_I_top_0_f(I_top_0_f[47]),
    .Tile_X0Y48_A_I_top_1_t(I_top_1_t[47]),
    .Tile_X0Y48_A_I_top_1_f(I_top_1_f[47]),
    .Tile_X0Y49_A_I_top_0_t(I_top_0_t[48]),
    .Tile_X0Y49_A_I_top_0_f(I_top_0_f[48]),
    .Tile_X0Y49_A_I_top_1_t(I_top_1_t[48]),
    .Tile_X0Y49_A_I_top_1_f(I_top_1_f[48]),
    .Tile_X0Y50_A_I_top_0_t(I_top_0_t[49]),
    .Tile_X0Y50_A_I_top_0_f(I_top_0_f[49]),
    .Tile_X0Y50_A_I_top_1_t(I_top_1_t[49]),
    .Tile_X0Y50_A_I_top_1_f(I_top_1_f[49]),
    .Tile_X0Y51_A_I_top_0_t(I_top_0_t[50]),
    .Tile_X0Y51_A_I_top_0_f(I_top_0_f[50]),
    .Tile_X0Y51_A_I_top_1_t(I_top_1_t[50]),
    .Tile_X0Y51_A_I_top_1_f(I_top_1_f[50]),
    .Tile_X0Y52_A_I_top_0_t(I_top_0_t[51]),
    .Tile_X0Y52_A_I_top_0_f(I_top_0_f[51]),
    .Tile_X0Y52_A_I_top_1_t(I_top_1_t[51]),
    .Tile_X0Y52_A_I_top_1_f(I_top_1_f[51]),
    .Tile_X0Y53_A_I_top_0_t(I_top_0_t[52]),
    .Tile_X0Y53_A_I_top_0_f(I_top_0_f[52]),
    .Tile_X0Y53_A_I_top_1_t(I_top_1_t[52]),
    .Tile_X0Y53_A_I_top_1_f(I_top_1_f[52]),
    .Tile_X0Y54_A_I_top_0_t(I_top_0_t[53]),
    .Tile_X0Y54_A_I_top_0_f(I_top_0_f[53]),
    .Tile_X0Y54_A_I_top_1_t(I_top_1_t[53]),
    .Tile_X0Y54_A_I_top_1_f(I_top_1_f[53]),
    .Tile_X0Y55_A_I_top_0_t(I_top_0_t[54]),
    .Tile_X0Y55_A_I_top_0_f(I_top_0_f[54]),
    .Tile_X0Y55_A_I_top_1_t(I_top_1_t[54]),
    .Tile_X0Y55_A_I_top_1_f(I_top_1_f[54]),
    .Tile_X0Y56_A_I_top_0_t(I_top_0_t[55]),
    .Tile_X0Y56_A_I_top_0_f(I_top_0_f[55]),
    .Tile_X0Y56_A_I_top_1_t(I_top_1_t[55]),
    .Tile_X0Y56_A_I_top_1_f(I_top_1_f[55]),
    .Tile_X0Y57_A_I_top_0_t(I_top_0_t[56]),
    .Tile_X0Y57_A_I_top_0_f(I_top_0_f[56]),
    .Tile_X0Y57_A_I_top_1_t(I_top_1_t[56]),
    .Tile_X0Y57_A_I_top_1_f(I_top_1_f[56]),
    .Tile_X0Y58_A_I_top_0_t(I_top_0_t[57]),
    .Tile_X0Y58_A_I_top_0_f(I_top_0_f[57]),
    .Tile_X0Y58_A_I_top_1_t(I_top_1_t[57]),
    .Tile_X0Y58_A_I_top_1_f(I_top_1_f[57]),
    .Tile_X0Y59_A_I_top_0_t(I_top_0_t[58]),
    .Tile_X0Y59_A_I_top_0_f(I_top_0_f[58]),
    .Tile_X0Y59_A_I_top_1_t(I_top_1_t[58]),
    .Tile_X0Y59_A_I_top_1_f(I_top_1_f[58]),
    .Tile_X0Y60_A_I_top_0_t(I_top_0_t[59]),
    .Tile_X0Y60_A_I_top_0_f(I_top_0_f[59]),
    .Tile_X0Y60_A_I_top_1_t(I_top_1_t[59]),
    .Tile_X0Y60_A_I_top_1_f(I_top_1_f[59]),
    .Tile_X0Y1_A_T_top(T_top[0]),
    .Tile_X0Y2_A_T_top(T_top[1]),
    .Tile_X0Y3_A_T_top(T_top[2]),
    .Tile_X0Y4_A_T_top(T_top[3]),
    .Tile_X0Y5_A_T_top(T_top[4]),
    .Tile_X0Y6_A_T_top(T_top[5]),
    .Tile_X0Y7_A_T_top(T_top[6]),
    .Tile_X0Y8_A_T_top(T_top[7]),
    .Tile_X0Y9_A_T_top(T_top[8]),
    .Tile_X0Y10_A_T_top(T_top[9]),
    .Tile_X0Y11_A_T_top(T_top[10]),
    .Tile_X0Y12_A_T_top(T_top[11]),
    .Tile_X0Y13_A_T_top(T_top[12]),
    .Tile_X0Y14_A_T_top(T_top[13]),
    .Tile_X0Y15_A_T_top(T_top[14]),
    .Tile_X0Y16_A_T_top(T_top[15]),
    .Tile_X0Y17_A_T_top(T_top[16]),
    .Tile_X0Y18_A_T_top(T_top[17]),
    .Tile_X0Y19_A_T_top(T_top[18]),
    .Tile_X0Y20_A_T_top(T_top[19]),
    .Tile_X0Y21_A_T_top(T_top[20]),
    .Tile_X0Y22_A_T_top(T_top[21]),
    .Tile_X0Y23_A_T_top(T_top[22]),
    .Tile_X0Y24_A_T_top(T_top[23]),
    .Tile_X0Y25_A_T_top(T_top[24]),
    .Tile_X0Y26_A_T_top(T_top[25]),
    .Tile_X0Y27_A_T_top(T_top[26]),
    .Tile_X0Y28_A_T_top(T_top[27]),
    .Tile_X0Y29_A_T_top(T_top[28]),
    .Tile_X0Y30_A_T_top(T_top[29]),
    .Tile_X0Y31_A_T_top(T_top[30]),
    .Tile_X0Y32_A_T_top(T_top[31]),
    .Tile_X0Y33_A_T_top(T_top[32]),
    .Tile_X0Y34_A_T_top(T_top[33]),
    .Tile_X0Y35_A_T_top(T_top[34]),
    .Tile_X0Y36_A_T_top(T_top[35]),
    .Tile_X0Y37_A_T_top(T_top[36]),
    .Tile_X0Y38_A_T_top(T_top[37]),
    .Tile_X0Y39_A_T_top(T_top[38]),
    .Tile_X0Y40_A_T_top(T_top[39]),
    .Tile_X0Y41_A_T_top(T_top[40]),
    .Tile_X0Y42_A_T_top(T_top[41]),
    .Tile_X0Y43_A_T_top(T_top[42]),
    .Tile_X0Y44_A_T_top(T_top[43]),
    .Tile_X0Y45_A_T_top(T_top[44]),
    .Tile_X0Y46_A_T_top(T_top[45]),
    .Tile_X0Y47_A_T_top(T_top[46]),
    .Tile_X0Y48_A_T_top(T_top[47]),
    .Tile_X0Y49_A_T_top(T_top[48]),
    .Tile_X0Y50_A_T_top(T_top[49]),
    .Tile_X0Y51_A_T_top(T_top[50]),
    .Tile_X0Y52_A_T_top(T_top[51]),
    .Tile_X0Y53_A_T_top(T_top[52]),
    .Tile_X0Y54_A_T_top(T_top[53]),
    .Tile_X0Y55_A_T_top(T_top[54]),
    .Tile_X0Y56_A_T_top(T_top[55]),
    .Tile_X0Y57_A_T_top(T_top[56]),
    .Tile_X0Y58_A_T_top(T_top[57]),
    .Tile_X0Y59_A_T_top(T_top[58]),
    .Tile_X0Y60_A_T_top(T_top[59]),
    .Tile_X0Y1_A_O_top_0_t(O_top_0_t[0]),
    .Tile_X0Y1_A_O_top_0_f(O_top_0_f[0]),
    .Tile_X0Y1_A_O_top_1_t(O_top_1_t[0]),
    .Tile_X0Y1_A_O_top_1_f(O_top_1_f[0]),
    .Tile_X0Y2_A_O_top_0_t(O_top_0_t[1]),
    .Tile_X0Y2_A_O_top_0_f(O_top_0_f[1]),
    .Tile_X0Y2_A_O_top_1_t(O_top_1_t[1]),
    .Tile_X0Y2_A_O_top_1_f(O_top_1_f[1]),
    .Tile_X0Y3_A_O_top_0_t(O_top_0_t[2]),
    .Tile_X0Y3_A_O_top_0_f(O_top_0_f[2]),
    .Tile_X0Y3_A_O_top_1_t(O_top_1_t[2]),
    .Tile_X0Y3_A_O_top_1_f(O_top_1_f[2]),
    .Tile_X0Y4_A_O_top_0_t(O_top_0_t[3]),
    .Tile_X0Y4_A_O_top_0_f(O_top_0_f[3]),
    .Tile_X0Y4_A_O_top_1_t(O_top_1_t[3]),
    .Tile_X0Y4_A_O_top_1_f(O_top_1_f[3]),
    .Tile_X0Y5_A_O_top_0_t(O_top_0_t[4]),
    .Tile_X0Y5_A_O_top_0_f(O_top_0_f[4]),
    .Tile_X0Y5_A_O_top_1_t(O_top_1_t[4]),
    .Tile_X0Y5_A_O_top_1_f(O_top_1_f[4]),
    .Tile_X0Y6_A_O_top_0_t(O_top_0_t[5]),
    .Tile_X0Y6_A_O_top_0_f(O_top_0_f[5]),
    .Tile_X0Y6_A_O_top_1_t(O_top_1_t[5]),
    .Tile_X0Y6_A_O_top_1_f(O_top_1_f[5]),
    .Tile_X0Y7_A_O_top_0_t(O_top_0_t[6]),
    .Tile_X0Y7_A_O_top_0_f(O_top_0_f[6]),
    .Tile_X0Y7_A_O_top_1_t(O_top_1_t[6]),
    .Tile_X0Y7_A_O_top_1_f(O_top_1_f[6]),
    .Tile_X0Y8_A_O_top_0_t(O_top_0_t[7]),
    .Tile_X0Y8_A_O_top_0_f(O_top_0_f[7]),
    .Tile_X0Y8_A_O_top_1_t(O_top_1_t[7]),
    .Tile_X0Y8_A_O_top_1_f(O_top_1_f[7]),
    .Tile_X0Y9_A_O_top_0_t(O_top_0_t[8]),
    .Tile_X0Y9_A_O_top_0_f(O_top_0_f[8]),
    .Tile_X0Y9_A_O_top_1_t(O_top_1_t[8]),
    .Tile_X0Y9_A_O_top_1_f(O_top_1_f[8]),
    .Tile_X0Y10_A_O_top_0_t(O_top_0_t[9]),
    .Tile_X0Y10_A_O_top_0_f(O_top_0_f[9]),
    .Tile_X0Y10_A_O_top_1_t(O_top_1_t[9]),
    .Tile_X0Y10_A_O_top_1_f(O_top_1_f[9]),
    .Tile_X0Y11_A_O_top_0_t(O_top_0_t[10]),
    .Tile_X0Y11_A_O_top_0_f(O_top_0_f[10]),
    .Tile_X0Y11_A_O_top_1_t(O_top_1_t[10]),
    .Tile_X0Y11_A_O_top_1_f(O_top_1_f[10]),
    .Tile_X0Y12_A_O_top_0_t(O_top_0_t[11]),
    .Tile_X0Y12_A_O_top_0_f(O_top_0_f[11]),
    .Tile_X0Y12_A_O_top_1_t(O_top_1_t[11]),
    .Tile_X0Y12_A_O_top_1_f(O_top_1_f[11]),
    .Tile_X0Y13_A_O_top_0_t(O_top_0_t[12]),
    .Tile_X0Y13_A_O_top_0_f(O_top_0_f[12]),
    .Tile_X0Y13_A_O_top_1_t(O_top_1_t[12]),
    .Tile_X0Y13_A_O_top_1_f(O_top_1_f[12]),
    .Tile_X0Y14_A_O_top_0_t(O_top_0_t[13]),
    .Tile_X0Y14_A_O_top_0_f(O_top_0_f[13]),
    .Tile_X0Y14_A_O_top_1_t(O_top_1_t[13]),
    .Tile_X0Y14_A_O_top_1_f(O_top_1_f[13]),
    .Tile_X0Y15_A_O_top_0_t(O_top_0_t[14]),
    .Tile_X0Y15_A_O_top_0_f(O_top_0_f[14]),
    .Tile_X0Y15_A_O_top_1_t(O_top_1_t[14]),
    .Tile_X0Y15_A_O_top_1_f(O_top_1_f[14]),
    .Tile_X0Y16_A_O_top_0_t(O_top_0_t[15]),
    .Tile_X0Y16_A_O_top_0_f(O_top_0_f[15]),
    .Tile_X0Y16_A_O_top_1_t(O_top_1_t[15]),
    .Tile_X0Y16_A_O_top_1_f(O_top_1_f[15]),
    .Tile_X0Y17_A_O_top_0_t(O_top_0_t[16]),
    .Tile_X0Y17_A_O_top_0_f(O_top_0_f[16]),
    .Tile_X0Y17_A_O_top_1_t(O_top_1_t[16]),
    .Tile_X0Y17_A_O_top_1_f(O_top_1_f[16]),
    .Tile_X0Y18_A_O_top_0_t(O_top_0_t[17]),
    .Tile_X0Y18_A_O_top_0_f(O_top_0_f[17]),
    .Tile_X0Y18_A_O_top_1_t(O_top_1_t[17]),
    .Tile_X0Y18_A_O_top_1_f(O_top_1_f[17]),
    .Tile_X0Y19_A_O_top_0_t(O_top_0_t[18]),
    .Tile_X0Y19_A_O_top_0_f(O_top_0_f[18]),
    .Tile_X0Y19_A_O_top_1_t(O_top_1_t[18]),
    .Tile_X0Y19_A_O_top_1_f(O_top_1_f[18]),
    .Tile_X0Y20_A_O_top_0_t(O_top_0_t[19]),
    .Tile_X0Y20_A_O_top_0_f(O_top_0_f[19]),
    .Tile_X0Y20_A_O_top_1_t(O_top_1_t[19]),
    .Tile_X0Y20_A_O_top_1_f(O_top_1_f[19]),
    .Tile_X0Y21_A_O_top_0_t(O_top_0_t[20]),
    .Tile_X0Y21_A_O_top_0_f(O_top_0_f[20]),
    .Tile_X0Y21_A_O_top_1_t(O_top_1_t[20]),
    .Tile_X0Y21_A_O_top_1_f(O_top_1_f[20]),
    .Tile_X0Y22_A_O_top_0_t(O_top_0_t[21]),
    .Tile_X0Y22_A_O_top_0_f(O_top_0_f[21]),
    .Tile_X0Y22_A_O_top_1_t(O_top_1_t[21]),
    .Tile_X0Y22_A_O_top_1_f(O_top_1_f[21]),
    .Tile_X0Y23_A_O_top_0_t(O_top_0_t[22]),
    .Tile_X0Y23_A_O_top_0_f(O_top_0_f[22]),
    .Tile_X0Y23_A_O_top_1_t(O_top_1_t[22]),
    .Tile_X0Y23_A_O_top_1_f(O_top_1_f[22]),
    .Tile_X0Y24_A_O_top_0_t(O_top_0_t[23]),
    .Tile_X0Y24_A_O_top_0_f(O_top_0_f[23]),
    .Tile_X0Y24_A_O_top_1_t(O_top_1_t[23]),
    .Tile_X0Y24_A_O_top_1_f(O_top_1_f[23]),
    .Tile_X0Y25_A_O_top_0_t(O_top_0_t[24]),
    .Tile_X0Y25_A_O_top_0_f(O_top_0_f[24]),
    .Tile_X0Y25_A_O_top_1_t(O_top_1_t[24]),
    .Tile_X0Y25_A_O_top_1_f(O_top_1_f[24]),
    .Tile_X0Y26_A_O_top_0_t(O_top_0_t[25]),
    .Tile_X0Y26_A_O_top_0_f(O_top_0_f[25]),
    .Tile_X0Y26_A_O_top_1_t(O_top_1_t[25]),
    .Tile_X0Y26_A_O_top_1_f(O_top_1_f[25]),
    .Tile_X0Y27_A_O_top_0_t(O_top_0_t[26]),
    .Tile_X0Y27_A_O_top_0_f(O_top_0_f[26]),
    .Tile_X0Y27_A_O_top_1_t(O_top_1_t[26]),
    .Tile_X0Y27_A_O_top_1_f(O_top_1_f[26]),
    .Tile_X0Y28_A_O_top_0_t(O_top_0_t[27]),
    .Tile_X0Y28_A_O_top_0_f(O_top_0_f[27]),
    .Tile_X0Y28_A_O_top_1_t(O_top_1_t[27]),
    .Tile_X0Y28_A_O_top_1_f(O_top_1_f[27]),
    .Tile_X0Y29_A_O_top_0_t(O_top_0_t[28]),
    .Tile_X0Y29_A_O_top_0_f(O_top_0_f[28]),
    .Tile_X0Y29_A_O_top_1_t(O_top_1_t[28]),
    .Tile_X0Y29_A_O_top_1_f(O_top_1_f[28]),
    .Tile_X0Y30_A_O_top_0_t(O_top_0_t[29]),
    .Tile_X0Y30_A_O_top_0_f(O_top_0_f[29]),
    .Tile_X0Y30_A_O_top_1_t(O_top_1_t[29]),
    .Tile_X0Y30_A_O_top_1_f(O_top_1_f[29]),
    .Tile_X0Y31_A_O_top_0_t(O_top_0_t[30]),
    .Tile_X0Y31_A_O_top_0_f(O_top_0_f[30]),
    .Tile_X0Y31_A_O_top_1_t(O_top_1_t[30]),
    .Tile_X0Y31_A_O_top_1_f(O_top_1_f[30]),
    .Tile_X0Y32_A_O_top_0_t(O_top_0_t[31]),
    .Tile_X0Y32_A_O_top_0_f(O_top_0_f[31]),
    .Tile_X0Y32_A_O_top_1_t(O_top_1_t[31]),
    .Tile_X0Y32_A_O_top_1_f(O_top_1_f[31]),
    .Tile_X0Y33_A_O_top_0_t(O_top_0_t[32]),
    .Tile_X0Y33_A_O_top_0_f(O_top_0_f[32]),
    .Tile_X0Y33_A_O_top_1_t(O_top_1_t[32]),
    .Tile_X0Y33_A_O_top_1_f(O_top_1_f[32]),
    .Tile_X0Y34_A_O_top_0_t(O_top_0_t[33]),
    .Tile_X0Y34_A_O_top_0_f(O_top_0_f[33]),
    .Tile_X0Y34_A_O_top_1_t(O_top_1_t[33]),
    .Tile_X0Y34_A_O_top_1_f(O_top_1_f[33]),
    .Tile_X0Y35_A_O_top_0_t(O_top_0_t[34]),
    .Tile_X0Y35_A_O_top_0_f(O_top_0_f[34]),
    .Tile_X0Y35_A_O_top_1_t(O_top_1_t[34]),
    .Tile_X0Y35_A_O_top_1_f(O_top_1_f[34]),
    .Tile_X0Y36_A_O_top_0_t(O_top_0_t[35]),
    .Tile_X0Y36_A_O_top_0_f(O_top_0_f[35]),
    .Tile_X0Y36_A_O_top_1_t(O_top_1_t[35]),
    .Tile_X0Y36_A_O_top_1_f(O_top_1_f[35]),
    .Tile_X0Y37_A_O_top_0_t(O_top_0_t[36]),
    .Tile_X0Y37_A_O_top_0_f(O_top_0_f[36]),
    .Tile_X0Y37_A_O_top_1_t(O_top_1_t[36]),
    .Tile_X0Y37_A_O_top_1_f(O_top_1_f[36]),
    .Tile_X0Y38_A_O_top_0_t(O_top_0_t[37]),
    .Tile_X0Y38_A_O_top_0_f(O_top_0_f[37]),
    .Tile_X0Y38_A_O_top_1_t(O_top_1_t[37]),
    .Tile_X0Y38_A_O_top_1_f(O_top_1_f[37]),
    .Tile_X0Y39_A_O_top_0_t(O_top_0_t[38]),
    .Tile_X0Y39_A_O_top_0_f(O_top_0_f[38]),
    .Tile_X0Y39_A_O_top_1_t(O_top_1_t[38]),
    .Tile_X0Y39_A_O_top_1_f(O_top_1_f[38]),
    .Tile_X0Y40_A_O_top_0_t(O_top_0_t[39]),
    .Tile_X0Y40_A_O_top_0_f(O_top_0_f[39]),
    .Tile_X0Y40_A_O_top_1_t(O_top_1_t[39]),
    .Tile_X0Y40_A_O_top_1_f(O_top_1_f[39]),
    .Tile_X0Y41_A_O_top_0_t(O_top_0_t[40]),
    .Tile_X0Y41_A_O_top_0_f(O_top_0_f[40]),
    .Tile_X0Y41_A_O_top_1_t(O_top_1_t[40]),
    .Tile_X0Y41_A_O_top_1_f(O_top_1_f[40]),
    .Tile_X0Y42_A_O_top_0_t(O_top_0_t[41]),
    .Tile_X0Y42_A_O_top_0_f(O_top_0_f[41]),
    .Tile_X0Y42_A_O_top_1_t(O_top_1_t[41]),
    .Tile_X0Y42_A_O_top_1_f(O_top_1_f[41]),
    .Tile_X0Y43_A_O_top_0_t(O_top_0_t[42]),
    .Tile_X0Y43_A_O_top_0_f(O_top_0_f[42]),
    .Tile_X0Y43_A_O_top_1_t(O_top_1_t[42]),
    .Tile_X0Y43_A_O_top_1_f(O_top_1_f[42]),
    .Tile_X0Y44_A_O_top_0_t(O_top_0_t[43]),
    .Tile_X0Y44_A_O_top_0_f(O_top_0_f[43]),
    .Tile_X0Y44_A_O_top_1_t(O_top_1_t[43]),
    .Tile_X0Y44_A_O_top_1_f(O_top_1_f[43]),
    .Tile_X0Y45_A_O_top_0_t(O_top_0_t[44]),
    .Tile_X0Y45_A_O_top_0_f(O_top_0_f[44]),
    .Tile_X0Y45_A_O_top_1_t(O_top_1_t[44]),
    .Tile_X0Y45_A_O_top_1_f(O_top_1_f[44]),
    .Tile_X0Y46_A_O_top_0_t(O_top_0_t[45]),
    .Tile_X0Y46_A_O_top_0_f(O_top_0_f[45]),
    .Tile_X0Y46_A_O_top_1_t(O_top_1_t[45]),
    .Tile_X0Y46_A_O_top_1_f(O_top_1_f[45]),
    .Tile_X0Y47_A_O_top_0_t(O_top_0_t[46]),
    .Tile_X0Y47_A_O_top_0_f(O_top_0_f[46]),
    .Tile_X0Y47_A_O_top_1_t(O_top_1_t[46]),
    .Tile_X0Y47_A_O_top_1_f(O_top_1_f[46]),
    .Tile_X0Y48_A_O_top_0_t(O_top_0_t[47]),
    .Tile_X0Y48_A_O_top_0_f(O_top_0_f[47]),
    .Tile_X0Y48_A_O_top_1_t(O_top_1_t[47]),
    .Tile_X0Y48_A_O_top_1_f(O_top_1_f[47]),
    .Tile_X0Y49_A_O_top_0_t(O_top_0_t[48]),
    .Tile_X0Y49_A_O_top_0_f(O_top_0_f[48]),
    .Tile_X0Y49_A_O_top_1_t(O_top_1_t[48]),
    .Tile_X0Y49_A_O_top_1_f(O_top_1_f[48]),
    .Tile_X0Y50_A_O_top_0_t(O_top_0_t[49]),
    .Tile_X0Y50_A_O_top_0_f(O_top_0_f[49]),
    .Tile_X0Y50_A_O_top_1_t(O_top_1_t[49]),
    .Tile_X0Y50_A_O_top_1_f(O_top_1_f[49]),
    .Tile_X0Y51_A_O_top_0_t(O_top_0_t[50]),
    .Tile_X0Y51_A_O_top_0_f(O_top_0_f[50]),
    .Tile_X0Y51_A_O_top_1_t(O_top_1_t[50]),
    .Tile_X0Y51_A_O_top_1_f(O_top_1_f[50]),
    .Tile_X0Y52_A_O_top_0_t(O_top_0_t[51]),
    .Tile_X0Y52_A_O_top_0_f(O_top_0_f[51]),
    .Tile_X0Y52_A_O_top_1_t(O_top_1_t[51]),
    .Tile_X0Y52_A_O_top_1_f(O_top_1_f[51]),
    .Tile_X0Y53_A_O_top_0_t(O_top_0_t[52]),
    .Tile_X0Y53_A_O_top_0_f(O_top_0_f[52]),
    .Tile_X0Y53_A_O_top_1_t(O_top_1_t[52]),
    .Tile_X0Y53_A_O_top_1_f(O_top_1_f[52]),
    .Tile_X0Y54_A_O_top_0_t(O_top_0_t[53]),
    .Tile_X0Y54_A_O_top_0_f(O_top_0_f[53]),
    .Tile_X0Y54_A_O_top_1_t(O_top_1_t[53]),
    .Tile_X0Y54_A_O_top_1_f(O_top_1_f[53]),
    .Tile_X0Y55_A_O_top_0_t(O_top_0_t[54]),
    .Tile_X0Y55_A_O_top_0_f(O_top_0_f[54]),
    .Tile_X0Y55_A_O_top_1_t(O_top_1_t[54]),
    .Tile_X0Y55_A_O_top_1_f(O_top_1_f[54]),
    .Tile_X0Y56_A_O_top_0_t(O_top_0_t[55]),
    .Tile_X0Y56_A_O_top_0_f(O_top_0_f[55]),
    .Tile_X0Y56_A_O_top_1_t(O_top_1_t[55]),
    .Tile_X0Y56_A_O_top_1_f(O_top_1_f[55]),
    .Tile_X0Y57_A_O_top_0_t(O_top_0_t[56]),
    .Tile_X0Y57_A_O_top_0_f(O_top_0_f[56]),
    .Tile_X0Y57_A_O_top_1_t(O_top_1_t[56]),
    .Tile_X0Y57_A_O_top_1_f(O_top_1_f[56]),
    .Tile_X0Y58_A_O_top_0_t(O_top_0_t[57]),
    .Tile_X0Y58_A_O_top_0_f(O_top_0_f[57]),
    .Tile_X0Y58_A_O_top_1_t(O_top_1_t[57]),
    .Tile_X0Y58_A_O_top_1_f(O_top_1_f[57]),
    .Tile_X0Y59_A_O_top_0_t(O_top_0_t[58]),
    .Tile_X0Y59_A_O_top_0_f(O_top_0_f[58]),
    .Tile_X0Y59_A_O_top_1_t(O_top_1_t[58]),
    .Tile_X0Y59_A_O_top_1_f(O_top_1_f[58]),
    .Tile_X0Y60_A_O_top_0_t(O_top_0_t[59]),
    .Tile_X0Y60_A_O_top_0_f(O_top_0_f[59]),
    .Tile_X0Y60_A_O_top_1_t(O_top_1_t[59]),
    .Tile_X0Y60_A_O_top_1_f(O_top_1_f[59]),
    .Tile_X38Y1_A_I_top_0_t(ctrl_I_top_0_t[0]),
    .Tile_X38Y1_A_I_top_0_f(ctrl_I_top_0_f[0]),
    .Tile_X38Y1_A_T_top(ctrl_T_top[0]),
    .Tile_X38Y1_A_O_top_0_t(ctrl_O_top_0_t[0]),
    .Tile_X38Y1_A_O_top_0_f(ctrl_O_top_0_f[0]),
    .Tile_X38Y2_A_I_top_0_t(ctrl_I_top_0_t[1]),
    .Tile_X38Y2_A_I_top_0_f(ctrl_I_top_0_f[1]),
    .Tile_X38Y2_A_T_top(ctrl_T_top[1]),
    .Tile_X38Y2_A_O_top_0_t(ctrl_O_top_0_t[1]),
    .Tile_X38Y2_A_O_top_0_f(ctrl_O_top_0_f[1]),
    .Tile_X38Y3_A_I_top_0_t(ctrl_I_top_0_t[2]),
    .Tile_X38Y3_A_I_top_0_f(ctrl_I_top_0_f[2]),
    .Tile_X38Y3_A_T_top(ctrl_T_top[2]),
    .Tile_X38Y3_A_O_top_0_t(ctrl_O_top_0_t[2]),
    .Tile_X38Y3_A_O_top_0_f(ctrl_O_top_0_f[2]),
    .Tile_X38Y4_A_I_top_0_t(ctrl_I_top_0_t[3]),
    .Tile_X38Y4_A_I_top_0_f(ctrl_I_top_0_f[3]),
    .Tile_X38Y4_A_T_top(ctrl_T_top[3]),
    .Tile_X38Y4_A_O_top_0_t(ctrl_O_top_0_t[3]),
    .Tile_X38Y4_A_O_top_0_f(ctrl_O_top_0_f[3]),
    .Tile_X38Y5_A_I_top_0_t(ctrl_I_top_0_t[4]),
    .Tile_X38Y5_A_I_top_0_f(ctrl_I_top_0_f[4]),
    .Tile_X38Y5_A_T_top(ctrl_T_top[4]),
    .Tile_X38Y5_A_O_top_0_t(ctrl_O_top_0_t[4]),
    .Tile_X38Y5_A_O_top_0_f(ctrl_O_top_0_f[4]),
    .Tile_X38Y6_A_I_top_0_t(ctrl_I_top_0_t[5]),
    .Tile_X38Y6_A_I_top_0_f(ctrl_I_top_0_f[5]),
    .Tile_X38Y6_A_T_top(ctrl_T_top[5]),
    .Tile_X38Y6_A_O_top_0_t(ctrl_O_top_0_t[5]),
    .Tile_X38Y6_A_O_top_0_f(ctrl_O_top_0_f[5]),
    .Tile_X38Y7_A_I_top_0_t(ctrl_I_top_0_t[6]),
    .Tile_X38Y7_A_I_top_0_f(ctrl_I_top_0_f[6]),
    .Tile_X38Y7_A_T_top(ctrl_T_top[6]),
    .Tile_X38Y7_A_O_top_0_t(ctrl_O_top_0_t[6]),
    .Tile_X38Y7_A_O_top_0_f(ctrl_O_top_0_f[6]),
    .Tile_X38Y8_A_I_top_0_t(ctrl_I_top_0_t[7]),
    .Tile_X38Y8_A_I_top_0_f(ctrl_I_top_0_f[7]),
    .Tile_X38Y8_A_T_top(ctrl_T_top[7]),
    .Tile_X38Y8_A_O_top_0_t(ctrl_O_top_0_t[7]),
    .Tile_X38Y8_A_O_top_0_f(ctrl_O_top_0_f[7]),
    .Tile_X38Y9_A_I_top_0_t(ctrl_I_top_0_t[8]),
    .Tile_X38Y9_A_I_top_0_f(ctrl_I_top_0_f[8]),
    .Tile_X38Y9_A_T_top(ctrl_T_top[8]),
    .Tile_X38Y9_A_O_top_0_t(ctrl_O_top_0_t[8]),
    .Tile_X38Y9_A_O_top_0_f(ctrl_O_top_0_f[8]),
    .Tile_X38Y10_A_I_top_0_t(ctrl_I_top_0_t[9]),
    .Tile_X38Y10_A_I_top_0_f(ctrl_I_top_0_f[9]),
    .Tile_X38Y10_A_T_top(ctrl_T_top[9]),
    .Tile_X38Y10_A_O_top_0_t(ctrl_O_top_0_t[9]),
    .Tile_X38Y10_A_O_top_0_f(ctrl_O_top_0_f[9]),
    .Tile_X38Y11_A_I_top_0_t(ctrl_I_top_0_t[10]),
    .Tile_X38Y11_A_I_top_0_f(ctrl_I_top_0_f[10]),
    .Tile_X38Y11_A_T_top(ctrl_T_top[10]),
    .Tile_X38Y11_A_O_top_0_t(ctrl_O_top_0_t[10]),
    .Tile_X38Y11_A_O_top_0_f(ctrl_O_top_0_f[10]),
    .Tile_X38Y12_A_I_top_0_t(ctrl_I_top_0_t[11]),
    .Tile_X38Y12_A_I_top_0_f(ctrl_I_top_0_f[11]),
    .Tile_X38Y12_A_T_top(ctrl_T_top[11]),
    .Tile_X38Y12_A_O_top_0_t(ctrl_O_top_0_t[11]),
    .Tile_X38Y12_A_O_top_0_f(ctrl_O_top_0_f[11]),
    .Tile_X38Y13_A_I_top_0_t(ctrl_I_top_0_t[12]),
    .Tile_X38Y13_A_I_top_0_f(ctrl_I_top_0_f[12]),
    .Tile_X38Y13_A_T_top(ctrl_T_top[12]),
    .Tile_X38Y13_A_O_top_0_t(ctrl_O_top_0_t[12]),
    .Tile_X38Y13_A_O_top_0_f(ctrl_O_top_0_f[12]),
    .Tile_X38Y14_A_I_top_0_t(ctrl_I_top_0_t[13]),
    .Tile_X38Y14_A_I_top_0_f(ctrl_I_top_0_f[13]),
    .Tile_X38Y14_A_T_top(ctrl_T_top[13]),
    .Tile_X38Y14_A_O_top_0_t(ctrl_O_top_0_t[13]),
    .Tile_X38Y14_A_O_top_0_f(ctrl_O_top_0_f[13]),
    .Tile_X38Y15_A_I_top_0_t(ctrl_I_top_0_t[14]),
    .Tile_X38Y15_A_I_top_0_f(ctrl_I_top_0_f[14]),
    .Tile_X38Y15_A_T_top(ctrl_T_top[14]),
    .Tile_X38Y15_A_O_top_0_t(ctrl_O_top_0_t[14]),
    .Tile_X38Y15_A_O_top_0_f(ctrl_O_top_0_f[14]),
    .Tile_X38Y16_A_I_top_0_t(ctrl_I_top_0_t[15]),
    .Tile_X38Y16_A_I_top_0_f(ctrl_I_top_0_f[15]),
    .Tile_X38Y16_A_T_top(ctrl_T_top[15]),
    .Tile_X38Y16_A_O_top_0_t(ctrl_O_top_0_t[15]),
    .Tile_X38Y16_A_O_top_0_f(ctrl_O_top_0_f[15]),
    .Tile_X38Y17_A_I_top_0_t(ctrl_I_top_0_t[16]),
    .Tile_X38Y17_A_I_top_0_f(ctrl_I_top_0_f[16]),
    .Tile_X38Y17_A_T_top(ctrl_T_top[16]),
    .Tile_X38Y17_A_O_top_0_t(ctrl_O_top_0_t[16]),
    .Tile_X38Y17_A_O_top_0_f(ctrl_O_top_0_f[16]),
    .Tile_X38Y18_A_I_top_0_t(ctrl_I_top_0_t[17]),
    .Tile_X38Y18_A_I_top_0_f(ctrl_I_top_0_f[17]),
    .Tile_X38Y18_A_T_top(ctrl_T_top[17]),
    .Tile_X38Y18_A_O_top_0_t(ctrl_O_top_0_t[17]),
    .Tile_X38Y18_A_O_top_0_f(ctrl_O_top_0_f[17]),
    .Tile_X38Y19_A_I_top_0_t(ctrl_I_top_0_t[18]),
    .Tile_X38Y19_A_I_top_0_f(ctrl_I_top_0_f[18]),
    .Tile_X38Y19_A_T_top(ctrl_T_top[18]),
    .Tile_X38Y19_A_O_top_0_t(ctrl_O_top_0_t[18]),
    .Tile_X38Y19_A_O_top_0_f(ctrl_O_top_0_f[18]),
    .Tile_X38Y20_A_I_top_0_t(ctrl_I_top_0_t[19]),
    .Tile_X38Y20_A_I_top_0_f(ctrl_I_top_0_f[19]),
    .Tile_X38Y20_A_T_top(ctrl_T_top[19]),
    .Tile_X38Y20_A_O_top_0_t(ctrl_O_top_0_t[19]),
    .Tile_X38Y20_A_O_top_0_f(ctrl_O_top_0_f[19]),
    .Tile_X38Y21_A_I_top_0_t(ctrl_I_top_0_t[20]),
    .Tile_X38Y21_A_I_top_0_f(ctrl_I_top_0_f[20]),
    .Tile_X38Y21_A_T_top(ctrl_T_top[20]),
    .Tile_X38Y21_A_O_top_0_t(ctrl_O_top_0_t[20]),
    .Tile_X38Y21_A_O_top_0_f(ctrl_O_top_0_f[20]),
    .Tile_X38Y22_A_I_top_0_t(ctrl_I_top_0_t[21]),
    .Tile_X38Y22_A_I_top_0_f(ctrl_I_top_0_f[21]),
    .Tile_X38Y22_A_T_top(ctrl_T_top[21]),
    .Tile_X38Y22_A_O_top_0_t(ctrl_O_top_0_t[21]),
    .Tile_X38Y22_A_O_top_0_f(ctrl_O_top_0_f[21]),
    .Tile_X38Y23_A_I_top_0_t(ctrl_I_top_0_t[22]),
    .Tile_X38Y23_A_I_top_0_f(ctrl_I_top_0_f[22]),
    .Tile_X38Y23_A_T_top(ctrl_T_top[22]),
    .Tile_X38Y23_A_O_top_0_t(ctrl_O_top_0_t[22]),
    .Tile_X38Y23_A_O_top_0_f(ctrl_O_top_0_f[22]),
    .Tile_X38Y24_A_I_top_0_t(ctrl_I_top_0_t[23]),
    .Tile_X38Y24_A_I_top_0_f(ctrl_I_top_0_f[23]),
    .Tile_X38Y24_A_T_top(ctrl_T_top[23]),
    .Tile_X38Y24_A_O_top_0_t(ctrl_O_top_0_t[23]),
    .Tile_X38Y24_A_O_top_0_f(ctrl_O_top_0_f[23]),
    .Tile_X38Y25_A_I_top_0_t(ctrl_I_top_0_t[24]),
    .Tile_X38Y25_A_I_top_0_f(ctrl_I_top_0_f[24]),
    .Tile_X38Y25_A_T_top(ctrl_T_top[24]),
    .Tile_X38Y25_A_O_top_0_t(ctrl_O_top_0_t[24]),
    .Tile_X38Y25_A_O_top_0_f(ctrl_O_top_0_f[24]),
    .Tile_X38Y26_A_I_top_0_t(ctrl_I_top_0_t[25]),
    .Tile_X38Y26_A_I_top_0_f(ctrl_I_top_0_f[25]),
    .Tile_X38Y26_A_T_top(ctrl_T_top[25]),
    .Tile_X38Y26_A_O_top_0_t(ctrl_O_top_0_t[25]),
    .Tile_X38Y26_A_O_top_0_f(ctrl_O_top_0_f[25]),
    .Tile_X38Y27_A_I_top_0_t(ctrl_I_top_0_t[26]),
    .Tile_X38Y27_A_I_top_0_f(ctrl_I_top_0_f[26]),
    .Tile_X38Y27_A_T_top(ctrl_T_top[26]),
    .Tile_X38Y27_A_O_top_0_t(ctrl_O_top_0_t[26]),
    .Tile_X38Y27_A_O_top_0_f(ctrl_O_top_0_f[26]),
    .Tile_X38Y28_A_I_top_0_t(ctrl_I_top_0_t[27]),
    .Tile_X38Y28_A_I_top_0_f(ctrl_I_top_0_f[27]),
    .Tile_X38Y28_A_T_top(ctrl_T_top[27]),
    .Tile_X38Y28_A_O_top_0_t(ctrl_O_top_0_t[27]),
    .Tile_X38Y28_A_O_top_0_f(ctrl_O_top_0_f[27]),
    .Tile_X38Y29_A_I_top_0_t(ctrl_I_top_0_t[28]),
    .Tile_X38Y29_A_I_top_0_f(ctrl_I_top_0_f[28]),
    .Tile_X38Y29_A_T_top(ctrl_T_top[28]),
    .Tile_X38Y29_A_O_top_0_t(ctrl_O_top_0_t[28]),
    .Tile_X38Y29_A_O_top_0_f(ctrl_O_top_0_f[28]),
    .Tile_X38Y30_A_I_top_0_t(ctrl_I_top_0_t[29]),
    .Tile_X38Y30_A_I_top_0_f(ctrl_I_top_0_f[29]),
    .Tile_X38Y30_A_T_top(ctrl_T_top[29]),
    .Tile_X38Y30_A_O_top_0_t(ctrl_O_top_0_t[29]),
    .Tile_X38Y30_A_O_top_0_f(ctrl_O_top_0_f[29]),
    .Tile_X38Y31_A_I_top_0_t(ctrl_I_top_0_t[30]),
    .Tile_X38Y31_A_I_top_0_f(ctrl_I_top_0_f[30]),
    .Tile_X38Y31_A_T_top(ctrl_T_top[30]),
    .Tile_X38Y31_A_O_top_0_t(ctrl_O_top_0_t[30]),
    .Tile_X38Y31_A_O_top_0_f(ctrl_O_top_0_f[30]),
    .Tile_X38Y32_A_I_top_0_t(ctrl_I_top_0_t[31]),
    .Tile_X38Y32_A_I_top_0_f(ctrl_I_top_0_f[31]),
    .Tile_X38Y32_A_T_top(ctrl_T_top[31]),
    .Tile_X38Y32_A_O_top_0_t(ctrl_O_top_0_t[31]),
    .Tile_X38Y32_A_O_top_0_f(ctrl_O_top_0_f[31]),
    .Tile_X38Y33_A_I_top_0_t(ctrl_I_top_0_t[32]),
    .Tile_X38Y33_A_I_top_0_f(ctrl_I_top_0_f[32]),
    .Tile_X38Y33_A_T_top(ctrl_T_top[32]),
    .Tile_X38Y33_A_O_top_0_t(ctrl_O_top_0_t[32]),
    .Tile_X38Y33_A_O_top_0_f(ctrl_O_top_0_f[32]),
    .Tile_X38Y34_A_I_top_0_t(ctrl_I_top_0_t[33]),
    .Tile_X38Y34_A_I_top_0_f(ctrl_I_top_0_f[33]),
    .Tile_X38Y34_A_T_top(ctrl_T_top[33]),
    .Tile_X38Y34_A_O_top_0_t(ctrl_O_top_0_t[33]),
    .Tile_X38Y34_A_O_top_0_f(ctrl_O_top_0_f[33]),
    .Tile_X38Y35_A_I_top_0_t(ctrl_I_top_0_t[34]),
    .Tile_X38Y35_A_I_top_0_f(ctrl_I_top_0_f[34]),
    .Tile_X38Y35_A_T_top(ctrl_T_top[34]),
    .Tile_X38Y35_A_O_top_0_t(ctrl_O_top_0_t[34]),
    .Tile_X38Y35_A_O_top_0_f(ctrl_O_top_0_f[34]),
    .Tile_X38Y36_A_I_top_0_t(ctrl_I_top_0_t[35]),
    .Tile_X38Y36_A_I_top_0_f(ctrl_I_top_0_f[35]),
    .Tile_X38Y36_A_T_top(ctrl_T_top[35]),
    .Tile_X38Y36_A_O_top_0_t(ctrl_O_top_0_t[35]),
    .Tile_X38Y36_A_O_top_0_f(ctrl_O_top_0_f[35]),
    .Tile_X38Y37_A_I_top_0_t(ctrl_I_top_0_t[36]),
    .Tile_X38Y37_A_I_top_0_f(ctrl_I_top_0_f[36]),
    .Tile_X38Y37_A_T_top(ctrl_T_top[36]),
    .Tile_X38Y37_A_O_top_0_t(ctrl_O_top_0_t[36]),
    .Tile_X38Y37_A_O_top_0_f(ctrl_O_top_0_f[36]),
    .Tile_X38Y38_A_I_top_0_t(ctrl_I_top_0_t[37]),
    .Tile_X38Y38_A_I_top_0_f(ctrl_I_top_0_f[37]),
    .Tile_X38Y38_A_T_top(ctrl_T_top[37]),
    .Tile_X38Y38_A_O_top_0_t(ctrl_O_top_0_t[37]),
    .Tile_X38Y38_A_O_top_0_f(ctrl_O_top_0_f[37]),
    .Tile_X38Y39_A_I_top_0_t(ctrl_I_top_0_t[38]),
    .Tile_X38Y39_A_I_top_0_f(ctrl_I_top_0_f[38]),
    .Tile_X38Y39_A_T_top(ctrl_T_top[38]),
    .Tile_X38Y39_A_O_top_0_t(ctrl_O_top_0_t[38]),
    .Tile_X38Y39_A_O_top_0_f(ctrl_O_top_0_f[38]),
    .Tile_X38Y40_A_I_top_0_t(ctrl_I_top_0_t[39]),
    .Tile_X38Y40_A_I_top_0_f(ctrl_I_top_0_f[39]),
    .Tile_X38Y40_A_T_top(ctrl_T_top[39]),
    .Tile_X38Y40_A_O_top_0_t(ctrl_O_top_0_t[39]),
    .Tile_X38Y40_A_O_top_0_f(ctrl_O_top_0_f[39]),
    .Tile_X38Y41_A_I_top_0_t(ctrl_I_top_0_t[40]),
    .Tile_X38Y41_A_I_top_0_f(ctrl_I_top_0_f[40]),
    .Tile_X38Y41_A_T_top(ctrl_T_top[40]),
    .Tile_X38Y41_A_O_top_0_t(ctrl_O_top_0_t[40]),
    .Tile_X38Y41_A_O_top_0_f(ctrl_O_top_0_f[40]),
    .Tile_X38Y42_A_I_top_0_t(ctrl_I_top_0_t[41]),
    .Tile_X38Y42_A_I_top_0_f(ctrl_I_top_0_f[41]),
    .Tile_X38Y42_A_T_top(ctrl_T_top[41]),
    .Tile_X38Y42_A_O_top_0_t(ctrl_O_top_0_t[41]),
    .Tile_X38Y42_A_O_top_0_f(ctrl_O_top_0_f[41]),
    .Tile_X38Y43_A_I_top_0_t(ctrl_I_top_0_t[42]),
    .Tile_X38Y43_A_I_top_0_f(ctrl_I_top_0_f[42]),
    .Tile_X38Y43_A_T_top(ctrl_T_top[42]),
    .Tile_X38Y43_A_O_top_0_t(ctrl_O_top_0_t[42]),
    .Tile_X38Y43_A_O_top_0_f(ctrl_O_top_0_f[42]),
    .Tile_X38Y44_A_I_top_0_t(ctrl_I_top_0_t[43]),
    .Tile_X38Y44_A_I_top_0_f(ctrl_I_top_0_f[43]),
    .Tile_X38Y44_A_T_top(ctrl_T_top[43]),
    .Tile_X38Y44_A_O_top_0_t(ctrl_O_top_0_t[43]),
    .Tile_X38Y44_A_O_top_0_f(ctrl_O_top_0_f[43]),
    .Tile_X38Y45_A_I_top_0_t(ctrl_I_top_0_t[44]),
    .Tile_X38Y45_A_I_top_0_f(ctrl_I_top_0_f[44]),
    .Tile_X38Y45_A_T_top(ctrl_T_top[44]),
    .Tile_X38Y45_A_O_top_0_t(ctrl_O_top_0_t[44]),
    .Tile_X38Y45_A_O_top_0_f(ctrl_O_top_0_f[44]),
    .Tile_X38Y46_A_I_top_0_t(ctrl_I_top_0_t[45]),
    .Tile_X38Y46_A_I_top_0_f(ctrl_I_top_0_f[45]),
    .Tile_X38Y46_A_T_top(ctrl_T_top[45]),
    .Tile_X38Y46_A_O_top_0_t(ctrl_O_top_0_t[45]),
    .Tile_X38Y46_A_O_top_0_f(ctrl_O_top_0_f[45]),
    .Tile_X38Y47_A_I_top_0_t(ctrl_I_top_0_t[46]),
    .Tile_X38Y47_A_I_top_0_f(ctrl_I_top_0_f[46]),
    .Tile_X38Y47_A_T_top(ctrl_T_top[46]),
    .Tile_X38Y47_A_O_top_0_t(ctrl_O_top_0_t[46]),
    .Tile_X38Y47_A_O_top_0_f(ctrl_O_top_0_f[46]),
    .Tile_X38Y48_A_I_top_0_t(ctrl_I_top_0_t[47]),
    .Tile_X38Y48_A_I_top_0_f(ctrl_I_top_0_f[47]),
    .Tile_X38Y48_A_T_top(ctrl_T_top[47]),
    .Tile_X38Y48_A_O_top_0_t(ctrl_O_top_0_t[47]),
    .Tile_X38Y48_A_O_top_0_f(ctrl_O_top_0_f[47]),
    .Tile_X38Y49_A_I_top_0_t(ctrl_I_top_0_t[48]),
    .Tile_X38Y49_A_I_top_0_f(ctrl_I_top_0_f[48]),
    .Tile_X38Y49_A_T_top(ctrl_T_top[48]),
    .Tile_X38Y49_A_O_top_0_t(ctrl_O_top_0_t[48]),
    .Tile_X38Y49_A_O_top_0_f(ctrl_O_top_0_f[48]),
    .Tile_X38Y50_A_I_top_0_t(ctrl_I_top_0_t[49]),
    .Tile_X38Y50_A_I_top_0_f(ctrl_I_top_0_f[49]),
    .Tile_X38Y50_A_T_top(ctrl_T_top[49]),
    .Tile_X38Y50_A_O_top_0_t(ctrl_O_top_0_t[49]),
    .Tile_X38Y50_A_O_top_0_f(ctrl_O_top_0_f[49]),
    .Tile_X38Y51_A_I_top_0_t(ctrl_I_top_0_t[50]),
    .Tile_X38Y51_A_I_top_0_f(ctrl_I_top_0_f[50]),
    .Tile_X38Y51_A_T_top(ctrl_T_top[50]),
    .Tile_X38Y51_A_O_top_0_t(ctrl_O_top_0_t[50]),
    .Tile_X38Y51_A_O_top_0_f(ctrl_O_top_0_f[50]),
    .Tile_X38Y52_A_I_top_0_t(ctrl_I_top_0_t[51]),
    .Tile_X38Y52_A_I_top_0_f(ctrl_I_top_0_f[51]),
    .Tile_X38Y52_A_T_top(ctrl_T_top[51]),
    .Tile_X38Y52_A_O_top_0_t(ctrl_O_top_0_t[51]),
    .Tile_X38Y52_A_O_top_0_f(ctrl_O_top_0_f[51]),
    .Tile_X38Y53_A_I_top_0_t(ctrl_I_top_0_t[52]),
    .Tile_X38Y53_A_I_top_0_f(ctrl_I_top_0_f[52]),
    .Tile_X38Y53_A_T_top(ctrl_T_top[52]),
    .Tile_X38Y53_A_O_top_0_t(ctrl_O_top_0_t[52]),
    .Tile_X38Y53_A_O_top_0_f(ctrl_O_top_0_f[52]),
    .Tile_X38Y54_A_I_top_0_t(ctrl_I_top_0_t[53]),
    .Tile_X38Y54_A_I_top_0_f(ctrl_I_top_0_f[53]),
    .Tile_X38Y54_A_T_top(ctrl_T_top[53]),
    .Tile_X38Y54_A_O_top_0_t(ctrl_O_top_0_t[53]),
    .Tile_X38Y54_A_O_top_0_f(ctrl_O_top_0_f[53]),
    .Tile_X38Y55_A_I_top_0_t(ctrl_I_top_0_t[54]),
    .Tile_X38Y55_A_I_top_0_f(ctrl_I_top_0_f[54]),
    .Tile_X38Y55_A_T_top(ctrl_T_top[54]),
    .Tile_X38Y55_A_O_top_0_t(ctrl_O_top_0_t[54]),
    .Tile_X38Y55_A_O_top_0_f(ctrl_O_top_0_f[54]),
    .Tile_X38Y56_A_I_top_0_t(ctrl_I_top_0_t[55]),
    .Tile_X38Y56_A_I_top_0_f(ctrl_I_top_0_f[55]),
    .Tile_X38Y56_A_T_top(ctrl_T_top[55]),
    .Tile_X38Y56_A_O_top_0_t(ctrl_O_top_0_t[55]),
    .Tile_X38Y56_A_O_top_0_f(ctrl_O_top_0_f[55]),
    .Tile_X38Y57_A_I_top_0_t(ctrl_I_top_0_t[56]),
    .Tile_X38Y57_A_I_top_0_f(ctrl_I_top_0_f[56]),
    .Tile_X38Y57_A_T_top(ctrl_T_top[56]),
    .Tile_X38Y57_A_O_top_0_t(ctrl_O_top_0_t[56]),
    .Tile_X38Y57_A_O_top_0_f(ctrl_O_top_0_f[56]),
    .Tile_X38Y58_A_I_top_0_t(ctrl_I_top_0_t[57]),
    .Tile_X38Y58_A_I_top_0_f(ctrl_I_top_0_f[57]),
    .Tile_X38Y58_A_T_top(ctrl_T_top[57]),
    .Tile_X38Y58_A_O_top_0_t(ctrl_O_top_0_t[57]),
    .Tile_X38Y58_A_O_top_0_f(ctrl_O_top_0_f[57]),
    .Tile_X38Y59_A_I_top_0_t(ctrl_I_top_0_t[58]),
    .Tile_X38Y59_A_I_top_0_f(ctrl_I_top_0_f[58]),
    .Tile_X38Y59_A_T_top(ctrl_T_top[58]),
    .Tile_X38Y59_A_O_top_0_t(ctrl_O_top_0_t[58]),
    .Tile_X38Y59_A_O_top_0_f(ctrl_O_top_0_f[58]),
    .Tile_X38Y60_A_I_top_0_t(ctrl_I_top_0_t[59]),
    .Tile_X38Y60_A_I_top_0_f(ctrl_I_top_0_f[59]),
    .Tile_X38Y60_A_T_top(ctrl_T_top[59]),
    .Tile_X38Y60_A_O_top_0_t(ctrl_O_top_0_t[59]),
    .Tile_X38Y60_A_O_top_0_f(ctrl_O_top_0_f[59]),
    .rst(rst),
    .Tile_X0Y1_A_config_C_bit0(A_config_C[239]),
    .Tile_X0Y1_A_config_C_bit1(A_config_C[238]),
    .Tile_X0Y1_A_config_C_bit2(A_config_C[237]),
    .Tile_X0Y1_A_config_C_bit3(A_config_C[236]),
    .Tile_X0Y2_A_config_C_bit0(A_config_C[235]),
    .Tile_X0Y2_A_config_C_bit1(A_config_C[234]),
    .Tile_X0Y2_A_config_C_bit2(A_config_C[233]),
    .Tile_X0Y2_A_config_C_bit3(A_config_C[232]),
    .Tile_X0Y3_A_config_C_bit0(A_config_C[231]),
    .Tile_X0Y3_A_config_C_bit1(A_config_C[230]),
    .Tile_X0Y3_A_config_C_bit2(A_config_C[229]),
    .Tile_X0Y3_A_config_C_bit3(A_config_C[228]),
    .Tile_X0Y4_A_config_C_bit0(A_config_C[227]),
    .Tile_X0Y4_A_config_C_bit1(A_config_C[226]),
    .Tile_X0Y4_A_config_C_bit2(A_config_C[225]),
    .Tile_X0Y4_A_config_C_bit3(A_config_C[224]),
    .Tile_X0Y5_A_config_C_bit0(A_config_C[223]),
    .Tile_X0Y5_A_config_C_bit1(A_config_C[222]),
    .Tile_X0Y5_A_config_C_bit2(A_config_C[221]),
    .Tile_X0Y5_A_config_C_bit3(A_config_C[220]),
    .Tile_X0Y6_A_config_C_bit0(A_config_C[219]),
    .Tile_X0Y6_A_config_C_bit1(A_config_C[218]),
    .Tile_X0Y6_A_config_C_bit2(A_config_C[217]),
    .Tile_X0Y6_A_config_C_bit3(A_config_C[216]),
    .Tile_X0Y7_A_config_C_bit0(A_config_C[215]),
    .Tile_X0Y7_A_config_C_bit1(A_config_C[214]),
    .Tile_X0Y7_A_config_C_bit2(A_config_C[213]),
    .Tile_X0Y7_A_config_C_bit3(A_config_C[212]),
    .Tile_X0Y8_A_config_C_bit0(A_config_C[211]),
    .Tile_X0Y8_A_config_C_bit1(A_config_C[210]),
    .Tile_X0Y8_A_config_C_bit2(A_config_C[209]),
    .Tile_X0Y8_A_config_C_bit3(A_config_C[208]),
    .Tile_X0Y9_A_config_C_bit0(A_config_C[207]),
    .Tile_X0Y9_A_config_C_bit1(A_config_C[206]),
    .Tile_X0Y9_A_config_C_bit2(A_config_C[205]),
    .Tile_X0Y9_A_config_C_bit3(A_config_C[204]),
    .Tile_X0Y10_A_config_C_bit0(A_config_C[203]),
    .Tile_X0Y10_A_config_C_bit1(A_config_C[202]),
    .Tile_X0Y10_A_config_C_bit2(A_config_C[201]),
    .Tile_X0Y10_A_config_C_bit3(A_config_C[200]),
    .Tile_X0Y11_A_config_C_bit0(A_config_C[199]),
    .Tile_X0Y11_A_config_C_bit1(A_config_C[198]),
    .Tile_X0Y11_A_config_C_bit2(A_config_C[197]),
    .Tile_X0Y11_A_config_C_bit3(A_config_C[196]),
    .Tile_X0Y12_A_config_C_bit0(A_config_C[195]),
    .Tile_X0Y12_A_config_C_bit1(A_config_C[194]),
    .Tile_X0Y12_A_config_C_bit2(A_config_C[193]),
    .Tile_X0Y12_A_config_C_bit3(A_config_C[192]),
    .Tile_X0Y13_A_config_C_bit0(A_config_C[191]),
    .Tile_X0Y13_A_config_C_bit1(A_config_C[190]),
    .Tile_X0Y13_A_config_C_bit2(A_config_C[189]),
    .Tile_X0Y13_A_config_C_bit3(A_config_C[188]),
    .Tile_X0Y14_A_config_C_bit0(A_config_C[187]),
    .Tile_X0Y14_A_config_C_bit1(A_config_C[186]),
    .Tile_X0Y14_A_config_C_bit2(A_config_C[185]),
    .Tile_X0Y14_A_config_C_bit3(A_config_C[184]),
    .Tile_X0Y15_A_config_C_bit0(A_config_C[183]),
    .Tile_X0Y15_A_config_C_bit1(A_config_C[182]),
    .Tile_X0Y15_A_config_C_bit2(A_config_C[181]),
    .Tile_X0Y15_A_config_C_bit3(A_config_C[180]),
    .Tile_X0Y16_A_config_C_bit0(A_config_C[179]),
    .Tile_X0Y16_A_config_C_bit1(A_config_C[178]),
    .Tile_X0Y16_A_config_C_bit2(A_config_C[177]),
    .Tile_X0Y16_A_config_C_bit3(A_config_C[176]),
    .Tile_X0Y17_A_config_C_bit0(A_config_C[175]),
    .Tile_X0Y17_A_config_C_bit1(A_config_C[174]),
    .Tile_X0Y17_A_config_C_bit2(A_config_C[173]),
    .Tile_X0Y17_A_config_C_bit3(A_config_C[172]),
    .Tile_X0Y18_A_config_C_bit0(A_config_C[171]),
    .Tile_X0Y18_A_config_C_bit1(A_config_C[170]),
    .Tile_X0Y18_A_config_C_bit2(A_config_C[169]),
    .Tile_X0Y18_A_config_C_bit3(A_config_C[168]),
    .Tile_X0Y19_A_config_C_bit0(A_config_C[167]),
    .Tile_X0Y19_A_config_C_bit1(A_config_C[166]),
    .Tile_X0Y19_A_config_C_bit2(A_config_C[165]),
    .Tile_X0Y19_A_config_C_bit3(A_config_C[164]),
    .Tile_X0Y20_A_config_C_bit0(A_config_C[163]),
    .Tile_X0Y20_A_config_C_bit1(A_config_C[162]),
    .Tile_X0Y20_A_config_C_bit2(A_config_C[161]),
    .Tile_X0Y20_A_config_C_bit3(A_config_C[160]),
    .Tile_X0Y21_A_config_C_bit0(A_config_C[159]),
    .Tile_X0Y21_A_config_C_bit1(A_config_C[158]),
    .Tile_X0Y21_A_config_C_bit2(A_config_C[157]),
    .Tile_X0Y21_A_config_C_bit3(A_config_C[156]),
    .Tile_X0Y22_A_config_C_bit0(A_config_C[155]),
    .Tile_X0Y22_A_config_C_bit1(A_config_C[154]),
    .Tile_X0Y22_A_config_C_bit2(A_config_C[153]),
    .Tile_X0Y22_A_config_C_bit3(A_config_C[152]),
    .Tile_X0Y23_A_config_C_bit0(A_config_C[151]),
    .Tile_X0Y23_A_config_C_bit1(A_config_C[150]),
    .Tile_X0Y23_A_config_C_bit2(A_config_C[149]),
    .Tile_X0Y23_A_config_C_bit3(A_config_C[148]),
    .Tile_X0Y24_A_config_C_bit0(A_config_C[147]),
    .Tile_X0Y24_A_config_C_bit1(A_config_C[146]),
    .Tile_X0Y24_A_config_C_bit2(A_config_C[145]),
    .Tile_X0Y24_A_config_C_bit3(A_config_C[144]),
    .Tile_X0Y25_A_config_C_bit0(A_config_C[143]),
    .Tile_X0Y25_A_config_C_bit1(A_config_C[142]),
    .Tile_X0Y25_A_config_C_bit2(A_config_C[141]),
    .Tile_X0Y25_A_config_C_bit3(A_config_C[140]),
    .Tile_X0Y26_A_config_C_bit0(A_config_C[139]),
    .Tile_X0Y26_A_config_C_bit1(A_config_C[138]),
    .Tile_X0Y26_A_config_C_bit2(A_config_C[137]),
    .Tile_X0Y26_A_config_C_bit3(A_config_C[136]),
    .Tile_X0Y27_A_config_C_bit0(A_config_C[135]),
    .Tile_X0Y27_A_config_C_bit1(A_config_C[134]),
    .Tile_X0Y27_A_config_C_bit2(A_config_C[133]),
    .Tile_X0Y27_A_config_C_bit3(A_config_C[132]),
    .Tile_X0Y28_A_config_C_bit0(A_config_C[131]),
    .Tile_X0Y28_A_config_C_bit1(A_config_C[130]),
    .Tile_X0Y28_A_config_C_bit2(A_config_C[129]),
    .Tile_X0Y28_A_config_C_bit3(A_config_C[128]),
    .Tile_X0Y29_A_config_C_bit0(A_config_C[127]),
    .Tile_X0Y29_A_config_C_bit1(A_config_C[126]),
    .Tile_X0Y29_A_config_C_bit2(A_config_C[125]),
    .Tile_X0Y29_A_config_C_bit3(A_config_C[124]),
    .Tile_X0Y30_A_config_C_bit0(A_config_C[123]),
    .Tile_X0Y30_A_config_C_bit1(A_config_C[122]),
    .Tile_X0Y30_A_config_C_bit2(A_config_C[121]),
    .Tile_X0Y30_A_config_C_bit3(A_config_C[120]),
    .Tile_X0Y31_A_config_C_bit0(A_config_C[119]),
    .Tile_X0Y31_A_config_C_bit1(A_config_C[118]),
    .Tile_X0Y31_A_config_C_bit2(A_config_C[117]),
    .Tile_X0Y31_A_config_C_bit3(A_config_C[116]),
    .Tile_X0Y32_A_config_C_bit0(A_config_C[115]),
    .Tile_X0Y32_A_config_C_bit1(A_config_C[114]),
    .Tile_X0Y32_A_config_C_bit2(A_config_C[113]),
    .Tile_X0Y32_A_config_C_bit3(A_config_C[112]),
    .Tile_X0Y33_A_config_C_bit0(A_config_C[111]),
    .Tile_X0Y33_A_config_C_bit1(A_config_C[110]),
    .Tile_X0Y33_A_config_C_bit2(A_config_C[109]),
    .Tile_X0Y33_A_config_C_bit3(A_config_C[108]),
    .Tile_X0Y34_A_config_C_bit0(A_config_C[107]),
    .Tile_X0Y34_A_config_C_bit1(A_config_C[106]),
    .Tile_X0Y34_A_config_C_bit2(A_config_C[105]),
    .Tile_X0Y34_A_config_C_bit3(A_config_C[104]),
    .Tile_X0Y35_A_config_C_bit0(A_config_C[103]),
    .Tile_X0Y35_A_config_C_bit1(A_config_C[102]),
    .Tile_X0Y35_A_config_C_bit2(A_config_C[101]),
    .Tile_X0Y35_A_config_C_bit3(A_config_C[100]),
    .Tile_X0Y36_A_config_C_bit0(A_config_C[99]),
    .Tile_X0Y36_A_config_C_bit1(A_config_C[98]),
    .Tile_X0Y36_A_config_C_bit2(A_config_C[97]),
    .Tile_X0Y36_A_config_C_bit3(A_config_C[96]),
    .Tile_X0Y37_A_config_C_bit0(A_config_C[95]),
    .Tile_X0Y37_A_config_C_bit1(A_config_C[94]),
    .Tile_X0Y37_A_config_C_bit2(A_config_C[93]),
    .Tile_X0Y37_A_config_C_bit3(A_config_C[92]),
    .Tile_X0Y38_A_config_C_bit0(A_config_C[91]),
    .Tile_X0Y38_A_config_C_bit1(A_config_C[90]),
    .Tile_X0Y38_A_config_C_bit2(A_config_C[89]),
    .Tile_X0Y38_A_config_C_bit3(A_config_C[88]),
    .Tile_X0Y39_A_config_C_bit0(A_config_C[87]),
    .Tile_X0Y39_A_config_C_bit1(A_config_C[86]),
    .Tile_X0Y39_A_config_C_bit2(A_config_C[85]),
    .Tile_X0Y39_A_config_C_bit3(A_config_C[84]),
    .Tile_X0Y40_A_config_C_bit0(A_config_C[83]),
    .Tile_X0Y40_A_config_C_bit1(A_config_C[82]),
    .Tile_X0Y40_A_config_C_bit2(A_config_C[81]),
    .Tile_X0Y40_A_config_C_bit3(A_config_C[80]),
    .Tile_X0Y41_A_config_C_bit0(A_config_C[79]),
    .Tile_X0Y41_A_config_C_bit1(A_config_C[78]),
    .Tile_X0Y41_A_config_C_bit2(A_config_C[77]),
    .Tile_X0Y41_A_config_C_bit3(A_config_C[76]),
    .Tile_X0Y42_A_config_C_bit0(A_config_C[75]),
    .Tile_X0Y42_A_config_C_bit1(A_config_C[74]),
    .Tile_X0Y42_A_config_C_bit2(A_config_C[73]),
    .Tile_X0Y42_A_config_C_bit3(A_config_C[72]),
    .Tile_X0Y43_A_config_C_bit0(A_config_C[71]),
    .Tile_X0Y43_A_config_C_bit1(A_config_C[70]),
    .Tile_X0Y43_A_config_C_bit2(A_config_C[69]),
    .Tile_X0Y43_A_config_C_bit3(A_config_C[68]),
    .Tile_X0Y44_A_config_C_bit0(A_config_C[67]),
    .Tile_X0Y44_A_config_C_bit1(A_config_C[66]),
    .Tile_X0Y44_A_config_C_bit2(A_config_C[65]),
    .Tile_X0Y44_A_config_C_bit3(A_config_C[64]),
    .Tile_X0Y45_A_config_C_bit0(A_config_C[63]),
    .Tile_X0Y45_A_config_C_bit1(A_config_C[62]),
    .Tile_X0Y45_A_config_C_bit2(A_config_C[61]),
    .Tile_X0Y45_A_config_C_bit3(A_config_C[60]),
    .Tile_X0Y46_A_config_C_bit0(A_config_C[59]),
    .Tile_X0Y46_A_config_C_bit1(A_config_C[58]),
    .Tile_X0Y46_A_config_C_bit2(A_config_C[57]),
    .Tile_X0Y46_A_config_C_bit3(A_config_C[56]),
    .Tile_X0Y47_A_config_C_bit0(A_config_C[55]),
    .Tile_X0Y47_A_config_C_bit1(A_config_C[54]),
    .Tile_X0Y47_A_config_C_bit2(A_config_C[53]),
    .Tile_X0Y47_A_config_C_bit3(A_config_C[52]),
    .Tile_X0Y48_A_config_C_bit0(A_config_C[51]),
    .Tile_X0Y48_A_config_C_bit1(A_config_C[50]),
    .Tile_X0Y48_A_config_C_bit2(A_config_C[49]),
    .Tile_X0Y48_A_config_C_bit3(A_config_C[48]),
    .Tile_X0Y49_A_config_C_bit0(A_config_C[47]),
    .Tile_X0Y49_A_config_C_bit1(A_config_C[46]),
    .Tile_X0Y49_A_config_C_bit2(A_config_C[45]),
    .Tile_X0Y49_A_config_C_bit3(A_config_C[44]),
    .Tile_X0Y50_A_config_C_bit0(A_config_C[43]),
    .Tile_X0Y50_A_config_C_bit1(A_config_C[42]),
    .Tile_X0Y50_A_config_C_bit2(A_config_C[41]),
    .Tile_X0Y50_A_config_C_bit3(A_config_C[40]),
    .Tile_X0Y51_A_config_C_bit0(A_config_C[39]),
    .Tile_X0Y51_A_config_C_bit1(A_config_C[38]),
    .Tile_X0Y51_A_config_C_bit2(A_config_C[37]),
    .Tile_X0Y51_A_config_C_bit3(A_config_C[36]),
    .Tile_X0Y52_A_config_C_bit0(A_config_C[35]),
    .Tile_X0Y52_A_config_C_bit1(A_config_C[34]),
    .Tile_X0Y52_A_config_C_bit2(A_config_C[33]),
    .Tile_X0Y52_A_config_C_bit3(A_config_C[32]),
    .Tile_X0Y53_A_config_C_bit0(A_config_C[31]),
    .Tile_X0Y53_A_config_C_bit1(A_config_C[30]),
    .Tile_X0Y53_A_config_C_bit2(A_config_C[29]),
    .Tile_X0Y53_A_config_C_bit3(A_config_C[28]),
    .Tile_X0Y54_A_config_C_bit0(A_config_C[27]),
    .Tile_X0Y54_A_config_C_bit1(A_config_C[26]),
    .Tile_X0Y54_A_config_C_bit2(A_config_C[25]),
    .Tile_X0Y54_A_config_C_bit3(A_config_C[24]),
    .Tile_X0Y55_A_config_C_bit0(A_config_C[23]),
    .Tile_X0Y55_A_config_C_bit1(A_config_C[22]),
    .Tile_X0Y55_A_config_C_bit2(A_config_C[21]),
    .Tile_X0Y55_A_config_C_bit3(A_config_C[20]),
    .Tile_X0Y56_A_config_C_bit0(A_config_C[19]),
    .Tile_X0Y56_A_config_C_bit1(A_config_C[18]),
    .Tile_X0Y56_A_config_C_bit2(A_config_C[17]),
    .Tile_X0Y56_A_config_C_bit3(A_config_C[16]),
    .Tile_X0Y57_A_config_C_bit0(A_config_C[15]),
    .Tile_X0Y57_A_config_C_bit1(A_config_C[14]),
    .Tile_X0Y57_A_config_C_bit2(A_config_C[13]),
    .Tile_X0Y57_A_config_C_bit3(A_config_C[12]),
    .Tile_X0Y58_A_config_C_bit0(A_config_C[11]),
    .Tile_X0Y58_A_config_C_bit1(A_config_C[10]),
    .Tile_X0Y58_A_config_C_bit2(A_config_C[9]),
    .Tile_X0Y58_A_config_C_bit3(A_config_C[8]),
    .Tile_X0Y59_A_config_C_bit0(A_config_C[7]),
    .Tile_X0Y59_A_config_C_bit1(A_config_C[6]),
    .Tile_X0Y59_A_config_C_bit2(A_config_C[5]),
    .Tile_X0Y59_A_config_C_bit3(A_config_C[4]),
    .Tile_X0Y60_A_config_C_bit0(A_config_C[3]),
    .Tile_X0Y60_A_config_C_bit1(A_config_C[2]),
    .Tile_X0Y60_A_config_C_bit2(A_config_C[1]),
    .Tile_X0Y60_A_config_C_bit3(A_config_C[0]),
    .Tile_X0Y1_B_config_C_bit0(B_config_C[239]),
    .Tile_X0Y1_B_config_C_bit1(B_config_C[238]),
    .Tile_X0Y1_B_config_C_bit2(B_config_C[237]),
    .Tile_X0Y1_B_config_C_bit3(B_config_C[236]),
    .Tile_X0Y2_B_config_C_bit0(B_config_C[235]),
    .Tile_X0Y2_B_config_C_bit1(B_config_C[234]),
    .Tile_X0Y2_B_config_C_bit2(B_config_C[233]),
    .Tile_X0Y2_B_config_C_bit3(B_config_C[232]),
    .Tile_X0Y3_B_config_C_bit0(B_config_C[231]),
    .Tile_X0Y3_B_config_C_bit1(B_config_C[230]),
    .Tile_X0Y3_B_config_C_bit2(B_config_C[229]),
    .Tile_X0Y3_B_config_C_bit3(B_config_C[228]),
    .Tile_X0Y4_B_config_C_bit0(B_config_C[227]),
    .Tile_X0Y4_B_config_C_bit1(B_config_C[226]),
    .Tile_X0Y4_B_config_C_bit2(B_config_C[225]),
    .Tile_X0Y4_B_config_C_bit3(B_config_C[224]),
    .Tile_X0Y5_B_config_C_bit0(B_config_C[223]),
    .Tile_X0Y5_B_config_C_bit1(B_config_C[222]),
    .Tile_X0Y5_B_config_C_bit2(B_config_C[221]),
    .Tile_X0Y5_B_config_C_bit3(B_config_C[220]),
    .Tile_X0Y6_B_config_C_bit0(B_config_C[219]),
    .Tile_X0Y6_B_config_C_bit1(B_config_C[218]),
    .Tile_X0Y6_B_config_C_bit2(B_config_C[217]),
    .Tile_X0Y6_B_config_C_bit3(B_config_C[216]),
    .Tile_X0Y7_B_config_C_bit0(B_config_C[215]),
    .Tile_X0Y7_B_config_C_bit1(B_config_C[214]),
    .Tile_X0Y7_B_config_C_bit2(B_config_C[213]),
    .Tile_X0Y7_B_config_C_bit3(B_config_C[212]),
    .Tile_X0Y8_B_config_C_bit0(B_config_C[211]),
    .Tile_X0Y8_B_config_C_bit1(B_config_C[210]),
    .Tile_X0Y8_B_config_C_bit2(B_config_C[209]),
    .Tile_X0Y8_B_config_C_bit3(B_config_C[208]),
    .Tile_X0Y9_B_config_C_bit0(B_config_C[207]),
    .Tile_X0Y9_B_config_C_bit1(B_config_C[206]),
    .Tile_X0Y9_B_config_C_bit2(B_config_C[205]),
    .Tile_X0Y9_B_config_C_bit3(B_config_C[204]),
    .Tile_X0Y10_B_config_C_bit0(B_config_C[203]),
    .Tile_X0Y10_B_config_C_bit1(B_config_C[202]),
    .Tile_X0Y10_B_config_C_bit2(B_config_C[201]),
    .Tile_X0Y10_B_config_C_bit3(B_config_C[200]),
    .Tile_X0Y11_B_config_C_bit0(B_config_C[199]),
    .Tile_X0Y11_B_config_C_bit1(B_config_C[198]),
    .Tile_X0Y11_B_config_C_bit2(B_config_C[197]),
    .Tile_X0Y11_B_config_C_bit3(B_config_C[196]),
    .Tile_X0Y12_B_config_C_bit0(B_config_C[195]),
    .Tile_X0Y12_B_config_C_bit1(B_config_C[194]),
    .Tile_X0Y12_B_config_C_bit2(B_config_C[193]),
    .Tile_X0Y12_B_config_C_bit3(B_config_C[192]),
    .Tile_X0Y13_B_config_C_bit0(B_config_C[191]),
    .Tile_X0Y13_B_config_C_bit1(B_config_C[190]),
    .Tile_X0Y13_B_config_C_bit2(B_config_C[189]),
    .Tile_X0Y13_B_config_C_bit3(B_config_C[188]),
    .Tile_X0Y14_B_config_C_bit0(B_config_C[187]),
    .Tile_X0Y14_B_config_C_bit1(B_config_C[186]),
    .Tile_X0Y14_B_config_C_bit2(B_config_C[185]),
    .Tile_X0Y14_B_config_C_bit3(B_config_C[184]),
    .Tile_X0Y15_B_config_C_bit0(B_config_C[183]),
    .Tile_X0Y15_B_config_C_bit1(B_config_C[182]),
    .Tile_X0Y15_B_config_C_bit2(B_config_C[181]),
    .Tile_X0Y15_B_config_C_bit3(B_config_C[180]),
    .Tile_X0Y16_B_config_C_bit0(B_config_C[179]),
    .Tile_X0Y16_B_config_C_bit1(B_config_C[178]),
    .Tile_X0Y16_B_config_C_bit2(B_config_C[177]),
    .Tile_X0Y16_B_config_C_bit3(B_config_C[176]),
    .Tile_X0Y17_B_config_C_bit0(B_config_C[175]),
    .Tile_X0Y17_B_config_C_bit1(B_config_C[174]),
    .Tile_X0Y17_B_config_C_bit2(B_config_C[173]),
    .Tile_X0Y17_B_config_C_bit3(B_config_C[172]),
    .Tile_X0Y18_B_config_C_bit0(B_config_C[171]),
    .Tile_X0Y18_B_config_C_bit1(B_config_C[170]),
    .Tile_X0Y18_B_config_C_bit2(B_config_C[169]),
    .Tile_X0Y18_B_config_C_bit3(B_config_C[168]),
    .Tile_X0Y19_B_config_C_bit0(B_config_C[167]),
    .Tile_X0Y19_B_config_C_bit1(B_config_C[166]),
    .Tile_X0Y19_B_config_C_bit2(B_config_C[165]),
    .Tile_X0Y19_B_config_C_bit3(B_config_C[164]),
    .Tile_X0Y20_B_config_C_bit0(B_config_C[163]),
    .Tile_X0Y20_B_config_C_bit1(B_config_C[162]),
    .Tile_X0Y20_B_config_C_bit2(B_config_C[161]),
    .Tile_X0Y20_B_config_C_bit3(B_config_C[160]),
    .Tile_X0Y21_B_config_C_bit0(B_config_C[159]),
    .Tile_X0Y21_B_config_C_bit1(B_config_C[158]),
    .Tile_X0Y21_B_config_C_bit2(B_config_C[157]),
    .Tile_X0Y21_B_config_C_bit3(B_config_C[156]),
    .Tile_X0Y22_B_config_C_bit0(B_config_C[155]),
    .Tile_X0Y22_B_config_C_bit1(B_config_C[154]),
    .Tile_X0Y22_B_config_C_bit2(B_config_C[153]),
    .Tile_X0Y22_B_config_C_bit3(B_config_C[152]),
    .Tile_X0Y23_B_config_C_bit0(B_config_C[151]),
    .Tile_X0Y23_B_config_C_bit1(B_config_C[150]),
    .Tile_X0Y23_B_config_C_bit2(B_config_C[149]),
    .Tile_X0Y23_B_config_C_bit3(B_config_C[148]),
    .Tile_X0Y24_B_config_C_bit0(B_config_C[147]),
    .Tile_X0Y24_B_config_C_bit1(B_config_C[146]),
    .Tile_X0Y24_B_config_C_bit2(B_config_C[145]),
    .Tile_X0Y24_B_config_C_bit3(B_config_C[144]),
    .Tile_X0Y25_B_config_C_bit0(B_config_C[143]),
    .Tile_X0Y25_B_config_C_bit1(B_config_C[142]),
    .Tile_X0Y25_B_config_C_bit2(B_config_C[141]),
    .Tile_X0Y25_B_config_C_bit3(B_config_C[140]),
    .Tile_X0Y26_B_config_C_bit0(B_config_C[139]),
    .Tile_X0Y26_B_config_C_bit1(B_config_C[138]),
    .Tile_X0Y26_B_config_C_bit2(B_config_C[137]),
    .Tile_X0Y26_B_config_C_bit3(B_config_C[136]),
    .Tile_X0Y27_B_config_C_bit0(B_config_C[135]),
    .Tile_X0Y27_B_config_C_bit1(B_config_C[134]),
    .Tile_X0Y27_B_config_C_bit2(B_config_C[133]),
    .Tile_X0Y27_B_config_C_bit3(B_config_C[132]),
    .Tile_X0Y28_B_config_C_bit0(B_config_C[131]),
    .Tile_X0Y28_B_config_C_bit1(B_config_C[130]),
    .Tile_X0Y28_B_config_C_bit2(B_config_C[129]),
    .Tile_X0Y28_B_config_C_bit3(B_config_C[128]),
    .Tile_X0Y29_B_config_C_bit0(B_config_C[127]),
    .Tile_X0Y29_B_config_C_bit1(B_config_C[126]),
    .Tile_X0Y29_B_config_C_bit2(B_config_C[125]),
    .Tile_X0Y29_B_config_C_bit3(B_config_C[124]),
    .Tile_X0Y30_B_config_C_bit0(B_config_C[123]),
    .Tile_X0Y30_B_config_C_bit1(B_config_C[122]),
    .Tile_X0Y30_B_config_C_bit2(B_config_C[121]),
    .Tile_X0Y30_B_config_C_bit3(B_config_C[120]),
    .Tile_X0Y31_B_config_C_bit0(B_config_C[119]),
    .Tile_X0Y31_B_config_C_bit1(B_config_C[118]),
    .Tile_X0Y31_B_config_C_bit2(B_config_C[117]),
    .Tile_X0Y31_B_config_C_bit3(B_config_C[116]),
    .Tile_X0Y32_B_config_C_bit0(B_config_C[115]),
    .Tile_X0Y32_B_config_C_bit1(B_config_C[114]),
    .Tile_X0Y32_B_config_C_bit2(B_config_C[113]),
    .Tile_X0Y32_B_config_C_bit3(B_config_C[112]),
    .Tile_X0Y33_B_config_C_bit0(B_config_C[111]),
    .Tile_X0Y33_B_config_C_bit1(B_config_C[110]),
    .Tile_X0Y33_B_config_C_bit2(B_config_C[109]),
    .Tile_X0Y33_B_config_C_bit3(B_config_C[108]),
    .Tile_X0Y34_B_config_C_bit0(B_config_C[107]),
    .Tile_X0Y34_B_config_C_bit1(B_config_C[106]),
    .Tile_X0Y34_B_config_C_bit2(B_config_C[105]),
    .Tile_X0Y34_B_config_C_bit3(B_config_C[104]),
    .Tile_X0Y35_B_config_C_bit0(B_config_C[103]),
    .Tile_X0Y35_B_config_C_bit1(B_config_C[102]),
    .Tile_X0Y35_B_config_C_bit2(B_config_C[101]),
    .Tile_X0Y35_B_config_C_bit3(B_config_C[100]),
    .Tile_X0Y36_B_config_C_bit0(B_config_C[99]),
    .Tile_X0Y36_B_config_C_bit1(B_config_C[98]),
    .Tile_X0Y36_B_config_C_bit2(B_config_C[97]),
    .Tile_X0Y36_B_config_C_bit3(B_config_C[96]),
    .Tile_X0Y37_B_config_C_bit0(B_config_C[95]),
    .Tile_X0Y37_B_config_C_bit1(B_config_C[94]),
    .Tile_X0Y37_B_config_C_bit2(B_config_C[93]),
    .Tile_X0Y37_B_config_C_bit3(B_config_C[92]),
    .Tile_X0Y38_B_config_C_bit0(B_config_C[91]),
    .Tile_X0Y38_B_config_C_bit1(B_config_C[90]),
    .Tile_X0Y38_B_config_C_bit2(B_config_C[89]),
    .Tile_X0Y38_B_config_C_bit3(B_config_C[88]),
    .Tile_X0Y39_B_config_C_bit0(B_config_C[87]),
    .Tile_X0Y39_B_config_C_bit1(B_config_C[86]),
    .Tile_X0Y39_B_config_C_bit2(B_config_C[85]),
    .Tile_X0Y39_B_config_C_bit3(B_config_C[84]),
    .Tile_X0Y40_B_config_C_bit0(B_config_C[83]),
    .Tile_X0Y40_B_config_C_bit1(B_config_C[82]),
    .Tile_X0Y40_B_config_C_bit2(B_config_C[81]),
    .Tile_X0Y40_B_config_C_bit3(B_config_C[80]),
    .Tile_X0Y41_B_config_C_bit0(B_config_C[79]),
    .Tile_X0Y41_B_config_C_bit1(B_config_C[78]),
    .Tile_X0Y41_B_config_C_bit2(B_config_C[77]),
    .Tile_X0Y41_B_config_C_bit3(B_config_C[76]),
    .Tile_X0Y42_B_config_C_bit0(B_config_C[75]),
    .Tile_X0Y42_B_config_C_bit1(B_config_C[74]),
    .Tile_X0Y42_B_config_C_bit2(B_config_C[73]),
    .Tile_X0Y42_B_config_C_bit3(B_config_C[72]),
    .Tile_X0Y43_B_config_C_bit0(B_config_C[71]),
    .Tile_X0Y43_B_config_C_bit1(B_config_C[70]),
    .Tile_X0Y43_B_config_C_bit2(B_config_C[69]),
    .Tile_X0Y43_B_config_C_bit3(B_config_C[68]),
    .Tile_X0Y44_B_config_C_bit0(B_config_C[67]),
    .Tile_X0Y44_B_config_C_bit1(B_config_C[66]),
    .Tile_X0Y44_B_config_C_bit2(B_config_C[65]),
    .Tile_X0Y44_B_config_C_bit3(B_config_C[64]),
    .Tile_X0Y45_B_config_C_bit0(B_config_C[63]),
    .Tile_X0Y45_B_config_C_bit1(B_config_C[62]),
    .Tile_X0Y45_B_config_C_bit2(B_config_C[61]),
    .Tile_X0Y45_B_config_C_bit3(B_config_C[60]),
    .Tile_X0Y46_B_config_C_bit0(B_config_C[59]),
    .Tile_X0Y46_B_config_C_bit1(B_config_C[58]),
    .Tile_X0Y46_B_config_C_bit2(B_config_C[57]),
    .Tile_X0Y46_B_config_C_bit3(B_config_C[56]),
    .Tile_X0Y47_B_config_C_bit0(B_config_C[55]),
    .Tile_X0Y47_B_config_C_bit1(B_config_C[54]),
    .Tile_X0Y47_B_config_C_bit2(B_config_C[53]),
    .Tile_X0Y47_B_config_C_bit3(B_config_C[52]),
    .Tile_X0Y48_B_config_C_bit0(B_config_C[51]),
    .Tile_X0Y48_B_config_C_bit1(B_config_C[50]),
    .Tile_X0Y48_B_config_C_bit2(B_config_C[49]),
    .Tile_X0Y48_B_config_C_bit3(B_config_C[48]),
    .Tile_X0Y49_B_config_C_bit0(B_config_C[47]),
    .Tile_X0Y49_B_config_C_bit1(B_config_C[46]),
    .Tile_X0Y49_B_config_C_bit2(B_config_C[45]),
    .Tile_X0Y49_B_config_C_bit3(B_config_C[44]),
    .Tile_X0Y50_B_config_C_bit0(B_config_C[43]),
    .Tile_X0Y50_B_config_C_bit1(B_config_C[42]),
    .Tile_X0Y50_B_config_C_bit2(B_config_C[41]),
    .Tile_X0Y50_B_config_C_bit3(B_config_C[40]),
    .Tile_X0Y51_B_config_C_bit0(B_config_C[39]),
    .Tile_X0Y51_B_config_C_bit1(B_config_C[38]),
    .Tile_X0Y51_B_config_C_bit2(B_config_C[37]),
    .Tile_X0Y51_B_config_C_bit3(B_config_C[36]),
    .Tile_X0Y52_B_config_C_bit0(B_config_C[35]),
    .Tile_X0Y52_B_config_C_bit1(B_config_C[34]),
    .Tile_X0Y52_B_config_C_bit2(B_config_C[33]),
    .Tile_X0Y52_B_config_C_bit3(B_config_C[32]),
    .Tile_X0Y53_B_config_C_bit0(B_config_C[31]),
    .Tile_X0Y53_B_config_C_bit1(B_config_C[30]),
    .Tile_X0Y53_B_config_C_bit2(B_config_C[29]),
    .Tile_X0Y53_B_config_C_bit3(B_config_C[28]),
    .Tile_X0Y54_B_config_C_bit0(B_config_C[27]),
    .Tile_X0Y54_B_config_C_bit1(B_config_C[26]),
    .Tile_X0Y54_B_config_C_bit2(B_config_C[25]),
    .Tile_X0Y54_B_config_C_bit3(B_config_C[24]),
    .Tile_X0Y55_B_config_C_bit0(B_config_C[23]),
    .Tile_X0Y55_B_config_C_bit1(B_config_C[22]),
    .Tile_X0Y55_B_config_C_bit2(B_config_C[21]),
    .Tile_X0Y55_B_config_C_bit3(B_config_C[20]),
    .Tile_X0Y56_B_config_C_bit0(B_config_C[19]),
    .Tile_X0Y56_B_config_C_bit1(B_config_C[18]),
    .Tile_X0Y56_B_config_C_bit2(B_config_C[17]),
    .Tile_X0Y56_B_config_C_bit3(B_config_C[16]),
    .Tile_X0Y57_B_config_C_bit0(B_config_C[15]),
    .Tile_X0Y57_B_config_C_bit1(B_config_C[14]),
    .Tile_X0Y57_B_config_C_bit2(B_config_C[13]),
    .Tile_X0Y57_B_config_C_bit3(B_config_C[12]),
    .Tile_X0Y58_B_config_C_bit0(B_config_C[11]),
    .Tile_X0Y58_B_config_C_bit1(B_config_C[10]),
    .Tile_X0Y58_B_config_C_bit2(B_config_C[9]),
    .Tile_X0Y58_B_config_C_bit3(B_config_C[8]),
    .Tile_X0Y59_B_config_C_bit0(B_config_C[7]),
    .Tile_X0Y59_B_config_C_bit1(B_config_C[6]),
    .Tile_X0Y59_B_config_C_bit2(B_config_C[5]),
    .Tile_X0Y59_B_config_C_bit3(B_config_C[4]),
    .Tile_X0Y60_B_config_C_bit0(B_config_C[3]),
    .Tile_X0Y60_B_config_C_bit1(B_config_C[2]),
    .Tile_X0Y60_B_config_C_bit2(B_config_C[1]),
    .Tile_X0Y60_B_config_C_bit3(B_config_C[0]),
    .UserCLK(CLK),
    .FrameData(FrameData),
    .FrameStrobe(FrameSelect)
);


fault_detector  #(.Nm1(59), .Nm2(59), .Nctrl(59)) DR_check (
    .CLK(CLK),
    .rst(rst),
    .prech1(prech1),
    .prech2(prech2),
    .f_m1(F_masked1_top),
    .f_m2(F_masked2_top),
    .f_ctrl(F_ctrl_top),
    .f_detected(f_detected)
);

prech_signal_module prech_signal_module_i (
    .rst(rst),
    .CLK(CLK),
    .prech1(prech1),
    .prech2(prech2)
);

Trivium_DRP  #(.output_bits(1500)) Trivium_DRP_i (
    .clk(CLK),
    .rst(prng_rst),
    .prech1(prech1),
    .key_t(key_t),
    .key_f(key_f),
    .iv_t(iv_t),
    .iv_f(iv_f),
    .stream_out_t(R_t_top),
    .stream_out_f(R_f_top)
);

assign FrameData = {32'h12345678,FrameRegister,32'h12345678};
endmodule