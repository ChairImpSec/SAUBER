/* modified netlist. Source: module SkinnyTop in file /mnt/c/Users/amirm/Desktop/Papers_in_progress/SAUBER/Design for our FPGA/9-Skinny64_64_round_based_encryption_PortParallel/4-AGEMA/SkinnyTop.v */
/* 0 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 1 register stage(s) in total */

module SkinnyTop_SAUBER_Pipeline_d1 (Plaintext, Key, rst, Ciphertext, done);
    input [63:0] Plaintext ;
    input [63:0] Key ;
    input rst ;
    output [63:0] Ciphertext ;
    output done ;
    wire PlaintextMUX_MUXInst_0_U1_Y ;
    wire PlaintextMUX_MUXInst_0_U1_X ;
    wire PlaintextMUX_MUXInst_1_U1_Y ;
    wire PlaintextMUX_MUXInst_1_U1_X ;
    wire PlaintextMUX_MUXInst_2_U1_Y ;
    wire PlaintextMUX_MUXInst_2_U1_X ;
    wire PlaintextMUX_MUXInst_3_U1_Y ;
    wire PlaintextMUX_MUXInst_3_U1_X ;
    wire PlaintextMUX_MUXInst_4_U1_Y ;
    wire PlaintextMUX_MUXInst_4_U1_X ;
    wire PlaintextMUX_MUXInst_5_U1_Y ;
    wire PlaintextMUX_MUXInst_5_U1_X ;
    wire PlaintextMUX_MUXInst_6_U1_Y ;
    wire PlaintextMUX_MUXInst_6_U1_X ;
    wire PlaintextMUX_MUXInst_7_U1_Y ;
    wire PlaintextMUX_MUXInst_7_U1_X ;
    wire PlaintextMUX_MUXInst_8_U1_Y ;
    wire PlaintextMUX_MUXInst_8_U1_X ;
    wire PlaintextMUX_MUXInst_9_U1_Y ;
    wire PlaintextMUX_MUXInst_9_U1_X ;
    wire PlaintextMUX_MUXInst_10_U1_Y ;
    wire PlaintextMUX_MUXInst_10_U1_X ;
    wire PlaintextMUX_MUXInst_11_U1_Y ;
    wire PlaintextMUX_MUXInst_11_U1_X ;
    wire PlaintextMUX_MUXInst_12_U1_Y ;
    wire PlaintextMUX_MUXInst_12_U1_X ;
    wire PlaintextMUX_MUXInst_13_U1_Y ;
    wire PlaintextMUX_MUXInst_13_U1_X ;
    wire PlaintextMUX_MUXInst_14_U1_Y ;
    wire PlaintextMUX_MUXInst_14_U1_X ;
    wire PlaintextMUX_MUXInst_15_U1_Y ;
    wire PlaintextMUX_MUXInst_15_U1_X ;
    wire PlaintextMUX_MUXInst_16_U1_Y ;
    wire PlaintextMUX_MUXInst_16_U1_X ;
    wire PlaintextMUX_MUXInst_17_U1_Y ;
    wire PlaintextMUX_MUXInst_17_U1_X ;
    wire PlaintextMUX_MUXInst_18_U1_Y ;
    wire PlaintextMUX_MUXInst_18_U1_X ;
    wire PlaintextMUX_MUXInst_19_U1_Y ;
    wire PlaintextMUX_MUXInst_19_U1_X ;
    wire PlaintextMUX_MUXInst_20_U1_Y ;
    wire PlaintextMUX_MUXInst_20_U1_X ;
    wire PlaintextMUX_MUXInst_21_U1_Y ;
    wire PlaintextMUX_MUXInst_21_U1_X ;
    wire PlaintextMUX_MUXInst_22_U1_Y ;
    wire PlaintextMUX_MUXInst_22_U1_X ;
    wire PlaintextMUX_MUXInst_23_U1_Y ;
    wire PlaintextMUX_MUXInst_23_U1_X ;
    wire PlaintextMUX_MUXInst_24_U1_Y ;
    wire PlaintextMUX_MUXInst_24_U1_X ;
    wire PlaintextMUX_MUXInst_25_U1_Y ;
    wire PlaintextMUX_MUXInst_25_U1_X ;
    wire PlaintextMUX_MUXInst_26_U1_Y ;
    wire PlaintextMUX_MUXInst_26_U1_X ;
    wire PlaintextMUX_MUXInst_27_U1_Y ;
    wire PlaintextMUX_MUXInst_27_U1_X ;
    wire PlaintextMUX_MUXInst_28_U1_Y ;
    wire PlaintextMUX_MUXInst_28_U1_X ;
    wire PlaintextMUX_MUXInst_29_U1_Y ;
    wire PlaintextMUX_MUXInst_29_U1_X ;
    wire PlaintextMUX_MUXInst_30_U1_Y ;
    wire PlaintextMUX_MUXInst_30_U1_X ;
    wire PlaintextMUX_MUXInst_31_U1_Y ;
    wire PlaintextMUX_MUXInst_31_U1_X ;
    wire PlaintextMUX_MUXInst_32_U1_Y ;
    wire PlaintextMUX_MUXInst_32_U1_X ;
    wire PlaintextMUX_MUXInst_33_U1_Y ;
    wire PlaintextMUX_MUXInst_33_U1_X ;
    wire PlaintextMUX_MUXInst_34_U1_Y ;
    wire PlaintextMUX_MUXInst_34_U1_X ;
    wire PlaintextMUX_MUXInst_35_U1_Y ;
    wire PlaintextMUX_MUXInst_35_U1_X ;
    wire PlaintextMUX_MUXInst_36_U1_Y ;
    wire PlaintextMUX_MUXInst_36_U1_X ;
    wire PlaintextMUX_MUXInst_37_U1_Y ;
    wire PlaintextMUX_MUXInst_37_U1_X ;
    wire PlaintextMUX_MUXInst_38_U1_Y ;
    wire PlaintextMUX_MUXInst_38_U1_X ;
    wire PlaintextMUX_MUXInst_39_U1_Y ;
    wire PlaintextMUX_MUXInst_39_U1_X ;
    wire PlaintextMUX_MUXInst_40_U1_Y ;
    wire PlaintextMUX_MUXInst_40_U1_X ;
    wire PlaintextMUX_MUXInst_41_U1_Y ;
    wire PlaintextMUX_MUXInst_41_U1_X ;
    wire PlaintextMUX_MUXInst_42_U1_Y ;
    wire PlaintextMUX_MUXInst_42_U1_X ;
    wire PlaintextMUX_MUXInst_43_U1_Y ;
    wire PlaintextMUX_MUXInst_43_U1_X ;
    wire PlaintextMUX_MUXInst_44_U1_Y ;
    wire PlaintextMUX_MUXInst_44_U1_X ;
    wire PlaintextMUX_MUXInst_45_U1_Y ;
    wire PlaintextMUX_MUXInst_45_U1_X ;
    wire PlaintextMUX_MUXInst_46_U1_Y ;
    wire PlaintextMUX_MUXInst_46_U1_X ;
    wire PlaintextMUX_MUXInst_47_U1_Y ;
    wire PlaintextMUX_MUXInst_47_U1_X ;
    wire PlaintextMUX_MUXInst_48_U1_Y ;
    wire PlaintextMUX_MUXInst_48_U1_X ;
    wire PlaintextMUX_MUXInst_49_U1_Y ;
    wire PlaintextMUX_MUXInst_49_U1_X ;
    wire PlaintextMUX_MUXInst_50_U1_Y ;
    wire PlaintextMUX_MUXInst_50_U1_X ;
    wire PlaintextMUX_MUXInst_51_U1_Y ;
    wire PlaintextMUX_MUXInst_51_U1_X ;
    wire PlaintextMUX_MUXInst_52_U1_Y ;
    wire PlaintextMUX_MUXInst_52_U1_X ;
    wire PlaintextMUX_MUXInst_53_U1_Y ;
    wire PlaintextMUX_MUXInst_53_U1_X ;
    wire PlaintextMUX_MUXInst_54_U1_Y ;
    wire PlaintextMUX_MUXInst_54_U1_X ;
    wire PlaintextMUX_MUXInst_55_U1_Y ;
    wire PlaintextMUX_MUXInst_55_U1_X ;
    wire PlaintextMUX_MUXInst_56_U1_Y ;
    wire PlaintextMUX_MUXInst_56_U1_X ;
    wire PlaintextMUX_MUXInst_57_U1_Y ;
    wire PlaintextMUX_MUXInst_57_U1_X ;
    wire PlaintextMUX_MUXInst_58_U1_Y ;
    wire PlaintextMUX_MUXInst_58_U1_X ;
    wire PlaintextMUX_MUXInst_59_U1_Y ;
    wire PlaintextMUX_MUXInst_59_U1_X ;
    wire PlaintextMUX_MUXInst_60_U1_Y ;
    wire PlaintextMUX_MUXInst_60_U1_X ;
    wire PlaintextMUX_MUXInst_61_U1_Y ;
    wire PlaintextMUX_MUXInst_61_U1_X ;
    wire PlaintextMUX_MUXInst_62_U1_Y ;
    wire PlaintextMUX_MUXInst_62_U1_X ;
    wire PlaintextMUX_MUXInst_63_U1_Y ;
    wire PlaintextMUX_MUXInst_63_U1_X ;
    wire SubCellInst_SboxInst_0_L3 ;
    wire SubCellInst_SboxInst_0_YY_3 ;
    wire SubCellInst_SboxInst_0_L2 ;
    wire SubCellInst_SboxInst_0_T3 ;
    wire SubCellInst_SboxInst_0_Q7 ;
    wire SubCellInst_SboxInst_0_L1 ;
    wire SubCellInst_SboxInst_0_Q6 ;
    wire SubCellInst_SboxInst_0_L0 ;
    wire SubCellInst_SboxInst_0_T2 ;
    wire SubCellInst_SboxInst_0_Q4 ;
    wire SubCellInst_SboxInst_0_T1 ;
    wire SubCellInst_SboxInst_0_Q2 ;
    wire SubCellInst_SboxInst_0_T0 ;
    wire SubCellInst_SboxInst_0_Q1 ;
    wire SubCellInst_SboxInst_0_Q0 ;
    wire SubCellInst_SboxInst_1_L3 ;
    wire SubCellInst_SboxInst_1_YY_3 ;
    wire SubCellInst_SboxInst_1_L2 ;
    wire SubCellInst_SboxInst_1_T3 ;
    wire SubCellInst_SboxInst_1_Q7 ;
    wire SubCellInst_SboxInst_1_L1 ;
    wire SubCellInst_SboxInst_1_Q6 ;
    wire SubCellInst_SboxInst_1_L0 ;
    wire SubCellInst_SboxInst_1_T2 ;
    wire SubCellInst_SboxInst_1_Q4 ;
    wire SubCellInst_SboxInst_1_T1 ;
    wire SubCellInst_SboxInst_1_Q2 ;
    wire SubCellInst_SboxInst_1_T0 ;
    wire SubCellInst_SboxInst_1_Q1 ;
    wire SubCellInst_SboxInst_1_Q0 ;
    wire SubCellInst_SboxInst_2_L3 ;
    wire SubCellInst_SboxInst_2_YY_3 ;
    wire SubCellInst_SboxInst_2_L2 ;
    wire SubCellInst_SboxInst_2_T3 ;
    wire SubCellInst_SboxInst_2_Q7 ;
    wire SubCellInst_SboxInst_2_L1 ;
    wire SubCellInst_SboxInst_2_Q6 ;
    wire SubCellInst_SboxInst_2_L0 ;
    wire SubCellInst_SboxInst_2_T2 ;
    wire SubCellInst_SboxInst_2_Q4 ;
    wire SubCellInst_SboxInst_2_T1 ;
    wire SubCellInst_SboxInst_2_Q2 ;
    wire SubCellInst_SboxInst_2_T0 ;
    wire SubCellInst_SboxInst_2_Q1 ;
    wire SubCellInst_SboxInst_2_Q0 ;
    wire SubCellInst_SboxInst_3_L3 ;
    wire SubCellInst_SboxInst_3_YY_3 ;
    wire SubCellInst_SboxInst_3_L2 ;
    wire SubCellInst_SboxInst_3_T3 ;
    wire SubCellInst_SboxInst_3_Q7 ;
    wire SubCellInst_SboxInst_3_L1 ;
    wire SubCellInst_SboxInst_3_Q6 ;
    wire SubCellInst_SboxInst_3_L0 ;
    wire SubCellInst_SboxInst_3_T2 ;
    wire SubCellInst_SboxInst_3_Q4 ;
    wire SubCellInst_SboxInst_3_T1 ;
    wire SubCellInst_SboxInst_3_Q2 ;
    wire SubCellInst_SboxInst_3_T0 ;
    wire SubCellInst_SboxInst_3_Q1 ;
    wire SubCellInst_SboxInst_3_Q0 ;
    wire SubCellInst_SboxInst_4_L3 ;
    wire SubCellInst_SboxInst_4_YY_3 ;
    wire SubCellInst_SboxInst_4_L2 ;
    wire SubCellInst_SboxInst_4_T3 ;
    wire SubCellInst_SboxInst_4_Q7 ;
    wire SubCellInst_SboxInst_4_L1 ;
    wire SubCellInst_SboxInst_4_Q6 ;
    wire SubCellInst_SboxInst_4_L0 ;
    wire SubCellInst_SboxInst_4_T2 ;
    wire SubCellInst_SboxInst_4_Q4 ;
    wire SubCellInst_SboxInst_4_T1 ;
    wire SubCellInst_SboxInst_4_Q2 ;
    wire SubCellInst_SboxInst_4_T0 ;
    wire SubCellInst_SboxInst_4_Q1 ;
    wire SubCellInst_SboxInst_4_Q0 ;
    wire SubCellInst_SboxInst_5_L3 ;
    wire SubCellInst_SboxInst_5_YY_3 ;
    wire SubCellInst_SboxInst_5_L2 ;
    wire SubCellInst_SboxInst_5_T3 ;
    wire SubCellInst_SboxInst_5_Q7 ;
    wire SubCellInst_SboxInst_5_L1 ;
    wire SubCellInst_SboxInst_5_Q6 ;
    wire SubCellInst_SboxInst_5_L0 ;
    wire SubCellInst_SboxInst_5_T2 ;
    wire SubCellInst_SboxInst_5_Q4 ;
    wire SubCellInst_SboxInst_5_T1 ;
    wire SubCellInst_SboxInst_5_Q2 ;
    wire SubCellInst_SboxInst_5_T0 ;
    wire SubCellInst_SboxInst_5_Q1 ;
    wire SubCellInst_SboxInst_5_Q0 ;
    wire SubCellInst_SboxInst_6_L3 ;
    wire SubCellInst_SboxInst_6_YY_3 ;
    wire SubCellInst_SboxInst_6_L2 ;
    wire SubCellInst_SboxInst_6_T3 ;
    wire SubCellInst_SboxInst_6_Q7 ;
    wire SubCellInst_SboxInst_6_L1 ;
    wire SubCellInst_SboxInst_6_Q6 ;
    wire SubCellInst_SboxInst_6_L0 ;
    wire SubCellInst_SboxInst_6_T2 ;
    wire SubCellInst_SboxInst_6_Q4 ;
    wire SubCellInst_SboxInst_6_T1 ;
    wire SubCellInst_SboxInst_6_Q2 ;
    wire SubCellInst_SboxInst_6_T0 ;
    wire SubCellInst_SboxInst_6_Q1 ;
    wire SubCellInst_SboxInst_6_Q0 ;
    wire SubCellInst_SboxInst_7_L3 ;
    wire SubCellInst_SboxInst_7_YY_3 ;
    wire SubCellInst_SboxInst_7_L2 ;
    wire SubCellInst_SboxInst_7_T3 ;
    wire SubCellInst_SboxInst_7_Q7 ;
    wire SubCellInst_SboxInst_7_L1 ;
    wire SubCellInst_SboxInst_7_Q6 ;
    wire SubCellInst_SboxInst_7_L0 ;
    wire SubCellInst_SboxInst_7_T2 ;
    wire SubCellInst_SboxInst_7_Q4 ;
    wire SubCellInst_SboxInst_7_T1 ;
    wire SubCellInst_SboxInst_7_Q2 ;
    wire SubCellInst_SboxInst_7_T0 ;
    wire SubCellInst_SboxInst_7_Q1 ;
    wire SubCellInst_SboxInst_7_Q0 ;
    wire SubCellInst_SboxInst_8_L3 ;
    wire SubCellInst_SboxInst_8_YY_3 ;
    wire SubCellInst_SboxInst_8_L2 ;
    wire SubCellInst_SboxInst_8_T3 ;
    wire SubCellInst_SboxInst_8_Q7 ;
    wire SubCellInst_SboxInst_8_L1 ;
    wire SubCellInst_SboxInst_8_Q6 ;
    wire SubCellInst_SboxInst_8_L0 ;
    wire SubCellInst_SboxInst_8_T2 ;
    wire SubCellInst_SboxInst_8_Q4 ;
    wire SubCellInst_SboxInst_8_T1 ;
    wire SubCellInst_SboxInst_8_Q2 ;
    wire SubCellInst_SboxInst_8_T0 ;
    wire SubCellInst_SboxInst_8_Q1 ;
    wire SubCellInst_SboxInst_8_Q0 ;
    wire SubCellInst_SboxInst_9_L3 ;
    wire SubCellInst_SboxInst_9_YY_3 ;
    wire SubCellInst_SboxInst_9_L2 ;
    wire SubCellInst_SboxInst_9_T3 ;
    wire SubCellInst_SboxInst_9_Q7 ;
    wire SubCellInst_SboxInst_9_L1 ;
    wire SubCellInst_SboxInst_9_Q6 ;
    wire SubCellInst_SboxInst_9_L0 ;
    wire SubCellInst_SboxInst_9_T2 ;
    wire SubCellInst_SboxInst_9_Q4 ;
    wire SubCellInst_SboxInst_9_T1 ;
    wire SubCellInst_SboxInst_9_Q2 ;
    wire SubCellInst_SboxInst_9_T0 ;
    wire SubCellInst_SboxInst_9_Q1 ;
    wire SubCellInst_SboxInst_9_Q0 ;
    wire SubCellInst_SboxInst_10_L3 ;
    wire SubCellInst_SboxInst_10_YY_3 ;
    wire SubCellInst_SboxInst_10_L2 ;
    wire SubCellInst_SboxInst_10_T3 ;
    wire SubCellInst_SboxInst_10_Q7 ;
    wire SubCellInst_SboxInst_10_L1 ;
    wire SubCellInst_SboxInst_10_Q6 ;
    wire SubCellInst_SboxInst_10_L0 ;
    wire SubCellInst_SboxInst_10_T2 ;
    wire SubCellInst_SboxInst_10_Q4 ;
    wire SubCellInst_SboxInst_10_T1 ;
    wire SubCellInst_SboxInst_10_Q2 ;
    wire SubCellInst_SboxInst_10_T0 ;
    wire SubCellInst_SboxInst_10_Q1 ;
    wire SubCellInst_SboxInst_10_Q0 ;
    wire SubCellInst_SboxInst_11_L3 ;
    wire SubCellInst_SboxInst_11_YY_3 ;
    wire SubCellInst_SboxInst_11_L2 ;
    wire SubCellInst_SboxInst_11_T3 ;
    wire SubCellInst_SboxInst_11_Q7 ;
    wire SubCellInst_SboxInst_11_L1 ;
    wire SubCellInst_SboxInst_11_Q6 ;
    wire SubCellInst_SboxInst_11_L0 ;
    wire SubCellInst_SboxInst_11_T2 ;
    wire SubCellInst_SboxInst_11_Q4 ;
    wire SubCellInst_SboxInst_11_T1 ;
    wire SubCellInst_SboxInst_11_Q2 ;
    wire SubCellInst_SboxInst_11_T0 ;
    wire SubCellInst_SboxInst_11_Q1 ;
    wire SubCellInst_SboxInst_11_Q0 ;
    wire SubCellInst_SboxInst_12_L3 ;
    wire SubCellInst_SboxInst_12_YY_3 ;
    wire SubCellInst_SboxInst_12_L2 ;
    wire SubCellInst_SboxInst_12_T3 ;
    wire SubCellInst_SboxInst_12_Q7 ;
    wire SubCellInst_SboxInst_12_L1 ;
    wire SubCellInst_SboxInst_12_Q6 ;
    wire SubCellInst_SboxInst_12_L0 ;
    wire SubCellInst_SboxInst_12_T2 ;
    wire SubCellInst_SboxInst_12_Q4 ;
    wire SubCellInst_SboxInst_12_T1 ;
    wire SubCellInst_SboxInst_12_Q2 ;
    wire SubCellInst_SboxInst_12_T0 ;
    wire SubCellInst_SboxInst_12_Q1 ;
    wire SubCellInst_SboxInst_12_Q0 ;
    wire SubCellInst_SboxInst_13_L3 ;
    wire SubCellInst_SboxInst_13_YY_3 ;
    wire SubCellInst_SboxInst_13_L2 ;
    wire SubCellInst_SboxInst_13_T3 ;
    wire SubCellInst_SboxInst_13_Q7 ;
    wire SubCellInst_SboxInst_13_L1 ;
    wire SubCellInst_SboxInst_13_Q6 ;
    wire SubCellInst_SboxInst_13_L0 ;
    wire SubCellInst_SboxInst_13_T2 ;
    wire SubCellInst_SboxInst_13_Q4 ;
    wire SubCellInst_SboxInst_13_T1 ;
    wire SubCellInst_SboxInst_13_Q2 ;
    wire SubCellInst_SboxInst_13_T0 ;
    wire SubCellInst_SboxInst_13_Q1 ;
    wire SubCellInst_SboxInst_13_Q0 ;
    wire SubCellInst_SboxInst_14_L3 ;
    wire SubCellInst_SboxInst_14_YY_3 ;
    wire SubCellInst_SboxInst_14_L2 ;
    wire SubCellInst_SboxInst_14_T3 ;
    wire SubCellInst_SboxInst_14_Q7 ;
    wire SubCellInst_SboxInst_14_L1 ;
    wire SubCellInst_SboxInst_14_Q6 ;
    wire SubCellInst_SboxInst_14_L0 ;
    wire SubCellInst_SboxInst_14_T2 ;
    wire SubCellInst_SboxInst_14_Q4 ;
    wire SubCellInst_SboxInst_14_T1 ;
    wire SubCellInst_SboxInst_14_Q2 ;
    wire SubCellInst_SboxInst_14_T0 ;
    wire SubCellInst_SboxInst_14_Q1 ;
    wire SubCellInst_SboxInst_14_Q0 ;
    wire SubCellInst_SboxInst_15_L3 ;
    wire SubCellInst_SboxInst_15_YY_3 ;
    wire SubCellInst_SboxInst_15_L2 ;
    wire SubCellInst_SboxInst_15_T3 ;
    wire SubCellInst_SboxInst_15_Q7 ;
    wire SubCellInst_SboxInst_15_L1 ;
    wire SubCellInst_SboxInst_15_Q6 ;
    wire SubCellInst_SboxInst_15_L0 ;
    wire SubCellInst_SboxInst_15_T2 ;
    wire SubCellInst_SboxInst_15_Q4 ;
    wire SubCellInst_SboxInst_15_T1 ;
    wire SubCellInst_SboxInst_15_Q2 ;
    wire SubCellInst_SboxInst_15_T0 ;
    wire SubCellInst_SboxInst_15_Q1 ;
    wire SubCellInst_SboxInst_15_Q0 ;
    wire MCInst_MCR0_XORInst_0_0_n1 ;
    wire MCInst_MCR0_XORInst_0_1_n1 ;
    wire MCInst_MCR0_XORInst_0_2_n1 ;
    wire MCInst_MCR0_XORInst_0_3_n1 ;
    wire MCInst_MCR0_XORInst_1_0_n1 ;
    wire MCInst_MCR0_XORInst_1_1_n1 ;
    wire MCInst_MCR0_XORInst_1_2_n1 ;
    wire MCInst_MCR0_XORInst_1_3_n1 ;
    wire MCInst_MCR0_XORInst_2_0_n1 ;
    wire MCInst_MCR0_XORInst_2_1_n1 ;
    wire MCInst_MCR0_XORInst_2_2_n1 ;
    wire MCInst_MCR0_XORInst_2_3_n1 ;
    wire MCInst_MCR0_XORInst_3_0_n1 ;
    wire MCInst_MCR0_XORInst_3_1_n1 ;
    wire MCInst_MCR0_XORInst_3_2_n1 ;
    wire MCInst_MCR0_XORInst_3_3_n1 ;
    wire TweakeyGeneration_KEYMUX_MUXInst_0_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_0_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_1_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_1_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_2_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_2_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_3_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_3_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_4_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_4_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_5_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_5_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_6_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_6_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_7_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_7_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_8_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_8_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_9_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_9_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_10_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_10_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_11_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_11_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_12_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_12_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_13_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_13_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_14_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_14_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_15_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_15_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_16_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_16_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_17_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_17_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_18_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_18_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_19_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_19_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_20_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_20_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_21_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_21_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_22_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_22_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_23_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_23_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_24_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_24_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_25_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_25_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_26_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_26_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_27_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_27_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_28_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_28_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_29_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_29_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_30_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_30_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_31_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_31_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_32_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_32_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_33_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_33_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_34_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_34_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_35_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_35_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_36_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_36_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_37_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_37_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_38_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_38_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_39_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_39_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_40_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_40_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_41_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_41_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_42_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_42_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_43_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_43_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_44_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_44_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_45_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_45_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_46_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_46_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_47_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_47_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_48_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_48_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_49_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_49_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_50_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_50_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_51_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_51_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_52_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_52_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_53_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_53_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_54_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_54_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_55_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_55_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_56_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_56_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_57_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_57_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_58_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_58_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_59_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_59_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_60_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_60_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_61_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_61_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_62_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_62_U1_X ;
    wire TweakeyGeneration_KEYMUX_MUXInst_63_U1_Y ;
    wire TweakeyGeneration_KEYMUX_MUXInst_63_U1_X ;
    wire FSMUpdateInst_StateUpdateInst_0_n3 ;
    wire FSMUpdateInst_StateUpdateInst_0_n2 ;
    wire FSMUpdateInst_StateUpdateInst_0_n1 ;
    wire FSMUpdateInst_StateUpdateInst_0_n4 ;
    wire FSMUpdateInst_StateUpdateInst_0_U7_Y ;
    wire FSMUpdateInst_StateUpdateInst_0_U7_X ;
    wire FSMUpdateInst_StateUpdateInst_2_n4 ;
    wire FSMUpdateInst_StateUpdateInst_2_n3 ;
    wire FSMUpdateInst_StateUpdateInst_2_n2 ;
    wire FSMUpdateInst_StateUpdateInst_2_n1 ;
    wire FSMUpdateInst_StateUpdateInst_5_n4 ;
    wire FSMUpdateInst_StateUpdateInst_5_n3 ;
    wire FSMUpdateInst_StateUpdateInst_5_n2 ;
    wire FSMUpdateInst_StateUpdateInst_5_n1 ;
    wire FSMSignalsInst_doneInst_n5 ;
    wire FSMSignalsInst_doneInst_n4 ;
    wire FSMSignalsInst_doneInst_n3 ;
    wire FSMSignalsInst_doneInst_n2 ;
    wire [63:0] MCOutput ;
    wire [61:29] SubCellOutput ;
    wire [5:1] FSM ;
    wire [63:32] AddRoundConstantOutput ;
    wire [47:0] ShiftRowsOutput ;
    wire [5:0] FSMUpdate ;
    wire [1:0] SubCellInst_SboxInst_0_YY ;
    wire [2:1] SubCellInst_SboxInst_0_XX ;
    wire [1:0] SubCellInst_SboxInst_1_YY ;
    wire [2:1] SubCellInst_SboxInst_1_XX ;
    wire [1:0] SubCellInst_SboxInst_2_YY ;
    wire [2:1] SubCellInst_SboxInst_2_XX ;
    wire [1:0] SubCellInst_SboxInst_3_YY ;
    wire [2:1] SubCellInst_SboxInst_3_XX ;
    wire [1:0] SubCellInst_SboxInst_4_YY ;
    wire [2:1] SubCellInst_SboxInst_4_XX ;
    wire [1:0] SubCellInst_SboxInst_5_YY ;
    wire [2:1] SubCellInst_SboxInst_5_XX ;
    wire [1:0] SubCellInst_SboxInst_6_YY ;
    wire [2:1] SubCellInst_SboxInst_6_XX ;
    wire [1:0] SubCellInst_SboxInst_7_YY ;
    wire [2:1] SubCellInst_SboxInst_7_XX ;
    wire [1:0] SubCellInst_SboxInst_8_YY ;
    wire [2:1] SubCellInst_SboxInst_8_XX ;
    wire [1:0] SubCellInst_SboxInst_9_YY ;
    wire [2:1] SubCellInst_SboxInst_9_XX ;
    wire [1:0] SubCellInst_SboxInst_10_YY ;
    wire [2:1] SubCellInst_SboxInst_10_XX ;
    wire [1:0] SubCellInst_SboxInst_11_YY ;
    wire [2:1] SubCellInst_SboxInst_11_XX ;
    wire [1:0] SubCellInst_SboxInst_12_YY ;
    wire [2:1] SubCellInst_SboxInst_12_XX ;
    wire [1:0] SubCellInst_SboxInst_13_YY ;
    wire [2:1] SubCellInst_SboxInst_13_XX ;
    wire [1:0] SubCellInst_SboxInst_14_YY ;
    wire [2:1] SubCellInst_SboxInst_14_XX ;
    wire [1:0] SubCellInst_SboxInst_15_YY ;
    wire [2:1] SubCellInst_SboxInst_15_XX ;
    wire [63:0] TweakeyGeneration_key_Feedback ;

    /* cells in depth 0 */
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_0_U1_XOR1_U1 ( .A0_t (MCOutput[0]), .B0_t (Plaintext[0]), .Z0_t (PlaintextMUX_MUXInst_0_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_0_U1_AND1_U1 ( .A0_t (rst), .B0_t (PlaintextMUX_MUXInst_0_U1_X), .Z0_t (PlaintextMUX_MUXInst_0_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_0_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_0_U1_Y), .B0_t (MCOutput[0]), .Z0_t (Ciphertext[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_1_U1_XOR1_U1 ( .A0_t (MCOutput[1]), .B0_t (Plaintext[1]), .Z0_t (PlaintextMUX_MUXInst_1_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_1_U1_AND1_U1 ( .A0_t (rst), .B0_t (PlaintextMUX_MUXInst_1_U1_X), .Z0_t (PlaintextMUX_MUXInst_1_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_1_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_1_U1_Y), .B0_t (MCOutput[1]), .Z0_t (Ciphertext[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_2_U1_XOR1_U1 ( .A0_t (MCOutput[2]), .B0_t (Plaintext[2]), .Z0_t (PlaintextMUX_MUXInst_2_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_2_U1_AND1_U1 ( .A0_t (rst), .B0_t (PlaintextMUX_MUXInst_2_U1_X), .Z0_t (PlaintextMUX_MUXInst_2_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_2_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_2_U1_Y), .B0_t (MCOutput[2]), .Z0_t (Ciphertext[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_3_U1_XOR1_U1 ( .A0_t (MCOutput[3]), .B0_t (Plaintext[3]), .Z0_t (PlaintextMUX_MUXInst_3_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_3_U1_AND1_U1 ( .A0_t (rst), .B0_t (PlaintextMUX_MUXInst_3_U1_X), .Z0_t (PlaintextMUX_MUXInst_3_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_3_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_3_U1_Y), .B0_t (MCOutput[3]), .Z0_t (Ciphertext[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_4_U1_XOR1_U1 ( .A0_t (MCOutput[4]), .B0_t (Plaintext[4]), .Z0_t (PlaintextMUX_MUXInst_4_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_4_U1_AND1_U1 ( .A0_t (rst), .B0_t (PlaintextMUX_MUXInst_4_U1_X), .Z0_t (PlaintextMUX_MUXInst_4_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_4_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_4_U1_Y), .B0_t (MCOutput[4]), .Z0_t (Ciphertext[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_5_U1_XOR1_U1 ( .A0_t (MCOutput[5]), .B0_t (Plaintext[5]), .Z0_t (PlaintextMUX_MUXInst_5_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_5_U1_AND1_U1 ( .A0_t (rst), .B0_t (PlaintextMUX_MUXInst_5_U1_X), .Z0_t (PlaintextMUX_MUXInst_5_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_5_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_5_U1_Y), .B0_t (MCOutput[5]), .Z0_t (Ciphertext[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_6_U1_XOR1_U1 ( .A0_t (MCOutput[6]), .B0_t (Plaintext[6]), .Z0_t (PlaintextMUX_MUXInst_6_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_6_U1_AND1_U1 ( .A0_t (rst), .B0_t (PlaintextMUX_MUXInst_6_U1_X), .Z0_t (PlaintextMUX_MUXInst_6_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_6_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_6_U1_Y), .B0_t (MCOutput[6]), .Z0_t (Ciphertext[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_7_U1_XOR1_U1 ( .A0_t (MCOutput[7]), .B0_t (Plaintext[7]), .Z0_t (PlaintextMUX_MUXInst_7_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_7_U1_AND1_U1 ( .A0_t (rst), .B0_t (PlaintextMUX_MUXInst_7_U1_X), .Z0_t (PlaintextMUX_MUXInst_7_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_7_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_7_U1_Y), .B0_t (MCOutput[7]), .Z0_t (Ciphertext[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_8_U1_XOR1_U1 ( .A0_t (MCOutput[8]), .B0_t (Plaintext[8]), .Z0_t (PlaintextMUX_MUXInst_8_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_8_U1_AND1_U1 ( .A0_t (rst), .B0_t (PlaintextMUX_MUXInst_8_U1_X), .Z0_t (PlaintextMUX_MUXInst_8_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_8_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_8_U1_Y), .B0_t (MCOutput[8]), .Z0_t (Ciphertext[8]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_9_U1_XOR1_U1 ( .A0_t (MCOutput[9]), .B0_t (Plaintext[9]), .Z0_t (PlaintextMUX_MUXInst_9_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_9_U1_AND1_U1 ( .A0_t (rst), .B0_t (PlaintextMUX_MUXInst_9_U1_X), .Z0_t (PlaintextMUX_MUXInst_9_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_9_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_9_U1_Y), .B0_t (MCOutput[9]), .Z0_t (Ciphertext[9]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_10_U1_XOR1_U1 ( .A0_t (MCOutput[10]), .B0_t (Plaintext[10]), .Z0_t (PlaintextMUX_MUXInst_10_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_10_U1_AND1_U1 ( .A0_t (rst), .B0_t (PlaintextMUX_MUXInst_10_U1_X), .Z0_t (PlaintextMUX_MUXInst_10_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_10_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_10_U1_Y), .B0_t (MCOutput[10]), .Z0_t (Ciphertext[10]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_11_U1_XOR1_U1 ( .A0_t (MCOutput[11]), .B0_t (Plaintext[11]), .Z0_t (PlaintextMUX_MUXInst_11_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_11_U1_AND1_U1 ( .A0_t (rst), .B0_t (PlaintextMUX_MUXInst_11_U1_X), .Z0_t (PlaintextMUX_MUXInst_11_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_11_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_11_U1_Y), .B0_t (MCOutput[11]), .Z0_t (Ciphertext[11]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_12_U1_XOR1_U1 ( .A0_t (MCOutput[12]), .B0_t (Plaintext[12]), .Z0_t (PlaintextMUX_MUXInst_12_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_12_U1_AND1_U1 ( .A0_t (rst), .B0_t (PlaintextMUX_MUXInst_12_U1_X), .Z0_t (PlaintextMUX_MUXInst_12_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_12_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_12_U1_Y), .B0_t (MCOutput[12]), .Z0_t (Ciphertext[12]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_13_U1_XOR1_U1 ( .A0_t (MCOutput[13]), .B0_t (Plaintext[13]), .Z0_t (PlaintextMUX_MUXInst_13_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_13_U1_AND1_U1 ( .A0_t (rst), .B0_t (PlaintextMUX_MUXInst_13_U1_X), .Z0_t (PlaintextMUX_MUXInst_13_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_13_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_13_U1_Y), .B0_t (MCOutput[13]), .Z0_t (Ciphertext[13]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_14_U1_XOR1_U1 ( .A0_t (MCOutput[14]), .B0_t (Plaintext[14]), .Z0_t (PlaintextMUX_MUXInst_14_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_14_U1_AND1_U1 ( .A0_t (rst), .B0_t (PlaintextMUX_MUXInst_14_U1_X), .Z0_t (PlaintextMUX_MUXInst_14_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_14_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_14_U1_Y), .B0_t (MCOutput[14]), .Z0_t (Ciphertext[14]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_15_U1_XOR1_U1 ( .A0_t (MCOutput[15]), .B0_t (Plaintext[15]), .Z0_t (PlaintextMUX_MUXInst_15_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_15_U1_AND1_U1 ( .A0_t (rst), .B0_t (PlaintextMUX_MUXInst_15_U1_X), .Z0_t (PlaintextMUX_MUXInst_15_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_15_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_15_U1_Y), .B0_t (MCOutput[15]), .Z0_t (Ciphertext[15]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_16_U1_XOR1_U1 ( .A0_t (MCOutput[16]), .B0_t (Plaintext[16]), .Z0_t (PlaintextMUX_MUXInst_16_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_16_U1_AND1_U1 ( .A0_t (rst), .B0_t (PlaintextMUX_MUXInst_16_U1_X), .Z0_t (PlaintextMUX_MUXInst_16_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_16_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_16_U1_Y), .B0_t (MCOutput[16]), .Z0_t (Ciphertext[16]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_17_U1_XOR1_U1 ( .A0_t (MCOutput[17]), .B0_t (Plaintext[17]), .Z0_t (PlaintextMUX_MUXInst_17_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_17_U1_AND1_U1 ( .A0_t (rst), .B0_t (PlaintextMUX_MUXInst_17_U1_X), .Z0_t (PlaintextMUX_MUXInst_17_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_17_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_17_U1_Y), .B0_t (MCOutput[17]), .Z0_t (Ciphertext[17]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_18_U1_XOR1_U1 ( .A0_t (MCOutput[18]), .B0_t (Plaintext[18]), .Z0_t (PlaintextMUX_MUXInst_18_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_18_U1_AND1_U1 ( .A0_t (rst), .B0_t (PlaintextMUX_MUXInst_18_U1_X), .Z0_t (PlaintextMUX_MUXInst_18_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_18_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_18_U1_Y), .B0_t (MCOutput[18]), .Z0_t (Ciphertext[18]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_19_U1_XOR1_U1 ( .A0_t (MCOutput[19]), .B0_t (Plaintext[19]), .Z0_t (PlaintextMUX_MUXInst_19_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_19_U1_AND1_U1 ( .A0_t (rst), .B0_t (PlaintextMUX_MUXInst_19_U1_X), .Z0_t (PlaintextMUX_MUXInst_19_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_19_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_19_U1_Y), .B0_t (MCOutput[19]), .Z0_t (Ciphertext[19]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_20_U1_XOR1_U1 ( .A0_t (MCOutput[20]), .B0_t (Plaintext[20]), .Z0_t (PlaintextMUX_MUXInst_20_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_20_U1_AND1_U1 ( .A0_t (rst), .B0_t (PlaintextMUX_MUXInst_20_U1_X), .Z0_t (PlaintextMUX_MUXInst_20_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_20_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_20_U1_Y), .B0_t (MCOutput[20]), .Z0_t (Ciphertext[20]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_21_U1_XOR1_U1 ( .A0_t (MCOutput[21]), .B0_t (Plaintext[21]), .Z0_t (PlaintextMUX_MUXInst_21_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_21_U1_AND1_U1 ( .A0_t (rst), .B0_t (PlaintextMUX_MUXInst_21_U1_X), .Z0_t (PlaintextMUX_MUXInst_21_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_21_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_21_U1_Y), .B0_t (MCOutput[21]), .Z0_t (Ciphertext[21]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_22_U1_XOR1_U1 ( .A0_t (MCOutput[22]), .B0_t (Plaintext[22]), .Z0_t (PlaintextMUX_MUXInst_22_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_22_U1_AND1_U1 ( .A0_t (rst), .B0_t (PlaintextMUX_MUXInst_22_U1_X), .Z0_t (PlaintextMUX_MUXInst_22_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_22_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_22_U1_Y), .B0_t (MCOutput[22]), .Z0_t (Ciphertext[22]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_23_U1_XOR1_U1 ( .A0_t (MCOutput[23]), .B0_t (Plaintext[23]), .Z0_t (PlaintextMUX_MUXInst_23_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_23_U1_AND1_U1 ( .A0_t (rst), .B0_t (PlaintextMUX_MUXInst_23_U1_X), .Z0_t (PlaintextMUX_MUXInst_23_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_23_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_23_U1_Y), .B0_t (MCOutput[23]), .Z0_t (Ciphertext[23]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_24_U1_XOR1_U1 ( .A0_t (MCOutput[24]), .B0_t (Plaintext[24]), .Z0_t (PlaintextMUX_MUXInst_24_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_24_U1_AND1_U1 ( .A0_t (rst), .B0_t (PlaintextMUX_MUXInst_24_U1_X), .Z0_t (PlaintextMUX_MUXInst_24_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_24_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_24_U1_Y), .B0_t (MCOutput[24]), .Z0_t (Ciphertext[24]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_25_U1_XOR1_U1 ( .A0_t (MCOutput[25]), .B0_t (Plaintext[25]), .Z0_t (PlaintextMUX_MUXInst_25_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_25_U1_AND1_U1 ( .A0_t (rst), .B0_t (PlaintextMUX_MUXInst_25_U1_X), .Z0_t (PlaintextMUX_MUXInst_25_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_25_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_25_U1_Y), .B0_t (MCOutput[25]), .Z0_t (Ciphertext[25]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_26_U1_XOR1_U1 ( .A0_t (MCOutput[26]), .B0_t (Plaintext[26]), .Z0_t (PlaintextMUX_MUXInst_26_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_26_U1_AND1_U1 ( .A0_t (rst), .B0_t (PlaintextMUX_MUXInst_26_U1_X), .Z0_t (PlaintextMUX_MUXInst_26_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_26_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_26_U1_Y), .B0_t (MCOutput[26]), .Z0_t (Ciphertext[26]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_27_U1_XOR1_U1 ( .A0_t (MCOutput[27]), .B0_t (Plaintext[27]), .Z0_t (PlaintextMUX_MUXInst_27_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_27_U1_AND1_U1 ( .A0_t (rst), .B0_t (PlaintextMUX_MUXInst_27_U1_X), .Z0_t (PlaintextMUX_MUXInst_27_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_27_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_27_U1_Y), .B0_t (MCOutput[27]), .Z0_t (Ciphertext[27]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_28_U1_XOR1_U1 ( .A0_t (MCOutput[28]), .B0_t (Plaintext[28]), .Z0_t (PlaintextMUX_MUXInst_28_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_28_U1_AND1_U1 ( .A0_t (rst), .B0_t (PlaintextMUX_MUXInst_28_U1_X), .Z0_t (PlaintextMUX_MUXInst_28_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_28_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_28_U1_Y), .B0_t (MCOutput[28]), .Z0_t (Ciphertext[28]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_29_U1_XOR1_U1 ( .A0_t (MCOutput[29]), .B0_t (Plaintext[29]), .Z0_t (PlaintextMUX_MUXInst_29_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_29_U1_AND1_U1 ( .A0_t (rst), .B0_t (PlaintextMUX_MUXInst_29_U1_X), .Z0_t (PlaintextMUX_MUXInst_29_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_29_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_29_U1_Y), .B0_t (MCOutput[29]), .Z0_t (Ciphertext[29]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_30_U1_XOR1_U1 ( .A0_t (MCOutput[30]), .B0_t (Plaintext[30]), .Z0_t (PlaintextMUX_MUXInst_30_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_30_U1_AND1_U1 ( .A0_t (rst), .B0_t (PlaintextMUX_MUXInst_30_U1_X), .Z0_t (PlaintextMUX_MUXInst_30_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_30_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_30_U1_Y), .B0_t (MCOutput[30]), .Z0_t (Ciphertext[30]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_31_U1_XOR1_U1 ( .A0_t (MCOutput[31]), .B0_t (Plaintext[31]), .Z0_t (PlaintextMUX_MUXInst_31_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_31_U1_AND1_U1 ( .A0_t (rst), .B0_t (PlaintextMUX_MUXInst_31_U1_X), .Z0_t (PlaintextMUX_MUXInst_31_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_31_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_31_U1_Y), .B0_t (MCOutput[31]), .Z0_t (Ciphertext[31]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_32_U1_XOR1_U1 ( .A0_t (MCOutput[32]), .B0_t (Plaintext[32]), .Z0_t (PlaintextMUX_MUXInst_32_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_32_U1_AND1_U1 ( .A0_t (rst), .B0_t (PlaintextMUX_MUXInst_32_U1_X), .Z0_t (PlaintextMUX_MUXInst_32_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_32_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_32_U1_Y), .B0_t (MCOutput[32]), .Z0_t (Ciphertext[32]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_33_U1_XOR1_U1 ( .A0_t (MCOutput[33]), .B0_t (Plaintext[33]), .Z0_t (PlaintextMUX_MUXInst_33_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_33_U1_AND1_U1 ( .A0_t (rst), .B0_t (PlaintextMUX_MUXInst_33_U1_X), .Z0_t (PlaintextMUX_MUXInst_33_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_33_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_33_U1_Y), .B0_t (MCOutput[33]), .Z0_t (Ciphertext[33]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_34_U1_XOR1_U1 ( .A0_t (MCOutput[34]), .B0_t (Plaintext[34]), .Z0_t (PlaintextMUX_MUXInst_34_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_34_U1_AND1_U1 ( .A0_t (rst), .B0_t (PlaintextMUX_MUXInst_34_U1_X), .Z0_t (PlaintextMUX_MUXInst_34_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_34_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_34_U1_Y), .B0_t (MCOutput[34]), .Z0_t (Ciphertext[34]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_35_U1_XOR1_U1 ( .A0_t (MCOutput[35]), .B0_t (Plaintext[35]), .Z0_t (PlaintextMUX_MUXInst_35_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_35_U1_AND1_U1 ( .A0_t (rst), .B0_t (PlaintextMUX_MUXInst_35_U1_X), .Z0_t (PlaintextMUX_MUXInst_35_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_35_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_35_U1_Y), .B0_t (MCOutput[35]), .Z0_t (Ciphertext[35]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_36_U1_XOR1_U1 ( .A0_t (MCOutput[36]), .B0_t (Plaintext[36]), .Z0_t (PlaintextMUX_MUXInst_36_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_36_U1_AND1_U1 ( .A0_t (rst), .B0_t (PlaintextMUX_MUXInst_36_U1_X), .Z0_t (PlaintextMUX_MUXInst_36_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_36_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_36_U1_Y), .B0_t (MCOutput[36]), .Z0_t (Ciphertext[36]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_37_U1_XOR1_U1 ( .A0_t (MCOutput[37]), .B0_t (Plaintext[37]), .Z0_t (PlaintextMUX_MUXInst_37_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_37_U1_AND1_U1 ( .A0_t (rst), .B0_t (PlaintextMUX_MUXInst_37_U1_X), .Z0_t (PlaintextMUX_MUXInst_37_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_37_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_37_U1_Y), .B0_t (MCOutput[37]), .Z0_t (Ciphertext[37]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_38_U1_XOR1_U1 ( .A0_t (MCOutput[38]), .B0_t (Plaintext[38]), .Z0_t (PlaintextMUX_MUXInst_38_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_38_U1_AND1_U1 ( .A0_t (rst), .B0_t (PlaintextMUX_MUXInst_38_U1_X), .Z0_t (PlaintextMUX_MUXInst_38_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_38_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_38_U1_Y), .B0_t (MCOutput[38]), .Z0_t (Ciphertext[38]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_39_U1_XOR1_U1 ( .A0_t (MCOutput[39]), .B0_t (Plaintext[39]), .Z0_t (PlaintextMUX_MUXInst_39_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_39_U1_AND1_U1 ( .A0_t (rst), .B0_t (PlaintextMUX_MUXInst_39_U1_X), .Z0_t (PlaintextMUX_MUXInst_39_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_39_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_39_U1_Y), .B0_t (MCOutput[39]), .Z0_t (Ciphertext[39]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_40_U1_XOR1_U1 ( .A0_t (MCOutput[40]), .B0_t (Plaintext[40]), .Z0_t (PlaintextMUX_MUXInst_40_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_40_U1_AND1_U1 ( .A0_t (rst), .B0_t (PlaintextMUX_MUXInst_40_U1_X), .Z0_t (PlaintextMUX_MUXInst_40_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_40_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_40_U1_Y), .B0_t (MCOutput[40]), .Z0_t (Ciphertext[40]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_41_U1_XOR1_U1 ( .A0_t (MCOutput[41]), .B0_t (Plaintext[41]), .Z0_t (PlaintextMUX_MUXInst_41_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_41_U1_AND1_U1 ( .A0_t (rst), .B0_t (PlaintextMUX_MUXInst_41_U1_X), .Z0_t (PlaintextMUX_MUXInst_41_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_41_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_41_U1_Y), .B0_t (MCOutput[41]), .Z0_t (Ciphertext[41]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_42_U1_XOR1_U1 ( .A0_t (MCOutput[42]), .B0_t (Plaintext[42]), .Z0_t (PlaintextMUX_MUXInst_42_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_42_U1_AND1_U1 ( .A0_t (rst), .B0_t (PlaintextMUX_MUXInst_42_U1_X), .Z0_t (PlaintextMUX_MUXInst_42_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_42_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_42_U1_Y), .B0_t (MCOutput[42]), .Z0_t (Ciphertext[42]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_43_U1_XOR1_U1 ( .A0_t (MCOutput[43]), .B0_t (Plaintext[43]), .Z0_t (PlaintextMUX_MUXInst_43_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_43_U1_AND1_U1 ( .A0_t (rst), .B0_t (PlaintextMUX_MUXInst_43_U1_X), .Z0_t (PlaintextMUX_MUXInst_43_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_43_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_43_U1_Y), .B0_t (MCOutput[43]), .Z0_t (Ciphertext[43]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_44_U1_XOR1_U1 ( .A0_t (MCOutput[44]), .B0_t (Plaintext[44]), .Z0_t (PlaintextMUX_MUXInst_44_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_44_U1_AND1_U1 ( .A0_t (rst), .B0_t (PlaintextMUX_MUXInst_44_U1_X), .Z0_t (PlaintextMUX_MUXInst_44_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_44_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_44_U1_Y), .B0_t (MCOutput[44]), .Z0_t (Ciphertext[44]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_45_U1_XOR1_U1 ( .A0_t (MCOutput[45]), .B0_t (Plaintext[45]), .Z0_t (PlaintextMUX_MUXInst_45_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_45_U1_AND1_U1 ( .A0_t (rst), .B0_t (PlaintextMUX_MUXInst_45_U1_X), .Z0_t (PlaintextMUX_MUXInst_45_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_45_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_45_U1_Y), .B0_t (MCOutput[45]), .Z0_t (Ciphertext[45]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_46_U1_XOR1_U1 ( .A0_t (MCOutput[46]), .B0_t (Plaintext[46]), .Z0_t (PlaintextMUX_MUXInst_46_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_46_U1_AND1_U1 ( .A0_t (rst), .B0_t (PlaintextMUX_MUXInst_46_U1_X), .Z0_t (PlaintextMUX_MUXInst_46_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_46_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_46_U1_Y), .B0_t (MCOutput[46]), .Z0_t (Ciphertext[46]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_47_U1_XOR1_U1 ( .A0_t (MCOutput[47]), .B0_t (Plaintext[47]), .Z0_t (PlaintextMUX_MUXInst_47_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_47_U1_AND1_U1 ( .A0_t (rst), .B0_t (PlaintextMUX_MUXInst_47_U1_X), .Z0_t (PlaintextMUX_MUXInst_47_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_47_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_47_U1_Y), .B0_t (MCOutput[47]), .Z0_t (Ciphertext[47]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_48_U1_XOR1_U1 ( .A0_t (MCOutput[48]), .B0_t (Plaintext[48]), .Z0_t (PlaintextMUX_MUXInst_48_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_48_U1_AND1_U1 ( .A0_t (rst), .B0_t (PlaintextMUX_MUXInst_48_U1_X), .Z0_t (PlaintextMUX_MUXInst_48_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_48_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_48_U1_Y), .B0_t (MCOutput[48]), .Z0_t (Ciphertext[48]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_49_U1_XOR1_U1 ( .A0_t (MCOutput[49]), .B0_t (Plaintext[49]), .Z0_t (PlaintextMUX_MUXInst_49_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_49_U1_AND1_U1 ( .A0_t (rst), .B0_t (PlaintextMUX_MUXInst_49_U1_X), .Z0_t (PlaintextMUX_MUXInst_49_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_49_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_49_U1_Y), .B0_t (MCOutput[49]), .Z0_t (Ciphertext[49]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_50_U1_XOR1_U1 ( .A0_t (MCOutput[50]), .B0_t (Plaintext[50]), .Z0_t (PlaintextMUX_MUXInst_50_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_50_U1_AND1_U1 ( .A0_t (rst), .B0_t (PlaintextMUX_MUXInst_50_U1_X), .Z0_t (PlaintextMUX_MUXInst_50_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_50_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_50_U1_Y), .B0_t (MCOutput[50]), .Z0_t (Ciphertext[50]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_51_U1_XOR1_U1 ( .A0_t (MCOutput[51]), .B0_t (Plaintext[51]), .Z0_t (PlaintextMUX_MUXInst_51_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_51_U1_AND1_U1 ( .A0_t (rst), .B0_t (PlaintextMUX_MUXInst_51_U1_X), .Z0_t (PlaintextMUX_MUXInst_51_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_51_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_51_U1_Y), .B0_t (MCOutput[51]), .Z0_t (Ciphertext[51]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_52_U1_XOR1_U1 ( .A0_t (MCOutput[52]), .B0_t (Plaintext[52]), .Z0_t (PlaintextMUX_MUXInst_52_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_52_U1_AND1_U1 ( .A0_t (rst), .B0_t (PlaintextMUX_MUXInst_52_U1_X), .Z0_t (PlaintextMUX_MUXInst_52_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_52_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_52_U1_Y), .B0_t (MCOutput[52]), .Z0_t (Ciphertext[52]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_53_U1_XOR1_U1 ( .A0_t (MCOutput[53]), .B0_t (Plaintext[53]), .Z0_t (PlaintextMUX_MUXInst_53_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_53_U1_AND1_U1 ( .A0_t (rst), .B0_t (PlaintextMUX_MUXInst_53_U1_X), .Z0_t (PlaintextMUX_MUXInst_53_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_53_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_53_U1_Y), .B0_t (MCOutput[53]), .Z0_t (Ciphertext[53]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_54_U1_XOR1_U1 ( .A0_t (MCOutput[54]), .B0_t (Plaintext[54]), .Z0_t (PlaintextMUX_MUXInst_54_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_54_U1_AND1_U1 ( .A0_t (rst), .B0_t (PlaintextMUX_MUXInst_54_U1_X), .Z0_t (PlaintextMUX_MUXInst_54_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_54_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_54_U1_Y), .B0_t (MCOutput[54]), .Z0_t (Ciphertext[54]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_55_U1_XOR1_U1 ( .A0_t (MCOutput[55]), .B0_t (Plaintext[55]), .Z0_t (PlaintextMUX_MUXInst_55_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_55_U1_AND1_U1 ( .A0_t (rst), .B0_t (PlaintextMUX_MUXInst_55_U1_X), .Z0_t (PlaintextMUX_MUXInst_55_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_55_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_55_U1_Y), .B0_t (MCOutput[55]), .Z0_t (Ciphertext[55]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_56_U1_XOR1_U1 ( .A0_t (MCOutput[56]), .B0_t (Plaintext[56]), .Z0_t (PlaintextMUX_MUXInst_56_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_56_U1_AND1_U1 ( .A0_t (rst), .B0_t (PlaintextMUX_MUXInst_56_U1_X), .Z0_t (PlaintextMUX_MUXInst_56_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_56_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_56_U1_Y), .B0_t (MCOutput[56]), .Z0_t (Ciphertext[56]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_57_U1_XOR1_U1 ( .A0_t (MCOutput[57]), .B0_t (Plaintext[57]), .Z0_t (PlaintextMUX_MUXInst_57_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_57_U1_AND1_U1 ( .A0_t (rst), .B0_t (PlaintextMUX_MUXInst_57_U1_X), .Z0_t (PlaintextMUX_MUXInst_57_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_57_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_57_U1_Y), .B0_t (MCOutput[57]), .Z0_t (Ciphertext[57]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_58_U1_XOR1_U1 ( .A0_t (MCOutput[58]), .B0_t (Plaintext[58]), .Z0_t (PlaintextMUX_MUXInst_58_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_58_U1_AND1_U1 ( .A0_t (rst), .B0_t (PlaintextMUX_MUXInst_58_U1_X), .Z0_t (PlaintextMUX_MUXInst_58_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_58_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_58_U1_Y), .B0_t (MCOutput[58]), .Z0_t (Ciphertext[58]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_59_U1_XOR1_U1 ( .A0_t (MCOutput[59]), .B0_t (Plaintext[59]), .Z0_t (PlaintextMUX_MUXInst_59_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_59_U1_AND1_U1 ( .A0_t (rst), .B0_t (PlaintextMUX_MUXInst_59_U1_X), .Z0_t (PlaintextMUX_MUXInst_59_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_59_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_59_U1_Y), .B0_t (MCOutput[59]), .Z0_t (Ciphertext[59]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_60_U1_XOR1_U1 ( .A0_t (MCOutput[60]), .B0_t (Plaintext[60]), .Z0_t (PlaintextMUX_MUXInst_60_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_60_U1_AND1_U1 ( .A0_t (rst), .B0_t (PlaintextMUX_MUXInst_60_U1_X), .Z0_t (PlaintextMUX_MUXInst_60_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_60_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_60_U1_Y), .B0_t (MCOutput[60]), .Z0_t (Ciphertext[60]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_61_U1_XOR1_U1 ( .A0_t (MCOutput[61]), .B0_t (Plaintext[61]), .Z0_t (PlaintextMUX_MUXInst_61_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_61_U1_AND1_U1 ( .A0_t (rst), .B0_t (PlaintextMUX_MUXInst_61_U1_X), .Z0_t (PlaintextMUX_MUXInst_61_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_61_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_61_U1_Y), .B0_t (MCOutput[61]), .Z0_t (Ciphertext[61]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_62_U1_XOR1_U1 ( .A0_t (MCOutput[62]), .B0_t (Plaintext[62]), .Z0_t (PlaintextMUX_MUXInst_62_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_62_U1_AND1_U1 ( .A0_t (rst), .B0_t (PlaintextMUX_MUXInst_62_U1_X), .Z0_t (PlaintextMUX_MUXInst_62_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_62_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_62_U1_Y), .B0_t (MCOutput[62]), .Z0_t (Ciphertext[62]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_63_U1_XOR1_U1 ( .A0_t (MCOutput[63]), .B0_t (Plaintext[63]), .Z0_t (PlaintextMUX_MUXInst_63_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) PlaintextMUX_MUXInst_63_U1_AND1_U1 ( .A0_t (rst), .B0_t (PlaintextMUX_MUXInst_63_U1_X), .Z0_t (PlaintextMUX_MUXInst_63_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) PlaintextMUX_MUXInst_63_U1_XOR2_U1 ( .A0_t (PlaintextMUX_MUXInst_63_U1_Y), .B0_t (MCOutput[63]), .Z0_t (Ciphertext[63]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_0_XOR_i1_U1 ( .A0_t (Ciphertext[2]), .B0_t (Ciphertext[3]), .Z0_t (SubCellInst_SboxInst_0_XX[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_0_XOR_i2_U1 ( .A0_t (Ciphertext[0]), .B0_t (Ciphertext[2]), .Z0_t (SubCellInst_SboxInst_0_XX[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_0_XOR0_U1 ( .A0_t (Ciphertext[1]), .B0_t (SubCellInst_SboxInst_0_XX[2]), .Z0_t (SubCellInst_SboxInst_0_Q0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_0_XOR1_U1 ( .A0_t (Ciphertext[1]), .B0_t (SubCellInst_SboxInst_0_XX[1]), .Z0_t (SubCellInst_SboxInst_0_Q1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_0_AND1_U1 ( .A0_t (Ciphertext[2]), .B0_t (SubCellInst_SboxInst_0_Q1), .Z0_t (SubCellInst_SboxInst_0_T0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_0_XOR2_U1 ( .A0_t (SubCellInst_SboxInst_0_Q0), .B0_t (SubCellInst_SboxInst_0_T0), .Z0_t (SubCellInst_SboxInst_0_Q2) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_0_AND2_U1 ( .A0_t (Ciphertext[1]), .B0_t (SubCellInst_SboxInst_0_Q2), .Z0_t (SubCellInst_SboxInst_0_T1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_0_XOR3_U1 ( .A0_t (Ciphertext[1]), .B0_t (Ciphertext[2]), .Z0_t (SubCellInst_SboxInst_0_Q4) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_0_AND3_U1 ( .A0_t (Ciphertext[2]), .B0_t (SubCellInst_SboxInst_0_Q4), .Z0_t (SubCellInst_SboxInst_0_T2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_0_XOR4_U1 ( .A0_t (SubCellInst_SboxInst_0_T1), .B0_t (SubCellInst_SboxInst_0_T2), .Z0_t (SubCellInst_SboxInst_0_L0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_0_XOR5_U1 ( .A0_t (SubCellInst_SboxInst_0_XX[2]), .B0_t (Ciphertext[2]), .Z0_t (SubCellInst_SboxInst_0_Q6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_0_XOR6_U1 ( .A0_t (SubCellInst_SboxInst_0_Q1), .B0_t (SubCellInst_SboxInst_0_Q6), .Z0_t (SubCellInst_SboxInst_0_L1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_0_XOR7_U1 ( .A0_t (SubCellInst_SboxInst_0_L1), .B0_t (SubCellInst_SboxInst_0_T2), .Z0_t (SubCellInst_SboxInst_0_Q7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_0_AND4_U1 ( .A0_t (SubCellInst_SboxInst_0_Q6), .B0_t (SubCellInst_SboxInst_0_Q7), .Z0_t (SubCellInst_SboxInst_0_T3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_0_XOR8_U1 ( .A0_t (Ciphertext[1]), .B0_t (Ciphertext[2]), .Z0_t (SubCellInst_SboxInst_0_L2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_0_XOR9_U1 ( .A0_t (SubCellInst_SboxInst_0_L0), .B0_t (SubCellInst_SboxInst_0_L2), .Z0_t (SubCellInst_SboxInst_0_YY_3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_0_XOR10_U1 ( .A0_t (SubCellInst_SboxInst_0_L0), .B0_t (SubCellInst_SboxInst_0_T3), .Z0_t (ShiftRowsOutput[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_0_XOR11_U1 ( .A0_t (SubCellInst_SboxInst_0_XX[2]), .B0_t (SubCellInst_SboxInst_0_T0), .Z0_t (SubCellInst_SboxInst_0_L3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_0_XOR12_U1 ( .A0_t (SubCellInst_SboxInst_0_L3), .B0_t (SubCellInst_SboxInst_0_T2), .Z0_t (SubCellInst_SboxInst_0_YY[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_0_XOR13_U1 ( .A0_t (SubCellInst_SboxInst_0_XX[1]), .B0_t (SubCellInst_SboxInst_0_T2), .Z0_t (SubCellInst_SboxInst_0_YY[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_0_XOR_o1_U1 ( .A0_t (SubCellInst_SboxInst_0_YY[1]), .B0_t (SubCellInst_SboxInst_0_YY_3), .Z0_t (ShiftRowsOutput[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_1_XOR_i1_U1 ( .A0_t (Ciphertext[6]), .B0_t (Ciphertext[7]), .Z0_t (SubCellInst_SboxInst_1_XX[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_1_XOR_i2_U1 ( .A0_t (Ciphertext[4]), .B0_t (Ciphertext[6]), .Z0_t (SubCellInst_SboxInst_1_XX[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_1_XOR0_U1 ( .A0_t (Ciphertext[5]), .B0_t (SubCellInst_SboxInst_1_XX[2]), .Z0_t (SubCellInst_SboxInst_1_Q0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_1_XOR1_U1 ( .A0_t (Ciphertext[5]), .B0_t (SubCellInst_SboxInst_1_XX[1]), .Z0_t (SubCellInst_SboxInst_1_Q1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_1_AND1_U1 ( .A0_t (Ciphertext[6]), .B0_t (SubCellInst_SboxInst_1_Q1), .Z0_t (SubCellInst_SboxInst_1_T0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_1_XOR2_U1 ( .A0_t (SubCellInst_SboxInst_1_Q0), .B0_t (SubCellInst_SboxInst_1_T0), .Z0_t (SubCellInst_SboxInst_1_Q2) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_1_AND2_U1 ( .A0_t (Ciphertext[5]), .B0_t (SubCellInst_SboxInst_1_Q2), .Z0_t (SubCellInst_SboxInst_1_T1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_1_XOR3_U1 ( .A0_t (Ciphertext[5]), .B0_t (Ciphertext[6]), .Z0_t (SubCellInst_SboxInst_1_Q4) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_1_AND3_U1 ( .A0_t (Ciphertext[6]), .B0_t (SubCellInst_SboxInst_1_Q4), .Z0_t (SubCellInst_SboxInst_1_T2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_1_XOR4_U1 ( .A0_t (SubCellInst_SboxInst_1_T1), .B0_t (SubCellInst_SboxInst_1_T2), .Z0_t (SubCellInst_SboxInst_1_L0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_1_XOR5_U1 ( .A0_t (SubCellInst_SboxInst_1_XX[2]), .B0_t (Ciphertext[6]), .Z0_t (SubCellInst_SboxInst_1_Q6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_1_XOR6_U1 ( .A0_t (SubCellInst_SboxInst_1_Q1), .B0_t (SubCellInst_SboxInst_1_Q6), .Z0_t (SubCellInst_SboxInst_1_L1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_1_XOR7_U1 ( .A0_t (SubCellInst_SboxInst_1_L1), .B0_t (SubCellInst_SboxInst_1_T2), .Z0_t (SubCellInst_SboxInst_1_Q7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_1_AND4_U1 ( .A0_t (SubCellInst_SboxInst_1_Q6), .B0_t (SubCellInst_SboxInst_1_Q7), .Z0_t (SubCellInst_SboxInst_1_T3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_1_XOR8_U1 ( .A0_t (Ciphertext[5]), .B0_t (Ciphertext[6]), .Z0_t (SubCellInst_SboxInst_1_L2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_1_XOR9_U1 ( .A0_t (SubCellInst_SboxInst_1_L0), .B0_t (SubCellInst_SboxInst_1_L2), .Z0_t (SubCellInst_SboxInst_1_YY_3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_1_XOR10_U1 ( .A0_t (SubCellInst_SboxInst_1_L0), .B0_t (SubCellInst_SboxInst_1_T3), .Z0_t (ShiftRowsOutput[8]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_1_XOR11_U1 ( .A0_t (SubCellInst_SboxInst_1_XX[2]), .B0_t (SubCellInst_SboxInst_1_T0), .Z0_t (SubCellInst_SboxInst_1_L3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_1_XOR12_U1 ( .A0_t (SubCellInst_SboxInst_1_L3), .B0_t (SubCellInst_SboxInst_1_T2), .Z0_t (SubCellInst_SboxInst_1_YY[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_1_XOR13_U1 ( .A0_t (SubCellInst_SboxInst_1_XX[1]), .B0_t (SubCellInst_SboxInst_1_T2), .Z0_t (SubCellInst_SboxInst_1_YY[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_1_XOR_o1_U1 ( .A0_t (SubCellInst_SboxInst_1_YY[1]), .B0_t (SubCellInst_SboxInst_1_YY_3), .Z0_t (ShiftRowsOutput[9]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_2_XOR_i1_U1 ( .A0_t (Ciphertext[10]), .B0_t (Ciphertext[11]), .Z0_t (SubCellInst_SboxInst_2_XX[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_2_XOR_i2_U1 ( .A0_t (Ciphertext[8]), .B0_t (Ciphertext[10]), .Z0_t (SubCellInst_SboxInst_2_XX[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_2_XOR0_U1 ( .A0_t (Ciphertext[9]), .B0_t (SubCellInst_SboxInst_2_XX[2]), .Z0_t (SubCellInst_SboxInst_2_Q0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_2_XOR1_U1 ( .A0_t (Ciphertext[9]), .B0_t (SubCellInst_SboxInst_2_XX[1]), .Z0_t (SubCellInst_SboxInst_2_Q1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_2_AND1_U1 ( .A0_t (Ciphertext[10]), .B0_t (SubCellInst_SboxInst_2_Q1), .Z0_t (SubCellInst_SboxInst_2_T0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_2_XOR2_U1 ( .A0_t (SubCellInst_SboxInst_2_Q0), .B0_t (SubCellInst_SboxInst_2_T0), .Z0_t (SubCellInst_SboxInst_2_Q2) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_2_AND2_U1 ( .A0_t (Ciphertext[9]), .B0_t (SubCellInst_SboxInst_2_Q2), .Z0_t (SubCellInst_SboxInst_2_T1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_2_XOR3_U1 ( .A0_t (Ciphertext[9]), .B0_t (Ciphertext[10]), .Z0_t (SubCellInst_SboxInst_2_Q4) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_2_AND3_U1 ( .A0_t (Ciphertext[10]), .B0_t (SubCellInst_SboxInst_2_Q4), .Z0_t (SubCellInst_SboxInst_2_T2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_2_XOR4_U1 ( .A0_t (SubCellInst_SboxInst_2_T1), .B0_t (SubCellInst_SboxInst_2_T2), .Z0_t (SubCellInst_SboxInst_2_L0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_2_XOR5_U1 ( .A0_t (SubCellInst_SboxInst_2_XX[2]), .B0_t (Ciphertext[10]), .Z0_t (SubCellInst_SboxInst_2_Q6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_2_XOR6_U1 ( .A0_t (SubCellInst_SboxInst_2_Q1), .B0_t (SubCellInst_SboxInst_2_Q6), .Z0_t (SubCellInst_SboxInst_2_L1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_2_XOR7_U1 ( .A0_t (SubCellInst_SboxInst_2_L1), .B0_t (SubCellInst_SboxInst_2_T2), .Z0_t (SubCellInst_SboxInst_2_Q7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_2_AND4_U1 ( .A0_t (SubCellInst_SboxInst_2_Q6), .B0_t (SubCellInst_SboxInst_2_Q7), .Z0_t (SubCellInst_SboxInst_2_T3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_2_XOR8_U1 ( .A0_t (Ciphertext[9]), .B0_t (Ciphertext[10]), .Z0_t (SubCellInst_SboxInst_2_L2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_2_XOR9_U1 ( .A0_t (SubCellInst_SboxInst_2_L0), .B0_t (SubCellInst_SboxInst_2_L2), .Z0_t (SubCellInst_SboxInst_2_YY_3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_2_XOR10_U1 ( .A0_t (SubCellInst_SboxInst_2_L0), .B0_t (SubCellInst_SboxInst_2_T3), .Z0_t (ShiftRowsOutput[12]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_2_XOR11_U1 ( .A0_t (SubCellInst_SboxInst_2_XX[2]), .B0_t (SubCellInst_SboxInst_2_T0), .Z0_t (SubCellInst_SboxInst_2_L3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_2_XOR12_U1 ( .A0_t (SubCellInst_SboxInst_2_L3), .B0_t (SubCellInst_SboxInst_2_T2), .Z0_t (SubCellInst_SboxInst_2_YY[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_2_XOR13_U1 ( .A0_t (SubCellInst_SboxInst_2_XX[1]), .B0_t (SubCellInst_SboxInst_2_T2), .Z0_t (SubCellInst_SboxInst_2_YY[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_2_XOR_o1_U1 ( .A0_t (SubCellInst_SboxInst_2_YY[1]), .B0_t (SubCellInst_SboxInst_2_YY_3), .Z0_t (ShiftRowsOutput[13]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_3_XOR_i1_U1 ( .A0_t (Ciphertext[14]), .B0_t (Ciphertext[15]), .Z0_t (SubCellInst_SboxInst_3_XX[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_3_XOR_i2_U1 ( .A0_t (Ciphertext[12]), .B0_t (Ciphertext[14]), .Z0_t (SubCellInst_SboxInst_3_XX[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_3_XOR0_U1 ( .A0_t (Ciphertext[13]), .B0_t (SubCellInst_SboxInst_3_XX[2]), .Z0_t (SubCellInst_SboxInst_3_Q0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_3_XOR1_U1 ( .A0_t (Ciphertext[13]), .B0_t (SubCellInst_SboxInst_3_XX[1]), .Z0_t (SubCellInst_SboxInst_3_Q1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_3_AND1_U1 ( .A0_t (Ciphertext[14]), .B0_t (SubCellInst_SboxInst_3_Q1), .Z0_t (SubCellInst_SboxInst_3_T0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_3_XOR2_U1 ( .A0_t (SubCellInst_SboxInst_3_Q0), .B0_t (SubCellInst_SboxInst_3_T0), .Z0_t (SubCellInst_SboxInst_3_Q2) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_3_AND2_U1 ( .A0_t (Ciphertext[13]), .B0_t (SubCellInst_SboxInst_3_Q2), .Z0_t (SubCellInst_SboxInst_3_T1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_3_XOR3_U1 ( .A0_t (Ciphertext[13]), .B0_t (Ciphertext[14]), .Z0_t (SubCellInst_SboxInst_3_Q4) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_3_AND3_U1 ( .A0_t (Ciphertext[14]), .B0_t (SubCellInst_SboxInst_3_Q4), .Z0_t (SubCellInst_SboxInst_3_T2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_3_XOR4_U1 ( .A0_t (SubCellInst_SboxInst_3_T1), .B0_t (SubCellInst_SboxInst_3_T2), .Z0_t (SubCellInst_SboxInst_3_L0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_3_XOR5_U1 ( .A0_t (SubCellInst_SboxInst_3_XX[2]), .B0_t (Ciphertext[14]), .Z0_t (SubCellInst_SboxInst_3_Q6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_3_XOR6_U1 ( .A0_t (SubCellInst_SboxInst_3_Q1), .B0_t (SubCellInst_SboxInst_3_Q6), .Z0_t (SubCellInst_SboxInst_3_L1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_3_XOR7_U1 ( .A0_t (SubCellInst_SboxInst_3_L1), .B0_t (SubCellInst_SboxInst_3_T2), .Z0_t (SubCellInst_SboxInst_3_Q7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_3_AND4_U1 ( .A0_t (SubCellInst_SboxInst_3_Q6), .B0_t (SubCellInst_SboxInst_3_Q7), .Z0_t (SubCellInst_SboxInst_3_T3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_3_XOR8_U1 ( .A0_t (Ciphertext[13]), .B0_t (Ciphertext[14]), .Z0_t (SubCellInst_SboxInst_3_L2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_3_XOR9_U1 ( .A0_t (SubCellInst_SboxInst_3_L0), .B0_t (SubCellInst_SboxInst_3_L2), .Z0_t (SubCellInst_SboxInst_3_YY_3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_3_XOR10_U1 ( .A0_t (SubCellInst_SboxInst_3_L0), .B0_t (SubCellInst_SboxInst_3_T3), .Z0_t (ShiftRowsOutput[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_3_XOR11_U1 ( .A0_t (SubCellInst_SboxInst_3_XX[2]), .B0_t (SubCellInst_SboxInst_3_T0), .Z0_t (SubCellInst_SboxInst_3_L3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_3_XOR12_U1 ( .A0_t (SubCellInst_SboxInst_3_L3), .B0_t (SubCellInst_SboxInst_3_T2), .Z0_t (SubCellInst_SboxInst_3_YY[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_3_XOR13_U1 ( .A0_t (SubCellInst_SboxInst_3_XX[1]), .B0_t (SubCellInst_SboxInst_3_T2), .Z0_t (SubCellInst_SboxInst_3_YY[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_3_XOR_o1_U1 ( .A0_t (SubCellInst_SboxInst_3_YY[1]), .B0_t (SubCellInst_SboxInst_3_YY_3), .Z0_t (ShiftRowsOutput[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_4_XOR_i1_U1 ( .A0_t (Ciphertext[18]), .B0_t (Ciphertext[19]), .Z0_t (SubCellInst_SboxInst_4_XX[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_4_XOR_i2_U1 ( .A0_t (Ciphertext[16]), .B0_t (Ciphertext[18]), .Z0_t (SubCellInst_SboxInst_4_XX[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_4_XOR0_U1 ( .A0_t (Ciphertext[17]), .B0_t (SubCellInst_SboxInst_4_XX[2]), .Z0_t (SubCellInst_SboxInst_4_Q0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_4_XOR1_U1 ( .A0_t (Ciphertext[17]), .B0_t (SubCellInst_SboxInst_4_XX[1]), .Z0_t (SubCellInst_SboxInst_4_Q1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_4_AND1_U1 ( .A0_t (Ciphertext[18]), .B0_t (SubCellInst_SboxInst_4_Q1), .Z0_t (SubCellInst_SboxInst_4_T0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_4_XOR2_U1 ( .A0_t (SubCellInst_SboxInst_4_Q0), .B0_t (SubCellInst_SboxInst_4_T0), .Z0_t (SubCellInst_SboxInst_4_Q2) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_4_AND2_U1 ( .A0_t (Ciphertext[17]), .B0_t (SubCellInst_SboxInst_4_Q2), .Z0_t (SubCellInst_SboxInst_4_T1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_4_XOR3_U1 ( .A0_t (Ciphertext[17]), .B0_t (Ciphertext[18]), .Z0_t (SubCellInst_SboxInst_4_Q4) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_4_AND3_U1 ( .A0_t (Ciphertext[18]), .B0_t (SubCellInst_SboxInst_4_Q4), .Z0_t (SubCellInst_SboxInst_4_T2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_4_XOR4_U1 ( .A0_t (SubCellInst_SboxInst_4_T1), .B0_t (SubCellInst_SboxInst_4_T2), .Z0_t (SubCellInst_SboxInst_4_L0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_4_XOR5_U1 ( .A0_t (SubCellInst_SboxInst_4_XX[2]), .B0_t (Ciphertext[18]), .Z0_t (SubCellInst_SboxInst_4_Q6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_4_XOR6_U1 ( .A0_t (SubCellInst_SboxInst_4_Q1), .B0_t (SubCellInst_SboxInst_4_Q6), .Z0_t (SubCellInst_SboxInst_4_L1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_4_XOR7_U1 ( .A0_t (SubCellInst_SboxInst_4_L1), .B0_t (SubCellInst_SboxInst_4_T2), .Z0_t (SubCellInst_SboxInst_4_Q7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_4_AND4_U1 ( .A0_t (SubCellInst_SboxInst_4_Q6), .B0_t (SubCellInst_SboxInst_4_Q7), .Z0_t (SubCellInst_SboxInst_4_T3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_4_XOR8_U1 ( .A0_t (Ciphertext[17]), .B0_t (Ciphertext[18]), .Z0_t (SubCellInst_SboxInst_4_L2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_4_XOR9_U1 ( .A0_t (SubCellInst_SboxInst_4_L0), .B0_t (SubCellInst_SboxInst_4_L2), .Z0_t (SubCellInst_SboxInst_4_YY_3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_4_XOR10_U1 ( .A0_t (SubCellInst_SboxInst_4_L0), .B0_t (SubCellInst_SboxInst_4_T3), .Z0_t (ShiftRowsOutput[24]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_4_XOR11_U1 ( .A0_t (SubCellInst_SboxInst_4_XX[2]), .B0_t (SubCellInst_SboxInst_4_T0), .Z0_t (SubCellInst_SboxInst_4_L3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_4_XOR12_U1 ( .A0_t (SubCellInst_SboxInst_4_L3), .B0_t (SubCellInst_SboxInst_4_T2), .Z0_t (SubCellInst_SboxInst_4_YY[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_4_XOR13_U1 ( .A0_t (SubCellInst_SboxInst_4_XX[1]), .B0_t (SubCellInst_SboxInst_4_T2), .Z0_t (SubCellInst_SboxInst_4_YY[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_4_XOR_o1_U1 ( .A0_t (SubCellInst_SboxInst_4_YY[1]), .B0_t (SubCellInst_SboxInst_4_YY_3), .Z0_t (ShiftRowsOutput[25]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_5_XOR_i1_U1 ( .A0_t (Ciphertext[22]), .B0_t (Ciphertext[23]), .Z0_t (SubCellInst_SboxInst_5_XX[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_5_XOR_i2_U1 ( .A0_t (Ciphertext[20]), .B0_t (Ciphertext[22]), .Z0_t (SubCellInst_SboxInst_5_XX[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_5_XOR0_U1 ( .A0_t (Ciphertext[21]), .B0_t (SubCellInst_SboxInst_5_XX[2]), .Z0_t (SubCellInst_SboxInst_5_Q0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_5_XOR1_U1 ( .A0_t (Ciphertext[21]), .B0_t (SubCellInst_SboxInst_5_XX[1]), .Z0_t (SubCellInst_SboxInst_5_Q1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_5_AND1_U1 ( .A0_t (Ciphertext[22]), .B0_t (SubCellInst_SboxInst_5_Q1), .Z0_t (SubCellInst_SboxInst_5_T0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_5_XOR2_U1 ( .A0_t (SubCellInst_SboxInst_5_Q0), .B0_t (SubCellInst_SboxInst_5_T0), .Z0_t (SubCellInst_SboxInst_5_Q2) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_5_AND2_U1 ( .A0_t (Ciphertext[21]), .B0_t (SubCellInst_SboxInst_5_Q2), .Z0_t (SubCellInst_SboxInst_5_T1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_5_XOR3_U1 ( .A0_t (Ciphertext[21]), .B0_t (Ciphertext[22]), .Z0_t (SubCellInst_SboxInst_5_Q4) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_5_AND3_U1 ( .A0_t (Ciphertext[22]), .B0_t (SubCellInst_SboxInst_5_Q4), .Z0_t (SubCellInst_SboxInst_5_T2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_5_XOR4_U1 ( .A0_t (SubCellInst_SboxInst_5_T1), .B0_t (SubCellInst_SboxInst_5_T2), .Z0_t (SubCellInst_SboxInst_5_L0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_5_XOR5_U1 ( .A0_t (SubCellInst_SboxInst_5_XX[2]), .B0_t (Ciphertext[22]), .Z0_t (SubCellInst_SboxInst_5_Q6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_5_XOR6_U1 ( .A0_t (SubCellInst_SboxInst_5_Q1), .B0_t (SubCellInst_SboxInst_5_Q6), .Z0_t (SubCellInst_SboxInst_5_L1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_5_XOR7_U1 ( .A0_t (SubCellInst_SboxInst_5_L1), .B0_t (SubCellInst_SboxInst_5_T2), .Z0_t (SubCellInst_SboxInst_5_Q7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_5_AND4_U1 ( .A0_t (SubCellInst_SboxInst_5_Q6), .B0_t (SubCellInst_SboxInst_5_Q7), .Z0_t (SubCellInst_SboxInst_5_T3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_5_XOR8_U1 ( .A0_t (Ciphertext[21]), .B0_t (Ciphertext[22]), .Z0_t (SubCellInst_SboxInst_5_L2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_5_XOR9_U1 ( .A0_t (SubCellInst_SboxInst_5_L0), .B0_t (SubCellInst_SboxInst_5_L2), .Z0_t (SubCellInst_SboxInst_5_YY_3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_5_XOR10_U1 ( .A0_t (SubCellInst_SboxInst_5_L0), .B0_t (SubCellInst_SboxInst_5_T3), .Z0_t (ShiftRowsOutput[28]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_5_XOR11_U1 ( .A0_t (SubCellInst_SboxInst_5_XX[2]), .B0_t (SubCellInst_SboxInst_5_T0), .Z0_t (SubCellInst_SboxInst_5_L3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_5_XOR12_U1 ( .A0_t (SubCellInst_SboxInst_5_L3), .B0_t (SubCellInst_SboxInst_5_T2), .Z0_t (SubCellInst_SboxInst_5_YY[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_5_XOR13_U1 ( .A0_t (SubCellInst_SboxInst_5_XX[1]), .B0_t (SubCellInst_SboxInst_5_T2), .Z0_t (SubCellInst_SboxInst_5_YY[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_5_XOR_o1_U1 ( .A0_t (SubCellInst_SboxInst_5_YY[1]), .B0_t (SubCellInst_SboxInst_5_YY_3), .Z0_t (ShiftRowsOutput[29]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_6_XOR_i1_U1 ( .A0_t (Ciphertext[26]), .B0_t (Ciphertext[27]), .Z0_t (SubCellInst_SboxInst_6_XX[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_6_XOR_i2_U1 ( .A0_t (Ciphertext[24]), .B0_t (Ciphertext[26]), .Z0_t (SubCellInst_SboxInst_6_XX[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_6_XOR0_U1 ( .A0_t (Ciphertext[25]), .B0_t (SubCellInst_SboxInst_6_XX[2]), .Z0_t (SubCellInst_SboxInst_6_Q0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_6_XOR1_U1 ( .A0_t (Ciphertext[25]), .B0_t (SubCellInst_SboxInst_6_XX[1]), .Z0_t (SubCellInst_SboxInst_6_Q1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_6_AND1_U1 ( .A0_t (Ciphertext[26]), .B0_t (SubCellInst_SboxInst_6_Q1), .Z0_t (SubCellInst_SboxInst_6_T0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_6_XOR2_U1 ( .A0_t (SubCellInst_SboxInst_6_Q0), .B0_t (SubCellInst_SboxInst_6_T0), .Z0_t (SubCellInst_SboxInst_6_Q2) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_6_AND2_U1 ( .A0_t (Ciphertext[25]), .B0_t (SubCellInst_SboxInst_6_Q2), .Z0_t (SubCellInst_SboxInst_6_T1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_6_XOR3_U1 ( .A0_t (Ciphertext[25]), .B0_t (Ciphertext[26]), .Z0_t (SubCellInst_SboxInst_6_Q4) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_6_AND3_U1 ( .A0_t (Ciphertext[26]), .B0_t (SubCellInst_SboxInst_6_Q4), .Z0_t (SubCellInst_SboxInst_6_T2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_6_XOR4_U1 ( .A0_t (SubCellInst_SboxInst_6_T1), .B0_t (SubCellInst_SboxInst_6_T2), .Z0_t (SubCellInst_SboxInst_6_L0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_6_XOR5_U1 ( .A0_t (SubCellInst_SboxInst_6_XX[2]), .B0_t (Ciphertext[26]), .Z0_t (SubCellInst_SboxInst_6_Q6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_6_XOR6_U1 ( .A0_t (SubCellInst_SboxInst_6_Q1), .B0_t (SubCellInst_SboxInst_6_Q6), .Z0_t (SubCellInst_SboxInst_6_L1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_6_XOR7_U1 ( .A0_t (SubCellInst_SboxInst_6_L1), .B0_t (SubCellInst_SboxInst_6_T2), .Z0_t (SubCellInst_SboxInst_6_Q7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_6_AND4_U1 ( .A0_t (SubCellInst_SboxInst_6_Q6), .B0_t (SubCellInst_SboxInst_6_Q7), .Z0_t (SubCellInst_SboxInst_6_T3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_6_XOR8_U1 ( .A0_t (Ciphertext[25]), .B0_t (Ciphertext[26]), .Z0_t (SubCellInst_SboxInst_6_L2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_6_XOR9_U1 ( .A0_t (SubCellInst_SboxInst_6_L0), .B0_t (SubCellInst_SboxInst_6_L2), .Z0_t (SubCellInst_SboxInst_6_YY_3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_6_XOR10_U1 ( .A0_t (SubCellInst_SboxInst_6_L0), .B0_t (SubCellInst_SboxInst_6_T3), .Z0_t (ShiftRowsOutput[16]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_6_XOR11_U1 ( .A0_t (SubCellInst_SboxInst_6_XX[2]), .B0_t (SubCellInst_SboxInst_6_T0), .Z0_t (SubCellInst_SboxInst_6_L3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_6_XOR12_U1 ( .A0_t (SubCellInst_SboxInst_6_L3), .B0_t (SubCellInst_SboxInst_6_T2), .Z0_t (SubCellInst_SboxInst_6_YY[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_6_XOR13_U1 ( .A0_t (SubCellInst_SboxInst_6_XX[1]), .B0_t (SubCellInst_SboxInst_6_T2), .Z0_t (SubCellInst_SboxInst_6_YY[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_6_XOR_o1_U1 ( .A0_t (SubCellInst_SboxInst_6_YY[1]), .B0_t (SubCellInst_SboxInst_6_YY_3), .Z0_t (ShiftRowsOutput[17]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_7_XOR_i1_U1 ( .A0_t (Ciphertext[30]), .B0_t (Ciphertext[31]), .Z0_t (SubCellInst_SboxInst_7_XX[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_7_XOR_i2_U1 ( .A0_t (Ciphertext[28]), .B0_t (Ciphertext[30]), .Z0_t (SubCellInst_SboxInst_7_XX[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_7_XOR0_U1 ( .A0_t (Ciphertext[29]), .B0_t (SubCellInst_SboxInst_7_XX[2]), .Z0_t (SubCellInst_SboxInst_7_Q0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_7_XOR1_U1 ( .A0_t (Ciphertext[29]), .B0_t (SubCellInst_SboxInst_7_XX[1]), .Z0_t (SubCellInst_SboxInst_7_Q1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_7_AND1_U1 ( .A0_t (Ciphertext[30]), .B0_t (SubCellInst_SboxInst_7_Q1), .Z0_t (SubCellInst_SboxInst_7_T0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_7_XOR2_U1 ( .A0_t (SubCellInst_SboxInst_7_Q0), .B0_t (SubCellInst_SboxInst_7_T0), .Z0_t (SubCellInst_SboxInst_7_Q2) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_7_AND2_U1 ( .A0_t (Ciphertext[29]), .B0_t (SubCellInst_SboxInst_7_Q2), .Z0_t (SubCellInst_SboxInst_7_T1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_7_XOR3_U1 ( .A0_t (Ciphertext[29]), .B0_t (Ciphertext[30]), .Z0_t (SubCellInst_SboxInst_7_Q4) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_7_AND3_U1 ( .A0_t (Ciphertext[30]), .B0_t (SubCellInst_SboxInst_7_Q4), .Z0_t (SubCellInst_SboxInst_7_T2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_7_XOR4_U1 ( .A0_t (SubCellInst_SboxInst_7_T1), .B0_t (SubCellInst_SboxInst_7_T2), .Z0_t (SubCellInst_SboxInst_7_L0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_7_XOR5_U1 ( .A0_t (SubCellInst_SboxInst_7_XX[2]), .B0_t (Ciphertext[30]), .Z0_t (SubCellInst_SboxInst_7_Q6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_7_XOR6_U1 ( .A0_t (SubCellInst_SboxInst_7_Q1), .B0_t (SubCellInst_SboxInst_7_Q6), .Z0_t (SubCellInst_SboxInst_7_L1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_7_XOR7_U1 ( .A0_t (SubCellInst_SboxInst_7_L1), .B0_t (SubCellInst_SboxInst_7_T2), .Z0_t (SubCellInst_SboxInst_7_Q7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_7_AND4_U1 ( .A0_t (SubCellInst_SboxInst_7_Q6), .B0_t (SubCellInst_SboxInst_7_Q7), .Z0_t (SubCellInst_SboxInst_7_T3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_7_XOR8_U1 ( .A0_t (Ciphertext[29]), .B0_t (Ciphertext[30]), .Z0_t (SubCellInst_SboxInst_7_L2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_7_XOR9_U1 ( .A0_t (SubCellInst_SboxInst_7_L0), .B0_t (SubCellInst_SboxInst_7_L2), .Z0_t (SubCellInst_SboxInst_7_YY_3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_7_XOR10_U1 ( .A0_t (SubCellInst_SboxInst_7_L0), .B0_t (SubCellInst_SboxInst_7_T3), .Z0_t (ShiftRowsOutput[20]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_7_XOR11_U1 ( .A0_t (SubCellInst_SboxInst_7_XX[2]), .B0_t (SubCellInst_SboxInst_7_T0), .Z0_t (SubCellInst_SboxInst_7_L3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_7_XOR12_U1 ( .A0_t (SubCellInst_SboxInst_7_L3), .B0_t (SubCellInst_SboxInst_7_T2), .Z0_t (SubCellInst_SboxInst_7_YY[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_7_XOR13_U1 ( .A0_t (SubCellInst_SboxInst_7_XX[1]), .B0_t (SubCellInst_SboxInst_7_T2), .Z0_t (SubCellInst_SboxInst_7_YY[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_7_XOR_o1_U1 ( .A0_t (SubCellInst_SboxInst_7_YY[1]), .B0_t (SubCellInst_SboxInst_7_YY_3), .Z0_t (SubCellOutput[29]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_8_XOR_i1_U1 ( .A0_t (Ciphertext[34]), .B0_t (Ciphertext[35]), .Z0_t (SubCellInst_SboxInst_8_XX[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_8_XOR_i2_U1 ( .A0_t (Ciphertext[32]), .B0_t (Ciphertext[34]), .Z0_t (SubCellInst_SboxInst_8_XX[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_8_XOR0_U1 ( .A0_t (Ciphertext[33]), .B0_t (SubCellInst_SboxInst_8_XX[2]), .Z0_t (SubCellInst_SboxInst_8_Q0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_8_XOR1_U1 ( .A0_t (Ciphertext[33]), .B0_t (SubCellInst_SboxInst_8_XX[1]), .Z0_t (SubCellInst_SboxInst_8_Q1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_8_AND1_U1 ( .A0_t (Ciphertext[34]), .B0_t (SubCellInst_SboxInst_8_Q1), .Z0_t (SubCellInst_SboxInst_8_T0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_8_XOR2_U1 ( .A0_t (SubCellInst_SboxInst_8_Q0), .B0_t (SubCellInst_SboxInst_8_T0), .Z0_t (SubCellInst_SboxInst_8_Q2) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_8_AND2_U1 ( .A0_t (Ciphertext[33]), .B0_t (SubCellInst_SboxInst_8_Q2), .Z0_t (SubCellInst_SboxInst_8_T1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_8_XOR3_U1 ( .A0_t (Ciphertext[33]), .B0_t (Ciphertext[34]), .Z0_t (SubCellInst_SboxInst_8_Q4) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_8_AND3_U1 ( .A0_t (Ciphertext[34]), .B0_t (SubCellInst_SboxInst_8_Q4), .Z0_t (SubCellInst_SboxInst_8_T2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_8_XOR4_U1 ( .A0_t (SubCellInst_SboxInst_8_T1), .B0_t (SubCellInst_SboxInst_8_T2), .Z0_t (SubCellInst_SboxInst_8_L0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_8_XOR5_U1 ( .A0_t (SubCellInst_SboxInst_8_XX[2]), .B0_t (Ciphertext[34]), .Z0_t (SubCellInst_SboxInst_8_Q6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_8_XOR6_U1 ( .A0_t (SubCellInst_SboxInst_8_Q1), .B0_t (SubCellInst_SboxInst_8_Q6), .Z0_t (SubCellInst_SboxInst_8_L1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_8_XOR7_U1 ( .A0_t (SubCellInst_SboxInst_8_L1), .B0_t (SubCellInst_SboxInst_8_T2), .Z0_t (SubCellInst_SboxInst_8_Q7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_8_AND4_U1 ( .A0_t (SubCellInst_SboxInst_8_Q6), .B0_t (SubCellInst_SboxInst_8_Q7), .Z0_t (SubCellInst_SboxInst_8_T3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_8_XOR8_U1 ( .A0_t (Ciphertext[33]), .B0_t (Ciphertext[34]), .Z0_t (SubCellInst_SboxInst_8_L2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_8_XOR9_U1 ( .A0_t (SubCellInst_SboxInst_8_L0), .B0_t (SubCellInst_SboxInst_8_L2), .Z0_t (SubCellInst_SboxInst_8_YY_3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_8_XOR10_U1 ( .A0_t (SubCellInst_SboxInst_8_L0), .B0_t (SubCellInst_SboxInst_8_T3), .Z0_t (AddRoundConstantOutput[32]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_8_XOR11_U1 ( .A0_t (SubCellInst_SboxInst_8_XX[2]), .B0_t (SubCellInst_SboxInst_8_T0), .Z0_t (SubCellInst_SboxInst_8_L3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_8_XOR12_U1 ( .A0_t (SubCellInst_SboxInst_8_L3), .B0_t (SubCellInst_SboxInst_8_T2), .Z0_t (SubCellInst_SboxInst_8_YY[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_8_XOR13_U1 ( .A0_t (SubCellInst_SboxInst_8_XX[1]), .B0_t (SubCellInst_SboxInst_8_T2), .Z0_t (SubCellInst_SboxInst_8_YY[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_8_XOR_o1_U1 ( .A0_t (SubCellInst_SboxInst_8_YY[1]), .B0_t (SubCellInst_SboxInst_8_YY_3), .Z0_t (AddRoundConstantOutput[33]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_9_XOR_i1_U1 ( .A0_t (Ciphertext[38]), .B0_t (Ciphertext[39]), .Z0_t (SubCellInst_SboxInst_9_XX[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_9_XOR_i2_U1 ( .A0_t (Ciphertext[36]), .B0_t (Ciphertext[38]), .Z0_t (SubCellInst_SboxInst_9_XX[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_9_XOR0_U1 ( .A0_t (Ciphertext[37]), .B0_t (SubCellInst_SboxInst_9_XX[2]), .Z0_t (SubCellInst_SboxInst_9_Q0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_9_XOR1_U1 ( .A0_t (Ciphertext[37]), .B0_t (SubCellInst_SboxInst_9_XX[1]), .Z0_t (SubCellInst_SboxInst_9_Q1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_9_AND1_U1 ( .A0_t (Ciphertext[38]), .B0_t (SubCellInst_SboxInst_9_Q1), .Z0_t (SubCellInst_SboxInst_9_T0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_9_XOR2_U1 ( .A0_t (SubCellInst_SboxInst_9_Q0), .B0_t (SubCellInst_SboxInst_9_T0), .Z0_t (SubCellInst_SboxInst_9_Q2) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_9_AND2_U1 ( .A0_t (Ciphertext[37]), .B0_t (SubCellInst_SboxInst_9_Q2), .Z0_t (SubCellInst_SboxInst_9_T1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_9_XOR3_U1 ( .A0_t (Ciphertext[37]), .B0_t (Ciphertext[38]), .Z0_t (SubCellInst_SboxInst_9_Q4) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_9_AND3_U1 ( .A0_t (Ciphertext[38]), .B0_t (SubCellInst_SboxInst_9_Q4), .Z0_t (SubCellInst_SboxInst_9_T2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_9_XOR4_U1 ( .A0_t (SubCellInst_SboxInst_9_T1), .B0_t (SubCellInst_SboxInst_9_T2), .Z0_t (SubCellInst_SboxInst_9_L0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_9_XOR5_U1 ( .A0_t (SubCellInst_SboxInst_9_XX[2]), .B0_t (Ciphertext[38]), .Z0_t (SubCellInst_SboxInst_9_Q6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_9_XOR6_U1 ( .A0_t (SubCellInst_SboxInst_9_Q1), .B0_t (SubCellInst_SboxInst_9_Q6), .Z0_t (SubCellInst_SboxInst_9_L1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_9_XOR7_U1 ( .A0_t (SubCellInst_SboxInst_9_L1), .B0_t (SubCellInst_SboxInst_9_T2), .Z0_t (SubCellInst_SboxInst_9_Q7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_9_AND4_U1 ( .A0_t (SubCellInst_SboxInst_9_Q6), .B0_t (SubCellInst_SboxInst_9_Q7), .Z0_t (SubCellInst_SboxInst_9_T3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_9_XOR8_U1 ( .A0_t (Ciphertext[37]), .B0_t (Ciphertext[38]), .Z0_t (SubCellInst_SboxInst_9_L2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_9_XOR9_U1 ( .A0_t (SubCellInst_SboxInst_9_L0), .B0_t (SubCellInst_SboxInst_9_L2), .Z0_t (SubCellInst_SboxInst_9_YY_3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_9_XOR10_U1 ( .A0_t (SubCellInst_SboxInst_9_L0), .B0_t (SubCellInst_SboxInst_9_T3), .Z0_t (AddRoundConstantOutput[36]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_9_XOR11_U1 ( .A0_t (SubCellInst_SboxInst_9_XX[2]), .B0_t (SubCellInst_SboxInst_9_T0), .Z0_t (SubCellInst_SboxInst_9_L3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_9_XOR12_U1 ( .A0_t (SubCellInst_SboxInst_9_L3), .B0_t (SubCellInst_SboxInst_9_T2), .Z0_t (SubCellInst_SboxInst_9_YY[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_9_XOR13_U1 ( .A0_t (SubCellInst_SboxInst_9_XX[1]), .B0_t (SubCellInst_SboxInst_9_T2), .Z0_t (SubCellInst_SboxInst_9_YY[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_9_XOR_o1_U1 ( .A0_t (SubCellInst_SboxInst_9_YY[1]), .B0_t (SubCellInst_SboxInst_9_YY_3), .Z0_t (AddRoundConstantOutput[37]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_10_XOR_i1_U1 ( .A0_t (Ciphertext[42]), .B0_t (Ciphertext[43]), .Z0_t (SubCellInst_SboxInst_10_XX[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_10_XOR_i2_U1 ( .A0_t (Ciphertext[40]), .B0_t (Ciphertext[42]), .Z0_t (SubCellInst_SboxInst_10_XX[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_10_XOR0_U1 ( .A0_t (Ciphertext[41]), .B0_t (SubCellInst_SboxInst_10_XX[2]), .Z0_t (SubCellInst_SboxInst_10_Q0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_10_XOR1_U1 ( .A0_t (Ciphertext[41]), .B0_t (SubCellInst_SboxInst_10_XX[1]), .Z0_t (SubCellInst_SboxInst_10_Q1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_10_AND1_U1 ( .A0_t (Ciphertext[42]), .B0_t (SubCellInst_SboxInst_10_Q1), .Z0_t (SubCellInst_SboxInst_10_T0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_10_XOR2_U1 ( .A0_t (SubCellInst_SboxInst_10_Q0), .B0_t (SubCellInst_SboxInst_10_T0), .Z0_t (SubCellInst_SboxInst_10_Q2) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_10_AND2_U1 ( .A0_t (Ciphertext[41]), .B0_t (SubCellInst_SboxInst_10_Q2), .Z0_t (SubCellInst_SboxInst_10_T1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_10_XOR3_U1 ( .A0_t (Ciphertext[41]), .B0_t (Ciphertext[42]), .Z0_t (SubCellInst_SboxInst_10_Q4) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_10_AND3_U1 ( .A0_t (Ciphertext[42]), .B0_t (SubCellInst_SboxInst_10_Q4), .Z0_t (SubCellInst_SboxInst_10_T2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_10_XOR4_U1 ( .A0_t (SubCellInst_SboxInst_10_T1), .B0_t (SubCellInst_SboxInst_10_T2), .Z0_t (SubCellInst_SboxInst_10_L0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_10_XOR5_U1 ( .A0_t (SubCellInst_SboxInst_10_XX[2]), .B0_t (Ciphertext[42]), .Z0_t (SubCellInst_SboxInst_10_Q6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_10_XOR6_U1 ( .A0_t (SubCellInst_SboxInst_10_Q1), .B0_t (SubCellInst_SboxInst_10_Q6), .Z0_t (SubCellInst_SboxInst_10_L1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_10_XOR7_U1 ( .A0_t (SubCellInst_SboxInst_10_L1), .B0_t (SubCellInst_SboxInst_10_T2), .Z0_t (SubCellInst_SboxInst_10_Q7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_10_AND4_U1 ( .A0_t (SubCellInst_SboxInst_10_Q6), .B0_t (SubCellInst_SboxInst_10_Q7), .Z0_t (SubCellInst_SboxInst_10_T3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_10_XOR8_U1 ( .A0_t (Ciphertext[41]), .B0_t (Ciphertext[42]), .Z0_t (SubCellInst_SboxInst_10_L2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_10_XOR9_U1 ( .A0_t (SubCellInst_SboxInst_10_L0), .B0_t (SubCellInst_SboxInst_10_L2), .Z0_t (SubCellInst_SboxInst_10_YY_3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_10_XOR10_U1 ( .A0_t (SubCellInst_SboxInst_10_L0), .B0_t (SubCellInst_SboxInst_10_T3), .Z0_t (AddRoundConstantOutput[40]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_10_XOR11_U1 ( .A0_t (SubCellInst_SboxInst_10_XX[2]), .B0_t (SubCellInst_SboxInst_10_T0), .Z0_t (SubCellInst_SboxInst_10_L3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_10_XOR12_U1 ( .A0_t (SubCellInst_SboxInst_10_L3), .B0_t (SubCellInst_SboxInst_10_T2), .Z0_t (SubCellInst_SboxInst_10_YY[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_10_XOR13_U1 ( .A0_t (SubCellInst_SboxInst_10_XX[1]), .B0_t (SubCellInst_SboxInst_10_T2), .Z0_t (SubCellInst_SboxInst_10_YY[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_10_XOR_o1_U1 ( .A0_t (SubCellInst_SboxInst_10_YY[1]), .B0_t (SubCellInst_SboxInst_10_YY_3), .Z0_t (AddRoundConstantOutput[41]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_11_XOR_i1_U1 ( .A0_t (Ciphertext[46]), .B0_t (Ciphertext[47]), .Z0_t (SubCellInst_SboxInst_11_XX[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_11_XOR_i2_U1 ( .A0_t (Ciphertext[44]), .B0_t (Ciphertext[46]), .Z0_t (SubCellInst_SboxInst_11_XX[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_11_XOR0_U1 ( .A0_t (Ciphertext[45]), .B0_t (SubCellInst_SboxInst_11_XX[2]), .Z0_t (SubCellInst_SboxInst_11_Q0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_11_XOR1_U1 ( .A0_t (Ciphertext[45]), .B0_t (SubCellInst_SboxInst_11_XX[1]), .Z0_t (SubCellInst_SboxInst_11_Q1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_11_AND1_U1 ( .A0_t (Ciphertext[46]), .B0_t (SubCellInst_SboxInst_11_Q1), .Z0_t (SubCellInst_SboxInst_11_T0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_11_XOR2_U1 ( .A0_t (SubCellInst_SboxInst_11_Q0), .B0_t (SubCellInst_SboxInst_11_T0), .Z0_t (SubCellInst_SboxInst_11_Q2) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_11_AND2_U1 ( .A0_t (Ciphertext[45]), .B0_t (SubCellInst_SboxInst_11_Q2), .Z0_t (SubCellInst_SboxInst_11_T1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_11_XOR3_U1 ( .A0_t (Ciphertext[45]), .B0_t (Ciphertext[46]), .Z0_t (SubCellInst_SboxInst_11_Q4) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_11_AND3_U1 ( .A0_t (Ciphertext[46]), .B0_t (SubCellInst_SboxInst_11_Q4), .Z0_t (SubCellInst_SboxInst_11_T2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_11_XOR4_U1 ( .A0_t (SubCellInst_SboxInst_11_T1), .B0_t (SubCellInst_SboxInst_11_T2), .Z0_t (SubCellInst_SboxInst_11_L0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_11_XOR5_U1 ( .A0_t (SubCellInst_SboxInst_11_XX[2]), .B0_t (Ciphertext[46]), .Z0_t (SubCellInst_SboxInst_11_Q6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_11_XOR6_U1 ( .A0_t (SubCellInst_SboxInst_11_Q1), .B0_t (SubCellInst_SboxInst_11_Q6), .Z0_t (SubCellInst_SboxInst_11_L1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_11_XOR7_U1 ( .A0_t (SubCellInst_SboxInst_11_L1), .B0_t (SubCellInst_SboxInst_11_T2), .Z0_t (SubCellInst_SboxInst_11_Q7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_11_AND4_U1 ( .A0_t (SubCellInst_SboxInst_11_Q6), .B0_t (SubCellInst_SboxInst_11_Q7), .Z0_t (SubCellInst_SboxInst_11_T3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_11_XOR8_U1 ( .A0_t (Ciphertext[45]), .B0_t (Ciphertext[46]), .Z0_t (SubCellInst_SboxInst_11_L2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_11_XOR9_U1 ( .A0_t (SubCellInst_SboxInst_11_L0), .B0_t (SubCellInst_SboxInst_11_L2), .Z0_t (SubCellInst_SboxInst_11_YY_3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_11_XOR10_U1 ( .A0_t (SubCellInst_SboxInst_11_L0), .B0_t (SubCellInst_SboxInst_11_T3), .Z0_t (SubCellOutput[44]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_11_XOR11_U1 ( .A0_t (SubCellInst_SboxInst_11_XX[2]), .B0_t (SubCellInst_SboxInst_11_T0), .Z0_t (SubCellInst_SboxInst_11_L3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_11_XOR12_U1 ( .A0_t (SubCellInst_SboxInst_11_L3), .B0_t (SubCellInst_SboxInst_11_T2), .Z0_t (SubCellInst_SboxInst_11_YY[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_11_XOR13_U1 ( .A0_t (SubCellInst_SboxInst_11_XX[1]), .B0_t (SubCellInst_SboxInst_11_T2), .Z0_t (SubCellInst_SboxInst_11_YY[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_11_XOR_o1_U1 ( .A0_t (SubCellInst_SboxInst_11_YY[1]), .B0_t (SubCellInst_SboxInst_11_YY_3), .Z0_t (SubCellOutput[45]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_12_XOR_i1_U1 ( .A0_t (Ciphertext[50]), .B0_t (Ciphertext[51]), .Z0_t (SubCellInst_SboxInst_12_XX[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_12_XOR_i2_U1 ( .A0_t (Ciphertext[48]), .B0_t (Ciphertext[50]), .Z0_t (SubCellInst_SboxInst_12_XX[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_12_XOR0_U1 ( .A0_t (Ciphertext[49]), .B0_t (SubCellInst_SboxInst_12_XX[2]), .Z0_t (SubCellInst_SboxInst_12_Q0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_12_XOR1_U1 ( .A0_t (Ciphertext[49]), .B0_t (SubCellInst_SboxInst_12_XX[1]), .Z0_t (SubCellInst_SboxInst_12_Q1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_12_AND1_U1 ( .A0_t (Ciphertext[50]), .B0_t (SubCellInst_SboxInst_12_Q1), .Z0_t (SubCellInst_SboxInst_12_T0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_12_XOR2_U1 ( .A0_t (SubCellInst_SboxInst_12_Q0), .B0_t (SubCellInst_SboxInst_12_T0), .Z0_t (SubCellInst_SboxInst_12_Q2) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_12_AND2_U1 ( .A0_t (Ciphertext[49]), .B0_t (SubCellInst_SboxInst_12_Q2), .Z0_t (SubCellInst_SboxInst_12_T1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_12_XOR3_U1 ( .A0_t (Ciphertext[49]), .B0_t (Ciphertext[50]), .Z0_t (SubCellInst_SboxInst_12_Q4) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_12_AND3_U1 ( .A0_t (Ciphertext[50]), .B0_t (SubCellInst_SboxInst_12_Q4), .Z0_t (SubCellInst_SboxInst_12_T2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_12_XOR4_U1 ( .A0_t (SubCellInst_SboxInst_12_T1), .B0_t (SubCellInst_SboxInst_12_T2), .Z0_t (SubCellInst_SboxInst_12_L0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_12_XOR5_U1 ( .A0_t (SubCellInst_SboxInst_12_XX[2]), .B0_t (Ciphertext[50]), .Z0_t (SubCellInst_SboxInst_12_Q6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_12_XOR6_U1 ( .A0_t (SubCellInst_SboxInst_12_Q1), .B0_t (SubCellInst_SboxInst_12_Q6), .Z0_t (SubCellInst_SboxInst_12_L1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_12_XOR7_U1 ( .A0_t (SubCellInst_SboxInst_12_L1), .B0_t (SubCellInst_SboxInst_12_T2), .Z0_t (SubCellInst_SboxInst_12_Q7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_12_AND4_U1 ( .A0_t (SubCellInst_SboxInst_12_Q6), .B0_t (SubCellInst_SboxInst_12_Q7), .Z0_t (SubCellInst_SboxInst_12_T3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_12_XOR8_U1 ( .A0_t (Ciphertext[49]), .B0_t (Ciphertext[50]), .Z0_t (SubCellInst_SboxInst_12_L2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_12_XOR9_U1 ( .A0_t (SubCellInst_SboxInst_12_L0), .B0_t (SubCellInst_SboxInst_12_L2), .Z0_t (SubCellInst_SboxInst_12_YY_3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_12_XOR10_U1 ( .A0_t (SubCellInst_SboxInst_12_L0), .B0_t (SubCellInst_SboxInst_12_T3), .Z0_t (AddRoundConstantOutput[48]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_12_XOR11_U1 ( .A0_t (SubCellInst_SboxInst_12_XX[2]), .B0_t (SubCellInst_SboxInst_12_T0), .Z0_t (SubCellInst_SboxInst_12_L3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_12_XOR12_U1 ( .A0_t (SubCellInst_SboxInst_12_L3), .B0_t (SubCellInst_SboxInst_12_T2), .Z0_t (SubCellInst_SboxInst_12_YY[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_12_XOR13_U1 ( .A0_t (SubCellInst_SboxInst_12_XX[1]), .B0_t (SubCellInst_SboxInst_12_T2), .Z0_t (SubCellInst_SboxInst_12_YY[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_12_XOR_o1_U1 ( .A0_t (SubCellInst_SboxInst_12_YY[1]), .B0_t (SubCellInst_SboxInst_12_YY_3), .Z0_t (AddRoundConstantOutput[49]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_13_XOR_i1_U1 ( .A0_t (Ciphertext[54]), .B0_t (Ciphertext[55]), .Z0_t (SubCellInst_SboxInst_13_XX[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_13_XOR_i2_U1 ( .A0_t (Ciphertext[52]), .B0_t (Ciphertext[54]), .Z0_t (SubCellInst_SboxInst_13_XX[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_13_XOR0_U1 ( .A0_t (Ciphertext[53]), .B0_t (SubCellInst_SboxInst_13_XX[2]), .Z0_t (SubCellInst_SboxInst_13_Q0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_13_XOR1_U1 ( .A0_t (Ciphertext[53]), .B0_t (SubCellInst_SboxInst_13_XX[1]), .Z0_t (SubCellInst_SboxInst_13_Q1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_13_AND1_U1 ( .A0_t (Ciphertext[54]), .B0_t (SubCellInst_SboxInst_13_Q1), .Z0_t (SubCellInst_SboxInst_13_T0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_13_XOR2_U1 ( .A0_t (SubCellInst_SboxInst_13_Q0), .B0_t (SubCellInst_SboxInst_13_T0), .Z0_t (SubCellInst_SboxInst_13_Q2) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_13_AND2_U1 ( .A0_t (Ciphertext[53]), .B0_t (SubCellInst_SboxInst_13_Q2), .Z0_t (SubCellInst_SboxInst_13_T1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_13_XOR3_U1 ( .A0_t (Ciphertext[53]), .B0_t (Ciphertext[54]), .Z0_t (SubCellInst_SboxInst_13_Q4) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_13_AND3_U1 ( .A0_t (Ciphertext[54]), .B0_t (SubCellInst_SboxInst_13_Q4), .Z0_t (SubCellInst_SboxInst_13_T2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_13_XOR4_U1 ( .A0_t (SubCellInst_SboxInst_13_T1), .B0_t (SubCellInst_SboxInst_13_T2), .Z0_t (SubCellInst_SboxInst_13_L0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_13_XOR5_U1 ( .A0_t (SubCellInst_SboxInst_13_XX[2]), .B0_t (Ciphertext[54]), .Z0_t (SubCellInst_SboxInst_13_Q6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_13_XOR6_U1 ( .A0_t (SubCellInst_SboxInst_13_Q1), .B0_t (SubCellInst_SboxInst_13_Q6), .Z0_t (SubCellInst_SboxInst_13_L1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_13_XOR7_U1 ( .A0_t (SubCellInst_SboxInst_13_L1), .B0_t (SubCellInst_SboxInst_13_T2), .Z0_t (SubCellInst_SboxInst_13_Q7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_13_AND4_U1 ( .A0_t (SubCellInst_SboxInst_13_Q6), .B0_t (SubCellInst_SboxInst_13_Q7), .Z0_t (SubCellInst_SboxInst_13_T3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_13_XOR8_U1 ( .A0_t (Ciphertext[53]), .B0_t (Ciphertext[54]), .Z0_t (SubCellInst_SboxInst_13_L2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_13_XOR9_U1 ( .A0_t (SubCellInst_SboxInst_13_L0), .B0_t (SubCellInst_SboxInst_13_L2), .Z0_t (SubCellInst_SboxInst_13_YY_3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_13_XOR10_U1 ( .A0_t (SubCellInst_SboxInst_13_L0), .B0_t (SubCellInst_SboxInst_13_T3), .Z0_t (AddRoundConstantOutput[52]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_13_XOR11_U1 ( .A0_t (SubCellInst_SboxInst_13_XX[2]), .B0_t (SubCellInst_SboxInst_13_T0), .Z0_t (SubCellInst_SboxInst_13_L3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_13_XOR12_U1 ( .A0_t (SubCellInst_SboxInst_13_L3), .B0_t (SubCellInst_SboxInst_13_T2), .Z0_t (SubCellInst_SboxInst_13_YY[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_13_XOR13_U1 ( .A0_t (SubCellInst_SboxInst_13_XX[1]), .B0_t (SubCellInst_SboxInst_13_T2), .Z0_t (SubCellInst_SboxInst_13_YY[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_13_XOR_o1_U1 ( .A0_t (SubCellInst_SboxInst_13_YY[1]), .B0_t (SubCellInst_SboxInst_13_YY_3), .Z0_t (AddRoundConstantOutput[53]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_14_XOR_i1_U1 ( .A0_t (Ciphertext[58]), .B0_t (Ciphertext[59]), .Z0_t (SubCellInst_SboxInst_14_XX[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_14_XOR_i2_U1 ( .A0_t (Ciphertext[56]), .B0_t (Ciphertext[58]), .Z0_t (SubCellInst_SboxInst_14_XX[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_14_XOR0_U1 ( .A0_t (Ciphertext[57]), .B0_t (SubCellInst_SboxInst_14_XX[2]), .Z0_t (SubCellInst_SboxInst_14_Q0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_14_XOR1_U1 ( .A0_t (Ciphertext[57]), .B0_t (SubCellInst_SboxInst_14_XX[1]), .Z0_t (SubCellInst_SboxInst_14_Q1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_14_AND1_U1 ( .A0_t (Ciphertext[58]), .B0_t (SubCellInst_SboxInst_14_Q1), .Z0_t (SubCellInst_SboxInst_14_T0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_14_XOR2_U1 ( .A0_t (SubCellInst_SboxInst_14_Q0), .B0_t (SubCellInst_SboxInst_14_T0), .Z0_t (SubCellInst_SboxInst_14_Q2) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_14_AND2_U1 ( .A0_t (Ciphertext[57]), .B0_t (SubCellInst_SboxInst_14_Q2), .Z0_t (SubCellInst_SboxInst_14_T1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_14_XOR3_U1 ( .A0_t (Ciphertext[57]), .B0_t (Ciphertext[58]), .Z0_t (SubCellInst_SboxInst_14_Q4) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_14_AND3_U1 ( .A0_t (Ciphertext[58]), .B0_t (SubCellInst_SboxInst_14_Q4), .Z0_t (SubCellInst_SboxInst_14_T2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_14_XOR4_U1 ( .A0_t (SubCellInst_SboxInst_14_T1), .B0_t (SubCellInst_SboxInst_14_T2), .Z0_t (SubCellInst_SboxInst_14_L0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_14_XOR5_U1 ( .A0_t (SubCellInst_SboxInst_14_XX[2]), .B0_t (Ciphertext[58]), .Z0_t (SubCellInst_SboxInst_14_Q6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_14_XOR6_U1 ( .A0_t (SubCellInst_SboxInst_14_Q1), .B0_t (SubCellInst_SboxInst_14_Q6), .Z0_t (SubCellInst_SboxInst_14_L1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_14_XOR7_U1 ( .A0_t (SubCellInst_SboxInst_14_L1), .B0_t (SubCellInst_SboxInst_14_T2), .Z0_t (SubCellInst_SboxInst_14_Q7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_14_AND4_U1 ( .A0_t (SubCellInst_SboxInst_14_Q6), .B0_t (SubCellInst_SboxInst_14_Q7), .Z0_t (SubCellInst_SboxInst_14_T3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_14_XOR8_U1 ( .A0_t (Ciphertext[57]), .B0_t (Ciphertext[58]), .Z0_t (SubCellInst_SboxInst_14_L2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_14_XOR9_U1 ( .A0_t (SubCellInst_SboxInst_14_L0), .B0_t (SubCellInst_SboxInst_14_L2), .Z0_t (SubCellInst_SboxInst_14_YY_3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_14_XOR10_U1 ( .A0_t (SubCellInst_SboxInst_14_L0), .B0_t (SubCellInst_SboxInst_14_T3), .Z0_t (AddRoundConstantOutput[56]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_14_XOR11_U1 ( .A0_t (SubCellInst_SboxInst_14_XX[2]), .B0_t (SubCellInst_SboxInst_14_T0), .Z0_t (SubCellInst_SboxInst_14_L3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_14_XOR12_U1 ( .A0_t (SubCellInst_SboxInst_14_L3), .B0_t (SubCellInst_SboxInst_14_T2), .Z0_t (SubCellInst_SboxInst_14_YY[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_14_XOR13_U1 ( .A0_t (SubCellInst_SboxInst_14_XX[1]), .B0_t (SubCellInst_SboxInst_14_T2), .Z0_t (SubCellInst_SboxInst_14_YY[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_14_XOR_o1_U1 ( .A0_t (SubCellInst_SboxInst_14_YY[1]), .B0_t (SubCellInst_SboxInst_14_YY_3), .Z0_t (AddRoundConstantOutput[57]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_15_XOR_i1_U1 ( .A0_t (Ciphertext[62]), .B0_t (Ciphertext[63]), .Z0_t (SubCellInst_SboxInst_15_XX[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_15_XOR_i2_U1 ( .A0_t (Ciphertext[60]), .B0_t (Ciphertext[62]), .Z0_t (SubCellInst_SboxInst_15_XX[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_15_XOR0_U1 ( .A0_t (Ciphertext[61]), .B0_t (SubCellInst_SboxInst_15_XX[2]), .Z0_t (SubCellInst_SboxInst_15_Q0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_15_XOR1_U1 ( .A0_t (Ciphertext[61]), .B0_t (SubCellInst_SboxInst_15_XX[1]), .Z0_t (SubCellInst_SboxInst_15_Q1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_15_AND1_U1 ( .A0_t (Ciphertext[62]), .B0_t (SubCellInst_SboxInst_15_Q1), .Z0_t (SubCellInst_SboxInst_15_T0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_15_XOR2_U1 ( .A0_t (SubCellInst_SboxInst_15_Q0), .B0_t (SubCellInst_SboxInst_15_T0), .Z0_t (SubCellInst_SboxInst_15_Q2) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_15_AND2_U1 ( .A0_t (Ciphertext[61]), .B0_t (SubCellInst_SboxInst_15_Q2), .Z0_t (SubCellInst_SboxInst_15_T1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_15_XOR3_U1 ( .A0_t (Ciphertext[61]), .B0_t (Ciphertext[62]), .Z0_t (SubCellInst_SboxInst_15_Q4) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_15_AND3_U1 ( .A0_t (Ciphertext[62]), .B0_t (SubCellInst_SboxInst_15_Q4), .Z0_t (SubCellInst_SboxInst_15_T2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_15_XOR4_U1 ( .A0_t (SubCellInst_SboxInst_15_T1), .B0_t (SubCellInst_SboxInst_15_T2), .Z0_t (SubCellInst_SboxInst_15_L0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_15_XOR5_U1 ( .A0_t (SubCellInst_SboxInst_15_XX[2]), .B0_t (Ciphertext[62]), .Z0_t (SubCellInst_SboxInst_15_Q6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_15_XOR6_U1 ( .A0_t (SubCellInst_SboxInst_15_Q1), .B0_t (SubCellInst_SboxInst_15_Q6), .Z0_t (SubCellInst_SboxInst_15_L1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_15_XOR7_U1 ( .A0_t (SubCellInst_SboxInst_15_L1), .B0_t (SubCellInst_SboxInst_15_T2), .Z0_t (SubCellInst_SboxInst_15_Q7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_15_AND4_U1 ( .A0_t (SubCellInst_SboxInst_15_Q6), .B0_t (SubCellInst_SboxInst_15_Q7), .Z0_t (SubCellInst_SboxInst_15_T3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_15_XOR8_U1 ( .A0_t (Ciphertext[61]), .B0_t (Ciphertext[62]), .Z0_t (SubCellInst_SboxInst_15_L2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_15_XOR9_U1 ( .A0_t (SubCellInst_SboxInst_15_L0), .B0_t (SubCellInst_SboxInst_15_L2), .Z0_t (SubCellInst_SboxInst_15_YY_3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_15_XOR10_U1 ( .A0_t (SubCellInst_SboxInst_15_L0), .B0_t (SubCellInst_SboxInst_15_T3), .Z0_t (SubCellOutput[60]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_15_XOR11_U1 ( .A0_t (SubCellInst_SboxInst_15_XX[2]), .B0_t (SubCellInst_SboxInst_15_T0), .Z0_t (SubCellInst_SboxInst_15_L3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_15_XOR12_U1 ( .A0_t (SubCellInst_SboxInst_15_L3), .B0_t (SubCellInst_SboxInst_15_T2), .Z0_t (SubCellInst_SboxInst_15_YY[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) SubCellInst_SboxInst_15_XOR13_U1 ( .A0_t (SubCellInst_SboxInst_15_XX[1]), .B0_t (SubCellInst_SboxInst_15_T2), .Z0_t (SubCellInst_SboxInst_15_YY[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) SubCellInst_SboxInst_15_XOR_o1_U1 ( .A0_t (SubCellInst_SboxInst_15_YY[1]), .B0_t (SubCellInst_SboxInst_15_YY_3), .Z0_t (SubCellOutput[61]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddConstXOR_AddConstXOR_XORInst_0_0_U1 ( .A0_t (SubCellOutput[60]), .B0_t (FSMUpdate[1]), .Z0_t (AddRoundConstantOutput[60]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddConstXOR_AddConstXOR_XORInst_0_1_U1 ( .A0_t (SubCellOutput[61]), .B0_t (FSM[1]), .Z0_t (AddRoundConstantOutput[61]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddConstXOR_AddConstXOR_XORInst_0_2_U1 ( .A0_t (SubCellInst_SboxInst_15_YY[0]), .B0_t (FSMUpdate[3]), .Z0_t (AddRoundConstantOutput[62]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddConstXOR_AddConstXOR_XORInst_0_3_U1 ( .A0_t (SubCellInst_SboxInst_15_YY[1]), .B0_t (FSMUpdate[4]), .Z0_t (AddRoundConstantOutput[63]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddConstXOR_AddConstXOR_XORInst_1_0_U1 ( .A0_t (SubCellOutput[44]), .B0_t (FSM[4]), .Z0_t (AddRoundConstantOutput[44]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddConstXOR_AddConstXOR_XORInst_1_1_U1 ( .A0_t (SubCellOutput[45]), .B0_t (FSM[5]), .Z0_t (AddRoundConstantOutput[45]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddRoundTweakeyXOR_XORInst_0_0_U1 ( .A0_t (AddRoundConstantOutput[32]), .B0_t (TweakeyGeneration_key_Feedback[0]), .Z0_t (ShiftRowsOutput[44]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddRoundTweakeyXOR_XORInst_0_1_U1 ( .A0_t (AddRoundConstantOutput[33]), .B0_t (TweakeyGeneration_key_Feedback[1]), .Z0_t (ShiftRowsOutput[45]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddRoundTweakeyXOR_XORInst_0_2_U1 ( .A0_t (SubCellInst_SboxInst_8_YY[0]), .B0_t (TweakeyGeneration_key_Feedback[2]), .Z0_t (ShiftRowsOutput[46]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddRoundTweakeyXOR_XORInst_0_3_U1 ( .A0_t (SubCellInst_SboxInst_8_YY[1]), .B0_t (TweakeyGeneration_key_Feedback[3]), .Z0_t (ShiftRowsOutput[47]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddRoundTweakeyXOR_XORInst_1_0_U1 ( .A0_t (AddRoundConstantOutput[36]), .B0_t (TweakeyGeneration_key_Feedback[4]), .Z0_t (ShiftRowsOutput[32]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddRoundTweakeyXOR_XORInst_1_1_U1 ( .A0_t (AddRoundConstantOutput[37]), .B0_t (TweakeyGeneration_key_Feedback[5]), .Z0_t (ShiftRowsOutput[33]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddRoundTweakeyXOR_XORInst_1_2_U1 ( .A0_t (SubCellInst_SboxInst_9_YY[0]), .B0_t (TweakeyGeneration_key_Feedback[6]), .Z0_t (ShiftRowsOutput[34]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddRoundTweakeyXOR_XORInst_1_3_U1 ( .A0_t (SubCellInst_SboxInst_9_YY[1]), .B0_t (TweakeyGeneration_key_Feedback[7]), .Z0_t (ShiftRowsOutput[35]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddRoundTweakeyXOR_XORInst_2_0_U1 ( .A0_t (AddRoundConstantOutput[40]), .B0_t (TweakeyGeneration_key_Feedback[8]), .Z0_t (ShiftRowsOutput[36]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddRoundTweakeyXOR_XORInst_2_1_U1 ( .A0_t (AddRoundConstantOutput[41]), .B0_t (TweakeyGeneration_key_Feedback[9]), .Z0_t (ShiftRowsOutput[37]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddRoundTweakeyXOR_XORInst_2_2_U1 ( .A0_t (SubCellInst_SboxInst_10_YY[0]), .B0_t (TweakeyGeneration_key_Feedback[10]), .Z0_t (ShiftRowsOutput[38]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddRoundTweakeyXOR_XORInst_2_3_U1 ( .A0_t (SubCellInst_SboxInst_10_YY[1]), .B0_t (TweakeyGeneration_key_Feedback[11]), .Z0_t (ShiftRowsOutput[39]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddRoundTweakeyXOR_XORInst_3_0_U1 ( .A0_t (AddRoundConstantOutput[44]), .B0_t (TweakeyGeneration_key_Feedback[12]), .Z0_t (ShiftRowsOutput[40]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddRoundTweakeyXOR_XORInst_3_1_U1 ( .A0_t (AddRoundConstantOutput[45]), .B0_t (TweakeyGeneration_key_Feedback[13]), .Z0_t (ShiftRowsOutput[41]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddRoundTweakeyXOR_XORInst_3_2_U1 ( .A0_t (SubCellInst_SboxInst_11_YY[0]), .B0_t (TweakeyGeneration_key_Feedback[14]), .Z0_t (ShiftRowsOutput[42]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddRoundTweakeyXOR_XORInst_3_3_U1 ( .A0_t (SubCellInst_SboxInst_11_YY[1]), .B0_t (TweakeyGeneration_key_Feedback[15]), .Z0_t (ShiftRowsOutput[43]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddRoundTweakeyXOR_XORInst_4_0_U1 ( .A0_t (AddRoundConstantOutput[48]), .B0_t (TweakeyGeneration_key_Feedback[16]), .Z0_t (MCOutput[32]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddRoundTweakeyXOR_XORInst_4_1_U1 ( .A0_t (AddRoundConstantOutput[49]), .B0_t (TweakeyGeneration_key_Feedback[17]), .Z0_t (MCOutput[33]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddRoundTweakeyXOR_XORInst_4_2_U1 ( .A0_t (SubCellInst_SboxInst_12_YY[0]), .B0_t (TweakeyGeneration_key_Feedback[18]), .Z0_t (MCOutput[34]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddRoundTweakeyXOR_XORInst_4_3_U1 ( .A0_t (SubCellInst_SboxInst_12_YY[1]), .B0_t (TweakeyGeneration_key_Feedback[19]), .Z0_t (MCOutput[35]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddRoundTweakeyXOR_XORInst_5_0_U1 ( .A0_t (AddRoundConstantOutput[52]), .B0_t (TweakeyGeneration_key_Feedback[20]), .Z0_t (MCOutput[36]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddRoundTweakeyXOR_XORInst_5_1_U1 ( .A0_t (AddRoundConstantOutput[53]), .B0_t (TweakeyGeneration_key_Feedback[21]), .Z0_t (MCOutput[37]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddRoundTweakeyXOR_XORInst_5_2_U1 ( .A0_t (SubCellInst_SboxInst_13_YY[0]), .B0_t (TweakeyGeneration_key_Feedback[22]), .Z0_t (MCOutput[38]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddRoundTweakeyXOR_XORInst_5_3_U1 ( .A0_t (SubCellInst_SboxInst_13_YY[1]), .B0_t (TweakeyGeneration_key_Feedback[23]), .Z0_t (MCOutput[39]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddRoundTweakeyXOR_XORInst_6_0_U1 ( .A0_t (AddRoundConstantOutput[56]), .B0_t (TweakeyGeneration_key_Feedback[24]), .Z0_t (MCOutput[40]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddRoundTweakeyXOR_XORInst_6_1_U1 ( .A0_t (AddRoundConstantOutput[57]), .B0_t (TweakeyGeneration_key_Feedback[25]), .Z0_t (MCOutput[41]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddRoundTweakeyXOR_XORInst_6_2_U1 ( .A0_t (SubCellInst_SboxInst_14_YY[0]), .B0_t (TweakeyGeneration_key_Feedback[26]), .Z0_t (MCOutput[42]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddRoundTweakeyXOR_XORInst_6_3_U1 ( .A0_t (SubCellInst_SboxInst_14_YY[1]), .B0_t (TweakeyGeneration_key_Feedback[27]), .Z0_t (MCOutput[43]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddRoundTweakeyXOR_XORInst_7_0_U1 ( .A0_t (AddRoundConstantOutput[60]), .B0_t (TweakeyGeneration_key_Feedback[28]), .Z0_t (MCOutput[44]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddRoundTweakeyXOR_XORInst_7_1_U1 ( .A0_t (AddRoundConstantOutput[61]), .B0_t (TweakeyGeneration_key_Feedback[29]), .Z0_t (MCOutput[45]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddRoundTweakeyXOR_XORInst_7_2_U1 ( .A0_t (AddRoundConstantOutput[62]), .B0_t (TweakeyGeneration_key_Feedback[30]), .Z0_t (MCOutput[46]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) AddRoundTweakeyXOR_XORInst_7_3_U1 ( .A0_t (AddRoundConstantOutput[63]), .B0_t (TweakeyGeneration_key_Feedback[31]), .Z0_t (MCOutput[47]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_MCR0_XORInst_0_0_U2 ( .A0_t (MCInst_MCR0_XORInst_0_0_n1), .B0_t (ShiftRowsOutput[0]), .Z0_t (MCOutput[48]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_MCR0_XORInst_0_0_U1 ( .A0_t (MCOutput[32]), .B0_t (ShiftRowsOutput[16]), .Z0_t (MCInst_MCR0_XORInst_0_0_n1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_MCR0_XORInst_0_1_U2 ( .A0_t (MCInst_MCR0_XORInst_0_1_n1), .B0_t (ShiftRowsOutput[1]), .Z0_t (MCOutput[49]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_MCR0_XORInst_0_1_U1 ( .A0_t (MCOutput[33]), .B0_t (ShiftRowsOutput[17]), .Z0_t (MCInst_MCR0_XORInst_0_1_n1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) MCInst_MCR0_XORInst_0_2_U2 ( .A0_t (MCInst_MCR0_XORInst_0_2_n1), .B0_t (SubCellInst_SboxInst_3_YY[0]), .Z0_t (MCOutput[50]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) MCInst_MCR0_XORInst_0_2_U1 ( .A0_t (MCOutput[34]), .B0_t (SubCellInst_SboxInst_6_YY[0]), .Z0_t (MCInst_MCR0_XORInst_0_2_n1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) MCInst_MCR0_XORInst_0_3_U2 ( .A0_t (MCInst_MCR0_XORInst_0_3_n1), .B0_t (SubCellInst_SboxInst_3_YY[1]), .Z0_t (MCOutput[51]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) MCInst_MCR0_XORInst_0_3_U1 ( .A0_t (MCOutput[35]), .B0_t (SubCellInst_SboxInst_6_YY[1]), .Z0_t (MCInst_MCR0_XORInst_0_3_n1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_MCR0_XORInst_1_0_U2 ( .A0_t (MCInst_MCR0_XORInst_1_0_n1), .B0_t (ShiftRowsOutput[4]), .Z0_t (MCOutput[52]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_MCR0_XORInst_1_0_U1 ( .A0_t (MCOutput[36]), .B0_t (ShiftRowsOutput[20]), .Z0_t (MCInst_MCR0_XORInst_1_0_n1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_MCR0_XORInst_1_1_U2 ( .A0_t (MCInst_MCR0_XORInst_1_1_n1), .B0_t (ShiftRowsOutput[5]), .Z0_t (MCOutput[53]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) MCInst_MCR0_XORInst_1_1_U1 ( .A0_t (MCOutput[37]), .B0_t (SubCellOutput[29]), .Z0_t (MCInst_MCR0_XORInst_1_1_n1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) MCInst_MCR0_XORInst_1_2_U2 ( .A0_t (MCInst_MCR0_XORInst_1_2_n1), .B0_t (SubCellInst_SboxInst_0_YY[0]), .Z0_t (MCOutput[54]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) MCInst_MCR0_XORInst_1_2_U1 ( .A0_t (MCOutput[38]), .B0_t (SubCellInst_SboxInst_7_YY[0]), .Z0_t (MCInst_MCR0_XORInst_1_2_n1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) MCInst_MCR0_XORInst_1_3_U2 ( .A0_t (MCInst_MCR0_XORInst_1_3_n1), .B0_t (SubCellInst_SboxInst_0_YY[1]), .Z0_t (MCOutput[55]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) MCInst_MCR0_XORInst_1_3_U1 ( .A0_t (MCOutput[39]), .B0_t (SubCellInst_SboxInst_7_YY[1]), .Z0_t (MCInst_MCR0_XORInst_1_3_n1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_MCR0_XORInst_2_0_U2 ( .A0_t (MCInst_MCR0_XORInst_2_0_n1), .B0_t (ShiftRowsOutput[8]), .Z0_t (MCOutput[56]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_MCR0_XORInst_2_0_U1 ( .A0_t (MCOutput[40]), .B0_t (ShiftRowsOutput[24]), .Z0_t (MCInst_MCR0_XORInst_2_0_n1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_MCR0_XORInst_2_1_U2 ( .A0_t (MCInst_MCR0_XORInst_2_1_n1), .B0_t (ShiftRowsOutput[9]), .Z0_t (MCOutput[57]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_MCR0_XORInst_2_1_U1 ( .A0_t (MCOutput[41]), .B0_t (ShiftRowsOutput[25]), .Z0_t (MCInst_MCR0_XORInst_2_1_n1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) MCInst_MCR0_XORInst_2_2_U2 ( .A0_t (MCInst_MCR0_XORInst_2_2_n1), .B0_t (SubCellInst_SboxInst_1_YY[0]), .Z0_t (MCOutput[58]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) MCInst_MCR0_XORInst_2_2_U1 ( .A0_t (MCOutput[42]), .B0_t (SubCellInst_SboxInst_4_YY[0]), .Z0_t (MCInst_MCR0_XORInst_2_2_n1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) MCInst_MCR0_XORInst_2_3_U2 ( .A0_t (MCInst_MCR0_XORInst_2_3_n1), .B0_t (SubCellInst_SboxInst_1_YY[1]), .Z0_t (MCOutput[59]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) MCInst_MCR0_XORInst_2_3_U1 ( .A0_t (MCOutput[43]), .B0_t (SubCellInst_SboxInst_4_YY[1]), .Z0_t (MCInst_MCR0_XORInst_2_3_n1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_MCR0_XORInst_3_0_U2 ( .A0_t (MCInst_MCR0_XORInst_3_0_n1), .B0_t (ShiftRowsOutput[12]), .Z0_t (MCOutput[60]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_MCR0_XORInst_3_0_U1 ( .A0_t (MCOutput[44]), .B0_t (ShiftRowsOutput[28]), .Z0_t (MCInst_MCR0_XORInst_3_0_n1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_MCR0_XORInst_3_1_U2 ( .A0_t (MCInst_MCR0_XORInst_3_1_n1), .B0_t (ShiftRowsOutput[13]), .Z0_t (MCOutput[61]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MCInst_MCR0_XORInst_3_1_U1 ( .A0_t (MCOutput[45]), .B0_t (ShiftRowsOutput[29]), .Z0_t (MCInst_MCR0_XORInst_3_1_n1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) MCInst_MCR0_XORInst_3_2_U2 ( .A0_t (MCInst_MCR0_XORInst_3_2_n1), .B0_t (SubCellInst_SboxInst_2_YY[0]), .Z0_t (MCOutput[62]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) MCInst_MCR0_XORInst_3_2_U1 ( .A0_t (MCOutput[46]), .B0_t (SubCellInst_SboxInst_5_YY[0]), .Z0_t (MCInst_MCR0_XORInst_3_2_n1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) MCInst_MCR0_XORInst_3_3_U2 ( .A0_t (MCInst_MCR0_XORInst_3_3_n1), .B0_t (SubCellInst_SboxInst_2_YY[1]), .Z0_t (MCOutput[63]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) MCInst_MCR0_XORInst_3_3_U1 ( .A0_t (MCOutput[47]), .B0_t (SubCellInst_SboxInst_5_YY[1]), .Z0_t (MCInst_MCR0_XORInst_3_3_n1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MCInst_MCR2_XORInst_0_0_U1 ( .A0_t (ShiftRowsOutput[32]), .B0_t (ShiftRowsOutput[16]), .Z0_t (MCOutput[16]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MCInst_MCR2_XORInst_0_1_U1 ( .A0_t (ShiftRowsOutput[33]), .B0_t (ShiftRowsOutput[17]), .Z0_t (MCOutput[17]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) MCInst_MCR2_XORInst_0_2_U1 ( .A0_t (ShiftRowsOutput[34]), .B0_t (SubCellInst_SboxInst_6_YY[0]), .Z0_t (MCOutput[18]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) MCInst_MCR2_XORInst_0_3_U1 ( .A0_t (ShiftRowsOutput[35]), .B0_t (SubCellInst_SboxInst_6_YY[1]), .Z0_t (MCOutput[19]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MCInst_MCR2_XORInst_1_0_U1 ( .A0_t (ShiftRowsOutput[36]), .B0_t (ShiftRowsOutput[20]), .Z0_t (MCOutput[20]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) MCInst_MCR2_XORInst_1_1_U1 ( .A0_t (ShiftRowsOutput[37]), .B0_t (SubCellOutput[29]), .Z0_t (MCOutput[21]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) MCInst_MCR2_XORInst_1_2_U1 ( .A0_t (ShiftRowsOutput[38]), .B0_t (SubCellInst_SboxInst_7_YY[0]), .Z0_t (MCOutput[22]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) MCInst_MCR2_XORInst_1_3_U1 ( .A0_t (ShiftRowsOutput[39]), .B0_t (SubCellInst_SboxInst_7_YY[1]), .Z0_t (MCOutput[23]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MCInst_MCR2_XORInst_2_0_U1 ( .A0_t (ShiftRowsOutput[40]), .B0_t (ShiftRowsOutput[24]), .Z0_t (MCOutput[24]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MCInst_MCR2_XORInst_2_1_U1 ( .A0_t (ShiftRowsOutput[41]), .B0_t (ShiftRowsOutput[25]), .Z0_t (MCOutput[25]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) MCInst_MCR2_XORInst_2_2_U1 ( .A0_t (ShiftRowsOutput[42]), .B0_t (SubCellInst_SboxInst_4_YY[0]), .Z0_t (MCOutput[26]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) MCInst_MCR2_XORInst_2_3_U1 ( .A0_t (ShiftRowsOutput[43]), .B0_t (SubCellInst_SboxInst_4_YY[1]), .Z0_t (MCOutput[27]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MCInst_MCR2_XORInst_3_0_U1 ( .A0_t (ShiftRowsOutput[44]), .B0_t (ShiftRowsOutput[28]), .Z0_t (MCOutput[28]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MCInst_MCR2_XORInst_3_1_U1 ( .A0_t (ShiftRowsOutput[45]), .B0_t (ShiftRowsOutput[29]), .Z0_t (MCOutput[29]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) MCInst_MCR2_XORInst_3_2_U1 ( .A0_t (ShiftRowsOutput[46]), .B0_t (SubCellInst_SboxInst_5_YY[0]), .Z0_t (MCOutput[30]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) MCInst_MCR2_XORInst_3_3_U1 ( .A0_t (ShiftRowsOutput[47]), .B0_t (SubCellInst_SboxInst_5_YY[1]), .Z0_t (MCOutput[31]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MCInst_MCR3_XORInst_0_0_U1 ( .A0_t (MCOutput[32]), .B0_t (ShiftRowsOutput[16]), .Z0_t (MCOutput[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MCInst_MCR3_XORInst_0_1_U1 ( .A0_t (MCOutput[33]), .B0_t (ShiftRowsOutput[17]), .Z0_t (MCOutput[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) MCInst_MCR3_XORInst_0_2_U1 ( .A0_t (MCOutput[34]), .B0_t (SubCellInst_SboxInst_6_YY[0]), .Z0_t (MCOutput[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) MCInst_MCR3_XORInst_0_3_U1 ( .A0_t (MCOutput[35]), .B0_t (SubCellInst_SboxInst_6_YY[1]), .Z0_t (MCOutput[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MCInst_MCR3_XORInst_1_0_U1 ( .A0_t (MCOutput[36]), .B0_t (ShiftRowsOutput[20]), .Z0_t (MCOutput[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) MCInst_MCR3_XORInst_1_1_U1 ( .A0_t (MCOutput[37]), .B0_t (SubCellOutput[29]), .Z0_t (MCOutput[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) MCInst_MCR3_XORInst_1_2_U1 ( .A0_t (MCOutput[38]), .B0_t (SubCellInst_SboxInst_7_YY[0]), .Z0_t (MCOutput[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) MCInst_MCR3_XORInst_1_3_U1 ( .A0_t (MCOutput[39]), .B0_t (SubCellInst_SboxInst_7_YY[1]), .Z0_t (MCOutput[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MCInst_MCR3_XORInst_2_0_U1 ( .A0_t (MCOutput[40]), .B0_t (ShiftRowsOutput[24]), .Z0_t (MCOutput[8]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MCInst_MCR3_XORInst_2_1_U1 ( .A0_t (MCOutput[41]), .B0_t (ShiftRowsOutput[25]), .Z0_t (MCOutput[9]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) MCInst_MCR3_XORInst_2_2_U1 ( .A0_t (MCOutput[42]), .B0_t (SubCellInst_SboxInst_4_YY[0]), .Z0_t (MCOutput[10]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) MCInst_MCR3_XORInst_2_3_U1 ( .A0_t (MCOutput[43]), .B0_t (SubCellInst_SboxInst_4_YY[1]), .Z0_t (MCOutput[11]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MCInst_MCR3_XORInst_3_0_U1 ( .A0_t (MCOutput[44]), .B0_t (ShiftRowsOutput[28]), .Z0_t (MCOutput[12]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MCInst_MCR3_XORInst_3_1_U1 ( .A0_t (MCOutput[45]), .B0_t (ShiftRowsOutput[29]), .Z0_t (MCOutput[13]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) MCInst_MCR3_XORInst_3_2_U1 ( .A0_t (MCOutput[46]), .B0_t (SubCellInst_SboxInst_5_YY[0]), .Z0_t (MCOutput[14]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) MCInst_MCR3_XORInst_3_3_U1 ( .A0_t (MCOutput[47]), .B0_t (SubCellInst_SboxInst_5_YY[1]), .Z0_t (MCOutput[15]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_0_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[0]), .B0_t (Key[0]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_0_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_0_U1_AND1_U1 ( .A0_t (rst), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_0_U1_X), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_0_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_0_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_0_U1_Y), .B0_t (TweakeyGeneration_key_Feedback[0]), .Z0_t (TweakeyGeneration_key_Feedback[56]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_1_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[1]), .B0_t (Key[1]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_1_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_1_U1_AND1_U1 ( .A0_t (rst), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_1_U1_X), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_1_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_1_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_1_U1_Y), .B0_t (TweakeyGeneration_key_Feedback[1]), .Z0_t (TweakeyGeneration_key_Feedback[57]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_2_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[2]), .B0_t (Key[2]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_2_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_2_U1_AND1_U1 ( .A0_t (rst), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_2_U1_X), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_2_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_2_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_2_U1_Y), .B0_t (TweakeyGeneration_key_Feedback[2]), .Z0_t (TweakeyGeneration_key_Feedback[58]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_3_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[3]), .B0_t (Key[3]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_3_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_3_U1_AND1_U1 ( .A0_t (rst), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_3_U1_X), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_3_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_3_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_3_U1_Y), .B0_t (TweakeyGeneration_key_Feedback[3]), .Z0_t (TweakeyGeneration_key_Feedback[59]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_4_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[4]), .B0_t (Key[4]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_4_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_4_U1_AND1_U1 ( .A0_t (rst), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_4_U1_X), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_4_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_4_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_4_U1_Y), .B0_t (TweakeyGeneration_key_Feedback[4]), .Z0_t (TweakeyGeneration_key_Feedback[40]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_5_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[5]), .B0_t (Key[5]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_5_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_5_U1_AND1_U1 ( .A0_t (rst), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_5_U1_X), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_5_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_5_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_5_U1_Y), .B0_t (TweakeyGeneration_key_Feedback[5]), .Z0_t (TweakeyGeneration_key_Feedback[41]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_6_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[6]), .B0_t (Key[6]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_6_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_6_U1_AND1_U1 ( .A0_t (rst), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_6_U1_X), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_6_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_6_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_6_U1_Y), .B0_t (TweakeyGeneration_key_Feedback[6]), .Z0_t (TweakeyGeneration_key_Feedback[42]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_7_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[7]), .B0_t (Key[7]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_7_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_7_U1_AND1_U1 ( .A0_t (rst), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_7_U1_X), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_7_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_7_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_7_U1_Y), .B0_t (TweakeyGeneration_key_Feedback[7]), .Z0_t (TweakeyGeneration_key_Feedback[43]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_8_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[8]), .B0_t (Key[8]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_8_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_8_U1_AND1_U1 ( .A0_t (rst), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_8_U1_X), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_8_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_8_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_8_U1_Y), .B0_t (TweakeyGeneration_key_Feedback[8]), .Z0_t (TweakeyGeneration_key_Feedback[48]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_9_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[9]), .B0_t (Key[9]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_9_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_9_U1_AND1_U1 ( .A0_t (rst), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_9_U1_X), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_9_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_9_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_9_U1_Y), .B0_t (TweakeyGeneration_key_Feedback[9]), .Z0_t (TweakeyGeneration_key_Feedback[49]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_10_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[10]), .B0_t (Key[10]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_10_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_10_U1_AND1_U1 ( .A0_t (rst), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_10_U1_X), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_10_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_10_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_10_U1_Y), .B0_t (TweakeyGeneration_key_Feedback[10]), .Z0_t (TweakeyGeneration_key_Feedback[50]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_11_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[11]), .B0_t (Key[11]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_11_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_11_U1_AND1_U1 ( .A0_t (rst), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_11_U1_X), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_11_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_11_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_11_U1_Y), .B0_t (TweakeyGeneration_key_Feedback[11]), .Z0_t (TweakeyGeneration_key_Feedback[51]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_12_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[12]), .B0_t (Key[12]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_12_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_12_U1_AND1_U1 ( .A0_t (rst), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_12_U1_X), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_12_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_12_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_12_U1_Y), .B0_t (TweakeyGeneration_key_Feedback[12]), .Z0_t (TweakeyGeneration_key_Feedback[36]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_13_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[13]), .B0_t (Key[13]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_13_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_13_U1_AND1_U1 ( .A0_t (rst), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_13_U1_X), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_13_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_13_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_13_U1_Y), .B0_t (TweakeyGeneration_key_Feedback[13]), .Z0_t (TweakeyGeneration_key_Feedback[37]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_14_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[14]), .B0_t (Key[14]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_14_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_14_U1_AND1_U1 ( .A0_t (rst), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_14_U1_X), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_14_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_14_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_14_U1_Y), .B0_t (TweakeyGeneration_key_Feedback[14]), .Z0_t (TweakeyGeneration_key_Feedback[38]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_15_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[15]), .B0_t (Key[15]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_15_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_15_U1_AND1_U1 ( .A0_t (rst), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_15_U1_X), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_15_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_15_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_15_U1_Y), .B0_t (TweakeyGeneration_key_Feedback[15]), .Z0_t (TweakeyGeneration_key_Feedback[39]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_16_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[16]), .B0_t (Key[16]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_16_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_16_U1_AND1_U1 ( .A0_t (rst), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_16_U1_X), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_16_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_16_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_16_U1_Y), .B0_t (TweakeyGeneration_key_Feedback[16]), .Z0_t (TweakeyGeneration_key_Feedback[32]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_17_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[17]), .B0_t (Key[17]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_17_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_17_U1_AND1_U1 ( .A0_t (rst), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_17_U1_X), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_17_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_17_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_17_U1_Y), .B0_t (TweakeyGeneration_key_Feedback[17]), .Z0_t (TweakeyGeneration_key_Feedback[33]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_18_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[18]), .B0_t (Key[18]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_18_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_18_U1_AND1_U1 ( .A0_t (rst), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_18_U1_X), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_18_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_18_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_18_U1_Y), .B0_t (TweakeyGeneration_key_Feedback[18]), .Z0_t (TweakeyGeneration_key_Feedback[34]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_19_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[19]), .B0_t (Key[19]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_19_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_19_U1_AND1_U1 ( .A0_t (rst), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_19_U1_X), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_19_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_19_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_19_U1_Y), .B0_t (TweakeyGeneration_key_Feedback[19]), .Z0_t (TweakeyGeneration_key_Feedback[35]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_20_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[20]), .B0_t (Key[20]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_20_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_20_U1_AND1_U1 ( .A0_t (rst), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_20_U1_X), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_20_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_20_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_20_U1_Y), .B0_t (TweakeyGeneration_key_Feedback[20]), .Z0_t (TweakeyGeneration_key_Feedback[44]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_21_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[21]), .B0_t (Key[21]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_21_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_21_U1_AND1_U1 ( .A0_t (rst), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_21_U1_X), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_21_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_21_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_21_U1_Y), .B0_t (TweakeyGeneration_key_Feedback[21]), .Z0_t (TweakeyGeneration_key_Feedback[45]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_22_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[22]), .B0_t (Key[22]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_22_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_22_U1_AND1_U1 ( .A0_t (rst), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_22_U1_X), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_22_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_22_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_22_U1_Y), .B0_t (TweakeyGeneration_key_Feedback[22]), .Z0_t (TweakeyGeneration_key_Feedback[46]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_23_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[23]), .B0_t (Key[23]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_23_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_23_U1_AND1_U1 ( .A0_t (rst), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_23_U1_X), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_23_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_23_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_23_U1_Y), .B0_t (TweakeyGeneration_key_Feedback[23]), .Z0_t (TweakeyGeneration_key_Feedback[47]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_24_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[24]), .B0_t (Key[24]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_24_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_24_U1_AND1_U1 ( .A0_t (rst), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_24_U1_X), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_24_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_24_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_24_U1_Y), .B0_t (TweakeyGeneration_key_Feedback[24]), .Z0_t (TweakeyGeneration_key_Feedback[60]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_25_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[25]), .B0_t (Key[25]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_25_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_25_U1_AND1_U1 ( .A0_t (rst), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_25_U1_X), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_25_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_25_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_25_U1_Y), .B0_t (TweakeyGeneration_key_Feedback[25]), .Z0_t (TweakeyGeneration_key_Feedback[61]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_26_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[26]), .B0_t (Key[26]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_26_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_26_U1_AND1_U1 ( .A0_t (rst), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_26_U1_X), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_26_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_26_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_26_U1_Y), .B0_t (TweakeyGeneration_key_Feedback[26]), .Z0_t (TweakeyGeneration_key_Feedback[62]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_27_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[27]), .B0_t (Key[27]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_27_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_27_U1_AND1_U1 ( .A0_t (rst), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_27_U1_X), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_27_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_27_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_27_U1_Y), .B0_t (TweakeyGeneration_key_Feedback[27]), .Z0_t (TweakeyGeneration_key_Feedback[63]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_28_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[28]), .B0_t (Key[28]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_28_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_28_U1_AND1_U1 ( .A0_t (rst), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_28_U1_X), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_28_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_28_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_28_U1_Y), .B0_t (TweakeyGeneration_key_Feedback[28]), .Z0_t (TweakeyGeneration_key_Feedback[52]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_29_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[29]), .B0_t (Key[29]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_29_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_29_U1_AND1_U1 ( .A0_t (rst), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_29_U1_X), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_29_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_29_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_29_U1_Y), .B0_t (TweakeyGeneration_key_Feedback[29]), .Z0_t (TweakeyGeneration_key_Feedback[53]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_30_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[30]), .B0_t (Key[30]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_30_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_30_U1_AND1_U1 ( .A0_t (rst), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_30_U1_X), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_30_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_30_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_30_U1_Y), .B0_t (TweakeyGeneration_key_Feedback[30]), .Z0_t (TweakeyGeneration_key_Feedback[54]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_31_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[31]), .B0_t (Key[31]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_31_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_31_U1_AND1_U1 ( .A0_t (rst), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_31_U1_X), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_31_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_31_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_31_U1_Y), .B0_t (TweakeyGeneration_key_Feedback[31]), .Z0_t (TweakeyGeneration_key_Feedback[55]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_32_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[32]), .B0_t (Key[32]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_32_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_32_U1_AND1_U1 ( .A0_t (rst), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_32_U1_X), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_32_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_32_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_32_U1_Y), .B0_t (TweakeyGeneration_key_Feedback[32]), .Z0_t (TweakeyGeneration_key_Feedback[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_33_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[33]), .B0_t (Key[33]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_33_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_33_U1_AND1_U1 ( .A0_t (rst), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_33_U1_X), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_33_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_33_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_33_U1_Y), .B0_t (TweakeyGeneration_key_Feedback[33]), .Z0_t (TweakeyGeneration_key_Feedback[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_34_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[34]), .B0_t (Key[34]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_34_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_34_U1_AND1_U1 ( .A0_t (rst), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_34_U1_X), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_34_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_34_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_34_U1_Y), .B0_t (TweakeyGeneration_key_Feedback[34]), .Z0_t (TweakeyGeneration_key_Feedback[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_35_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[35]), .B0_t (Key[35]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_35_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_35_U1_AND1_U1 ( .A0_t (rst), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_35_U1_X), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_35_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_35_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_35_U1_Y), .B0_t (TweakeyGeneration_key_Feedback[35]), .Z0_t (TweakeyGeneration_key_Feedback[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_36_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[36]), .B0_t (Key[36]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_36_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_36_U1_AND1_U1 ( .A0_t (rst), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_36_U1_X), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_36_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_36_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_36_U1_Y), .B0_t (TweakeyGeneration_key_Feedback[36]), .Z0_t (TweakeyGeneration_key_Feedback[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_37_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[37]), .B0_t (Key[37]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_37_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_37_U1_AND1_U1 ( .A0_t (rst), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_37_U1_X), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_37_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_37_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_37_U1_Y), .B0_t (TweakeyGeneration_key_Feedback[37]), .Z0_t (TweakeyGeneration_key_Feedback[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_38_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[38]), .B0_t (Key[38]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_38_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_38_U1_AND1_U1 ( .A0_t (rst), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_38_U1_X), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_38_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_38_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_38_U1_Y), .B0_t (TweakeyGeneration_key_Feedback[38]), .Z0_t (TweakeyGeneration_key_Feedback[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_39_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[39]), .B0_t (Key[39]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_39_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_39_U1_AND1_U1 ( .A0_t (rst), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_39_U1_X), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_39_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_39_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_39_U1_Y), .B0_t (TweakeyGeneration_key_Feedback[39]), .Z0_t (TweakeyGeneration_key_Feedback[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_40_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[40]), .B0_t (Key[40]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_40_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_40_U1_AND1_U1 ( .A0_t (rst), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_40_U1_X), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_40_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_40_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_40_U1_Y), .B0_t (TweakeyGeneration_key_Feedback[40]), .Z0_t (TweakeyGeneration_key_Feedback[8]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_41_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[41]), .B0_t (Key[41]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_41_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_41_U1_AND1_U1 ( .A0_t (rst), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_41_U1_X), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_41_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_41_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_41_U1_Y), .B0_t (TweakeyGeneration_key_Feedback[41]), .Z0_t (TweakeyGeneration_key_Feedback[9]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_42_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[42]), .B0_t (Key[42]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_42_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_42_U1_AND1_U1 ( .A0_t (rst), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_42_U1_X), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_42_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_42_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_42_U1_Y), .B0_t (TweakeyGeneration_key_Feedback[42]), .Z0_t (TweakeyGeneration_key_Feedback[10]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_43_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[43]), .B0_t (Key[43]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_43_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_43_U1_AND1_U1 ( .A0_t (rst), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_43_U1_X), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_43_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_43_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_43_U1_Y), .B0_t (TweakeyGeneration_key_Feedback[43]), .Z0_t (TweakeyGeneration_key_Feedback[11]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_44_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[44]), .B0_t (Key[44]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_44_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_44_U1_AND1_U1 ( .A0_t (rst), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_44_U1_X), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_44_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_44_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_44_U1_Y), .B0_t (TweakeyGeneration_key_Feedback[44]), .Z0_t (TweakeyGeneration_key_Feedback[12]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_45_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[45]), .B0_t (Key[45]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_45_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_45_U1_AND1_U1 ( .A0_t (rst), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_45_U1_X), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_45_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_45_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_45_U1_Y), .B0_t (TweakeyGeneration_key_Feedback[45]), .Z0_t (TweakeyGeneration_key_Feedback[13]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_46_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[46]), .B0_t (Key[46]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_46_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_46_U1_AND1_U1 ( .A0_t (rst), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_46_U1_X), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_46_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_46_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_46_U1_Y), .B0_t (TweakeyGeneration_key_Feedback[46]), .Z0_t (TweakeyGeneration_key_Feedback[14]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_47_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[47]), .B0_t (Key[47]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_47_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_47_U1_AND1_U1 ( .A0_t (rst), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_47_U1_X), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_47_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_47_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_47_U1_Y), .B0_t (TweakeyGeneration_key_Feedback[47]), .Z0_t (TweakeyGeneration_key_Feedback[15]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_48_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[48]), .B0_t (Key[48]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_48_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_48_U1_AND1_U1 ( .A0_t (rst), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_48_U1_X), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_48_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_48_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_48_U1_Y), .B0_t (TweakeyGeneration_key_Feedback[48]), .Z0_t (TweakeyGeneration_key_Feedback[16]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_49_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[49]), .B0_t (Key[49]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_49_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_49_U1_AND1_U1 ( .A0_t (rst), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_49_U1_X), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_49_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_49_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_49_U1_Y), .B0_t (TweakeyGeneration_key_Feedback[49]), .Z0_t (TweakeyGeneration_key_Feedback[17]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_50_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[50]), .B0_t (Key[50]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_50_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_50_U1_AND1_U1 ( .A0_t (rst), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_50_U1_X), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_50_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_50_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_50_U1_Y), .B0_t (TweakeyGeneration_key_Feedback[50]), .Z0_t (TweakeyGeneration_key_Feedback[18]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_51_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[51]), .B0_t (Key[51]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_51_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_51_U1_AND1_U1 ( .A0_t (rst), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_51_U1_X), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_51_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_51_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_51_U1_Y), .B0_t (TweakeyGeneration_key_Feedback[51]), .Z0_t (TweakeyGeneration_key_Feedback[19]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_52_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[52]), .B0_t (Key[52]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_52_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_52_U1_AND1_U1 ( .A0_t (rst), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_52_U1_X), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_52_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_52_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_52_U1_Y), .B0_t (TweakeyGeneration_key_Feedback[52]), .Z0_t (TweakeyGeneration_key_Feedback[20]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_53_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[53]), .B0_t (Key[53]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_53_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_53_U1_AND1_U1 ( .A0_t (rst), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_53_U1_X), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_53_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_53_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_53_U1_Y), .B0_t (TweakeyGeneration_key_Feedback[53]), .Z0_t (TweakeyGeneration_key_Feedback[21]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_54_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[54]), .B0_t (Key[54]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_54_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_54_U1_AND1_U1 ( .A0_t (rst), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_54_U1_X), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_54_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_54_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_54_U1_Y), .B0_t (TweakeyGeneration_key_Feedback[54]), .Z0_t (TweakeyGeneration_key_Feedback[22]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_55_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[55]), .B0_t (Key[55]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_55_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_55_U1_AND1_U1 ( .A0_t (rst), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_55_U1_X), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_55_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_55_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_55_U1_Y), .B0_t (TweakeyGeneration_key_Feedback[55]), .Z0_t (TweakeyGeneration_key_Feedback[23]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_56_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[56]), .B0_t (Key[56]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_56_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_56_U1_AND1_U1 ( .A0_t (rst), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_56_U1_X), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_56_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_56_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_56_U1_Y), .B0_t (TweakeyGeneration_key_Feedback[56]), .Z0_t (TweakeyGeneration_key_Feedback[24]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_57_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[57]), .B0_t (Key[57]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_57_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_57_U1_AND1_U1 ( .A0_t (rst), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_57_U1_X), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_57_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_57_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_57_U1_Y), .B0_t (TweakeyGeneration_key_Feedback[57]), .Z0_t (TweakeyGeneration_key_Feedback[25]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_58_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[58]), .B0_t (Key[58]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_58_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_58_U1_AND1_U1 ( .A0_t (rst), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_58_U1_X), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_58_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_58_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_58_U1_Y), .B0_t (TweakeyGeneration_key_Feedback[58]), .Z0_t (TweakeyGeneration_key_Feedback[26]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_59_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[59]), .B0_t (Key[59]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_59_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_59_U1_AND1_U1 ( .A0_t (rst), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_59_U1_X), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_59_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_59_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_59_U1_Y), .B0_t (TweakeyGeneration_key_Feedback[59]), .Z0_t (TweakeyGeneration_key_Feedback[27]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_60_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[60]), .B0_t (Key[60]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_60_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_60_U1_AND1_U1 ( .A0_t (rst), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_60_U1_X), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_60_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_60_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_60_U1_Y), .B0_t (TweakeyGeneration_key_Feedback[60]), .Z0_t (TweakeyGeneration_key_Feedback[28]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_61_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[61]), .B0_t (Key[61]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_61_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_61_U1_AND1_U1 ( .A0_t (rst), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_61_U1_X), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_61_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_61_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_61_U1_Y), .B0_t (TweakeyGeneration_key_Feedback[61]), .Z0_t (TweakeyGeneration_key_Feedback[29]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_62_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[62]), .B0_t (Key[62]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_62_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_62_U1_AND1_U1 ( .A0_t (rst), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_62_U1_X), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_62_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_62_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_62_U1_Y), .B0_t (TweakeyGeneration_key_Feedback[62]), .Z0_t (TweakeyGeneration_key_Feedback[30]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_63_U1_XOR1_U1 ( .A0_t (TweakeyGeneration_key_Feedback[63]), .B0_t (Key[63]), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_63_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) TweakeyGeneration_KEYMUX_MUXInst_63_U1_AND1_U1 ( .A0_t (rst), .B0_t (TweakeyGeneration_KEYMUX_MUXInst_63_U1_X), .Z0_t (TweakeyGeneration_KEYMUX_MUXInst_63_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) TweakeyGeneration_KEYMUX_MUXInst_63_U1_XOR2_U1 ( .A0_t (TweakeyGeneration_KEYMUX_MUXInst_63_U1_Y), .B0_t (TweakeyGeneration_key_Feedback[63]), .Z0_t (TweakeyGeneration_key_Feedback[31]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b1), .NL(1'b1)) FSMMUX_MUXInst_0_U1 ( .A0_t (FSMUpdate[0]), .B0_t (rst), .Z0_t (FSMUpdate[1]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) FSMMUX_MUXInst_1_U2 ( .A0_t (rst), .B0_t (FSMUpdate[1]), .Z0_t (FSM[1]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) FSMMUX_MUXInst_2_U2 ( .A0_t (rst), .B0_t (FSMUpdate[2]), .Z0_t (FSMUpdate[3]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) FSMMUX_MUXInst_3_U2 ( .A0_t (rst), .B0_t (FSMUpdate[3]), .Z0_t (FSMUpdate[4]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) FSMMUX_MUXInst_4_U2 ( .A0_t (rst), .B0_t (FSMUpdate[4]), .Z0_t (FSM[4]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) FSMMUX_MUXInst_5_U2 ( .A0_t (rst), .B0_t (FSMUpdate[5]), .Z0_t (FSM[5]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) FSMUpdateInst_StateUpdateInst_0_U4 ( .A0_t (FSM[5]), .B0_t (FSMUpdateInst_StateUpdateInst_0_n3), .Z0_t (FSMUpdateInst_StateUpdateInst_0_n4) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) FSMUpdateInst_StateUpdateInst_0_U3 ( .A0_t (FSMUpdateInst_StateUpdateInst_0_n2), .B0_t (FSMUpdateInst_StateUpdateInst_0_n1), .Z0_t (FSMUpdateInst_StateUpdateInst_0_n3) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) FSMUpdateInst_StateUpdateInst_0_U2 ( .A0_t (FSMUpdate[4]), .B0_t (FSMUpdate[3]), .Z0_t (FSMUpdateInst_StateUpdateInst_0_n1) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) FSMUpdateInst_StateUpdateInst_0_U1 ( .A0_t (FSMUpdate[1]), .B0_t (FSM[1]), .Z0_t (FSMUpdateInst_StateUpdateInst_0_n2) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) FSMUpdateInst_StateUpdateInst_0_U7_XOR1_U1 ( .A0_t (FSMUpdateInst_StateUpdateInst_0_n4), .B0_t (FSM[5]), .Z0_t (FSMUpdateInst_StateUpdateInst_0_U7_X) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) FSMUpdateInst_StateUpdateInst_0_U7_AND1_U1 ( .A0_t (FSM[4]), .B0_t (FSMUpdateInst_StateUpdateInst_0_U7_X), .Z0_t (FSMUpdateInst_StateUpdateInst_0_U7_Y) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) FSMUpdateInst_StateUpdateInst_0_U7_XOR2_U1 ( .A0_t (FSMUpdateInst_StateUpdateInst_0_U7_Y), .B0_t (FSMUpdateInst_StateUpdateInst_0_n4), .Z0_t (FSMUpdate[0]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) FSMUpdateInst_StateUpdateInst_2_U5 ( .A0_t (FSMUpdateInst_StateUpdateInst_2_n4), .B0_t (FSM[1]), .Z0_t (FSMUpdate[2]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) FSMUpdateInst_StateUpdateInst_2_U4 ( .A0_t (FSMUpdateInst_StateUpdateInst_2_n3), .B0_t (FSM[5]), .Z0_t (FSMUpdateInst_StateUpdateInst_2_n4) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) FSMUpdateInst_StateUpdateInst_2_U3 ( .A0_t (FSM[4]), .B0_t (FSMUpdateInst_StateUpdateInst_2_n2), .Z0_t (FSMUpdateInst_StateUpdateInst_2_n3) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) FSMUpdateInst_StateUpdateInst_2_U2 ( .A0_t (FSMUpdate[1]), .B0_t (FSMUpdateInst_StateUpdateInst_2_n1), .Z0_t (FSMUpdateInst_StateUpdateInst_2_n2) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) FSMUpdateInst_StateUpdateInst_2_U1 ( .A0_t (FSMUpdate[4]), .B0_t (FSMUpdate[3]), .Z0_t (FSMUpdateInst_StateUpdateInst_2_n1) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) FSMUpdateInst_StateUpdateInst_5_U5 ( .A0_t (FSM[4]), .B0_t (FSMUpdateInst_StateUpdateInst_5_n4), .Z0_t (FSMUpdate[5]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) FSMUpdateInst_StateUpdateInst_5_U4 ( .A0_t (FSMUpdate[4]), .B0_t (FSMUpdateInst_StateUpdateInst_5_n3), .Z0_t (FSMUpdateInst_StateUpdateInst_5_n4) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) FSMUpdateInst_StateUpdateInst_5_U3 ( .A0_t (FSM[5]), .B0_t (FSMUpdateInst_StateUpdateInst_5_n2), .Z0_t (FSMUpdateInst_StateUpdateInst_5_n3) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) FSMUpdateInst_StateUpdateInst_5_U2 ( .A0_t (FSMUpdate[3]), .B0_t (FSMUpdateInst_StateUpdateInst_5_n1), .Z0_t (FSMUpdateInst_StateUpdateInst_5_n2) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) FSMUpdateInst_StateUpdateInst_5_U1 ( .A0_t (FSMUpdate[1]), .B0_t (FSM[1]), .Z0_t (FSMUpdateInst_StateUpdateInst_5_n1) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) FSMSignalsInst_doneInst_U6 ( .A0_t (FSMSignalsInst_doneInst_n5), .B0_t (FSMSignalsInst_doneInst_n4), .Z0_t (done) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) FSMSignalsInst_doneInst_U5 ( .A0_t (FSM[4]), .B0_t (FSM[5]), .Z0_t (FSMSignalsInst_doneInst_n4) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) FSMSignalsInst_doneInst_U4 ( .A0_t (FSMSignalsInst_doneInst_n3), .B0_t (FSMSignalsInst_doneInst_n2), .Z0_t (FSMSignalsInst_doneInst_n5) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) FSMSignalsInst_doneInst_U3 ( .A0_t (FSMUpdate[4]), .B0_t (FSMUpdate[1]), .Z0_t (FSMSignalsInst_doneInst_n2) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) FSMSignalsInst_doneInst_U1 ( .A0_t (FSMUpdate[3]), .B0_t (FSM[1]), .Z0_t (FSMSignalsInst_doneInst_n3) ) ;

    /* register cells */
endmodule
