
module AES ( clk, start, port_in, port_out, done );
  input [7:0] port_in;
  output [7:0] port_out;
  input clk, start;
  output done;
  wire   start_done, n286, n287, notdone, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         RoundReg_n10, RoundReg_n9, RoundReg_n8, RoundReg_n7, RoundReg_n6,
         RoundReg_Inst_ff_SDE_0_next_state, RoundReg_Inst_ff_SDE_0_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_0_MUX_inst_X,
         RoundReg_Inst_ff_SDE_0_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_1_next_state, RoundReg_Inst_ff_SDE_1_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_1_MUX_inst_X,
         RoundReg_Inst_ff_SDE_1_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_2_next_state, RoundReg_Inst_ff_SDE_2_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_2_MUX_inst_X,
         RoundReg_Inst_ff_SDE_2_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_3_next_state, RoundReg_Inst_ff_SDE_3_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_3_MUX_inst_X,
         RoundReg_Inst_ff_SDE_3_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_4_next_state, RoundReg_Inst_ff_SDE_4_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_4_MUX_inst_X,
         RoundReg_Inst_ff_SDE_4_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_5_next_state, RoundReg_Inst_ff_SDE_5_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_5_MUX_inst_X,
         RoundReg_Inst_ff_SDE_5_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_6_next_state, RoundReg_Inst_ff_SDE_6_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_6_MUX_inst_X,
         RoundReg_Inst_ff_SDE_6_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_7_next_state, RoundReg_Inst_ff_SDE_7_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_7_MUX_inst_X,
         RoundReg_Inst_ff_SDE_7_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_8_next_state, RoundReg_Inst_ff_SDE_8_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_8_MUX_inst_X,
         RoundReg_Inst_ff_SDE_8_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_9_next_state, RoundReg_Inst_ff_SDE_9_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_9_MUX_inst_X,
         RoundReg_Inst_ff_SDE_9_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_10_next_state,
         RoundReg_Inst_ff_SDE_10_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_10_MUX_inst_X,
         RoundReg_Inst_ff_SDE_10_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_11_next_state,
         RoundReg_Inst_ff_SDE_11_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_11_MUX_inst_X,
         RoundReg_Inst_ff_SDE_11_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_12_next_state,
         RoundReg_Inst_ff_SDE_12_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_12_MUX_inst_X,
         RoundReg_Inst_ff_SDE_12_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_13_next_state,
         RoundReg_Inst_ff_SDE_13_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_13_MUX_inst_X,
         RoundReg_Inst_ff_SDE_13_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_14_next_state,
         RoundReg_Inst_ff_SDE_14_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_14_MUX_inst_X,
         RoundReg_Inst_ff_SDE_14_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_15_next_state,
         RoundReg_Inst_ff_SDE_15_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_15_MUX_inst_X,
         RoundReg_Inst_ff_SDE_15_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_16_next_state,
         RoundReg_Inst_ff_SDE_16_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_16_MUX_inst_X,
         RoundReg_Inst_ff_SDE_16_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_17_next_state,
         RoundReg_Inst_ff_SDE_17_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_17_MUX_inst_X,
         RoundReg_Inst_ff_SDE_17_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_18_next_state,
         RoundReg_Inst_ff_SDE_18_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_18_MUX_inst_X,
         RoundReg_Inst_ff_SDE_18_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_19_next_state,
         RoundReg_Inst_ff_SDE_19_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_19_MUX_inst_X,
         RoundReg_Inst_ff_SDE_19_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_20_next_state,
         RoundReg_Inst_ff_SDE_20_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_20_MUX_inst_X,
         RoundReg_Inst_ff_SDE_20_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_21_next_state,
         RoundReg_Inst_ff_SDE_21_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_21_MUX_inst_X,
         RoundReg_Inst_ff_SDE_21_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_22_next_state,
         RoundReg_Inst_ff_SDE_22_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_22_MUX_inst_X,
         RoundReg_Inst_ff_SDE_22_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_23_next_state,
         RoundReg_Inst_ff_SDE_23_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_23_MUX_inst_X,
         RoundReg_Inst_ff_SDE_23_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_24_next_state,
         RoundReg_Inst_ff_SDE_24_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_24_MUX_inst_X,
         RoundReg_Inst_ff_SDE_24_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_25_next_state,
         RoundReg_Inst_ff_SDE_25_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_25_MUX_inst_X,
         RoundReg_Inst_ff_SDE_25_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_26_next_state,
         RoundReg_Inst_ff_SDE_26_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_26_MUX_inst_X,
         RoundReg_Inst_ff_SDE_26_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_27_next_state,
         RoundReg_Inst_ff_SDE_27_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_27_MUX_inst_X,
         RoundReg_Inst_ff_SDE_27_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_28_next_state,
         RoundReg_Inst_ff_SDE_28_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_28_MUX_inst_X,
         RoundReg_Inst_ff_SDE_28_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_29_next_state,
         RoundReg_Inst_ff_SDE_29_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_29_MUX_inst_X,
         RoundReg_Inst_ff_SDE_29_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_30_next_state,
         RoundReg_Inst_ff_SDE_30_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_30_MUX_inst_X,
         RoundReg_Inst_ff_SDE_30_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_31_next_state,
         RoundReg_Inst_ff_SDE_31_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_31_MUX_inst_X,
         RoundReg_Inst_ff_SDE_31_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_32_next_state,
         RoundReg_Inst_ff_SDE_32_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_32_MUX_inst_X,
         RoundReg_Inst_ff_SDE_32_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_33_next_state,
         RoundReg_Inst_ff_SDE_33_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_33_MUX_inst_X,
         RoundReg_Inst_ff_SDE_33_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_34_next_state,
         RoundReg_Inst_ff_SDE_34_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_34_MUX_inst_X,
         RoundReg_Inst_ff_SDE_34_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_35_next_state,
         RoundReg_Inst_ff_SDE_35_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_35_MUX_inst_X,
         RoundReg_Inst_ff_SDE_35_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_36_next_state,
         RoundReg_Inst_ff_SDE_36_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_36_MUX_inst_X,
         RoundReg_Inst_ff_SDE_36_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_37_next_state,
         RoundReg_Inst_ff_SDE_37_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_37_MUX_inst_X,
         RoundReg_Inst_ff_SDE_37_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_38_next_state,
         RoundReg_Inst_ff_SDE_38_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_38_MUX_inst_X,
         RoundReg_Inst_ff_SDE_38_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_39_next_state,
         RoundReg_Inst_ff_SDE_39_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_39_MUX_inst_X,
         RoundReg_Inst_ff_SDE_39_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_40_next_state,
         RoundReg_Inst_ff_SDE_40_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_40_MUX_inst_X,
         RoundReg_Inst_ff_SDE_40_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_41_next_state,
         RoundReg_Inst_ff_SDE_41_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_41_MUX_inst_X,
         RoundReg_Inst_ff_SDE_41_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_42_next_state,
         RoundReg_Inst_ff_SDE_42_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_42_MUX_inst_X,
         RoundReg_Inst_ff_SDE_42_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_43_next_state,
         RoundReg_Inst_ff_SDE_43_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_43_MUX_inst_X,
         RoundReg_Inst_ff_SDE_43_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_44_next_state,
         RoundReg_Inst_ff_SDE_44_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_44_MUX_inst_X,
         RoundReg_Inst_ff_SDE_44_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_45_next_state,
         RoundReg_Inst_ff_SDE_45_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_45_MUX_inst_X,
         RoundReg_Inst_ff_SDE_45_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_46_next_state,
         RoundReg_Inst_ff_SDE_46_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_46_MUX_inst_X,
         RoundReg_Inst_ff_SDE_46_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_47_next_state,
         RoundReg_Inst_ff_SDE_47_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_47_MUX_inst_X,
         RoundReg_Inst_ff_SDE_47_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_48_next_state,
         RoundReg_Inst_ff_SDE_48_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_48_MUX_inst_X,
         RoundReg_Inst_ff_SDE_48_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_49_next_state,
         RoundReg_Inst_ff_SDE_49_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_49_MUX_inst_X,
         RoundReg_Inst_ff_SDE_49_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_50_next_state,
         RoundReg_Inst_ff_SDE_50_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_50_MUX_inst_X,
         RoundReg_Inst_ff_SDE_50_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_51_next_state,
         RoundReg_Inst_ff_SDE_51_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_51_MUX_inst_X,
         RoundReg_Inst_ff_SDE_51_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_52_next_state,
         RoundReg_Inst_ff_SDE_52_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_52_MUX_inst_X,
         RoundReg_Inst_ff_SDE_52_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_53_next_state,
         RoundReg_Inst_ff_SDE_53_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_53_MUX_inst_X,
         RoundReg_Inst_ff_SDE_53_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_54_next_state,
         RoundReg_Inst_ff_SDE_54_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_54_MUX_inst_X,
         RoundReg_Inst_ff_SDE_54_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_55_next_state,
         RoundReg_Inst_ff_SDE_55_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_55_MUX_inst_X,
         RoundReg_Inst_ff_SDE_55_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_56_next_state,
         RoundReg_Inst_ff_SDE_56_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_56_MUX_inst_X,
         RoundReg_Inst_ff_SDE_56_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_57_next_state,
         RoundReg_Inst_ff_SDE_57_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_57_MUX_inst_X,
         RoundReg_Inst_ff_SDE_57_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_58_next_state,
         RoundReg_Inst_ff_SDE_58_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_58_MUX_inst_X,
         RoundReg_Inst_ff_SDE_58_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_59_next_state,
         RoundReg_Inst_ff_SDE_59_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_59_MUX_inst_X,
         RoundReg_Inst_ff_SDE_59_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_60_next_state,
         RoundReg_Inst_ff_SDE_60_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_60_MUX_inst_X,
         RoundReg_Inst_ff_SDE_60_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_61_next_state,
         RoundReg_Inst_ff_SDE_61_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_61_MUX_inst_X,
         RoundReg_Inst_ff_SDE_61_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_62_next_state,
         RoundReg_Inst_ff_SDE_62_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_62_MUX_inst_X,
         RoundReg_Inst_ff_SDE_62_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_63_next_state,
         RoundReg_Inst_ff_SDE_63_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_63_MUX_inst_X,
         RoundReg_Inst_ff_SDE_63_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_64_next_state,
         RoundReg_Inst_ff_SDE_64_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_64_MUX_inst_X,
         RoundReg_Inst_ff_SDE_64_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_65_next_state,
         RoundReg_Inst_ff_SDE_65_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_65_MUX_inst_X,
         RoundReg_Inst_ff_SDE_65_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_66_next_state,
         RoundReg_Inst_ff_SDE_66_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_66_MUX_inst_X,
         RoundReg_Inst_ff_SDE_66_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_67_next_state,
         RoundReg_Inst_ff_SDE_67_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_67_MUX_inst_X,
         RoundReg_Inst_ff_SDE_67_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_68_next_state,
         RoundReg_Inst_ff_SDE_68_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_68_MUX_inst_X,
         RoundReg_Inst_ff_SDE_68_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_69_next_state,
         RoundReg_Inst_ff_SDE_69_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_69_MUX_inst_X,
         RoundReg_Inst_ff_SDE_69_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_70_next_state,
         RoundReg_Inst_ff_SDE_70_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_70_MUX_inst_X,
         RoundReg_Inst_ff_SDE_70_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_71_next_state,
         RoundReg_Inst_ff_SDE_71_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_71_MUX_inst_X,
         RoundReg_Inst_ff_SDE_71_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_72_next_state,
         RoundReg_Inst_ff_SDE_72_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_72_MUX_inst_X,
         RoundReg_Inst_ff_SDE_72_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_73_next_state,
         RoundReg_Inst_ff_SDE_73_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_73_MUX_inst_X,
         RoundReg_Inst_ff_SDE_73_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_74_next_state,
         RoundReg_Inst_ff_SDE_74_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_74_MUX_inst_X,
         RoundReg_Inst_ff_SDE_74_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_75_next_state,
         RoundReg_Inst_ff_SDE_75_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_75_MUX_inst_X,
         RoundReg_Inst_ff_SDE_75_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_76_next_state,
         RoundReg_Inst_ff_SDE_76_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_76_MUX_inst_X,
         RoundReg_Inst_ff_SDE_76_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_77_next_state,
         RoundReg_Inst_ff_SDE_77_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_77_MUX_inst_X,
         RoundReg_Inst_ff_SDE_77_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_78_next_state,
         RoundReg_Inst_ff_SDE_78_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_78_MUX_inst_X,
         RoundReg_Inst_ff_SDE_78_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_79_next_state,
         RoundReg_Inst_ff_SDE_79_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_79_MUX_inst_X,
         RoundReg_Inst_ff_SDE_79_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_80_next_state,
         RoundReg_Inst_ff_SDE_80_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_80_MUX_inst_X,
         RoundReg_Inst_ff_SDE_80_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_81_next_state,
         RoundReg_Inst_ff_SDE_81_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_81_MUX_inst_X,
         RoundReg_Inst_ff_SDE_81_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_82_next_state,
         RoundReg_Inst_ff_SDE_82_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_82_MUX_inst_X,
         RoundReg_Inst_ff_SDE_82_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_83_next_state,
         RoundReg_Inst_ff_SDE_83_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_83_MUX_inst_X,
         RoundReg_Inst_ff_SDE_83_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_84_next_state,
         RoundReg_Inst_ff_SDE_84_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_84_MUX_inst_X,
         RoundReg_Inst_ff_SDE_84_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_85_next_state,
         RoundReg_Inst_ff_SDE_85_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_85_MUX_inst_X,
         RoundReg_Inst_ff_SDE_85_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_86_next_state,
         RoundReg_Inst_ff_SDE_86_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_86_MUX_inst_X,
         RoundReg_Inst_ff_SDE_86_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_87_next_state,
         RoundReg_Inst_ff_SDE_87_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_87_MUX_inst_X,
         RoundReg_Inst_ff_SDE_87_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_88_next_state,
         RoundReg_Inst_ff_SDE_88_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_88_MUX_inst_X,
         RoundReg_Inst_ff_SDE_88_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_89_next_state,
         RoundReg_Inst_ff_SDE_89_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_89_MUX_inst_X,
         RoundReg_Inst_ff_SDE_89_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_90_next_state,
         RoundReg_Inst_ff_SDE_90_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_90_MUX_inst_X,
         RoundReg_Inst_ff_SDE_90_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_91_next_state,
         RoundReg_Inst_ff_SDE_91_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_91_MUX_inst_X,
         RoundReg_Inst_ff_SDE_91_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_92_next_state,
         RoundReg_Inst_ff_SDE_92_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_92_MUX_inst_X,
         RoundReg_Inst_ff_SDE_92_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_93_next_state,
         RoundReg_Inst_ff_SDE_93_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_93_MUX_inst_X,
         RoundReg_Inst_ff_SDE_93_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_94_next_state,
         RoundReg_Inst_ff_SDE_94_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_94_MUX_inst_X,
         RoundReg_Inst_ff_SDE_94_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_95_next_state,
         RoundReg_Inst_ff_SDE_95_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_95_MUX_inst_X,
         RoundReg_Inst_ff_SDE_95_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_96_next_state,
         RoundReg_Inst_ff_SDE_96_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_96_MUX_inst_X,
         RoundReg_Inst_ff_SDE_96_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_97_next_state,
         RoundReg_Inst_ff_SDE_97_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_97_MUX_inst_X,
         RoundReg_Inst_ff_SDE_97_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_98_next_state,
         RoundReg_Inst_ff_SDE_98_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_98_MUX_inst_X,
         RoundReg_Inst_ff_SDE_98_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_99_next_state,
         RoundReg_Inst_ff_SDE_99_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_99_MUX_inst_X,
         RoundReg_Inst_ff_SDE_99_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_100_next_state,
         RoundReg_Inst_ff_SDE_100_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_100_MUX_inst_X,
         RoundReg_Inst_ff_SDE_100_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_101_next_state,
         RoundReg_Inst_ff_SDE_101_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_101_MUX_inst_X,
         RoundReg_Inst_ff_SDE_101_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_102_next_state,
         RoundReg_Inst_ff_SDE_102_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_102_MUX_inst_X,
         RoundReg_Inst_ff_SDE_102_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_103_next_state,
         RoundReg_Inst_ff_SDE_103_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_103_MUX_inst_X,
         RoundReg_Inst_ff_SDE_103_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_104_next_state,
         RoundReg_Inst_ff_SDE_104_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_104_MUX_inst_X,
         RoundReg_Inst_ff_SDE_104_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_105_next_state,
         RoundReg_Inst_ff_SDE_105_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_105_MUX_inst_X,
         RoundReg_Inst_ff_SDE_105_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_106_next_state,
         RoundReg_Inst_ff_SDE_106_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_106_MUX_inst_X,
         RoundReg_Inst_ff_SDE_106_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_107_next_state,
         RoundReg_Inst_ff_SDE_107_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_107_MUX_inst_X,
         RoundReg_Inst_ff_SDE_107_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_108_next_state,
         RoundReg_Inst_ff_SDE_108_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_108_MUX_inst_X,
         RoundReg_Inst_ff_SDE_108_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_109_next_state,
         RoundReg_Inst_ff_SDE_109_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_109_MUX_inst_X,
         RoundReg_Inst_ff_SDE_109_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_110_next_state,
         RoundReg_Inst_ff_SDE_110_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_110_MUX_inst_X,
         RoundReg_Inst_ff_SDE_110_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_111_next_state,
         RoundReg_Inst_ff_SDE_111_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_111_MUX_inst_X,
         RoundReg_Inst_ff_SDE_111_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_112_next_state,
         RoundReg_Inst_ff_SDE_112_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_112_MUX_inst_X,
         RoundReg_Inst_ff_SDE_112_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_113_next_state,
         RoundReg_Inst_ff_SDE_113_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_113_MUX_inst_X,
         RoundReg_Inst_ff_SDE_113_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_114_next_state,
         RoundReg_Inst_ff_SDE_114_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_114_MUX_inst_X,
         RoundReg_Inst_ff_SDE_114_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_115_next_state,
         RoundReg_Inst_ff_SDE_115_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_115_MUX_inst_X,
         RoundReg_Inst_ff_SDE_115_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_116_next_state,
         RoundReg_Inst_ff_SDE_116_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_116_MUX_inst_X,
         RoundReg_Inst_ff_SDE_116_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_117_next_state,
         RoundReg_Inst_ff_SDE_117_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_117_MUX_inst_X,
         RoundReg_Inst_ff_SDE_117_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_118_next_state,
         RoundReg_Inst_ff_SDE_118_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_118_MUX_inst_X,
         RoundReg_Inst_ff_SDE_118_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_119_next_state,
         RoundReg_Inst_ff_SDE_119_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_119_MUX_inst_X,
         RoundReg_Inst_ff_SDE_119_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_120_next_state,
         RoundReg_Inst_ff_SDE_120_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_120_MUX_inst_X,
         RoundReg_Inst_ff_SDE_120_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_121_next_state,
         RoundReg_Inst_ff_SDE_121_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_121_MUX_inst_X,
         RoundReg_Inst_ff_SDE_121_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_122_next_state,
         RoundReg_Inst_ff_SDE_122_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_122_MUX_inst_X,
         RoundReg_Inst_ff_SDE_122_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_123_next_state,
         RoundReg_Inst_ff_SDE_123_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_123_MUX_inst_X,
         RoundReg_Inst_ff_SDE_123_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_124_next_state,
         RoundReg_Inst_ff_SDE_124_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_124_MUX_inst_X,
         RoundReg_Inst_ff_SDE_124_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_125_next_state,
         RoundReg_Inst_ff_SDE_125_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_125_MUX_inst_X,
         RoundReg_Inst_ff_SDE_125_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_126_next_state,
         RoundReg_Inst_ff_SDE_126_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_126_MUX_inst_X,
         RoundReg_Inst_ff_SDE_126_current_state_reg_QN,
         RoundReg_Inst_ff_SDE_127_next_state,
         RoundReg_Inst_ff_SDE_127_MUX_inst_Y,
         RoundReg_Inst_ff_SDE_127_MUX_inst_X,
         RoundReg_Inst_ff_SDE_127_current_state_reg_QN,
         SubBytesIns_Inst_Sbox_0_L29, SubBytesIns_Inst_Sbox_0_L28,
         SubBytesIns_Inst_Sbox_0_L27, SubBytesIns_Inst_Sbox_0_L26,
         SubBytesIns_Inst_Sbox_0_L25, SubBytesIns_Inst_Sbox_0_L24,
         SubBytesIns_Inst_Sbox_0_L23, SubBytesIns_Inst_Sbox_0_L22,
         SubBytesIns_Inst_Sbox_0_L21, SubBytesIns_Inst_Sbox_0_L20,
         SubBytesIns_Inst_Sbox_0_L19, SubBytesIns_Inst_Sbox_0_L18,
         SubBytesIns_Inst_Sbox_0_L17, SubBytesIns_Inst_Sbox_0_L16,
         SubBytesIns_Inst_Sbox_0_L15, SubBytesIns_Inst_Sbox_0_L14,
         SubBytesIns_Inst_Sbox_0_L13, SubBytesIns_Inst_Sbox_0_L12,
         SubBytesIns_Inst_Sbox_0_L11, SubBytesIns_Inst_Sbox_0_L10,
         SubBytesIns_Inst_Sbox_0_L9, SubBytesIns_Inst_Sbox_0_L8,
         SubBytesIns_Inst_Sbox_0_L7, SubBytesIns_Inst_Sbox_0_L6,
         SubBytesIns_Inst_Sbox_0_L5, SubBytesIns_Inst_Sbox_0_L4,
         SubBytesIns_Inst_Sbox_0_L3, SubBytesIns_Inst_Sbox_0_L2,
         SubBytesIns_Inst_Sbox_0_L1, SubBytesIns_Inst_Sbox_0_L0,
         SubBytesIns_Inst_Sbox_0_M63, SubBytesIns_Inst_Sbox_0_M62,
         SubBytesIns_Inst_Sbox_0_M61, SubBytesIns_Inst_Sbox_0_M60,
         SubBytesIns_Inst_Sbox_0_M59, SubBytesIns_Inst_Sbox_0_M58,
         SubBytesIns_Inst_Sbox_0_M57, SubBytesIns_Inst_Sbox_0_M56,
         SubBytesIns_Inst_Sbox_0_M55, SubBytesIns_Inst_Sbox_0_M54,
         SubBytesIns_Inst_Sbox_0_M53, SubBytesIns_Inst_Sbox_0_M52,
         SubBytesIns_Inst_Sbox_0_M51, SubBytesIns_Inst_Sbox_0_M50,
         SubBytesIns_Inst_Sbox_0_M49, SubBytesIns_Inst_Sbox_0_M48,
         SubBytesIns_Inst_Sbox_0_M47, SubBytesIns_Inst_Sbox_0_M46,
         SubBytesIns_Inst_Sbox_0_M45, SubBytesIns_Inst_Sbox_0_M44,
         SubBytesIns_Inst_Sbox_0_M43, SubBytesIns_Inst_Sbox_0_M42,
         SubBytesIns_Inst_Sbox_0_M41, SubBytesIns_Inst_Sbox_0_M40,
         SubBytesIns_Inst_Sbox_0_M39, SubBytesIns_Inst_Sbox_0_M38,
         SubBytesIns_Inst_Sbox_0_M37, SubBytesIns_Inst_Sbox_0_M36,
         SubBytesIns_Inst_Sbox_0_M35, SubBytesIns_Inst_Sbox_0_M34,
         SubBytesIns_Inst_Sbox_0_M33, SubBytesIns_Inst_Sbox_0_M32,
         SubBytesIns_Inst_Sbox_0_M31, SubBytesIns_Inst_Sbox_0_M30,
         SubBytesIns_Inst_Sbox_0_M29, SubBytesIns_Inst_Sbox_0_M28,
         SubBytesIns_Inst_Sbox_0_M27, SubBytesIns_Inst_Sbox_0_M26,
         SubBytesIns_Inst_Sbox_0_M25, SubBytesIns_Inst_Sbox_0_M24,
         SubBytesIns_Inst_Sbox_0_M23, SubBytesIns_Inst_Sbox_0_M22,
         SubBytesIns_Inst_Sbox_0_M21, SubBytesIns_Inst_Sbox_0_M20,
         SubBytesIns_Inst_Sbox_0_M19, SubBytesIns_Inst_Sbox_0_M18,
         SubBytesIns_Inst_Sbox_0_M17, SubBytesIns_Inst_Sbox_0_M16,
         SubBytesIns_Inst_Sbox_0_M15, SubBytesIns_Inst_Sbox_0_M14,
         SubBytesIns_Inst_Sbox_0_M13, SubBytesIns_Inst_Sbox_0_M12,
         SubBytesIns_Inst_Sbox_0_M11, SubBytesIns_Inst_Sbox_0_M10,
         SubBytesIns_Inst_Sbox_0_M9, SubBytesIns_Inst_Sbox_0_M8,
         SubBytesIns_Inst_Sbox_0_M7, SubBytesIns_Inst_Sbox_0_M6,
         SubBytesIns_Inst_Sbox_0_M5, SubBytesIns_Inst_Sbox_0_M4,
         SubBytesIns_Inst_Sbox_0_M3, SubBytesIns_Inst_Sbox_0_M2,
         SubBytesIns_Inst_Sbox_0_M1, SubBytesIns_Inst_Sbox_0_T27,
         SubBytesIns_Inst_Sbox_0_T26, SubBytesIns_Inst_Sbox_0_T25,
         SubBytesIns_Inst_Sbox_0_T24, SubBytesIns_Inst_Sbox_0_T23,
         SubBytesIns_Inst_Sbox_0_T22, SubBytesIns_Inst_Sbox_0_T21,
         SubBytesIns_Inst_Sbox_0_T20, SubBytesIns_Inst_Sbox_0_T19,
         SubBytesIns_Inst_Sbox_0_T18, SubBytesIns_Inst_Sbox_0_T17,
         SubBytesIns_Inst_Sbox_0_T16, SubBytesIns_Inst_Sbox_0_T15,
         SubBytesIns_Inst_Sbox_0_T14, SubBytesIns_Inst_Sbox_0_T13,
         SubBytesIns_Inst_Sbox_0_T12, SubBytesIns_Inst_Sbox_0_T11,
         SubBytesIns_Inst_Sbox_0_T10, SubBytesIns_Inst_Sbox_0_T9,
         SubBytesIns_Inst_Sbox_0_T8, SubBytesIns_Inst_Sbox_0_T7,
         SubBytesIns_Inst_Sbox_0_T6, SubBytesIns_Inst_Sbox_0_T5,
         SubBytesIns_Inst_Sbox_0_T4, SubBytesIns_Inst_Sbox_0_T3,
         SubBytesIns_Inst_Sbox_0_T2, SubBytesIns_Inst_Sbox_0_T1,
         SubBytesIns_Inst_Sbox_1_L29, SubBytesIns_Inst_Sbox_1_L28,
         SubBytesIns_Inst_Sbox_1_L27, SubBytesIns_Inst_Sbox_1_L26,
         SubBytesIns_Inst_Sbox_1_L25, SubBytesIns_Inst_Sbox_1_L24,
         SubBytesIns_Inst_Sbox_1_L23, SubBytesIns_Inst_Sbox_1_L22,
         SubBytesIns_Inst_Sbox_1_L21, SubBytesIns_Inst_Sbox_1_L20,
         SubBytesIns_Inst_Sbox_1_L19, SubBytesIns_Inst_Sbox_1_L18,
         SubBytesIns_Inst_Sbox_1_L17, SubBytesIns_Inst_Sbox_1_L16,
         SubBytesIns_Inst_Sbox_1_L15, SubBytesIns_Inst_Sbox_1_L14,
         SubBytesIns_Inst_Sbox_1_L13, SubBytesIns_Inst_Sbox_1_L12,
         SubBytesIns_Inst_Sbox_1_L11, SubBytesIns_Inst_Sbox_1_L10,
         SubBytesIns_Inst_Sbox_1_L9, SubBytesIns_Inst_Sbox_1_L8,
         SubBytesIns_Inst_Sbox_1_L7, SubBytesIns_Inst_Sbox_1_L6,
         SubBytesIns_Inst_Sbox_1_L5, SubBytesIns_Inst_Sbox_1_L4,
         SubBytesIns_Inst_Sbox_1_L3, SubBytesIns_Inst_Sbox_1_L2,
         SubBytesIns_Inst_Sbox_1_L1, SubBytesIns_Inst_Sbox_1_L0,
         SubBytesIns_Inst_Sbox_1_M63, SubBytesIns_Inst_Sbox_1_M62,
         SubBytesIns_Inst_Sbox_1_M61, SubBytesIns_Inst_Sbox_1_M60,
         SubBytesIns_Inst_Sbox_1_M59, SubBytesIns_Inst_Sbox_1_M58,
         SubBytesIns_Inst_Sbox_1_M57, SubBytesIns_Inst_Sbox_1_M56,
         SubBytesIns_Inst_Sbox_1_M55, SubBytesIns_Inst_Sbox_1_M54,
         SubBytesIns_Inst_Sbox_1_M53, SubBytesIns_Inst_Sbox_1_M52,
         SubBytesIns_Inst_Sbox_1_M51, SubBytesIns_Inst_Sbox_1_M50,
         SubBytesIns_Inst_Sbox_1_M49, SubBytesIns_Inst_Sbox_1_M48,
         SubBytesIns_Inst_Sbox_1_M47, SubBytesIns_Inst_Sbox_1_M46,
         SubBytesIns_Inst_Sbox_1_M45, SubBytesIns_Inst_Sbox_1_M44,
         SubBytesIns_Inst_Sbox_1_M43, SubBytesIns_Inst_Sbox_1_M42,
         SubBytesIns_Inst_Sbox_1_M41, SubBytesIns_Inst_Sbox_1_M40,
         SubBytesIns_Inst_Sbox_1_M39, SubBytesIns_Inst_Sbox_1_M38,
         SubBytesIns_Inst_Sbox_1_M37, SubBytesIns_Inst_Sbox_1_M36,
         SubBytesIns_Inst_Sbox_1_M35, SubBytesIns_Inst_Sbox_1_M34,
         SubBytesIns_Inst_Sbox_1_M33, SubBytesIns_Inst_Sbox_1_M32,
         SubBytesIns_Inst_Sbox_1_M31, SubBytesIns_Inst_Sbox_1_M30,
         SubBytesIns_Inst_Sbox_1_M29, SubBytesIns_Inst_Sbox_1_M28,
         SubBytesIns_Inst_Sbox_1_M27, SubBytesIns_Inst_Sbox_1_M26,
         SubBytesIns_Inst_Sbox_1_M25, SubBytesIns_Inst_Sbox_1_M24,
         SubBytesIns_Inst_Sbox_1_M23, SubBytesIns_Inst_Sbox_1_M22,
         SubBytesIns_Inst_Sbox_1_M21, SubBytesIns_Inst_Sbox_1_M20,
         SubBytesIns_Inst_Sbox_1_M19, SubBytesIns_Inst_Sbox_1_M18,
         SubBytesIns_Inst_Sbox_1_M17, SubBytesIns_Inst_Sbox_1_M16,
         SubBytesIns_Inst_Sbox_1_M15, SubBytesIns_Inst_Sbox_1_M14,
         SubBytesIns_Inst_Sbox_1_M13, SubBytesIns_Inst_Sbox_1_M12,
         SubBytesIns_Inst_Sbox_1_M11, SubBytesIns_Inst_Sbox_1_M10,
         SubBytesIns_Inst_Sbox_1_M9, SubBytesIns_Inst_Sbox_1_M8,
         SubBytesIns_Inst_Sbox_1_M7, SubBytesIns_Inst_Sbox_1_M6,
         SubBytesIns_Inst_Sbox_1_M5, SubBytesIns_Inst_Sbox_1_M4,
         SubBytesIns_Inst_Sbox_1_M3, SubBytesIns_Inst_Sbox_1_M2,
         SubBytesIns_Inst_Sbox_1_M1, SubBytesIns_Inst_Sbox_1_T27,
         SubBytesIns_Inst_Sbox_1_T26, SubBytesIns_Inst_Sbox_1_T25,
         SubBytesIns_Inst_Sbox_1_T24, SubBytesIns_Inst_Sbox_1_T23,
         SubBytesIns_Inst_Sbox_1_T22, SubBytesIns_Inst_Sbox_1_T21,
         SubBytesIns_Inst_Sbox_1_T20, SubBytesIns_Inst_Sbox_1_T19,
         SubBytesIns_Inst_Sbox_1_T18, SubBytesIns_Inst_Sbox_1_T17,
         SubBytesIns_Inst_Sbox_1_T16, SubBytesIns_Inst_Sbox_1_T15,
         SubBytesIns_Inst_Sbox_1_T14, SubBytesIns_Inst_Sbox_1_T13,
         SubBytesIns_Inst_Sbox_1_T12, SubBytesIns_Inst_Sbox_1_T11,
         SubBytesIns_Inst_Sbox_1_T10, SubBytesIns_Inst_Sbox_1_T9,
         SubBytesIns_Inst_Sbox_1_T8, SubBytesIns_Inst_Sbox_1_T7,
         SubBytesIns_Inst_Sbox_1_T6, SubBytesIns_Inst_Sbox_1_T5,
         SubBytesIns_Inst_Sbox_1_T4, SubBytesIns_Inst_Sbox_1_T3,
         SubBytesIns_Inst_Sbox_1_T2, SubBytesIns_Inst_Sbox_1_T1,
         SubBytesIns_Inst_Sbox_2_L29, SubBytesIns_Inst_Sbox_2_L28,
         SubBytesIns_Inst_Sbox_2_L27, SubBytesIns_Inst_Sbox_2_L26,
         SubBytesIns_Inst_Sbox_2_L25, SubBytesIns_Inst_Sbox_2_L24,
         SubBytesIns_Inst_Sbox_2_L23, SubBytesIns_Inst_Sbox_2_L22,
         SubBytesIns_Inst_Sbox_2_L21, SubBytesIns_Inst_Sbox_2_L20,
         SubBytesIns_Inst_Sbox_2_L19, SubBytesIns_Inst_Sbox_2_L18,
         SubBytesIns_Inst_Sbox_2_L17, SubBytesIns_Inst_Sbox_2_L16,
         SubBytesIns_Inst_Sbox_2_L15, SubBytesIns_Inst_Sbox_2_L14,
         SubBytesIns_Inst_Sbox_2_L13, SubBytesIns_Inst_Sbox_2_L12,
         SubBytesIns_Inst_Sbox_2_L11, SubBytesIns_Inst_Sbox_2_L10,
         SubBytesIns_Inst_Sbox_2_L9, SubBytesIns_Inst_Sbox_2_L8,
         SubBytesIns_Inst_Sbox_2_L7, SubBytesIns_Inst_Sbox_2_L6,
         SubBytesIns_Inst_Sbox_2_L5, SubBytesIns_Inst_Sbox_2_L4,
         SubBytesIns_Inst_Sbox_2_L3, SubBytesIns_Inst_Sbox_2_L2,
         SubBytesIns_Inst_Sbox_2_L1, SubBytesIns_Inst_Sbox_2_L0,
         SubBytesIns_Inst_Sbox_2_M63, SubBytesIns_Inst_Sbox_2_M62,
         SubBytesIns_Inst_Sbox_2_M61, SubBytesIns_Inst_Sbox_2_M60,
         SubBytesIns_Inst_Sbox_2_M59, SubBytesIns_Inst_Sbox_2_M58,
         SubBytesIns_Inst_Sbox_2_M57, SubBytesIns_Inst_Sbox_2_M56,
         SubBytesIns_Inst_Sbox_2_M55, SubBytesIns_Inst_Sbox_2_M54,
         SubBytesIns_Inst_Sbox_2_M53, SubBytesIns_Inst_Sbox_2_M52,
         SubBytesIns_Inst_Sbox_2_M51, SubBytesIns_Inst_Sbox_2_M50,
         SubBytesIns_Inst_Sbox_2_M49, SubBytesIns_Inst_Sbox_2_M48,
         SubBytesIns_Inst_Sbox_2_M47, SubBytesIns_Inst_Sbox_2_M46,
         SubBytesIns_Inst_Sbox_2_M45, SubBytesIns_Inst_Sbox_2_M44,
         SubBytesIns_Inst_Sbox_2_M43, SubBytesIns_Inst_Sbox_2_M42,
         SubBytesIns_Inst_Sbox_2_M41, SubBytesIns_Inst_Sbox_2_M40,
         SubBytesIns_Inst_Sbox_2_M39, SubBytesIns_Inst_Sbox_2_M38,
         SubBytesIns_Inst_Sbox_2_M37, SubBytesIns_Inst_Sbox_2_M36,
         SubBytesIns_Inst_Sbox_2_M35, SubBytesIns_Inst_Sbox_2_M34,
         SubBytesIns_Inst_Sbox_2_M33, SubBytesIns_Inst_Sbox_2_M32,
         SubBytesIns_Inst_Sbox_2_M31, SubBytesIns_Inst_Sbox_2_M30,
         SubBytesIns_Inst_Sbox_2_M29, SubBytesIns_Inst_Sbox_2_M28,
         SubBytesIns_Inst_Sbox_2_M27, SubBytesIns_Inst_Sbox_2_M26,
         SubBytesIns_Inst_Sbox_2_M25, SubBytesIns_Inst_Sbox_2_M24,
         SubBytesIns_Inst_Sbox_2_M23, SubBytesIns_Inst_Sbox_2_M22,
         SubBytesIns_Inst_Sbox_2_M21, SubBytesIns_Inst_Sbox_2_M20,
         SubBytesIns_Inst_Sbox_2_M19, SubBytesIns_Inst_Sbox_2_M18,
         SubBytesIns_Inst_Sbox_2_M17, SubBytesIns_Inst_Sbox_2_M16,
         SubBytesIns_Inst_Sbox_2_M15, SubBytesIns_Inst_Sbox_2_M14,
         SubBytesIns_Inst_Sbox_2_M13, SubBytesIns_Inst_Sbox_2_M12,
         SubBytesIns_Inst_Sbox_2_M11, SubBytesIns_Inst_Sbox_2_M10,
         SubBytesIns_Inst_Sbox_2_M9, SubBytesIns_Inst_Sbox_2_M8,
         SubBytesIns_Inst_Sbox_2_M7, SubBytesIns_Inst_Sbox_2_M6,
         SubBytesIns_Inst_Sbox_2_M5, SubBytesIns_Inst_Sbox_2_M4,
         SubBytesIns_Inst_Sbox_2_M3, SubBytesIns_Inst_Sbox_2_M2,
         SubBytesIns_Inst_Sbox_2_M1, SubBytesIns_Inst_Sbox_2_T27,
         SubBytesIns_Inst_Sbox_2_T26, SubBytesIns_Inst_Sbox_2_T25,
         SubBytesIns_Inst_Sbox_2_T24, SubBytesIns_Inst_Sbox_2_T23,
         SubBytesIns_Inst_Sbox_2_T22, SubBytesIns_Inst_Sbox_2_T21,
         SubBytesIns_Inst_Sbox_2_T20, SubBytesIns_Inst_Sbox_2_T19,
         SubBytesIns_Inst_Sbox_2_T18, SubBytesIns_Inst_Sbox_2_T17,
         SubBytesIns_Inst_Sbox_2_T16, SubBytesIns_Inst_Sbox_2_T15,
         SubBytesIns_Inst_Sbox_2_T14, SubBytesIns_Inst_Sbox_2_T13,
         SubBytesIns_Inst_Sbox_2_T12, SubBytesIns_Inst_Sbox_2_T11,
         SubBytesIns_Inst_Sbox_2_T10, SubBytesIns_Inst_Sbox_2_T9,
         SubBytesIns_Inst_Sbox_2_T8, SubBytesIns_Inst_Sbox_2_T7,
         SubBytesIns_Inst_Sbox_2_T6, SubBytesIns_Inst_Sbox_2_T5,
         SubBytesIns_Inst_Sbox_2_T4, SubBytesIns_Inst_Sbox_2_T3,
         SubBytesIns_Inst_Sbox_2_T2, SubBytesIns_Inst_Sbox_2_T1,
         SubBytesIns_Inst_Sbox_3_L29, SubBytesIns_Inst_Sbox_3_L28,
         SubBytesIns_Inst_Sbox_3_L27, SubBytesIns_Inst_Sbox_3_L26,
         SubBytesIns_Inst_Sbox_3_L25, SubBytesIns_Inst_Sbox_3_L24,
         SubBytesIns_Inst_Sbox_3_L23, SubBytesIns_Inst_Sbox_3_L22,
         SubBytesIns_Inst_Sbox_3_L21, SubBytesIns_Inst_Sbox_3_L20,
         SubBytesIns_Inst_Sbox_3_L19, SubBytesIns_Inst_Sbox_3_L18,
         SubBytesIns_Inst_Sbox_3_L17, SubBytesIns_Inst_Sbox_3_L16,
         SubBytesIns_Inst_Sbox_3_L15, SubBytesIns_Inst_Sbox_3_L14,
         SubBytesIns_Inst_Sbox_3_L13, SubBytesIns_Inst_Sbox_3_L12,
         SubBytesIns_Inst_Sbox_3_L11, SubBytesIns_Inst_Sbox_3_L10,
         SubBytesIns_Inst_Sbox_3_L9, SubBytesIns_Inst_Sbox_3_L8,
         SubBytesIns_Inst_Sbox_3_L7, SubBytesIns_Inst_Sbox_3_L6,
         SubBytesIns_Inst_Sbox_3_L5, SubBytesIns_Inst_Sbox_3_L4,
         SubBytesIns_Inst_Sbox_3_L3, SubBytesIns_Inst_Sbox_3_L2,
         SubBytesIns_Inst_Sbox_3_L1, SubBytesIns_Inst_Sbox_3_L0,
         SubBytesIns_Inst_Sbox_3_M63, SubBytesIns_Inst_Sbox_3_M62,
         SubBytesIns_Inst_Sbox_3_M61, SubBytesIns_Inst_Sbox_3_M60,
         SubBytesIns_Inst_Sbox_3_M59, SubBytesIns_Inst_Sbox_3_M58,
         SubBytesIns_Inst_Sbox_3_M57, SubBytesIns_Inst_Sbox_3_M56,
         SubBytesIns_Inst_Sbox_3_M55, SubBytesIns_Inst_Sbox_3_M54,
         SubBytesIns_Inst_Sbox_3_M53, SubBytesIns_Inst_Sbox_3_M52,
         SubBytesIns_Inst_Sbox_3_M51, SubBytesIns_Inst_Sbox_3_M50,
         SubBytesIns_Inst_Sbox_3_M49, SubBytesIns_Inst_Sbox_3_M48,
         SubBytesIns_Inst_Sbox_3_M47, SubBytesIns_Inst_Sbox_3_M46,
         SubBytesIns_Inst_Sbox_3_M45, SubBytesIns_Inst_Sbox_3_M44,
         SubBytesIns_Inst_Sbox_3_M43, SubBytesIns_Inst_Sbox_3_M42,
         SubBytesIns_Inst_Sbox_3_M41, SubBytesIns_Inst_Sbox_3_M40,
         SubBytesIns_Inst_Sbox_3_M39, SubBytesIns_Inst_Sbox_3_M38,
         SubBytesIns_Inst_Sbox_3_M37, SubBytesIns_Inst_Sbox_3_M36,
         SubBytesIns_Inst_Sbox_3_M35, SubBytesIns_Inst_Sbox_3_M34,
         SubBytesIns_Inst_Sbox_3_M33, SubBytesIns_Inst_Sbox_3_M32,
         SubBytesIns_Inst_Sbox_3_M31, SubBytesIns_Inst_Sbox_3_M30,
         SubBytesIns_Inst_Sbox_3_M29, SubBytesIns_Inst_Sbox_3_M28,
         SubBytesIns_Inst_Sbox_3_M27, SubBytesIns_Inst_Sbox_3_M26,
         SubBytesIns_Inst_Sbox_3_M25, SubBytesIns_Inst_Sbox_3_M24,
         SubBytesIns_Inst_Sbox_3_M23, SubBytesIns_Inst_Sbox_3_M22,
         SubBytesIns_Inst_Sbox_3_M21, SubBytesIns_Inst_Sbox_3_M20,
         SubBytesIns_Inst_Sbox_3_M19, SubBytesIns_Inst_Sbox_3_M18,
         SubBytesIns_Inst_Sbox_3_M17, SubBytesIns_Inst_Sbox_3_M16,
         SubBytesIns_Inst_Sbox_3_M15, SubBytesIns_Inst_Sbox_3_M14,
         SubBytesIns_Inst_Sbox_3_M13, SubBytesIns_Inst_Sbox_3_M12,
         SubBytesIns_Inst_Sbox_3_M11, SubBytesIns_Inst_Sbox_3_M10,
         SubBytesIns_Inst_Sbox_3_M9, SubBytesIns_Inst_Sbox_3_M8,
         SubBytesIns_Inst_Sbox_3_M7, SubBytesIns_Inst_Sbox_3_M6,
         SubBytesIns_Inst_Sbox_3_M5, SubBytesIns_Inst_Sbox_3_M4,
         SubBytesIns_Inst_Sbox_3_M3, SubBytesIns_Inst_Sbox_3_M2,
         SubBytesIns_Inst_Sbox_3_M1, SubBytesIns_Inst_Sbox_3_T27,
         SubBytesIns_Inst_Sbox_3_T26, SubBytesIns_Inst_Sbox_3_T25,
         SubBytesIns_Inst_Sbox_3_T24, SubBytesIns_Inst_Sbox_3_T23,
         SubBytesIns_Inst_Sbox_3_T22, SubBytesIns_Inst_Sbox_3_T21,
         SubBytesIns_Inst_Sbox_3_T20, SubBytesIns_Inst_Sbox_3_T19,
         SubBytesIns_Inst_Sbox_3_T18, SubBytesIns_Inst_Sbox_3_T17,
         SubBytesIns_Inst_Sbox_3_T16, SubBytesIns_Inst_Sbox_3_T15,
         SubBytesIns_Inst_Sbox_3_T14, SubBytesIns_Inst_Sbox_3_T13,
         SubBytesIns_Inst_Sbox_3_T12, SubBytesIns_Inst_Sbox_3_T11,
         SubBytesIns_Inst_Sbox_3_T10, SubBytesIns_Inst_Sbox_3_T9,
         SubBytesIns_Inst_Sbox_3_T8, SubBytesIns_Inst_Sbox_3_T7,
         SubBytesIns_Inst_Sbox_3_T6, SubBytesIns_Inst_Sbox_3_T5,
         SubBytesIns_Inst_Sbox_3_T4, SubBytesIns_Inst_Sbox_3_T3,
         SubBytesIns_Inst_Sbox_3_T2, SubBytesIns_Inst_Sbox_3_T1,
         SubBytesIns_Inst_Sbox_4_L29, SubBytesIns_Inst_Sbox_4_L28,
         SubBytesIns_Inst_Sbox_4_L27, SubBytesIns_Inst_Sbox_4_L26,
         SubBytesIns_Inst_Sbox_4_L25, SubBytesIns_Inst_Sbox_4_L24,
         SubBytesIns_Inst_Sbox_4_L23, SubBytesIns_Inst_Sbox_4_L22,
         SubBytesIns_Inst_Sbox_4_L21, SubBytesIns_Inst_Sbox_4_L20,
         SubBytesIns_Inst_Sbox_4_L19, SubBytesIns_Inst_Sbox_4_L18,
         SubBytesIns_Inst_Sbox_4_L17, SubBytesIns_Inst_Sbox_4_L16,
         SubBytesIns_Inst_Sbox_4_L15, SubBytesIns_Inst_Sbox_4_L14,
         SubBytesIns_Inst_Sbox_4_L13, SubBytesIns_Inst_Sbox_4_L12,
         SubBytesIns_Inst_Sbox_4_L11, SubBytesIns_Inst_Sbox_4_L10,
         SubBytesIns_Inst_Sbox_4_L9, SubBytesIns_Inst_Sbox_4_L8,
         SubBytesIns_Inst_Sbox_4_L7, SubBytesIns_Inst_Sbox_4_L6,
         SubBytesIns_Inst_Sbox_4_L5, SubBytesIns_Inst_Sbox_4_L4,
         SubBytesIns_Inst_Sbox_4_L3, SubBytesIns_Inst_Sbox_4_L2,
         SubBytesIns_Inst_Sbox_4_L1, SubBytesIns_Inst_Sbox_4_L0,
         SubBytesIns_Inst_Sbox_4_M63, SubBytesIns_Inst_Sbox_4_M62,
         SubBytesIns_Inst_Sbox_4_M61, SubBytesIns_Inst_Sbox_4_M60,
         SubBytesIns_Inst_Sbox_4_M59, SubBytesIns_Inst_Sbox_4_M58,
         SubBytesIns_Inst_Sbox_4_M57, SubBytesIns_Inst_Sbox_4_M56,
         SubBytesIns_Inst_Sbox_4_M55, SubBytesIns_Inst_Sbox_4_M54,
         SubBytesIns_Inst_Sbox_4_M53, SubBytesIns_Inst_Sbox_4_M52,
         SubBytesIns_Inst_Sbox_4_M51, SubBytesIns_Inst_Sbox_4_M50,
         SubBytesIns_Inst_Sbox_4_M49, SubBytesIns_Inst_Sbox_4_M48,
         SubBytesIns_Inst_Sbox_4_M47, SubBytesIns_Inst_Sbox_4_M46,
         SubBytesIns_Inst_Sbox_4_M45, SubBytesIns_Inst_Sbox_4_M44,
         SubBytesIns_Inst_Sbox_4_M43, SubBytesIns_Inst_Sbox_4_M42,
         SubBytesIns_Inst_Sbox_4_M41, SubBytesIns_Inst_Sbox_4_M40,
         SubBytesIns_Inst_Sbox_4_M39, SubBytesIns_Inst_Sbox_4_M38,
         SubBytesIns_Inst_Sbox_4_M37, SubBytesIns_Inst_Sbox_4_M36,
         SubBytesIns_Inst_Sbox_4_M35, SubBytesIns_Inst_Sbox_4_M34,
         SubBytesIns_Inst_Sbox_4_M33, SubBytesIns_Inst_Sbox_4_M32,
         SubBytesIns_Inst_Sbox_4_M31, SubBytesIns_Inst_Sbox_4_M30,
         SubBytesIns_Inst_Sbox_4_M29, SubBytesIns_Inst_Sbox_4_M28,
         SubBytesIns_Inst_Sbox_4_M27, SubBytesIns_Inst_Sbox_4_M26,
         SubBytesIns_Inst_Sbox_4_M25, SubBytesIns_Inst_Sbox_4_M24,
         SubBytesIns_Inst_Sbox_4_M23, SubBytesIns_Inst_Sbox_4_M22,
         SubBytesIns_Inst_Sbox_4_M21, SubBytesIns_Inst_Sbox_4_M20,
         SubBytesIns_Inst_Sbox_4_M19, SubBytesIns_Inst_Sbox_4_M18,
         SubBytesIns_Inst_Sbox_4_M17, SubBytesIns_Inst_Sbox_4_M16,
         SubBytesIns_Inst_Sbox_4_M15, SubBytesIns_Inst_Sbox_4_M14,
         SubBytesIns_Inst_Sbox_4_M13, SubBytesIns_Inst_Sbox_4_M12,
         SubBytesIns_Inst_Sbox_4_M11, SubBytesIns_Inst_Sbox_4_M10,
         SubBytesIns_Inst_Sbox_4_M9, SubBytesIns_Inst_Sbox_4_M8,
         SubBytesIns_Inst_Sbox_4_M7, SubBytesIns_Inst_Sbox_4_M6,
         SubBytesIns_Inst_Sbox_4_M5, SubBytesIns_Inst_Sbox_4_M4,
         SubBytesIns_Inst_Sbox_4_M3, SubBytesIns_Inst_Sbox_4_M2,
         SubBytesIns_Inst_Sbox_4_M1, SubBytesIns_Inst_Sbox_4_T27,
         SubBytesIns_Inst_Sbox_4_T26, SubBytesIns_Inst_Sbox_4_T25,
         SubBytesIns_Inst_Sbox_4_T24, SubBytesIns_Inst_Sbox_4_T23,
         SubBytesIns_Inst_Sbox_4_T22, SubBytesIns_Inst_Sbox_4_T21,
         SubBytesIns_Inst_Sbox_4_T20, SubBytesIns_Inst_Sbox_4_T19,
         SubBytesIns_Inst_Sbox_4_T18, SubBytesIns_Inst_Sbox_4_T17,
         SubBytesIns_Inst_Sbox_4_T16, SubBytesIns_Inst_Sbox_4_T15,
         SubBytesIns_Inst_Sbox_4_T14, SubBytesIns_Inst_Sbox_4_T13,
         SubBytesIns_Inst_Sbox_4_T12, SubBytesIns_Inst_Sbox_4_T11,
         SubBytesIns_Inst_Sbox_4_T10, SubBytesIns_Inst_Sbox_4_T9,
         SubBytesIns_Inst_Sbox_4_T8, SubBytesIns_Inst_Sbox_4_T7,
         SubBytesIns_Inst_Sbox_4_T6, SubBytesIns_Inst_Sbox_4_T5,
         SubBytesIns_Inst_Sbox_4_T4, SubBytesIns_Inst_Sbox_4_T3,
         SubBytesIns_Inst_Sbox_4_T2, SubBytesIns_Inst_Sbox_4_T1,
         SubBytesIns_Inst_Sbox_5_L29, SubBytesIns_Inst_Sbox_5_L28,
         SubBytesIns_Inst_Sbox_5_L27, SubBytesIns_Inst_Sbox_5_L26,
         SubBytesIns_Inst_Sbox_5_L25, SubBytesIns_Inst_Sbox_5_L24,
         SubBytesIns_Inst_Sbox_5_L23, SubBytesIns_Inst_Sbox_5_L22,
         SubBytesIns_Inst_Sbox_5_L21, SubBytesIns_Inst_Sbox_5_L20,
         SubBytesIns_Inst_Sbox_5_L19, SubBytesIns_Inst_Sbox_5_L18,
         SubBytesIns_Inst_Sbox_5_L17, SubBytesIns_Inst_Sbox_5_L16,
         SubBytesIns_Inst_Sbox_5_L15, SubBytesIns_Inst_Sbox_5_L14,
         SubBytesIns_Inst_Sbox_5_L13, SubBytesIns_Inst_Sbox_5_L12,
         SubBytesIns_Inst_Sbox_5_L11, SubBytesIns_Inst_Sbox_5_L10,
         SubBytesIns_Inst_Sbox_5_L9, SubBytesIns_Inst_Sbox_5_L8,
         SubBytesIns_Inst_Sbox_5_L7, SubBytesIns_Inst_Sbox_5_L6,
         SubBytesIns_Inst_Sbox_5_L5, SubBytesIns_Inst_Sbox_5_L4,
         SubBytesIns_Inst_Sbox_5_L3, SubBytesIns_Inst_Sbox_5_L2,
         SubBytesIns_Inst_Sbox_5_L1, SubBytesIns_Inst_Sbox_5_L0,
         SubBytesIns_Inst_Sbox_5_M63, SubBytesIns_Inst_Sbox_5_M62,
         SubBytesIns_Inst_Sbox_5_M61, SubBytesIns_Inst_Sbox_5_M60,
         SubBytesIns_Inst_Sbox_5_M59, SubBytesIns_Inst_Sbox_5_M58,
         SubBytesIns_Inst_Sbox_5_M57, SubBytesIns_Inst_Sbox_5_M56,
         SubBytesIns_Inst_Sbox_5_M55, SubBytesIns_Inst_Sbox_5_M54,
         SubBytesIns_Inst_Sbox_5_M53, SubBytesIns_Inst_Sbox_5_M52,
         SubBytesIns_Inst_Sbox_5_M51, SubBytesIns_Inst_Sbox_5_M50,
         SubBytesIns_Inst_Sbox_5_M49, SubBytesIns_Inst_Sbox_5_M48,
         SubBytesIns_Inst_Sbox_5_M47, SubBytesIns_Inst_Sbox_5_M46,
         SubBytesIns_Inst_Sbox_5_M45, SubBytesIns_Inst_Sbox_5_M44,
         SubBytesIns_Inst_Sbox_5_M43, SubBytesIns_Inst_Sbox_5_M42,
         SubBytesIns_Inst_Sbox_5_M41, SubBytesIns_Inst_Sbox_5_M40,
         SubBytesIns_Inst_Sbox_5_M39, SubBytesIns_Inst_Sbox_5_M38,
         SubBytesIns_Inst_Sbox_5_M37, SubBytesIns_Inst_Sbox_5_M36,
         SubBytesIns_Inst_Sbox_5_M35, SubBytesIns_Inst_Sbox_5_M34,
         SubBytesIns_Inst_Sbox_5_M33, SubBytesIns_Inst_Sbox_5_M32,
         SubBytesIns_Inst_Sbox_5_M31, SubBytesIns_Inst_Sbox_5_M30,
         SubBytesIns_Inst_Sbox_5_M29, SubBytesIns_Inst_Sbox_5_M28,
         SubBytesIns_Inst_Sbox_5_M27, SubBytesIns_Inst_Sbox_5_M26,
         SubBytesIns_Inst_Sbox_5_M25, SubBytesIns_Inst_Sbox_5_M24,
         SubBytesIns_Inst_Sbox_5_M23, SubBytesIns_Inst_Sbox_5_M22,
         SubBytesIns_Inst_Sbox_5_M21, SubBytesIns_Inst_Sbox_5_M20,
         SubBytesIns_Inst_Sbox_5_M19, SubBytesIns_Inst_Sbox_5_M18,
         SubBytesIns_Inst_Sbox_5_M17, SubBytesIns_Inst_Sbox_5_M16,
         SubBytesIns_Inst_Sbox_5_M15, SubBytesIns_Inst_Sbox_5_M14,
         SubBytesIns_Inst_Sbox_5_M13, SubBytesIns_Inst_Sbox_5_M12,
         SubBytesIns_Inst_Sbox_5_M11, SubBytesIns_Inst_Sbox_5_M10,
         SubBytesIns_Inst_Sbox_5_M9, SubBytesIns_Inst_Sbox_5_M8,
         SubBytesIns_Inst_Sbox_5_M7, SubBytesIns_Inst_Sbox_5_M6,
         SubBytesIns_Inst_Sbox_5_M5, SubBytesIns_Inst_Sbox_5_M4,
         SubBytesIns_Inst_Sbox_5_M3, SubBytesIns_Inst_Sbox_5_M2,
         SubBytesIns_Inst_Sbox_5_M1, SubBytesIns_Inst_Sbox_5_T27,
         SubBytesIns_Inst_Sbox_5_T26, SubBytesIns_Inst_Sbox_5_T25,
         SubBytesIns_Inst_Sbox_5_T24, SubBytesIns_Inst_Sbox_5_T23,
         SubBytesIns_Inst_Sbox_5_T22, SubBytesIns_Inst_Sbox_5_T21,
         SubBytesIns_Inst_Sbox_5_T20, SubBytesIns_Inst_Sbox_5_T19,
         SubBytesIns_Inst_Sbox_5_T18, SubBytesIns_Inst_Sbox_5_T17,
         SubBytesIns_Inst_Sbox_5_T16, SubBytesIns_Inst_Sbox_5_T15,
         SubBytesIns_Inst_Sbox_5_T14, SubBytesIns_Inst_Sbox_5_T13,
         SubBytesIns_Inst_Sbox_5_T12, SubBytesIns_Inst_Sbox_5_T11,
         SubBytesIns_Inst_Sbox_5_T10, SubBytesIns_Inst_Sbox_5_T9,
         SubBytesIns_Inst_Sbox_5_T8, SubBytesIns_Inst_Sbox_5_T7,
         SubBytesIns_Inst_Sbox_5_T6, SubBytesIns_Inst_Sbox_5_T5,
         SubBytesIns_Inst_Sbox_5_T4, SubBytesIns_Inst_Sbox_5_T3,
         SubBytesIns_Inst_Sbox_5_T2, SubBytesIns_Inst_Sbox_5_T1,
         SubBytesIns_Inst_Sbox_6_L29, SubBytesIns_Inst_Sbox_6_L28,
         SubBytesIns_Inst_Sbox_6_L27, SubBytesIns_Inst_Sbox_6_L26,
         SubBytesIns_Inst_Sbox_6_L25, SubBytesIns_Inst_Sbox_6_L24,
         SubBytesIns_Inst_Sbox_6_L23, SubBytesIns_Inst_Sbox_6_L22,
         SubBytesIns_Inst_Sbox_6_L21, SubBytesIns_Inst_Sbox_6_L20,
         SubBytesIns_Inst_Sbox_6_L19, SubBytesIns_Inst_Sbox_6_L18,
         SubBytesIns_Inst_Sbox_6_L17, SubBytesIns_Inst_Sbox_6_L16,
         SubBytesIns_Inst_Sbox_6_L15, SubBytesIns_Inst_Sbox_6_L14,
         SubBytesIns_Inst_Sbox_6_L13, SubBytesIns_Inst_Sbox_6_L12,
         SubBytesIns_Inst_Sbox_6_L11, SubBytesIns_Inst_Sbox_6_L10,
         SubBytesIns_Inst_Sbox_6_L9, SubBytesIns_Inst_Sbox_6_L8,
         SubBytesIns_Inst_Sbox_6_L7, SubBytesIns_Inst_Sbox_6_L6,
         SubBytesIns_Inst_Sbox_6_L5, SubBytesIns_Inst_Sbox_6_L4,
         SubBytesIns_Inst_Sbox_6_L3, SubBytesIns_Inst_Sbox_6_L2,
         SubBytesIns_Inst_Sbox_6_L1, SubBytesIns_Inst_Sbox_6_L0,
         SubBytesIns_Inst_Sbox_6_M63, SubBytesIns_Inst_Sbox_6_M62,
         SubBytesIns_Inst_Sbox_6_M61, SubBytesIns_Inst_Sbox_6_M60,
         SubBytesIns_Inst_Sbox_6_M59, SubBytesIns_Inst_Sbox_6_M58,
         SubBytesIns_Inst_Sbox_6_M57, SubBytesIns_Inst_Sbox_6_M56,
         SubBytesIns_Inst_Sbox_6_M55, SubBytesIns_Inst_Sbox_6_M54,
         SubBytesIns_Inst_Sbox_6_M53, SubBytesIns_Inst_Sbox_6_M52,
         SubBytesIns_Inst_Sbox_6_M51, SubBytesIns_Inst_Sbox_6_M50,
         SubBytesIns_Inst_Sbox_6_M49, SubBytesIns_Inst_Sbox_6_M48,
         SubBytesIns_Inst_Sbox_6_M47, SubBytesIns_Inst_Sbox_6_M46,
         SubBytesIns_Inst_Sbox_6_M45, SubBytesIns_Inst_Sbox_6_M44,
         SubBytesIns_Inst_Sbox_6_M43, SubBytesIns_Inst_Sbox_6_M42,
         SubBytesIns_Inst_Sbox_6_M41, SubBytesIns_Inst_Sbox_6_M40,
         SubBytesIns_Inst_Sbox_6_M39, SubBytesIns_Inst_Sbox_6_M38,
         SubBytesIns_Inst_Sbox_6_M37, SubBytesIns_Inst_Sbox_6_M36,
         SubBytesIns_Inst_Sbox_6_M35, SubBytesIns_Inst_Sbox_6_M34,
         SubBytesIns_Inst_Sbox_6_M33, SubBytesIns_Inst_Sbox_6_M32,
         SubBytesIns_Inst_Sbox_6_M31, SubBytesIns_Inst_Sbox_6_M30,
         SubBytesIns_Inst_Sbox_6_M29, SubBytesIns_Inst_Sbox_6_M28,
         SubBytesIns_Inst_Sbox_6_M27, SubBytesIns_Inst_Sbox_6_M26,
         SubBytesIns_Inst_Sbox_6_M25, SubBytesIns_Inst_Sbox_6_M24,
         SubBytesIns_Inst_Sbox_6_M23, SubBytesIns_Inst_Sbox_6_M22,
         SubBytesIns_Inst_Sbox_6_M21, SubBytesIns_Inst_Sbox_6_M20,
         SubBytesIns_Inst_Sbox_6_M19, SubBytesIns_Inst_Sbox_6_M18,
         SubBytesIns_Inst_Sbox_6_M17, SubBytesIns_Inst_Sbox_6_M16,
         SubBytesIns_Inst_Sbox_6_M15, SubBytesIns_Inst_Sbox_6_M14,
         SubBytesIns_Inst_Sbox_6_M13, SubBytesIns_Inst_Sbox_6_M12,
         SubBytesIns_Inst_Sbox_6_M11, SubBytesIns_Inst_Sbox_6_M10,
         SubBytesIns_Inst_Sbox_6_M9, SubBytesIns_Inst_Sbox_6_M8,
         SubBytesIns_Inst_Sbox_6_M7, SubBytesIns_Inst_Sbox_6_M6,
         SubBytesIns_Inst_Sbox_6_M5, SubBytesIns_Inst_Sbox_6_M4,
         SubBytesIns_Inst_Sbox_6_M3, SubBytesIns_Inst_Sbox_6_M2,
         SubBytesIns_Inst_Sbox_6_M1, SubBytesIns_Inst_Sbox_6_T27,
         SubBytesIns_Inst_Sbox_6_T26, SubBytesIns_Inst_Sbox_6_T25,
         SubBytesIns_Inst_Sbox_6_T24, SubBytesIns_Inst_Sbox_6_T23,
         SubBytesIns_Inst_Sbox_6_T22, SubBytesIns_Inst_Sbox_6_T21,
         SubBytesIns_Inst_Sbox_6_T20, SubBytesIns_Inst_Sbox_6_T19,
         SubBytesIns_Inst_Sbox_6_T18, SubBytesIns_Inst_Sbox_6_T17,
         SubBytesIns_Inst_Sbox_6_T16, SubBytesIns_Inst_Sbox_6_T15,
         SubBytesIns_Inst_Sbox_6_T14, SubBytesIns_Inst_Sbox_6_T13,
         SubBytesIns_Inst_Sbox_6_T12, SubBytesIns_Inst_Sbox_6_T11,
         SubBytesIns_Inst_Sbox_6_T10, SubBytesIns_Inst_Sbox_6_T9,
         SubBytesIns_Inst_Sbox_6_T8, SubBytesIns_Inst_Sbox_6_T7,
         SubBytesIns_Inst_Sbox_6_T6, SubBytesIns_Inst_Sbox_6_T5,
         SubBytesIns_Inst_Sbox_6_T4, SubBytesIns_Inst_Sbox_6_T3,
         SubBytesIns_Inst_Sbox_6_T2, SubBytesIns_Inst_Sbox_6_T1,
         SubBytesIns_Inst_Sbox_7_L29, SubBytesIns_Inst_Sbox_7_L28,
         SubBytesIns_Inst_Sbox_7_L27, SubBytesIns_Inst_Sbox_7_L26,
         SubBytesIns_Inst_Sbox_7_L25, SubBytesIns_Inst_Sbox_7_L24,
         SubBytesIns_Inst_Sbox_7_L23, SubBytesIns_Inst_Sbox_7_L22,
         SubBytesIns_Inst_Sbox_7_L21, SubBytesIns_Inst_Sbox_7_L20,
         SubBytesIns_Inst_Sbox_7_L19, SubBytesIns_Inst_Sbox_7_L18,
         SubBytesIns_Inst_Sbox_7_L17, SubBytesIns_Inst_Sbox_7_L16,
         SubBytesIns_Inst_Sbox_7_L15, SubBytesIns_Inst_Sbox_7_L14,
         SubBytesIns_Inst_Sbox_7_L13, SubBytesIns_Inst_Sbox_7_L12,
         SubBytesIns_Inst_Sbox_7_L11, SubBytesIns_Inst_Sbox_7_L10,
         SubBytesIns_Inst_Sbox_7_L9, SubBytesIns_Inst_Sbox_7_L8,
         SubBytesIns_Inst_Sbox_7_L7, SubBytesIns_Inst_Sbox_7_L6,
         SubBytesIns_Inst_Sbox_7_L5, SubBytesIns_Inst_Sbox_7_L4,
         SubBytesIns_Inst_Sbox_7_L3, SubBytesIns_Inst_Sbox_7_L2,
         SubBytesIns_Inst_Sbox_7_L1, SubBytesIns_Inst_Sbox_7_L0,
         SubBytesIns_Inst_Sbox_7_M63, SubBytesIns_Inst_Sbox_7_M62,
         SubBytesIns_Inst_Sbox_7_M61, SubBytesIns_Inst_Sbox_7_M60,
         SubBytesIns_Inst_Sbox_7_M59, SubBytesIns_Inst_Sbox_7_M58,
         SubBytesIns_Inst_Sbox_7_M57, SubBytesIns_Inst_Sbox_7_M56,
         SubBytesIns_Inst_Sbox_7_M55, SubBytesIns_Inst_Sbox_7_M54,
         SubBytesIns_Inst_Sbox_7_M53, SubBytesIns_Inst_Sbox_7_M52,
         SubBytesIns_Inst_Sbox_7_M51, SubBytesIns_Inst_Sbox_7_M50,
         SubBytesIns_Inst_Sbox_7_M49, SubBytesIns_Inst_Sbox_7_M48,
         SubBytesIns_Inst_Sbox_7_M47, SubBytesIns_Inst_Sbox_7_M46,
         SubBytesIns_Inst_Sbox_7_M45, SubBytesIns_Inst_Sbox_7_M44,
         SubBytesIns_Inst_Sbox_7_M43, SubBytesIns_Inst_Sbox_7_M42,
         SubBytesIns_Inst_Sbox_7_M41, SubBytesIns_Inst_Sbox_7_M40,
         SubBytesIns_Inst_Sbox_7_M39, SubBytesIns_Inst_Sbox_7_M38,
         SubBytesIns_Inst_Sbox_7_M37, SubBytesIns_Inst_Sbox_7_M36,
         SubBytesIns_Inst_Sbox_7_M35, SubBytesIns_Inst_Sbox_7_M34,
         SubBytesIns_Inst_Sbox_7_M33, SubBytesIns_Inst_Sbox_7_M32,
         SubBytesIns_Inst_Sbox_7_M31, SubBytesIns_Inst_Sbox_7_M30,
         SubBytesIns_Inst_Sbox_7_M29, SubBytesIns_Inst_Sbox_7_M28,
         SubBytesIns_Inst_Sbox_7_M27, SubBytesIns_Inst_Sbox_7_M26,
         SubBytesIns_Inst_Sbox_7_M25, SubBytesIns_Inst_Sbox_7_M24,
         SubBytesIns_Inst_Sbox_7_M23, SubBytesIns_Inst_Sbox_7_M22,
         SubBytesIns_Inst_Sbox_7_M21, SubBytesIns_Inst_Sbox_7_M20,
         SubBytesIns_Inst_Sbox_7_M19, SubBytesIns_Inst_Sbox_7_M18,
         SubBytesIns_Inst_Sbox_7_M17, SubBytesIns_Inst_Sbox_7_M16,
         SubBytesIns_Inst_Sbox_7_M15, SubBytesIns_Inst_Sbox_7_M14,
         SubBytesIns_Inst_Sbox_7_M13, SubBytesIns_Inst_Sbox_7_M12,
         SubBytesIns_Inst_Sbox_7_M11, SubBytesIns_Inst_Sbox_7_M10,
         SubBytesIns_Inst_Sbox_7_M9, SubBytesIns_Inst_Sbox_7_M8,
         SubBytesIns_Inst_Sbox_7_M7, SubBytesIns_Inst_Sbox_7_M6,
         SubBytesIns_Inst_Sbox_7_M5, SubBytesIns_Inst_Sbox_7_M4,
         SubBytesIns_Inst_Sbox_7_M3, SubBytesIns_Inst_Sbox_7_M2,
         SubBytesIns_Inst_Sbox_7_M1, SubBytesIns_Inst_Sbox_7_T27,
         SubBytesIns_Inst_Sbox_7_T26, SubBytesIns_Inst_Sbox_7_T25,
         SubBytesIns_Inst_Sbox_7_T24, SubBytesIns_Inst_Sbox_7_T23,
         SubBytesIns_Inst_Sbox_7_T22, SubBytesIns_Inst_Sbox_7_T21,
         SubBytesIns_Inst_Sbox_7_T20, SubBytesIns_Inst_Sbox_7_T19,
         SubBytesIns_Inst_Sbox_7_T18, SubBytesIns_Inst_Sbox_7_T17,
         SubBytesIns_Inst_Sbox_7_T16, SubBytesIns_Inst_Sbox_7_T15,
         SubBytesIns_Inst_Sbox_7_T14, SubBytesIns_Inst_Sbox_7_T13,
         SubBytesIns_Inst_Sbox_7_T12, SubBytesIns_Inst_Sbox_7_T11,
         SubBytesIns_Inst_Sbox_7_T10, SubBytesIns_Inst_Sbox_7_T9,
         SubBytesIns_Inst_Sbox_7_T8, SubBytesIns_Inst_Sbox_7_T7,
         SubBytesIns_Inst_Sbox_7_T6, SubBytesIns_Inst_Sbox_7_T5,
         SubBytesIns_Inst_Sbox_7_T4, SubBytesIns_Inst_Sbox_7_T3,
         SubBytesIns_Inst_Sbox_7_T2, SubBytesIns_Inst_Sbox_7_T1,
         SubBytesIns_Inst_Sbox_8_L29, SubBytesIns_Inst_Sbox_8_L28,
         SubBytesIns_Inst_Sbox_8_L27, SubBytesIns_Inst_Sbox_8_L26,
         SubBytesIns_Inst_Sbox_8_L25, SubBytesIns_Inst_Sbox_8_L24,
         SubBytesIns_Inst_Sbox_8_L23, SubBytesIns_Inst_Sbox_8_L22,
         SubBytesIns_Inst_Sbox_8_L21, SubBytesIns_Inst_Sbox_8_L20,
         SubBytesIns_Inst_Sbox_8_L19, SubBytesIns_Inst_Sbox_8_L18,
         SubBytesIns_Inst_Sbox_8_L17, SubBytesIns_Inst_Sbox_8_L16,
         SubBytesIns_Inst_Sbox_8_L15, SubBytesIns_Inst_Sbox_8_L14,
         SubBytesIns_Inst_Sbox_8_L13, SubBytesIns_Inst_Sbox_8_L12,
         SubBytesIns_Inst_Sbox_8_L11, SubBytesIns_Inst_Sbox_8_L10,
         SubBytesIns_Inst_Sbox_8_L9, SubBytesIns_Inst_Sbox_8_L8,
         SubBytesIns_Inst_Sbox_8_L7, SubBytesIns_Inst_Sbox_8_L6,
         SubBytesIns_Inst_Sbox_8_L5, SubBytesIns_Inst_Sbox_8_L4,
         SubBytesIns_Inst_Sbox_8_L3, SubBytesIns_Inst_Sbox_8_L2,
         SubBytesIns_Inst_Sbox_8_L1, SubBytesIns_Inst_Sbox_8_L0,
         SubBytesIns_Inst_Sbox_8_M63, SubBytesIns_Inst_Sbox_8_M62,
         SubBytesIns_Inst_Sbox_8_M61, SubBytesIns_Inst_Sbox_8_M60,
         SubBytesIns_Inst_Sbox_8_M59, SubBytesIns_Inst_Sbox_8_M58,
         SubBytesIns_Inst_Sbox_8_M57, SubBytesIns_Inst_Sbox_8_M56,
         SubBytesIns_Inst_Sbox_8_M55, SubBytesIns_Inst_Sbox_8_M54,
         SubBytesIns_Inst_Sbox_8_M53, SubBytesIns_Inst_Sbox_8_M52,
         SubBytesIns_Inst_Sbox_8_M51, SubBytesIns_Inst_Sbox_8_M50,
         SubBytesIns_Inst_Sbox_8_M49, SubBytesIns_Inst_Sbox_8_M48,
         SubBytesIns_Inst_Sbox_8_M47, SubBytesIns_Inst_Sbox_8_M46,
         SubBytesIns_Inst_Sbox_8_M45, SubBytesIns_Inst_Sbox_8_M44,
         SubBytesIns_Inst_Sbox_8_M43, SubBytesIns_Inst_Sbox_8_M42,
         SubBytesIns_Inst_Sbox_8_M41, SubBytesIns_Inst_Sbox_8_M40,
         SubBytesIns_Inst_Sbox_8_M39, SubBytesIns_Inst_Sbox_8_M38,
         SubBytesIns_Inst_Sbox_8_M37, SubBytesIns_Inst_Sbox_8_M36,
         SubBytesIns_Inst_Sbox_8_M35, SubBytesIns_Inst_Sbox_8_M34,
         SubBytesIns_Inst_Sbox_8_M33, SubBytesIns_Inst_Sbox_8_M32,
         SubBytesIns_Inst_Sbox_8_M31, SubBytesIns_Inst_Sbox_8_M30,
         SubBytesIns_Inst_Sbox_8_M29, SubBytesIns_Inst_Sbox_8_M28,
         SubBytesIns_Inst_Sbox_8_M27, SubBytesIns_Inst_Sbox_8_M26,
         SubBytesIns_Inst_Sbox_8_M25, SubBytesIns_Inst_Sbox_8_M24,
         SubBytesIns_Inst_Sbox_8_M23, SubBytesIns_Inst_Sbox_8_M22,
         SubBytesIns_Inst_Sbox_8_M21, SubBytesIns_Inst_Sbox_8_M20,
         SubBytesIns_Inst_Sbox_8_M19, SubBytesIns_Inst_Sbox_8_M18,
         SubBytesIns_Inst_Sbox_8_M17, SubBytesIns_Inst_Sbox_8_M16,
         SubBytesIns_Inst_Sbox_8_M15, SubBytesIns_Inst_Sbox_8_M14,
         SubBytesIns_Inst_Sbox_8_M13, SubBytesIns_Inst_Sbox_8_M12,
         SubBytesIns_Inst_Sbox_8_M11, SubBytesIns_Inst_Sbox_8_M10,
         SubBytesIns_Inst_Sbox_8_M9, SubBytesIns_Inst_Sbox_8_M8,
         SubBytesIns_Inst_Sbox_8_M7, SubBytesIns_Inst_Sbox_8_M6,
         SubBytesIns_Inst_Sbox_8_M5, SubBytesIns_Inst_Sbox_8_M4,
         SubBytesIns_Inst_Sbox_8_M3, SubBytesIns_Inst_Sbox_8_M2,
         SubBytesIns_Inst_Sbox_8_M1, SubBytesIns_Inst_Sbox_8_T27,
         SubBytesIns_Inst_Sbox_8_T26, SubBytesIns_Inst_Sbox_8_T25,
         SubBytesIns_Inst_Sbox_8_T24, SubBytesIns_Inst_Sbox_8_T23,
         SubBytesIns_Inst_Sbox_8_T22, SubBytesIns_Inst_Sbox_8_T21,
         SubBytesIns_Inst_Sbox_8_T20, SubBytesIns_Inst_Sbox_8_T19,
         SubBytesIns_Inst_Sbox_8_T18, SubBytesIns_Inst_Sbox_8_T17,
         SubBytesIns_Inst_Sbox_8_T16, SubBytesIns_Inst_Sbox_8_T15,
         SubBytesIns_Inst_Sbox_8_T14, SubBytesIns_Inst_Sbox_8_T13,
         SubBytesIns_Inst_Sbox_8_T12, SubBytesIns_Inst_Sbox_8_T11,
         SubBytesIns_Inst_Sbox_8_T10, SubBytesIns_Inst_Sbox_8_T9,
         SubBytesIns_Inst_Sbox_8_T8, SubBytesIns_Inst_Sbox_8_T7,
         SubBytesIns_Inst_Sbox_8_T6, SubBytesIns_Inst_Sbox_8_T5,
         SubBytesIns_Inst_Sbox_8_T4, SubBytesIns_Inst_Sbox_8_T3,
         SubBytesIns_Inst_Sbox_8_T2, SubBytesIns_Inst_Sbox_8_T1,
         SubBytesIns_Inst_Sbox_9_L29, SubBytesIns_Inst_Sbox_9_L28,
         SubBytesIns_Inst_Sbox_9_L27, SubBytesIns_Inst_Sbox_9_L26,
         SubBytesIns_Inst_Sbox_9_L25, SubBytesIns_Inst_Sbox_9_L24,
         SubBytesIns_Inst_Sbox_9_L23, SubBytesIns_Inst_Sbox_9_L22,
         SubBytesIns_Inst_Sbox_9_L21, SubBytesIns_Inst_Sbox_9_L20,
         SubBytesIns_Inst_Sbox_9_L19, SubBytesIns_Inst_Sbox_9_L18,
         SubBytesIns_Inst_Sbox_9_L17, SubBytesIns_Inst_Sbox_9_L16,
         SubBytesIns_Inst_Sbox_9_L15, SubBytesIns_Inst_Sbox_9_L14,
         SubBytesIns_Inst_Sbox_9_L13, SubBytesIns_Inst_Sbox_9_L12,
         SubBytesIns_Inst_Sbox_9_L11, SubBytesIns_Inst_Sbox_9_L10,
         SubBytesIns_Inst_Sbox_9_L9, SubBytesIns_Inst_Sbox_9_L8,
         SubBytesIns_Inst_Sbox_9_L7, SubBytesIns_Inst_Sbox_9_L6,
         SubBytesIns_Inst_Sbox_9_L5, SubBytesIns_Inst_Sbox_9_L4,
         SubBytesIns_Inst_Sbox_9_L3, SubBytesIns_Inst_Sbox_9_L2,
         SubBytesIns_Inst_Sbox_9_L1, SubBytesIns_Inst_Sbox_9_L0,
         SubBytesIns_Inst_Sbox_9_M63, SubBytesIns_Inst_Sbox_9_M62,
         SubBytesIns_Inst_Sbox_9_M61, SubBytesIns_Inst_Sbox_9_M60,
         SubBytesIns_Inst_Sbox_9_M59, SubBytesIns_Inst_Sbox_9_M58,
         SubBytesIns_Inst_Sbox_9_M57, SubBytesIns_Inst_Sbox_9_M56,
         SubBytesIns_Inst_Sbox_9_M55, SubBytesIns_Inst_Sbox_9_M54,
         SubBytesIns_Inst_Sbox_9_M53, SubBytesIns_Inst_Sbox_9_M52,
         SubBytesIns_Inst_Sbox_9_M51, SubBytesIns_Inst_Sbox_9_M50,
         SubBytesIns_Inst_Sbox_9_M49, SubBytesIns_Inst_Sbox_9_M48,
         SubBytesIns_Inst_Sbox_9_M47, SubBytesIns_Inst_Sbox_9_M46,
         SubBytesIns_Inst_Sbox_9_M45, SubBytesIns_Inst_Sbox_9_M44,
         SubBytesIns_Inst_Sbox_9_M43, SubBytesIns_Inst_Sbox_9_M42,
         SubBytesIns_Inst_Sbox_9_M41, SubBytesIns_Inst_Sbox_9_M40,
         SubBytesIns_Inst_Sbox_9_M39, SubBytesIns_Inst_Sbox_9_M38,
         SubBytesIns_Inst_Sbox_9_M37, SubBytesIns_Inst_Sbox_9_M36,
         SubBytesIns_Inst_Sbox_9_M35, SubBytesIns_Inst_Sbox_9_M34,
         SubBytesIns_Inst_Sbox_9_M33, SubBytesIns_Inst_Sbox_9_M32,
         SubBytesIns_Inst_Sbox_9_M31, SubBytesIns_Inst_Sbox_9_M30,
         SubBytesIns_Inst_Sbox_9_M29, SubBytesIns_Inst_Sbox_9_M28,
         SubBytesIns_Inst_Sbox_9_M27, SubBytesIns_Inst_Sbox_9_M26,
         SubBytesIns_Inst_Sbox_9_M25, SubBytesIns_Inst_Sbox_9_M24,
         SubBytesIns_Inst_Sbox_9_M23, SubBytesIns_Inst_Sbox_9_M22,
         SubBytesIns_Inst_Sbox_9_M21, SubBytesIns_Inst_Sbox_9_M20,
         SubBytesIns_Inst_Sbox_9_M19, SubBytesIns_Inst_Sbox_9_M18,
         SubBytesIns_Inst_Sbox_9_M17, SubBytesIns_Inst_Sbox_9_M16,
         SubBytesIns_Inst_Sbox_9_M15, SubBytesIns_Inst_Sbox_9_M14,
         SubBytesIns_Inst_Sbox_9_M13, SubBytesIns_Inst_Sbox_9_M12,
         SubBytesIns_Inst_Sbox_9_M11, SubBytesIns_Inst_Sbox_9_M10,
         SubBytesIns_Inst_Sbox_9_M9, SubBytesIns_Inst_Sbox_9_M8,
         SubBytesIns_Inst_Sbox_9_M7, SubBytesIns_Inst_Sbox_9_M6,
         SubBytesIns_Inst_Sbox_9_M5, SubBytesIns_Inst_Sbox_9_M4,
         SubBytesIns_Inst_Sbox_9_M3, SubBytesIns_Inst_Sbox_9_M2,
         SubBytesIns_Inst_Sbox_9_M1, SubBytesIns_Inst_Sbox_9_T27,
         SubBytesIns_Inst_Sbox_9_T26, SubBytesIns_Inst_Sbox_9_T25,
         SubBytesIns_Inst_Sbox_9_T24, SubBytesIns_Inst_Sbox_9_T23,
         SubBytesIns_Inst_Sbox_9_T22, SubBytesIns_Inst_Sbox_9_T21,
         SubBytesIns_Inst_Sbox_9_T20, SubBytesIns_Inst_Sbox_9_T19,
         SubBytesIns_Inst_Sbox_9_T18, SubBytesIns_Inst_Sbox_9_T17,
         SubBytesIns_Inst_Sbox_9_T16, SubBytesIns_Inst_Sbox_9_T15,
         SubBytesIns_Inst_Sbox_9_T14, SubBytesIns_Inst_Sbox_9_T13,
         SubBytesIns_Inst_Sbox_9_T12, SubBytesIns_Inst_Sbox_9_T11,
         SubBytesIns_Inst_Sbox_9_T10, SubBytesIns_Inst_Sbox_9_T9,
         SubBytesIns_Inst_Sbox_9_T8, SubBytesIns_Inst_Sbox_9_T7,
         SubBytesIns_Inst_Sbox_9_T6, SubBytesIns_Inst_Sbox_9_T5,
         SubBytesIns_Inst_Sbox_9_T4, SubBytesIns_Inst_Sbox_9_T3,
         SubBytesIns_Inst_Sbox_9_T2, SubBytesIns_Inst_Sbox_9_T1,
         SubBytesIns_Inst_Sbox_10_L29, SubBytesIns_Inst_Sbox_10_L28,
         SubBytesIns_Inst_Sbox_10_L27, SubBytesIns_Inst_Sbox_10_L26,
         SubBytesIns_Inst_Sbox_10_L25, SubBytesIns_Inst_Sbox_10_L24,
         SubBytesIns_Inst_Sbox_10_L23, SubBytesIns_Inst_Sbox_10_L22,
         SubBytesIns_Inst_Sbox_10_L21, SubBytesIns_Inst_Sbox_10_L20,
         SubBytesIns_Inst_Sbox_10_L19, SubBytesIns_Inst_Sbox_10_L18,
         SubBytesIns_Inst_Sbox_10_L17, SubBytesIns_Inst_Sbox_10_L16,
         SubBytesIns_Inst_Sbox_10_L15, SubBytesIns_Inst_Sbox_10_L14,
         SubBytesIns_Inst_Sbox_10_L13, SubBytesIns_Inst_Sbox_10_L12,
         SubBytesIns_Inst_Sbox_10_L11, SubBytesIns_Inst_Sbox_10_L10,
         SubBytesIns_Inst_Sbox_10_L9, SubBytesIns_Inst_Sbox_10_L8,
         SubBytesIns_Inst_Sbox_10_L7, SubBytesIns_Inst_Sbox_10_L6,
         SubBytesIns_Inst_Sbox_10_L5, SubBytesIns_Inst_Sbox_10_L4,
         SubBytesIns_Inst_Sbox_10_L3, SubBytesIns_Inst_Sbox_10_L2,
         SubBytesIns_Inst_Sbox_10_L1, SubBytesIns_Inst_Sbox_10_L0,
         SubBytesIns_Inst_Sbox_10_M63, SubBytesIns_Inst_Sbox_10_M62,
         SubBytesIns_Inst_Sbox_10_M61, SubBytesIns_Inst_Sbox_10_M60,
         SubBytesIns_Inst_Sbox_10_M59, SubBytesIns_Inst_Sbox_10_M58,
         SubBytesIns_Inst_Sbox_10_M57, SubBytesIns_Inst_Sbox_10_M56,
         SubBytesIns_Inst_Sbox_10_M55, SubBytesIns_Inst_Sbox_10_M54,
         SubBytesIns_Inst_Sbox_10_M53, SubBytesIns_Inst_Sbox_10_M52,
         SubBytesIns_Inst_Sbox_10_M51, SubBytesIns_Inst_Sbox_10_M50,
         SubBytesIns_Inst_Sbox_10_M49, SubBytesIns_Inst_Sbox_10_M48,
         SubBytesIns_Inst_Sbox_10_M47, SubBytesIns_Inst_Sbox_10_M46,
         SubBytesIns_Inst_Sbox_10_M45, SubBytesIns_Inst_Sbox_10_M44,
         SubBytesIns_Inst_Sbox_10_M43, SubBytesIns_Inst_Sbox_10_M42,
         SubBytesIns_Inst_Sbox_10_M41, SubBytesIns_Inst_Sbox_10_M40,
         SubBytesIns_Inst_Sbox_10_M39, SubBytesIns_Inst_Sbox_10_M38,
         SubBytesIns_Inst_Sbox_10_M37, SubBytesIns_Inst_Sbox_10_M36,
         SubBytesIns_Inst_Sbox_10_M35, SubBytesIns_Inst_Sbox_10_M34,
         SubBytesIns_Inst_Sbox_10_M33, SubBytesIns_Inst_Sbox_10_M32,
         SubBytesIns_Inst_Sbox_10_M31, SubBytesIns_Inst_Sbox_10_M30,
         SubBytesIns_Inst_Sbox_10_M29, SubBytesIns_Inst_Sbox_10_M28,
         SubBytesIns_Inst_Sbox_10_M27, SubBytesIns_Inst_Sbox_10_M26,
         SubBytesIns_Inst_Sbox_10_M25, SubBytesIns_Inst_Sbox_10_M24,
         SubBytesIns_Inst_Sbox_10_M23, SubBytesIns_Inst_Sbox_10_M22,
         SubBytesIns_Inst_Sbox_10_M21, SubBytesIns_Inst_Sbox_10_M20,
         SubBytesIns_Inst_Sbox_10_M19, SubBytesIns_Inst_Sbox_10_M18,
         SubBytesIns_Inst_Sbox_10_M17, SubBytesIns_Inst_Sbox_10_M16,
         SubBytesIns_Inst_Sbox_10_M15, SubBytesIns_Inst_Sbox_10_M14,
         SubBytesIns_Inst_Sbox_10_M13, SubBytesIns_Inst_Sbox_10_M12,
         SubBytesIns_Inst_Sbox_10_M11, SubBytesIns_Inst_Sbox_10_M10,
         SubBytesIns_Inst_Sbox_10_M9, SubBytesIns_Inst_Sbox_10_M8,
         SubBytesIns_Inst_Sbox_10_M7, SubBytesIns_Inst_Sbox_10_M6,
         SubBytesIns_Inst_Sbox_10_M5, SubBytesIns_Inst_Sbox_10_M4,
         SubBytesIns_Inst_Sbox_10_M3, SubBytesIns_Inst_Sbox_10_M2,
         SubBytesIns_Inst_Sbox_10_M1, SubBytesIns_Inst_Sbox_10_T27,
         SubBytesIns_Inst_Sbox_10_T26, SubBytesIns_Inst_Sbox_10_T25,
         SubBytesIns_Inst_Sbox_10_T24, SubBytesIns_Inst_Sbox_10_T23,
         SubBytesIns_Inst_Sbox_10_T22, SubBytesIns_Inst_Sbox_10_T21,
         SubBytesIns_Inst_Sbox_10_T20, SubBytesIns_Inst_Sbox_10_T19,
         SubBytesIns_Inst_Sbox_10_T18, SubBytesIns_Inst_Sbox_10_T17,
         SubBytesIns_Inst_Sbox_10_T16, SubBytesIns_Inst_Sbox_10_T15,
         SubBytesIns_Inst_Sbox_10_T14, SubBytesIns_Inst_Sbox_10_T13,
         SubBytesIns_Inst_Sbox_10_T12, SubBytesIns_Inst_Sbox_10_T11,
         SubBytesIns_Inst_Sbox_10_T10, SubBytesIns_Inst_Sbox_10_T9,
         SubBytesIns_Inst_Sbox_10_T8, SubBytesIns_Inst_Sbox_10_T7,
         SubBytesIns_Inst_Sbox_10_T6, SubBytesIns_Inst_Sbox_10_T5,
         SubBytesIns_Inst_Sbox_10_T4, SubBytesIns_Inst_Sbox_10_T3,
         SubBytesIns_Inst_Sbox_10_T2, SubBytesIns_Inst_Sbox_10_T1,
         SubBytesIns_Inst_Sbox_11_L29, SubBytesIns_Inst_Sbox_11_L28,
         SubBytesIns_Inst_Sbox_11_L27, SubBytesIns_Inst_Sbox_11_L26,
         SubBytesIns_Inst_Sbox_11_L25, SubBytesIns_Inst_Sbox_11_L24,
         SubBytesIns_Inst_Sbox_11_L23, SubBytesIns_Inst_Sbox_11_L22,
         SubBytesIns_Inst_Sbox_11_L21, SubBytesIns_Inst_Sbox_11_L20,
         SubBytesIns_Inst_Sbox_11_L19, SubBytesIns_Inst_Sbox_11_L18,
         SubBytesIns_Inst_Sbox_11_L17, SubBytesIns_Inst_Sbox_11_L16,
         SubBytesIns_Inst_Sbox_11_L15, SubBytesIns_Inst_Sbox_11_L14,
         SubBytesIns_Inst_Sbox_11_L13, SubBytesIns_Inst_Sbox_11_L12,
         SubBytesIns_Inst_Sbox_11_L11, SubBytesIns_Inst_Sbox_11_L10,
         SubBytesIns_Inst_Sbox_11_L9, SubBytesIns_Inst_Sbox_11_L8,
         SubBytesIns_Inst_Sbox_11_L7, SubBytesIns_Inst_Sbox_11_L6,
         SubBytesIns_Inst_Sbox_11_L5, SubBytesIns_Inst_Sbox_11_L4,
         SubBytesIns_Inst_Sbox_11_L3, SubBytesIns_Inst_Sbox_11_L2,
         SubBytesIns_Inst_Sbox_11_L1, SubBytesIns_Inst_Sbox_11_L0,
         SubBytesIns_Inst_Sbox_11_M63, SubBytesIns_Inst_Sbox_11_M62,
         SubBytesIns_Inst_Sbox_11_M61, SubBytesIns_Inst_Sbox_11_M60,
         SubBytesIns_Inst_Sbox_11_M59, SubBytesIns_Inst_Sbox_11_M58,
         SubBytesIns_Inst_Sbox_11_M57, SubBytesIns_Inst_Sbox_11_M56,
         SubBytesIns_Inst_Sbox_11_M55, SubBytesIns_Inst_Sbox_11_M54,
         SubBytesIns_Inst_Sbox_11_M53, SubBytesIns_Inst_Sbox_11_M52,
         SubBytesIns_Inst_Sbox_11_M51, SubBytesIns_Inst_Sbox_11_M50,
         SubBytesIns_Inst_Sbox_11_M49, SubBytesIns_Inst_Sbox_11_M48,
         SubBytesIns_Inst_Sbox_11_M47, SubBytesIns_Inst_Sbox_11_M46,
         SubBytesIns_Inst_Sbox_11_M45, SubBytesIns_Inst_Sbox_11_M44,
         SubBytesIns_Inst_Sbox_11_M43, SubBytesIns_Inst_Sbox_11_M42,
         SubBytesIns_Inst_Sbox_11_M41, SubBytesIns_Inst_Sbox_11_M40,
         SubBytesIns_Inst_Sbox_11_M39, SubBytesIns_Inst_Sbox_11_M38,
         SubBytesIns_Inst_Sbox_11_M37, SubBytesIns_Inst_Sbox_11_M36,
         SubBytesIns_Inst_Sbox_11_M35, SubBytesIns_Inst_Sbox_11_M34,
         SubBytesIns_Inst_Sbox_11_M33, SubBytesIns_Inst_Sbox_11_M32,
         SubBytesIns_Inst_Sbox_11_M31, SubBytesIns_Inst_Sbox_11_M30,
         SubBytesIns_Inst_Sbox_11_M29, SubBytesIns_Inst_Sbox_11_M28,
         SubBytesIns_Inst_Sbox_11_M27, SubBytesIns_Inst_Sbox_11_M26,
         SubBytesIns_Inst_Sbox_11_M25, SubBytesIns_Inst_Sbox_11_M24,
         SubBytesIns_Inst_Sbox_11_M23, SubBytesIns_Inst_Sbox_11_M22,
         SubBytesIns_Inst_Sbox_11_M21, SubBytesIns_Inst_Sbox_11_M20,
         SubBytesIns_Inst_Sbox_11_M19, SubBytesIns_Inst_Sbox_11_M18,
         SubBytesIns_Inst_Sbox_11_M17, SubBytesIns_Inst_Sbox_11_M16,
         SubBytesIns_Inst_Sbox_11_M15, SubBytesIns_Inst_Sbox_11_M14,
         SubBytesIns_Inst_Sbox_11_M13, SubBytesIns_Inst_Sbox_11_M12,
         SubBytesIns_Inst_Sbox_11_M11, SubBytesIns_Inst_Sbox_11_M10,
         SubBytesIns_Inst_Sbox_11_M9, SubBytesIns_Inst_Sbox_11_M8,
         SubBytesIns_Inst_Sbox_11_M7, SubBytesIns_Inst_Sbox_11_M6,
         SubBytesIns_Inst_Sbox_11_M5, SubBytesIns_Inst_Sbox_11_M4,
         SubBytesIns_Inst_Sbox_11_M3, SubBytesIns_Inst_Sbox_11_M2,
         SubBytesIns_Inst_Sbox_11_M1, SubBytesIns_Inst_Sbox_11_T27,
         SubBytesIns_Inst_Sbox_11_T26, SubBytesIns_Inst_Sbox_11_T25,
         SubBytesIns_Inst_Sbox_11_T24, SubBytesIns_Inst_Sbox_11_T23,
         SubBytesIns_Inst_Sbox_11_T22, SubBytesIns_Inst_Sbox_11_T21,
         SubBytesIns_Inst_Sbox_11_T20, SubBytesIns_Inst_Sbox_11_T19,
         SubBytesIns_Inst_Sbox_11_T18, SubBytesIns_Inst_Sbox_11_T17,
         SubBytesIns_Inst_Sbox_11_T16, SubBytesIns_Inst_Sbox_11_T15,
         SubBytesIns_Inst_Sbox_11_T14, SubBytesIns_Inst_Sbox_11_T13,
         SubBytesIns_Inst_Sbox_11_T12, SubBytesIns_Inst_Sbox_11_T11,
         SubBytesIns_Inst_Sbox_11_T10, SubBytesIns_Inst_Sbox_11_T9,
         SubBytesIns_Inst_Sbox_11_T8, SubBytesIns_Inst_Sbox_11_T7,
         SubBytesIns_Inst_Sbox_11_T6, SubBytesIns_Inst_Sbox_11_T5,
         SubBytesIns_Inst_Sbox_11_T4, SubBytesIns_Inst_Sbox_11_T3,
         SubBytesIns_Inst_Sbox_11_T2, SubBytesIns_Inst_Sbox_11_T1,
         SubBytesIns_Inst_Sbox_12_L29, SubBytesIns_Inst_Sbox_12_L28,
         SubBytesIns_Inst_Sbox_12_L27, SubBytesIns_Inst_Sbox_12_L26,
         SubBytesIns_Inst_Sbox_12_L25, SubBytesIns_Inst_Sbox_12_L24,
         SubBytesIns_Inst_Sbox_12_L23, SubBytesIns_Inst_Sbox_12_L22,
         SubBytesIns_Inst_Sbox_12_L21, SubBytesIns_Inst_Sbox_12_L20,
         SubBytesIns_Inst_Sbox_12_L19, SubBytesIns_Inst_Sbox_12_L18,
         SubBytesIns_Inst_Sbox_12_L17, SubBytesIns_Inst_Sbox_12_L16,
         SubBytesIns_Inst_Sbox_12_L15, SubBytesIns_Inst_Sbox_12_L14,
         SubBytesIns_Inst_Sbox_12_L13, SubBytesIns_Inst_Sbox_12_L12,
         SubBytesIns_Inst_Sbox_12_L11, SubBytesIns_Inst_Sbox_12_L10,
         SubBytesIns_Inst_Sbox_12_L9, SubBytesIns_Inst_Sbox_12_L8,
         SubBytesIns_Inst_Sbox_12_L7, SubBytesIns_Inst_Sbox_12_L6,
         SubBytesIns_Inst_Sbox_12_L5, SubBytesIns_Inst_Sbox_12_L4,
         SubBytesIns_Inst_Sbox_12_L3, SubBytesIns_Inst_Sbox_12_L2,
         SubBytesIns_Inst_Sbox_12_L1, SubBytesIns_Inst_Sbox_12_L0,
         SubBytesIns_Inst_Sbox_12_M63, SubBytesIns_Inst_Sbox_12_M62,
         SubBytesIns_Inst_Sbox_12_M61, SubBytesIns_Inst_Sbox_12_M60,
         SubBytesIns_Inst_Sbox_12_M59, SubBytesIns_Inst_Sbox_12_M58,
         SubBytesIns_Inst_Sbox_12_M57, SubBytesIns_Inst_Sbox_12_M56,
         SubBytesIns_Inst_Sbox_12_M55, SubBytesIns_Inst_Sbox_12_M54,
         SubBytesIns_Inst_Sbox_12_M53, SubBytesIns_Inst_Sbox_12_M52,
         SubBytesIns_Inst_Sbox_12_M51, SubBytesIns_Inst_Sbox_12_M50,
         SubBytesIns_Inst_Sbox_12_M49, SubBytesIns_Inst_Sbox_12_M48,
         SubBytesIns_Inst_Sbox_12_M47, SubBytesIns_Inst_Sbox_12_M46,
         SubBytesIns_Inst_Sbox_12_M45, SubBytesIns_Inst_Sbox_12_M44,
         SubBytesIns_Inst_Sbox_12_M43, SubBytesIns_Inst_Sbox_12_M42,
         SubBytesIns_Inst_Sbox_12_M41, SubBytesIns_Inst_Sbox_12_M40,
         SubBytesIns_Inst_Sbox_12_M39, SubBytesIns_Inst_Sbox_12_M38,
         SubBytesIns_Inst_Sbox_12_M37, SubBytesIns_Inst_Sbox_12_M36,
         SubBytesIns_Inst_Sbox_12_M35, SubBytesIns_Inst_Sbox_12_M34,
         SubBytesIns_Inst_Sbox_12_M33, SubBytesIns_Inst_Sbox_12_M32,
         SubBytesIns_Inst_Sbox_12_M31, SubBytesIns_Inst_Sbox_12_M30,
         SubBytesIns_Inst_Sbox_12_M29, SubBytesIns_Inst_Sbox_12_M28,
         SubBytesIns_Inst_Sbox_12_M27, SubBytesIns_Inst_Sbox_12_M26,
         SubBytesIns_Inst_Sbox_12_M25, SubBytesIns_Inst_Sbox_12_M24,
         SubBytesIns_Inst_Sbox_12_M23, SubBytesIns_Inst_Sbox_12_M22,
         SubBytesIns_Inst_Sbox_12_M21, SubBytesIns_Inst_Sbox_12_M20,
         SubBytesIns_Inst_Sbox_12_M19, SubBytesIns_Inst_Sbox_12_M18,
         SubBytesIns_Inst_Sbox_12_M17, SubBytesIns_Inst_Sbox_12_M16,
         SubBytesIns_Inst_Sbox_12_M15, SubBytesIns_Inst_Sbox_12_M14,
         SubBytesIns_Inst_Sbox_12_M13, SubBytesIns_Inst_Sbox_12_M12,
         SubBytesIns_Inst_Sbox_12_M11, SubBytesIns_Inst_Sbox_12_M10,
         SubBytesIns_Inst_Sbox_12_M9, SubBytesIns_Inst_Sbox_12_M8,
         SubBytesIns_Inst_Sbox_12_M7, SubBytesIns_Inst_Sbox_12_M6,
         SubBytesIns_Inst_Sbox_12_M5, SubBytesIns_Inst_Sbox_12_M4,
         SubBytesIns_Inst_Sbox_12_M3, SubBytesIns_Inst_Sbox_12_M2,
         SubBytesIns_Inst_Sbox_12_M1, SubBytesIns_Inst_Sbox_12_T27,
         SubBytesIns_Inst_Sbox_12_T26, SubBytesIns_Inst_Sbox_12_T25,
         SubBytesIns_Inst_Sbox_12_T24, SubBytesIns_Inst_Sbox_12_T23,
         SubBytesIns_Inst_Sbox_12_T22, SubBytesIns_Inst_Sbox_12_T21,
         SubBytesIns_Inst_Sbox_12_T20, SubBytesIns_Inst_Sbox_12_T19,
         SubBytesIns_Inst_Sbox_12_T18, SubBytesIns_Inst_Sbox_12_T17,
         SubBytesIns_Inst_Sbox_12_T16, SubBytesIns_Inst_Sbox_12_T15,
         SubBytesIns_Inst_Sbox_12_T14, SubBytesIns_Inst_Sbox_12_T13,
         SubBytesIns_Inst_Sbox_12_T12, SubBytesIns_Inst_Sbox_12_T11,
         SubBytesIns_Inst_Sbox_12_T10, SubBytesIns_Inst_Sbox_12_T9,
         SubBytesIns_Inst_Sbox_12_T8, SubBytesIns_Inst_Sbox_12_T7,
         SubBytesIns_Inst_Sbox_12_T6, SubBytesIns_Inst_Sbox_12_T5,
         SubBytesIns_Inst_Sbox_12_T4, SubBytesIns_Inst_Sbox_12_T3,
         SubBytesIns_Inst_Sbox_12_T2, SubBytesIns_Inst_Sbox_12_T1,
         SubBytesIns_Inst_Sbox_13_L29, SubBytesIns_Inst_Sbox_13_L28,
         SubBytesIns_Inst_Sbox_13_L27, SubBytesIns_Inst_Sbox_13_L26,
         SubBytesIns_Inst_Sbox_13_L25, SubBytesIns_Inst_Sbox_13_L24,
         SubBytesIns_Inst_Sbox_13_L23, SubBytesIns_Inst_Sbox_13_L22,
         SubBytesIns_Inst_Sbox_13_L21, SubBytesIns_Inst_Sbox_13_L20,
         SubBytesIns_Inst_Sbox_13_L19, SubBytesIns_Inst_Sbox_13_L18,
         SubBytesIns_Inst_Sbox_13_L17, SubBytesIns_Inst_Sbox_13_L16,
         SubBytesIns_Inst_Sbox_13_L15, SubBytesIns_Inst_Sbox_13_L14,
         SubBytesIns_Inst_Sbox_13_L13, SubBytesIns_Inst_Sbox_13_L12,
         SubBytesIns_Inst_Sbox_13_L11, SubBytesIns_Inst_Sbox_13_L10,
         SubBytesIns_Inst_Sbox_13_L9, SubBytesIns_Inst_Sbox_13_L8,
         SubBytesIns_Inst_Sbox_13_L7, SubBytesIns_Inst_Sbox_13_L6,
         SubBytesIns_Inst_Sbox_13_L5, SubBytesIns_Inst_Sbox_13_L4,
         SubBytesIns_Inst_Sbox_13_L3, SubBytesIns_Inst_Sbox_13_L2,
         SubBytesIns_Inst_Sbox_13_L1, SubBytesIns_Inst_Sbox_13_L0,
         SubBytesIns_Inst_Sbox_13_M63, SubBytesIns_Inst_Sbox_13_M62,
         SubBytesIns_Inst_Sbox_13_M61, SubBytesIns_Inst_Sbox_13_M60,
         SubBytesIns_Inst_Sbox_13_M59, SubBytesIns_Inst_Sbox_13_M58,
         SubBytesIns_Inst_Sbox_13_M57, SubBytesIns_Inst_Sbox_13_M56,
         SubBytesIns_Inst_Sbox_13_M55, SubBytesIns_Inst_Sbox_13_M54,
         SubBytesIns_Inst_Sbox_13_M53, SubBytesIns_Inst_Sbox_13_M52,
         SubBytesIns_Inst_Sbox_13_M51, SubBytesIns_Inst_Sbox_13_M50,
         SubBytesIns_Inst_Sbox_13_M49, SubBytesIns_Inst_Sbox_13_M48,
         SubBytesIns_Inst_Sbox_13_M47, SubBytesIns_Inst_Sbox_13_M46,
         SubBytesIns_Inst_Sbox_13_M45, SubBytesIns_Inst_Sbox_13_M44,
         SubBytesIns_Inst_Sbox_13_M43, SubBytesIns_Inst_Sbox_13_M42,
         SubBytesIns_Inst_Sbox_13_M41, SubBytesIns_Inst_Sbox_13_M40,
         SubBytesIns_Inst_Sbox_13_M39, SubBytesIns_Inst_Sbox_13_M38,
         SubBytesIns_Inst_Sbox_13_M37, SubBytesIns_Inst_Sbox_13_M36,
         SubBytesIns_Inst_Sbox_13_M35, SubBytesIns_Inst_Sbox_13_M34,
         SubBytesIns_Inst_Sbox_13_M33, SubBytesIns_Inst_Sbox_13_M32,
         SubBytesIns_Inst_Sbox_13_M31, SubBytesIns_Inst_Sbox_13_M30,
         SubBytesIns_Inst_Sbox_13_M29, SubBytesIns_Inst_Sbox_13_M28,
         SubBytesIns_Inst_Sbox_13_M27, SubBytesIns_Inst_Sbox_13_M26,
         SubBytesIns_Inst_Sbox_13_M25, SubBytesIns_Inst_Sbox_13_M24,
         SubBytesIns_Inst_Sbox_13_M23, SubBytesIns_Inst_Sbox_13_M22,
         SubBytesIns_Inst_Sbox_13_M21, SubBytesIns_Inst_Sbox_13_M20,
         SubBytesIns_Inst_Sbox_13_M19, SubBytesIns_Inst_Sbox_13_M18,
         SubBytesIns_Inst_Sbox_13_M17, SubBytesIns_Inst_Sbox_13_M16,
         SubBytesIns_Inst_Sbox_13_M15, SubBytesIns_Inst_Sbox_13_M14,
         SubBytesIns_Inst_Sbox_13_M13, SubBytesIns_Inst_Sbox_13_M12,
         SubBytesIns_Inst_Sbox_13_M11, SubBytesIns_Inst_Sbox_13_M10,
         SubBytesIns_Inst_Sbox_13_M9, SubBytesIns_Inst_Sbox_13_M8,
         SubBytesIns_Inst_Sbox_13_M7, SubBytesIns_Inst_Sbox_13_M6,
         SubBytesIns_Inst_Sbox_13_M5, SubBytesIns_Inst_Sbox_13_M4,
         SubBytesIns_Inst_Sbox_13_M3, SubBytesIns_Inst_Sbox_13_M2,
         SubBytesIns_Inst_Sbox_13_M1, SubBytesIns_Inst_Sbox_13_T27,
         SubBytesIns_Inst_Sbox_13_T26, SubBytesIns_Inst_Sbox_13_T25,
         SubBytesIns_Inst_Sbox_13_T24, SubBytesIns_Inst_Sbox_13_T23,
         SubBytesIns_Inst_Sbox_13_T22, SubBytesIns_Inst_Sbox_13_T21,
         SubBytesIns_Inst_Sbox_13_T20, SubBytesIns_Inst_Sbox_13_T19,
         SubBytesIns_Inst_Sbox_13_T18, SubBytesIns_Inst_Sbox_13_T17,
         SubBytesIns_Inst_Sbox_13_T16, SubBytesIns_Inst_Sbox_13_T15,
         SubBytesIns_Inst_Sbox_13_T14, SubBytesIns_Inst_Sbox_13_T13,
         SubBytesIns_Inst_Sbox_13_T12, SubBytesIns_Inst_Sbox_13_T11,
         SubBytesIns_Inst_Sbox_13_T10, SubBytesIns_Inst_Sbox_13_T9,
         SubBytesIns_Inst_Sbox_13_T8, SubBytesIns_Inst_Sbox_13_T7,
         SubBytesIns_Inst_Sbox_13_T6, SubBytesIns_Inst_Sbox_13_T5,
         SubBytesIns_Inst_Sbox_13_T4, SubBytesIns_Inst_Sbox_13_T3,
         SubBytesIns_Inst_Sbox_13_T2, SubBytesIns_Inst_Sbox_13_T1,
         SubBytesIns_Inst_Sbox_14_L29, SubBytesIns_Inst_Sbox_14_L28,
         SubBytesIns_Inst_Sbox_14_L27, SubBytesIns_Inst_Sbox_14_L26,
         SubBytesIns_Inst_Sbox_14_L25, SubBytesIns_Inst_Sbox_14_L24,
         SubBytesIns_Inst_Sbox_14_L23, SubBytesIns_Inst_Sbox_14_L22,
         SubBytesIns_Inst_Sbox_14_L21, SubBytesIns_Inst_Sbox_14_L20,
         SubBytesIns_Inst_Sbox_14_L19, SubBytesIns_Inst_Sbox_14_L18,
         SubBytesIns_Inst_Sbox_14_L17, SubBytesIns_Inst_Sbox_14_L16,
         SubBytesIns_Inst_Sbox_14_L15, SubBytesIns_Inst_Sbox_14_L14,
         SubBytesIns_Inst_Sbox_14_L13, SubBytesIns_Inst_Sbox_14_L12,
         SubBytesIns_Inst_Sbox_14_L11, SubBytesIns_Inst_Sbox_14_L10,
         SubBytesIns_Inst_Sbox_14_L9, SubBytesIns_Inst_Sbox_14_L8,
         SubBytesIns_Inst_Sbox_14_L7, SubBytesIns_Inst_Sbox_14_L6,
         SubBytesIns_Inst_Sbox_14_L5, SubBytesIns_Inst_Sbox_14_L4,
         SubBytesIns_Inst_Sbox_14_L3, SubBytesIns_Inst_Sbox_14_L2,
         SubBytesIns_Inst_Sbox_14_L1, SubBytesIns_Inst_Sbox_14_L0,
         SubBytesIns_Inst_Sbox_14_M63, SubBytesIns_Inst_Sbox_14_M62,
         SubBytesIns_Inst_Sbox_14_M61, SubBytesIns_Inst_Sbox_14_M60,
         SubBytesIns_Inst_Sbox_14_M59, SubBytesIns_Inst_Sbox_14_M58,
         SubBytesIns_Inst_Sbox_14_M57, SubBytesIns_Inst_Sbox_14_M56,
         SubBytesIns_Inst_Sbox_14_M55, SubBytesIns_Inst_Sbox_14_M54,
         SubBytesIns_Inst_Sbox_14_M53, SubBytesIns_Inst_Sbox_14_M52,
         SubBytesIns_Inst_Sbox_14_M51, SubBytesIns_Inst_Sbox_14_M50,
         SubBytesIns_Inst_Sbox_14_M49, SubBytesIns_Inst_Sbox_14_M48,
         SubBytesIns_Inst_Sbox_14_M47, SubBytesIns_Inst_Sbox_14_M46,
         SubBytesIns_Inst_Sbox_14_M45, SubBytesIns_Inst_Sbox_14_M44,
         SubBytesIns_Inst_Sbox_14_M43, SubBytesIns_Inst_Sbox_14_M42,
         SubBytesIns_Inst_Sbox_14_M41, SubBytesIns_Inst_Sbox_14_M40,
         SubBytesIns_Inst_Sbox_14_M39, SubBytesIns_Inst_Sbox_14_M38,
         SubBytesIns_Inst_Sbox_14_M37, SubBytesIns_Inst_Sbox_14_M36,
         SubBytesIns_Inst_Sbox_14_M35, SubBytesIns_Inst_Sbox_14_M34,
         SubBytesIns_Inst_Sbox_14_M33, SubBytesIns_Inst_Sbox_14_M32,
         SubBytesIns_Inst_Sbox_14_M31, SubBytesIns_Inst_Sbox_14_M30,
         SubBytesIns_Inst_Sbox_14_M29, SubBytesIns_Inst_Sbox_14_M28,
         SubBytesIns_Inst_Sbox_14_M27, SubBytesIns_Inst_Sbox_14_M26,
         SubBytesIns_Inst_Sbox_14_M25, SubBytesIns_Inst_Sbox_14_M24,
         SubBytesIns_Inst_Sbox_14_M23, SubBytesIns_Inst_Sbox_14_M22,
         SubBytesIns_Inst_Sbox_14_M21, SubBytesIns_Inst_Sbox_14_M20,
         SubBytesIns_Inst_Sbox_14_M19, SubBytesIns_Inst_Sbox_14_M18,
         SubBytesIns_Inst_Sbox_14_M17, SubBytesIns_Inst_Sbox_14_M16,
         SubBytesIns_Inst_Sbox_14_M15, SubBytesIns_Inst_Sbox_14_M14,
         SubBytesIns_Inst_Sbox_14_M13, SubBytesIns_Inst_Sbox_14_M12,
         SubBytesIns_Inst_Sbox_14_M11, SubBytesIns_Inst_Sbox_14_M10,
         SubBytesIns_Inst_Sbox_14_M9, SubBytesIns_Inst_Sbox_14_M8,
         SubBytesIns_Inst_Sbox_14_M7, SubBytesIns_Inst_Sbox_14_M6,
         SubBytesIns_Inst_Sbox_14_M5, SubBytesIns_Inst_Sbox_14_M4,
         SubBytesIns_Inst_Sbox_14_M3, SubBytesIns_Inst_Sbox_14_M2,
         SubBytesIns_Inst_Sbox_14_M1, SubBytesIns_Inst_Sbox_14_T27,
         SubBytesIns_Inst_Sbox_14_T26, SubBytesIns_Inst_Sbox_14_T25,
         SubBytesIns_Inst_Sbox_14_T24, SubBytesIns_Inst_Sbox_14_T23,
         SubBytesIns_Inst_Sbox_14_T22, SubBytesIns_Inst_Sbox_14_T21,
         SubBytesIns_Inst_Sbox_14_T20, SubBytesIns_Inst_Sbox_14_T19,
         SubBytesIns_Inst_Sbox_14_T18, SubBytesIns_Inst_Sbox_14_T17,
         SubBytesIns_Inst_Sbox_14_T16, SubBytesIns_Inst_Sbox_14_T15,
         SubBytesIns_Inst_Sbox_14_T14, SubBytesIns_Inst_Sbox_14_T13,
         SubBytesIns_Inst_Sbox_14_T12, SubBytesIns_Inst_Sbox_14_T11,
         SubBytesIns_Inst_Sbox_14_T10, SubBytesIns_Inst_Sbox_14_T9,
         SubBytesIns_Inst_Sbox_14_T8, SubBytesIns_Inst_Sbox_14_T7,
         SubBytesIns_Inst_Sbox_14_T6, SubBytesIns_Inst_Sbox_14_T5,
         SubBytesIns_Inst_Sbox_14_T4, SubBytesIns_Inst_Sbox_14_T3,
         SubBytesIns_Inst_Sbox_14_T2, SubBytesIns_Inst_Sbox_14_T1,
         SubBytesIns_Inst_Sbox_15_L29, SubBytesIns_Inst_Sbox_15_L28,
         SubBytesIns_Inst_Sbox_15_L27, SubBytesIns_Inst_Sbox_15_L26,
         SubBytesIns_Inst_Sbox_15_L25, SubBytesIns_Inst_Sbox_15_L24,
         SubBytesIns_Inst_Sbox_15_L23, SubBytesIns_Inst_Sbox_15_L22,
         SubBytesIns_Inst_Sbox_15_L21, SubBytesIns_Inst_Sbox_15_L20,
         SubBytesIns_Inst_Sbox_15_L19, SubBytesIns_Inst_Sbox_15_L18,
         SubBytesIns_Inst_Sbox_15_L17, SubBytesIns_Inst_Sbox_15_L16,
         SubBytesIns_Inst_Sbox_15_L15, SubBytesIns_Inst_Sbox_15_L14,
         SubBytesIns_Inst_Sbox_15_L13, SubBytesIns_Inst_Sbox_15_L12,
         SubBytesIns_Inst_Sbox_15_L11, SubBytesIns_Inst_Sbox_15_L10,
         SubBytesIns_Inst_Sbox_15_L9, SubBytesIns_Inst_Sbox_15_L8,
         SubBytesIns_Inst_Sbox_15_L7, SubBytesIns_Inst_Sbox_15_L6,
         SubBytesIns_Inst_Sbox_15_L5, SubBytesIns_Inst_Sbox_15_L4,
         SubBytesIns_Inst_Sbox_15_L3, SubBytesIns_Inst_Sbox_15_L2,
         SubBytesIns_Inst_Sbox_15_L1, SubBytesIns_Inst_Sbox_15_L0,
         SubBytesIns_Inst_Sbox_15_M63, SubBytesIns_Inst_Sbox_15_M62,
         SubBytesIns_Inst_Sbox_15_M61, SubBytesIns_Inst_Sbox_15_M60,
         SubBytesIns_Inst_Sbox_15_M59, SubBytesIns_Inst_Sbox_15_M58,
         SubBytesIns_Inst_Sbox_15_M57, SubBytesIns_Inst_Sbox_15_M56,
         SubBytesIns_Inst_Sbox_15_M55, SubBytesIns_Inst_Sbox_15_M54,
         SubBytesIns_Inst_Sbox_15_M53, SubBytesIns_Inst_Sbox_15_M52,
         SubBytesIns_Inst_Sbox_15_M51, SubBytesIns_Inst_Sbox_15_M50,
         SubBytesIns_Inst_Sbox_15_M49, SubBytesIns_Inst_Sbox_15_M48,
         SubBytesIns_Inst_Sbox_15_M47, SubBytesIns_Inst_Sbox_15_M46,
         SubBytesIns_Inst_Sbox_15_M45, SubBytesIns_Inst_Sbox_15_M44,
         SubBytesIns_Inst_Sbox_15_M43, SubBytesIns_Inst_Sbox_15_M42,
         SubBytesIns_Inst_Sbox_15_M41, SubBytesIns_Inst_Sbox_15_M40,
         SubBytesIns_Inst_Sbox_15_M39, SubBytesIns_Inst_Sbox_15_M38,
         SubBytesIns_Inst_Sbox_15_M37, SubBytesIns_Inst_Sbox_15_M36,
         SubBytesIns_Inst_Sbox_15_M35, SubBytesIns_Inst_Sbox_15_M34,
         SubBytesIns_Inst_Sbox_15_M33, SubBytesIns_Inst_Sbox_15_M32,
         SubBytesIns_Inst_Sbox_15_M31, SubBytesIns_Inst_Sbox_15_M30,
         SubBytesIns_Inst_Sbox_15_M29, SubBytesIns_Inst_Sbox_15_M28,
         SubBytesIns_Inst_Sbox_15_M27, SubBytesIns_Inst_Sbox_15_M26,
         SubBytesIns_Inst_Sbox_15_M25, SubBytesIns_Inst_Sbox_15_M24,
         SubBytesIns_Inst_Sbox_15_M23, SubBytesIns_Inst_Sbox_15_M22,
         SubBytesIns_Inst_Sbox_15_M21, SubBytesIns_Inst_Sbox_15_M20,
         SubBytesIns_Inst_Sbox_15_M19, SubBytesIns_Inst_Sbox_15_M18,
         SubBytesIns_Inst_Sbox_15_M17, SubBytesIns_Inst_Sbox_15_M16,
         SubBytesIns_Inst_Sbox_15_M15, SubBytesIns_Inst_Sbox_15_M14,
         SubBytesIns_Inst_Sbox_15_M13, SubBytesIns_Inst_Sbox_15_M12,
         SubBytesIns_Inst_Sbox_15_M11, SubBytesIns_Inst_Sbox_15_M10,
         SubBytesIns_Inst_Sbox_15_M9, SubBytesIns_Inst_Sbox_15_M8,
         SubBytesIns_Inst_Sbox_15_M7, SubBytesIns_Inst_Sbox_15_M6,
         SubBytesIns_Inst_Sbox_15_M5, SubBytesIns_Inst_Sbox_15_M4,
         SubBytesIns_Inst_Sbox_15_M3, SubBytesIns_Inst_Sbox_15_M2,
         SubBytesIns_Inst_Sbox_15_M1, SubBytesIns_Inst_Sbox_15_T27,
         SubBytesIns_Inst_Sbox_15_T26, SubBytesIns_Inst_Sbox_15_T25,
         SubBytesIns_Inst_Sbox_15_T24, SubBytesIns_Inst_Sbox_15_T23,
         SubBytesIns_Inst_Sbox_15_T22, SubBytesIns_Inst_Sbox_15_T21,
         SubBytesIns_Inst_Sbox_15_T20, SubBytesIns_Inst_Sbox_15_T19,
         SubBytesIns_Inst_Sbox_15_T18, SubBytesIns_Inst_Sbox_15_T17,
         SubBytesIns_Inst_Sbox_15_T16, SubBytesIns_Inst_Sbox_15_T15,
         SubBytesIns_Inst_Sbox_15_T14, SubBytesIns_Inst_Sbox_15_T13,
         SubBytesIns_Inst_Sbox_15_T12, SubBytesIns_Inst_Sbox_15_T11,
         SubBytesIns_Inst_Sbox_15_T10, SubBytesIns_Inst_Sbox_15_T9,
         SubBytesIns_Inst_Sbox_15_T8, SubBytesIns_Inst_Sbox_15_T7,
         SubBytesIns_Inst_Sbox_15_T6, SubBytesIns_Inst_Sbox_15_T5,
         SubBytesIns_Inst_Sbox_15_T4, SubBytesIns_Inst_Sbox_15_T3,
         SubBytesIns_Inst_Sbox_15_T2, SubBytesIns_Inst_Sbox_15_T1,
         MixColumnsIns_MixOneColumnInst_0_n64,
         MixColumnsIns_MixOneColumnInst_0_n63,
         MixColumnsIns_MixOneColumnInst_0_n62,
         MixColumnsIns_MixOneColumnInst_0_n61,
         MixColumnsIns_MixOneColumnInst_0_n60,
         MixColumnsIns_MixOneColumnInst_0_n59,
         MixColumnsIns_MixOneColumnInst_0_n58,
         MixColumnsIns_MixOneColumnInst_0_n57,
         MixColumnsIns_MixOneColumnInst_0_n56,
         MixColumnsIns_MixOneColumnInst_0_n55,
         MixColumnsIns_MixOneColumnInst_0_n54,
         MixColumnsIns_MixOneColumnInst_0_n53,
         MixColumnsIns_MixOneColumnInst_0_n52,
         MixColumnsIns_MixOneColumnInst_0_n51,
         MixColumnsIns_MixOneColumnInst_0_n50,
         MixColumnsIns_MixOneColumnInst_0_n49,
         MixColumnsIns_MixOneColumnInst_0_n48,
         MixColumnsIns_MixOneColumnInst_0_n47,
         MixColumnsIns_MixOneColumnInst_0_n46,
         MixColumnsIns_MixOneColumnInst_0_n45,
         MixColumnsIns_MixOneColumnInst_0_n44,
         MixColumnsIns_MixOneColumnInst_0_n43,
         MixColumnsIns_MixOneColumnInst_0_n42,
         MixColumnsIns_MixOneColumnInst_0_n41,
         MixColumnsIns_MixOneColumnInst_0_n40,
         MixColumnsIns_MixOneColumnInst_0_n39,
         MixColumnsIns_MixOneColumnInst_0_n38,
         MixColumnsIns_MixOneColumnInst_0_n37,
         MixColumnsIns_MixOneColumnInst_0_n36,
         MixColumnsIns_MixOneColumnInst_0_n35,
         MixColumnsIns_MixOneColumnInst_0_n34,
         MixColumnsIns_MixOneColumnInst_0_n33,
         MixColumnsIns_MixOneColumnInst_0_n32,
         MixColumnsIns_MixOneColumnInst_0_n31,
         MixColumnsIns_MixOneColumnInst_0_n30,
         MixColumnsIns_MixOneColumnInst_0_n29,
         MixColumnsIns_MixOneColumnInst_0_n28,
         MixColumnsIns_MixOneColumnInst_0_n27,
         MixColumnsIns_MixOneColumnInst_0_n26,
         MixColumnsIns_MixOneColumnInst_0_n25,
         MixColumnsIns_MixOneColumnInst_0_n24,
         MixColumnsIns_MixOneColumnInst_0_n23,
         MixColumnsIns_MixOneColumnInst_0_n22,
         MixColumnsIns_MixOneColumnInst_0_n21,
         MixColumnsIns_MixOneColumnInst_0_n20,
         MixColumnsIns_MixOneColumnInst_0_n19,
         MixColumnsIns_MixOneColumnInst_0_n18,
         MixColumnsIns_MixOneColumnInst_0_n17,
         MixColumnsIns_MixOneColumnInst_0_n16,
         MixColumnsIns_MixOneColumnInst_0_n15,
         MixColumnsIns_MixOneColumnInst_0_n14,
         MixColumnsIns_MixOneColumnInst_0_n13,
         MixColumnsIns_MixOneColumnInst_0_n12,
         MixColumnsIns_MixOneColumnInst_0_n11,
         MixColumnsIns_MixOneColumnInst_0_n10,
         MixColumnsIns_MixOneColumnInst_0_n9,
         MixColumnsIns_MixOneColumnInst_0_n8,
         MixColumnsIns_MixOneColumnInst_0_n7,
         MixColumnsIns_MixOneColumnInst_0_n6,
         MixColumnsIns_MixOneColumnInst_0_n5,
         MixColumnsIns_MixOneColumnInst_0_n4,
         MixColumnsIns_MixOneColumnInst_0_n3,
         MixColumnsIns_MixOneColumnInst_0_n2,
         MixColumnsIns_MixOneColumnInst_0_n1,
         MixColumnsIns_MixOneColumnInst_1_n64,
         MixColumnsIns_MixOneColumnInst_1_n63,
         MixColumnsIns_MixOneColumnInst_1_n62,
         MixColumnsIns_MixOneColumnInst_1_n61,
         MixColumnsIns_MixOneColumnInst_1_n60,
         MixColumnsIns_MixOneColumnInst_1_n59,
         MixColumnsIns_MixOneColumnInst_1_n58,
         MixColumnsIns_MixOneColumnInst_1_n57,
         MixColumnsIns_MixOneColumnInst_1_n56,
         MixColumnsIns_MixOneColumnInst_1_n55,
         MixColumnsIns_MixOneColumnInst_1_n54,
         MixColumnsIns_MixOneColumnInst_1_n53,
         MixColumnsIns_MixOneColumnInst_1_n52,
         MixColumnsIns_MixOneColumnInst_1_n51,
         MixColumnsIns_MixOneColumnInst_1_n50,
         MixColumnsIns_MixOneColumnInst_1_n49,
         MixColumnsIns_MixOneColumnInst_1_n48,
         MixColumnsIns_MixOneColumnInst_1_n47,
         MixColumnsIns_MixOneColumnInst_1_n46,
         MixColumnsIns_MixOneColumnInst_1_n45,
         MixColumnsIns_MixOneColumnInst_1_n44,
         MixColumnsIns_MixOneColumnInst_1_n43,
         MixColumnsIns_MixOneColumnInst_1_n42,
         MixColumnsIns_MixOneColumnInst_1_n41,
         MixColumnsIns_MixOneColumnInst_1_n40,
         MixColumnsIns_MixOneColumnInst_1_n39,
         MixColumnsIns_MixOneColumnInst_1_n38,
         MixColumnsIns_MixOneColumnInst_1_n37,
         MixColumnsIns_MixOneColumnInst_1_n36,
         MixColumnsIns_MixOneColumnInst_1_n35,
         MixColumnsIns_MixOneColumnInst_1_n34,
         MixColumnsIns_MixOneColumnInst_1_n33,
         MixColumnsIns_MixOneColumnInst_1_n32,
         MixColumnsIns_MixOneColumnInst_1_n31,
         MixColumnsIns_MixOneColumnInst_1_n30,
         MixColumnsIns_MixOneColumnInst_1_n29,
         MixColumnsIns_MixOneColumnInst_1_n28,
         MixColumnsIns_MixOneColumnInst_1_n27,
         MixColumnsIns_MixOneColumnInst_1_n26,
         MixColumnsIns_MixOneColumnInst_1_n25,
         MixColumnsIns_MixOneColumnInst_1_n24,
         MixColumnsIns_MixOneColumnInst_1_n23,
         MixColumnsIns_MixOneColumnInst_1_n22,
         MixColumnsIns_MixOneColumnInst_1_n21,
         MixColumnsIns_MixOneColumnInst_1_n20,
         MixColumnsIns_MixOneColumnInst_1_n19,
         MixColumnsIns_MixOneColumnInst_1_n18,
         MixColumnsIns_MixOneColumnInst_1_n17,
         MixColumnsIns_MixOneColumnInst_1_n16,
         MixColumnsIns_MixOneColumnInst_1_n15,
         MixColumnsIns_MixOneColumnInst_1_n14,
         MixColumnsIns_MixOneColumnInst_1_n13,
         MixColumnsIns_MixOneColumnInst_1_n12,
         MixColumnsIns_MixOneColumnInst_1_n11,
         MixColumnsIns_MixOneColumnInst_1_n10,
         MixColumnsIns_MixOneColumnInst_1_n9,
         MixColumnsIns_MixOneColumnInst_1_n8,
         MixColumnsIns_MixOneColumnInst_1_n7,
         MixColumnsIns_MixOneColumnInst_1_n6,
         MixColumnsIns_MixOneColumnInst_1_n5,
         MixColumnsIns_MixOneColumnInst_1_n4,
         MixColumnsIns_MixOneColumnInst_1_n3,
         MixColumnsIns_MixOneColumnInst_1_n2,
         MixColumnsIns_MixOneColumnInst_1_n1,
         MixColumnsIns_MixOneColumnInst_2_n64,
         MixColumnsIns_MixOneColumnInst_2_n63,
         MixColumnsIns_MixOneColumnInst_2_n62,
         MixColumnsIns_MixOneColumnInst_2_n61,
         MixColumnsIns_MixOneColumnInst_2_n60,
         MixColumnsIns_MixOneColumnInst_2_n59,
         MixColumnsIns_MixOneColumnInst_2_n58,
         MixColumnsIns_MixOneColumnInst_2_n57,
         MixColumnsIns_MixOneColumnInst_2_n56,
         MixColumnsIns_MixOneColumnInst_2_n55,
         MixColumnsIns_MixOneColumnInst_2_n54,
         MixColumnsIns_MixOneColumnInst_2_n53,
         MixColumnsIns_MixOneColumnInst_2_n52,
         MixColumnsIns_MixOneColumnInst_2_n51,
         MixColumnsIns_MixOneColumnInst_2_n50,
         MixColumnsIns_MixOneColumnInst_2_n49,
         MixColumnsIns_MixOneColumnInst_2_n48,
         MixColumnsIns_MixOneColumnInst_2_n47,
         MixColumnsIns_MixOneColumnInst_2_n46,
         MixColumnsIns_MixOneColumnInst_2_n45,
         MixColumnsIns_MixOneColumnInst_2_n44,
         MixColumnsIns_MixOneColumnInst_2_n43,
         MixColumnsIns_MixOneColumnInst_2_n42,
         MixColumnsIns_MixOneColumnInst_2_n41,
         MixColumnsIns_MixOneColumnInst_2_n40,
         MixColumnsIns_MixOneColumnInst_2_n39,
         MixColumnsIns_MixOneColumnInst_2_n38,
         MixColumnsIns_MixOneColumnInst_2_n37,
         MixColumnsIns_MixOneColumnInst_2_n36,
         MixColumnsIns_MixOneColumnInst_2_n35,
         MixColumnsIns_MixOneColumnInst_2_n34,
         MixColumnsIns_MixOneColumnInst_2_n33,
         MixColumnsIns_MixOneColumnInst_2_n32,
         MixColumnsIns_MixOneColumnInst_2_n31,
         MixColumnsIns_MixOneColumnInst_2_n30,
         MixColumnsIns_MixOneColumnInst_2_n29,
         MixColumnsIns_MixOneColumnInst_2_n28,
         MixColumnsIns_MixOneColumnInst_2_n27,
         MixColumnsIns_MixOneColumnInst_2_n26,
         MixColumnsIns_MixOneColumnInst_2_n25,
         MixColumnsIns_MixOneColumnInst_2_n24,
         MixColumnsIns_MixOneColumnInst_2_n23,
         MixColumnsIns_MixOneColumnInst_2_n22,
         MixColumnsIns_MixOneColumnInst_2_n21,
         MixColumnsIns_MixOneColumnInst_2_n20,
         MixColumnsIns_MixOneColumnInst_2_n19,
         MixColumnsIns_MixOneColumnInst_2_n18,
         MixColumnsIns_MixOneColumnInst_2_n17,
         MixColumnsIns_MixOneColumnInst_2_n16,
         MixColumnsIns_MixOneColumnInst_2_n15,
         MixColumnsIns_MixOneColumnInst_2_n14,
         MixColumnsIns_MixOneColumnInst_2_n13,
         MixColumnsIns_MixOneColumnInst_2_n12,
         MixColumnsIns_MixOneColumnInst_2_n11,
         MixColumnsIns_MixOneColumnInst_2_n10,
         MixColumnsIns_MixOneColumnInst_2_n9,
         MixColumnsIns_MixOneColumnInst_2_n8,
         MixColumnsIns_MixOneColumnInst_2_n7,
         MixColumnsIns_MixOneColumnInst_2_n6,
         MixColumnsIns_MixOneColumnInst_2_n5,
         MixColumnsIns_MixOneColumnInst_2_n4,
         MixColumnsIns_MixOneColumnInst_2_n3,
         MixColumnsIns_MixOneColumnInst_2_n2,
         MixColumnsIns_MixOneColumnInst_2_n1,
         MixColumnsIns_MixOneColumnInst_3_n64,
         MixColumnsIns_MixOneColumnInst_3_n63,
         MixColumnsIns_MixOneColumnInst_3_n62,
         MixColumnsIns_MixOneColumnInst_3_n61,
         MixColumnsIns_MixOneColumnInst_3_n60,
         MixColumnsIns_MixOneColumnInst_3_n59,
         MixColumnsIns_MixOneColumnInst_3_n58,
         MixColumnsIns_MixOneColumnInst_3_n57,
         MixColumnsIns_MixOneColumnInst_3_n56,
         MixColumnsIns_MixOneColumnInst_3_n55,
         MixColumnsIns_MixOneColumnInst_3_n54,
         MixColumnsIns_MixOneColumnInst_3_n53,
         MixColumnsIns_MixOneColumnInst_3_n52,
         MixColumnsIns_MixOneColumnInst_3_n51,
         MixColumnsIns_MixOneColumnInst_3_n50,
         MixColumnsIns_MixOneColumnInst_3_n49,
         MixColumnsIns_MixOneColumnInst_3_n48,
         MixColumnsIns_MixOneColumnInst_3_n47,
         MixColumnsIns_MixOneColumnInst_3_n46,
         MixColumnsIns_MixOneColumnInst_3_n45,
         MixColumnsIns_MixOneColumnInst_3_n44,
         MixColumnsIns_MixOneColumnInst_3_n43,
         MixColumnsIns_MixOneColumnInst_3_n42,
         MixColumnsIns_MixOneColumnInst_3_n41,
         MixColumnsIns_MixOneColumnInst_3_n40,
         MixColumnsIns_MixOneColumnInst_3_n39,
         MixColumnsIns_MixOneColumnInst_3_n38,
         MixColumnsIns_MixOneColumnInst_3_n37,
         MixColumnsIns_MixOneColumnInst_3_n36,
         MixColumnsIns_MixOneColumnInst_3_n35,
         MixColumnsIns_MixOneColumnInst_3_n34,
         MixColumnsIns_MixOneColumnInst_3_n33,
         MixColumnsIns_MixOneColumnInst_3_n32,
         MixColumnsIns_MixOneColumnInst_3_n31,
         MixColumnsIns_MixOneColumnInst_3_n30,
         MixColumnsIns_MixOneColumnInst_3_n29,
         MixColumnsIns_MixOneColumnInst_3_n28,
         MixColumnsIns_MixOneColumnInst_3_n27,
         MixColumnsIns_MixOneColumnInst_3_n26,
         MixColumnsIns_MixOneColumnInst_3_n25,
         MixColumnsIns_MixOneColumnInst_3_n24,
         MixColumnsIns_MixOneColumnInst_3_n23,
         MixColumnsIns_MixOneColumnInst_3_n22,
         MixColumnsIns_MixOneColumnInst_3_n21,
         MixColumnsIns_MixOneColumnInst_3_n20,
         MixColumnsIns_MixOneColumnInst_3_n19,
         MixColumnsIns_MixOneColumnInst_3_n18,
         MixColumnsIns_MixOneColumnInst_3_n17,
         MixColumnsIns_MixOneColumnInst_3_n16,
         MixColumnsIns_MixOneColumnInst_3_n15,
         MixColumnsIns_MixOneColumnInst_3_n14,
         MixColumnsIns_MixOneColumnInst_3_n13,
         MixColumnsIns_MixOneColumnInst_3_n12,
         MixColumnsIns_MixOneColumnInst_3_n11,
         MixColumnsIns_MixOneColumnInst_3_n10,
         MixColumnsIns_MixOneColumnInst_3_n9,
         MixColumnsIns_MixOneColumnInst_3_n8,
         MixColumnsIns_MixOneColumnInst_3_n7,
         MixColumnsIns_MixOneColumnInst_3_n6,
         MixColumnsIns_MixOneColumnInst_3_n5,
         MixColumnsIns_MixOneColumnInst_3_n4,
         MixColumnsIns_MixOneColumnInst_3_n3,
         MixColumnsIns_MixOneColumnInst_3_n2,
         MixColumnsIns_MixOneColumnInst_3_n1, KeyReg_n10, KeyReg_n9, KeyReg_n8,
         KeyReg_n7, KeyReg_n6, KeyReg_Inst_ff_SDE_0_next_state,
         KeyReg_Inst_ff_SDE_0_MUX_inst_Y, KeyReg_Inst_ff_SDE_0_MUX_inst_X,
         KeyReg_Inst_ff_SDE_0_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_1_next_state, KeyReg_Inst_ff_SDE_1_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_1_MUX_inst_X,
         KeyReg_Inst_ff_SDE_1_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_2_next_state, KeyReg_Inst_ff_SDE_2_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_2_MUX_inst_X,
         KeyReg_Inst_ff_SDE_2_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_3_next_state, KeyReg_Inst_ff_SDE_3_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_3_MUX_inst_X,
         KeyReg_Inst_ff_SDE_3_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_4_next_state, KeyReg_Inst_ff_SDE_4_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_4_MUX_inst_X,
         KeyReg_Inst_ff_SDE_4_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_5_next_state, KeyReg_Inst_ff_SDE_5_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_5_MUX_inst_X,
         KeyReg_Inst_ff_SDE_5_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_6_next_state, KeyReg_Inst_ff_SDE_6_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_6_MUX_inst_X,
         KeyReg_Inst_ff_SDE_6_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_7_next_state, KeyReg_Inst_ff_SDE_7_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_7_MUX_inst_X,
         KeyReg_Inst_ff_SDE_7_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_8_next_state, KeyReg_Inst_ff_SDE_8_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_8_MUX_inst_X,
         KeyReg_Inst_ff_SDE_8_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_9_next_state, KeyReg_Inst_ff_SDE_9_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_9_MUX_inst_X,
         KeyReg_Inst_ff_SDE_9_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_10_next_state, KeyReg_Inst_ff_SDE_10_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_10_MUX_inst_X,
         KeyReg_Inst_ff_SDE_10_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_11_next_state, KeyReg_Inst_ff_SDE_11_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_11_MUX_inst_X,
         KeyReg_Inst_ff_SDE_11_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_12_next_state, KeyReg_Inst_ff_SDE_12_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_12_MUX_inst_X,
         KeyReg_Inst_ff_SDE_12_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_13_next_state, KeyReg_Inst_ff_SDE_13_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_13_MUX_inst_X,
         KeyReg_Inst_ff_SDE_13_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_14_next_state, KeyReg_Inst_ff_SDE_14_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_14_MUX_inst_X,
         KeyReg_Inst_ff_SDE_14_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_15_next_state, KeyReg_Inst_ff_SDE_15_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_15_MUX_inst_X,
         KeyReg_Inst_ff_SDE_15_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_16_next_state, KeyReg_Inst_ff_SDE_16_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_16_MUX_inst_X,
         KeyReg_Inst_ff_SDE_16_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_17_next_state, KeyReg_Inst_ff_SDE_17_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_17_MUX_inst_X,
         KeyReg_Inst_ff_SDE_17_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_18_next_state, KeyReg_Inst_ff_SDE_18_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_18_MUX_inst_X,
         KeyReg_Inst_ff_SDE_18_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_19_next_state, KeyReg_Inst_ff_SDE_19_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_19_MUX_inst_X,
         KeyReg_Inst_ff_SDE_19_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_20_next_state, KeyReg_Inst_ff_SDE_20_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_20_MUX_inst_X,
         KeyReg_Inst_ff_SDE_20_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_21_next_state, KeyReg_Inst_ff_SDE_21_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_21_MUX_inst_X,
         KeyReg_Inst_ff_SDE_21_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_22_next_state, KeyReg_Inst_ff_SDE_22_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_22_MUX_inst_X,
         KeyReg_Inst_ff_SDE_22_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_23_next_state, KeyReg_Inst_ff_SDE_23_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_23_MUX_inst_X,
         KeyReg_Inst_ff_SDE_23_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_24_next_state, KeyReg_Inst_ff_SDE_24_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_24_MUX_inst_X,
         KeyReg_Inst_ff_SDE_24_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_25_next_state, KeyReg_Inst_ff_SDE_25_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_25_MUX_inst_X,
         KeyReg_Inst_ff_SDE_25_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_26_next_state, KeyReg_Inst_ff_SDE_26_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_26_MUX_inst_X,
         KeyReg_Inst_ff_SDE_26_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_27_next_state, KeyReg_Inst_ff_SDE_27_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_27_MUX_inst_X,
         KeyReg_Inst_ff_SDE_27_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_28_next_state, KeyReg_Inst_ff_SDE_28_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_28_MUX_inst_X,
         KeyReg_Inst_ff_SDE_28_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_29_next_state, KeyReg_Inst_ff_SDE_29_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_29_MUX_inst_X,
         KeyReg_Inst_ff_SDE_29_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_30_next_state, KeyReg_Inst_ff_SDE_30_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_30_MUX_inst_X,
         KeyReg_Inst_ff_SDE_30_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_31_next_state, KeyReg_Inst_ff_SDE_31_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_31_MUX_inst_X,
         KeyReg_Inst_ff_SDE_31_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_32_next_state, KeyReg_Inst_ff_SDE_32_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_32_MUX_inst_X,
         KeyReg_Inst_ff_SDE_32_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_33_next_state, KeyReg_Inst_ff_SDE_33_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_33_MUX_inst_X,
         KeyReg_Inst_ff_SDE_33_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_34_next_state, KeyReg_Inst_ff_SDE_34_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_34_MUX_inst_X,
         KeyReg_Inst_ff_SDE_34_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_35_next_state, KeyReg_Inst_ff_SDE_35_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_35_MUX_inst_X,
         KeyReg_Inst_ff_SDE_35_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_36_next_state, KeyReg_Inst_ff_SDE_36_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_36_MUX_inst_X,
         KeyReg_Inst_ff_SDE_36_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_37_next_state, KeyReg_Inst_ff_SDE_37_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_37_MUX_inst_X,
         KeyReg_Inst_ff_SDE_37_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_38_next_state, KeyReg_Inst_ff_SDE_38_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_38_MUX_inst_X,
         KeyReg_Inst_ff_SDE_38_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_39_next_state, KeyReg_Inst_ff_SDE_39_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_39_MUX_inst_X,
         KeyReg_Inst_ff_SDE_39_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_40_next_state, KeyReg_Inst_ff_SDE_40_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_40_MUX_inst_X,
         KeyReg_Inst_ff_SDE_40_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_41_next_state, KeyReg_Inst_ff_SDE_41_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_41_MUX_inst_X,
         KeyReg_Inst_ff_SDE_41_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_42_next_state, KeyReg_Inst_ff_SDE_42_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_42_MUX_inst_X,
         KeyReg_Inst_ff_SDE_42_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_43_next_state, KeyReg_Inst_ff_SDE_43_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_43_MUX_inst_X,
         KeyReg_Inst_ff_SDE_43_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_44_next_state, KeyReg_Inst_ff_SDE_44_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_44_MUX_inst_X,
         KeyReg_Inst_ff_SDE_44_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_45_next_state, KeyReg_Inst_ff_SDE_45_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_45_MUX_inst_X,
         KeyReg_Inst_ff_SDE_45_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_46_next_state, KeyReg_Inst_ff_SDE_46_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_46_MUX_inst_X,
         KeyReg_Inst_ff_SDE_46_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_47_next_state, KeyReg_Inst_ff_SDE_47_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_47_MUX_inst_X,
         KeyReg_Inst_ff_SDE_47_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_48_next_state, KeyReg_Inst_ff_SDE_48_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_48_MUX_inst_X,
         KeyReg_Inst_ff_SDE_48_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_49_next_state, KeyReg_Inst_ff_SDE_49_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_49_MUX_inst_X,
         KeyReg_Inst_ff_SDE_49_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_50_next_state, KeyReg_Inst_ff_SDE_50_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_50_MUX_inst_X,
         KeyReg_Inst_ff_SDE_50_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_51_next_state, KeyReg_Inst_ff_SDE_51_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_51_MUX_inst_X,
         KeyReg_Inst_ff_SDE_51_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_52_next_state, KeyReg_Inst_ff_SDE_52_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_52_MUX_inst_X,
         KeyReg_Inst_ff_SDE_52_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_53_next_state, KeyReg_Inst_ff_SDE_53_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_53_MUX_inst_X,
         KeyReg_Inst_ff_SDE_53_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_54_next_state, KeyReg_Inst_ff_SDE_54_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_54_MUX_inst_X,
         KeyReg_Inst_ff_SDE_54_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_55_next_state, KeyReg_Inst_ff_SDE_55_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_55_MUX_inst_X,
         KeyReg_Inst_ff_SDE_55_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_56_next_state, KeyReg_Inst_ff_SDE_56_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_56_MUX_inst_X,
         KeyReg_Inst_ff_SDE_56_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_57_next_state, KeyReg_Inst_ff_SDE_57_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_57_MUX_inst_X,
         KeyReg_Inst_ff_SDE_57_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_58_next_state, KeyReg_Inst_ff_SDE_58_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_58_MUX_inst_X,
         KeyReg_Inst_ff_SDE_58_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_59_next_state, KeyReg_Inst_ff_SDE_59_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_59_MUX_inst_X,
         KeyReg_Inst_ff_SDE_59_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_60_next_state, KeyReg_Inst_ff_SDE_60_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_60_MUX_inst_X,
         KeyReg_Inst_ff_SDE_60_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_61_next_state, KeyReg_Inst_ff_SDE_61_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_61_MUX_inst_X,
         KeyReg_Inst_ff_SDE_61_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_62_next_state, KeyReg_Inst_ff_SDE_62_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_62_MUX_inst_X,
         KeyReg_Inst_ff_SDE_62_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_63_next_state, KeyReg_Inst_ff_SDE_63_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_63_MUX_inst_X,
         KeyReg_Inst_ff_SDE_63_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_64_next_state, KeyReg_Inst_ff_SDE_64_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_64_MUX_inst_X,
         KeyReg_Inst_ff_SDE_64_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_65_next_state, KeyReg_Inst_ff_SDE_65_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_65_MUX_inst_X,
         KeyReg_Inst_ff_SDE_65_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_66_next_state, KeyReg_Inst_ff_SDE_66_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_66_MUX_inst_X,
         KeyReg_Inst_ff_SDE_66_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_67_next_state, KeyReg_Inst_ff_SDE_67_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_67_MUX_inst_X,
         KeyReg_Inst_ff_SDE_67_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_68_next_state, KeyReg_Inst_ff_SDE_68_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_68_MUX_inst_X,
         KeyReg_Inst_ff_SDE_68_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_69_next_state, KeyReg_Inst_ff_SDE_69_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_69_MUX_inst_X,
         KeyReg_Inst_ff_SDE_69_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_70_next_state, KeyReg_Inst_ff_SDE_70_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_70_MUX_inst_X,
         KeyReg_Inst_ff_SDE_70_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_71_next_state, KeyReg_Inst_ff_SDE_71_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_71_MUX_inst_X,
         KeyReg_Inst_ff_SDE_71_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_72_next_state, KeyReg_Inst_ff_SDE_72_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_72_MUX_inst_X,
         KeyReg_Inst_ff_SDE_72_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_73_next_state, KeyReg_Inst_ff_SDE_73_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_73_MUX_inst_X,
         KeyReg_Inst_ff_SDE_73_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_74_next_state, KeyReg_Inst_ff_SDE_74_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_74_MUX_inst_X,
         KeyReg_Inst_ff_SDE_74_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_75_next_state, KeyReg_Inst_ff_SDE_75_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_75_MUX_inst_X,
         KeyReg_Inst_ff_SDE_75_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_76_next_state, KeyReg_Inst_ff_SDE_76_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_76_MUX_inst_X,
         KeyReg_Inst_ff_SDE_76_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_77_next_state, KeyReg_Inst_ff_SDE_77_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_77_MUX_inst_X,
         KeyReg_Inst_ff_SDE_77_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_78_next_state, KeyReg_Inst_ff_SDE_78_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_78_MUX_inst_X,
         KeyReg_Inst_ff_SDE_78_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_79_next_state, KeyReg_Inst_ff_SDE_79_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_79_MUX_inst_X,
         KeyReg_Inst_ff_SDE_79_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_80_next_state, KeyReg_Inst_ff_SDE_80_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_80_MUX_inst_X,
         KeyReg_Inst_ff_SDE_80_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_81_next_state, KeyReg_Inst_ff_SDE_81_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_81_MUX_inst_X,
         KeyReg_Inst_ff_SDE_81_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_82_next_state, KeyReg_Inst_ff_SDE_82_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_82_MUX_inst_X,
         KeyReg_Inst_ff_SDE_82_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_83_next_state, KeyReg_Inst_ff_SDE_83_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_83_MUX_inst_X,
         KeyReg_Inst_ff_SDE_83_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_84_next_state, KeyReg_Inst_ff_SDE_84_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_84_MUX_inst_X,
         KeyReg_Inst_ff_SDE_84_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_85_next_state, KeyReg_Inst_ff_SDE_85_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_85_MUX_inst_X,
         KeyReg_Inst_ff_SDE_85_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_86_next_state, KeyReg_Inst_ff_SDE_86_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_86_MUX_inst_X,
         KeyReg_Inst_ff_SDE_86_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_87_next_state, KeyReg_Inst_ff_SDE_87_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_87_MUX_inst_X,
         KeyReg_Inst_ff_SDE_87_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_88_next_state, KeyReg_Inst_ff_SDE_88_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_88_MUX_inst_X,
         KeyReg_Inst_ff_SDE_88_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_89_next_state, KeyReg_Inst_ff_SDE_89_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_89_MUX_inst_X,
         KeyReg_Inst_ff_SDE_89_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_90_next_state, KeyReg_Inst_ff_SDE_90_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_90_MUX_inst_X,
         KeyReg_Inst_ff_SDE_90_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_91_next_state, KeyReg_Inst_ff_SDE_91_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_91_MUX_inst_X,
         KeyReg_Inst_ff_SDE_91_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_92_next_state, KeyReg_Inst_ff_SDE_92_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_92_MUX_inst_X,
         KeyReg_Inst_ff_SDE_92_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_93_next_state, KeyReg_Inst_ff_SDE_93_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_93_MUX_inst_X,
         KeyReg_Inst_ff_SDE_93_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_94_next_state, KeyReg_Inst_ff_SDE_94_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_94_MUX_inst_X,
         KeyReg_Inst_ff_SDE_94_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_95_next_state, KeyReg_Inst_ff_SDE_95_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_95_MUX_inst_X,
         KeyReg_Inst_ff_SDE_95_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_96_next_state, KeyReg_Inst_ff_SDE_96_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_96_MUX_inst_X,
         KeyReg_Inst_ff_SDE_96_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_97_next_state, KeyReg_Inst_ff_SDE_97_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_97_MUX_inst_X,
         KeyReg_Inst_ff_SDE_97_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_98_next_state, KeyReg_Inst_ff_SDE_98_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_98_MUX_inst_X,
         KeyReg_Inst_ff_SDE_98_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_99_next_state, KeyReg_Inst_ff_SDE_99_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_99_MUX_inst_X,
         KeyReg_Inst_ff_SDE_99_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_100_next_state, KeyReg_Inst_ff_SDE_100_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_100_MUX_inst_X,
         KeyReg_Inst_ff_SDE_100_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_101_next_state, KeyReg_Inst_ff_SDE_101_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_101_MUX_inst_X,
         KeyReg_Inst_ff_SDE_101_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_102_next_state, KeyReg_Inst_ff_SDE_102_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_102_MUX_inst_X,
         KeyReg_Inst_ff_SDE_102_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_103_next_state, KeyReg_Inst_ff_SDE_103_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_103_MUX_inst_X,
         KeyReg_Inst_ff_SDE_103_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_104_next_state, KeyReg_Inst_ff_SDE_104_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_104_MUX_inst_X,
         KeyReg_Inst_ff_SDE_104_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_105_next_state, KeyReg_Inst_ff_SDE_105_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_105_MUX_inst_X,
         KeyReg_Inst_ff_SDE_105_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_106_next_state, KeyReg_Inst_ff_SDE_106_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_106_MUX_inst_X,
         KeyReg_Inst_ff_SDE_106_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_107_next_state, KeyReg_Inst_ff_SDE_107_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_107_MUX_inst_X,
         KeyReg_Inst_ff_SDE_107_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_108_next_state, KeyReg_Inst_ff_SDE_108_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_108_MUX_inst_X,
         KeyReg_Inst_ff_SDE_108_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_109_next_state, KeyReg_Inst_ff_SDE_109_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_109_MUX_inst_X,
         KeyReg_Inst_ff_SDE_109_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_110_next_state, KeyReg_Inst_ff_SDE_110_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_110_MUX_inst_X,
         KeyReg_Inst_ff_SDE_110_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_111_next_state, KeyReg_Inst_ff_SDE_111_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_111_MUX_inst_X,
         KeyReg_Inst_ff_SDE_111_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_112_next_state, KeyReg_Inst_ff_SDE_112_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_112_MUX_inst_X,
         KeyReg_Inst_ff_SDE_112_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_113_next_state, KeyReg_Inst_ff_SDE_113_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_113_MUX_inst_X,
         KeyReg_Inst_ff_SDE_113_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_114_next_state, KeyReg_Inst_ff_SDE_114_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_114_MUX_inst_X,
         KeyReg_Inst_ff_SDE_114_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_115_next_state, KeyReg_Inst_ff_SDE_115_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_115_MUX_inst_X,
         KeyReg_Inst_ff_SDE_115_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_116_next_state, KeyReg_Inst_ff_SDE_116_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_116_MUX_inst_X,
         KeyReg_Inst_ff_SDE_116_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_117_next_state, KeyReg_Inst_ff_SDE_117_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_117_MUX_inst_X,
         KeyReg_Inst_ff_SDE_117_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_118_next_state, KeyReg_Inst_ff_SDE_118_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_118_MUX_inst_X,
         KeyReg_Inst_ff_SDE_118_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_119_next_state, KeyReg_Inst_ff_SDE_119_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_119_MUX_inst_X,
         KeyReg_Inst_ff_SDE_119_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_120_next_state, KeyReg_Inst_ff_SDE_120_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_120_MUX_inst_X,
         KeyReg_Inst_ff_SDE_120_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_121_next_state, KeyReg_Inst_ff_SDE_121_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_121_MUX_inst_X,
         KeyReg_Inst_ff_SDE_121_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_122_next_state, KeyReg_Inst_ff_SDE_122_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_122_MUX_inst_X,
         KeyReg_Inst_ff_SDE_122_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_123_next_state, KeyReg_Inst_ff_SDE_123_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_123_MUX_inst_X,
         KeyReg_Inst_ff_SDE_123_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_124_next_state, KeyReg_Inst_ff_SDE_124_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_124_MUX_inst_X,
         KeyReg_Inst_ff_SDE_124_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_125_next_state, KeyReg_Inst_ff_SDE_125_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_125_MUX_inst_X,
         KeyReg_Inst_ff_SDE_125_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_126_next_state, KeyReg_Inst_ff_SDE_126_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_126_MUX_inst_X,
         KeyReg_Inst_ff_SDE_126_current_state_reg_QN,
         KeyReg_Inst_ff_SDE_127_next_state, KeyReg_Inst_ff_SDE_127_MUX_inst_Y,
         KeyReg_Inst_ff_SDE_127_MUX_inst_X,
         KeyReg_Inst_ff_SDE_127_current_state_reg_QN,
         KeyExpansionIns_KeySchedCoreInst_OutBytes_0__0_,
         KeyExpansionIns_KeySchedCoreInst_OutBytes_0__1_,
         KeyExpansionIns_KeySchedCoreInst_OutBytes_0__2_,
         KeyExpansionIns_KeySchedCoreInst_OutBytes_0__3_,
         KeyExpansionIns_KeySchedCoreInst_OutBytes_0__4_,
         KeyExpansionIns_KeySchedCoreInst_OutBytes_0__5_,
         KeyExpansionIns_KeySchedCoreInst_OutBytes_0__6_,
         KeyExpansionIns_KeySchedCoreInst_OutBytes_0__7_,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L29,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L28,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L27,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L26,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L25,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L24,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L23,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L22,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L21,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L20,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L19,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L18,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L17,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L16,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L15,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L14,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L13,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L12,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L11,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L10,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L9,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L8,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L7,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L6,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L5,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L4,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L3,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L2,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L1,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L0,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M63,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M62,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M61,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M60,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M59,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M58,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M57,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M56,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M55,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M54,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M53,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M52,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M51,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M50,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M49,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M48,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M47,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M46,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M45,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M44,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M43,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M42,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M41,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M40,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M39,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M38,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M37,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M36,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M35,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M34,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M33,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M32,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M31,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M30,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M29,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M28,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M27,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M26,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M25,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M24,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M23,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M22,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M21,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M20,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M19,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M18,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M17,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M16,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M15,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M14,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M13,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M12,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M11,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M10,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M9,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M8,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M7,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M6,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M5,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M4,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M3,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M2,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M1,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T27,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T26,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T25,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T24,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T23,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T22,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T21,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T20,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T19,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T18,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T17,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T16,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T15,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T14,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T13,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T12,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T11,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T10,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T9,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T8,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T7,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T5,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T4,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T3,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T2,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L29,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L28,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L27,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L26,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L25,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L24,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L23,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L22,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L21,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L20,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L19,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L18,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L17,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L16,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L15,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L14,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L13,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L12,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L11,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L10,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L9,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L8,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L7,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L6,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L5,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L4,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L3,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L2,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L1,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L0,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M63,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M62,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M61,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M60,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M59,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M58,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M57,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M56,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M55,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M54,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M53,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M52,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M51,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M50,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M49,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M48,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M47,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M46,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M45,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M44,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M43,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M42,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M41,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M40,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M39,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M38,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M37,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M36,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M35,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M34,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M33,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M32,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M31,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M30,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M29,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M28,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M27,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M26,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M25,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M24,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M23,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M22,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M21,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M20,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M19,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M18,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M17,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M16,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M15,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M14,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M13,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M12,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M11,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M10,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M9,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M8,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M7,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M6,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M5,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M4,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M3,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M2,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M1,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T27,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T26,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T25,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T24,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T23,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T22,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T21,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T20,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T19,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T18,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T17,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T16,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T15,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T14,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T13,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T12,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T11,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T10,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T9,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T8,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T7,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T5,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T4,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T3,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T2,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L29,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L28,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L27,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L26,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L25,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L24,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L23,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L22,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L21,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L20,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L19,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L18,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L17,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L16,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L15,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L14,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L13,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L12,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L11,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L10,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L9,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L8,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L7,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L6,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L5,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L4,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L3,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L2,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L1,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L0,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M63,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M62,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M61,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M60,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M59,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M58,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M57,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M56,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M55,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M54,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M53,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M52,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M51,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M50,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M49,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M48,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M47,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M46,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M45,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M44,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M43,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M42,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M41,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M40,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M39,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M38,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M37,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M36,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M35,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M34,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M33,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M32,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M31,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M30,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M29,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M28,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M27,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M26,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M25,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M24,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M23,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M22,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M21,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M20,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M19,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M18,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M17,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M16,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M15,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M14,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M13,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M12,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M11,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M10,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M9,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M8,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M7,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M6,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M5,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M4,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M3,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M2,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M1,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T27,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T26,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T25,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T24,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T23,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T22,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T21,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T20,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T19,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T18,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T17,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T16,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T15,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T14,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T13,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T12,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T11,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T10,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T9,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T8,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T7,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T5,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T4,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T3,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T2,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L29,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L28,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L27,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L26,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L25,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L24,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L23,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L22,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L21,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L20,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L19,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L18,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L17,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L16,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L15,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L14,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L13,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L12,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L11,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L10,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L9,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L8,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L7,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L6,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L5,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L4,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L3,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L2,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L1,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L0,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M63,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M62,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M61,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M60,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M59,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M58,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M57,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M56,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M55,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M54,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M53,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M52,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M51,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M50,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M49,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M48,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M47,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M46,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M45,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M44,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M43,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M42,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M41,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M40,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M39,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M38,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M37,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M36,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M35,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M34,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M33,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M32,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M31,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M30,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M29,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M28,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M27,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M26,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M25,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M24,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M23,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M22,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M21,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M20,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M19,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M18,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M17,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M16,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M15,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M14,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M13,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M12,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M11,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M10,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M9,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M8,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M7,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M6,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M5,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M4,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M3,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M2,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M1,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T27,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T26,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T25,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T24,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T23,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T22,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T21,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T20,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T19,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T18,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T17,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T16,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T15,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T14,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T13,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T12,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T11,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T10,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T9,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T8,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T7,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T5,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T4,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T3,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T2,
         KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1, RoundCounterIns_n8,
         RoundCounterIns_n7, RoundCounterIns_n6, RoundCounterIns_n5,
         RoundCounterIns_n4, RoundCounterIns_n3, RoundCounterIns_n2,
         RoundCounterIns_n24, RoundCounterIns_n25, RoundCounterIns_n1,
         RoundCounterIns_n26, RoundCounterIns_n27,
         RoundCounterIns_count_reg_0__QN, RoundCounterIns_count_reg_2__QN,
         RoundCounterIns_count_reg_3__QN;
  wire   [127:0] RoundOutput;
  wire   [127:8] state_shifted;
  wire   [127:120] RoundInput;
  wire   [119:0] SubBytesInput;
  wire   [123:0] MixColumnsInput;
  wire   [127:0] MixColumnsOutput;
  wire   [127:0] KeyExpansionOutput;
  wire   [127:8] key_shifted;
  wire   [127:120] RoundKey;
  wire   [5:0] Rcon;
  wire   [3:0] RoundCounter;
  wire   [31:0] MixColumnsIns_MixOneColumnInst_0_DoubleBytes;
  wire   [31:0] MixColumnsIns_MixOneColumnInst_1_DoubleBytes;
  wire   [31:0] MixColumnsIns_MixOneColumnInst_2_DoubleBytes;
  wire   [31:0] MixColumnsIns_MixOneColumnInst_3_DoubleBytes;
  wire   [31:0] KeyExpansionIns_tmp;

  INV_X8 U1092 ( .A(n845), .ZN(n579) );
  OR2_X1 U1093 ( .A1(start), .A2(done), .ZN(start_done) );
  INV_X1 U1094 ( .A(n579), .ZN(n574) );
  INV_X1 U1095 ( .A(n579), .ZN(n576) );
  INV_X1 U1096 ( .A(n579), .ZN(n575) );
  INV_X1 U1097 ( .A(n579), .ZN(n577) );
  INV_X1 U1098 ( .A(n579), .ZN(n578) );
  NAND2_X1 U1099 ( .A1(RoundCounter[0]), .A2(n587), .ZN(n845) );
  NOR2_X1 U1100 ( .A1(n852), .A2(n580), .ZN(n587) );
  INV_X1 U1101 ( .A(notdone), .ZN(done) );
  NAND2_X1 U1102 ( .A1(n854), .A2(n853), .ZN(notdone) );
  INV_X1 U1103 ( .A(RoundCounter[3]), .ZN(n852) );
  NOR2_X1 U1104 ( .A1(RoundCounter[2]), .A2(n584), .ZN(n854) );
  INV_X1 U1105 ( .A(RoundCounter[1]), .ZN(n584) );
  INV_X1 U1106 ( .A(RoundCounter[2]), .ZN(n851) );
  NOR2_X1 U1107 ( .A1(RoundCounter[0]), .A2(n852), .ZN(n853) );
  NAND2_X1 U1108 ( .A1(n851), .A2(n584), .ZN(n580) );
  NOR2_X1 U1109 ( .A1(RoundCounter[0]), .A2(n580), .ZN(Rcon[0]) );
  NOR2_X1 U1110 ( .A1(RoundCounter[0]), .A2(RoundCounter[3]), .ZN(n849) );
  NOR2_X1 U1111 ( .A1(n849), .A2(n580), .ZN(Rcon[1]) );
  NAND2_X1 U1112 ( .A1(n854), .A2(n849), .ZN(n581) );
  NAND2_X1 U1113 ( .A1(n578), .A2(n581), .ZN(Rcon[2]) );
  NAND2_X1 U1114 ( .A1(RoundCounter[0]), .A2(n852), .ZN(n589) );
  NOR2_X1 U1115 ( .A1(n584), .A2(n589), .ZN(n848) );
  NAND2_X1 U1116 ( .A1(n848), .A2(n851), .ZN(n583) );
  NAND2_X1 U1117 ( .A1(RoundCounter[3]), .A2(Rcon[0]), .ZN(n582) );
  NAND2_X1 U1118 ( .A1(n583), .A2(n582), .ZN(Rcon[3]) );
  INV_X1 U1119 ( .A(n849), .ZN(n585) );
  NAND2_X1 U1120 ( .A1(RoundCounter[2]), .A2(n584), .ZN(n588) );
  NOR2_X1 U1121 ( .A1(n585), .A2(n588), .ZN(n586) );
  OR2_X1 U1122 ( .A1(n587), .A2(n586), .ZN(Rcon[4]) );
  OR2_X1 U1123 ( .A1(n589), .A2(n588), .ZN(n590) );
  NAND2_X1 U1124 ( .A1(n578), .A2(n590), .ZN(Rcon[5]) );
  NAND2_X1 U1125 ( .A1(MixColumnsOutput[0]), .A2(n578), .ZN(n592) );
  NAND2_X1 U1126 ( .A1(n579), .A2(MixColumnsInput[0]), .ZN(n591) );
  NAND2_X1 U1127 ( .A1(n592), .A2(n591), .ZN(RoundOutput[0]) );
  NAND2_X1 U1128 ( .A1(MixColumnsOutput[100]), .A2(n578), .ZN(n594) );
  NAND2_X1 U1129 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[5]), .ZN(n593) );
  NAND2_X1 U1130 ( .A1(n594), .A2(n593), .ZN(RoundOutput[100]) );
  NAND2_X1 U1131 ( .A1(MixColumnsOutput[101]), .A2(n578), .ZN(n596) );
  NAND2_X1 U1132 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[6]), .ZN(n595) );
  NAND2_X1 U1133 ( .A1(n596), .A2(n595), .ZN(RoundOutput[101]) );
  NAND2_X1 U1134 ( .A1(MixColumnsOutput[102]), .A2(n578), .ZN(n598) );
  NAND2_X1 U1135 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[7]), .ZN(n597) );
  NAND2_X1 U1136 ( .A1(n598), .A2(n597), .ZN(RoundOutput[102]) );
  NAND2_X1 U1137 ( .A1(MixColumnsOutput[103]), .A2(n578), .ZN(n600) );
  NAND2_X1 U1138 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]), .ZN(n599) );
  NAND2_X1 U1139 ( .A1(n600), .A2(n599), .ZN(RoundOutput[103]) );
  NAND2_X1 U1140 ( .A1(MixColumnsOutput[104]), .A2(n578), .ZN(n602) );
  NAND2_X1 U1141 ( .A1(n579), .A2(MixColumnsInput[104]), .ZN(n601) );
  NAND2_X1 U1142 ( .A1(n602), .A2(n601), .ZN(RoundOutput[104]) );
  NAND2_X1 U1143 ( .A1(MixColumnsOutput[105]), .A2(n578), .ZN(n604) );
  NAND2_X1 U1144 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[10]), .ZN(n603) );
  NAND2_X1 U1145 ( .A1(n604), .A2(n603), .ZN(RoundOutput[105]) );
  NAND2_X1 U1146 ( .A1(MixColumnsOutput[106]), .A2(n578), .ZN(n606) );
  NAND2_X1 U1147 ( .A1(n579), .A2(MixColumnsInput[106]), .ZN(n605) );
  NAND2_X1 U1148 ( .A1(n606), .A2(n605), .ZN(RoundOutput[106]) );
  NAND2_X1 U1149 ( .A1(MixColumnsOutput[107]), .A2(n577), .ZN(n608) );
  NAND2_X1 U1150 ( .A1(n579), .A2(MixColumnsInput[107]), .ZN(n607) );
  NAND2_X1 U1151 ( .A1(n608), .A2(n607), .ZN(RoundOutput[107]) );
  NAND2_X1 U1152 ( .A1(MixColumnsOutput[108]), .A2(n577), .ZN(n610) );
  NAND2_X1 U1153 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[13]), .ZN(n609) );
  NAND2_X1 U1154 ( .A1(n610), .A2(n609), .ZN(RoundOutput[108]) );
  NAND2_X1 U1155 ( .A1(MixColumnsOutput[109]), .A2(n577), .ZN(n612) );
  NAND2_X1 U1156 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[14]), .ZN(n611) );
  NAND2_X1 U1157 ( .A1(n612), .A2(n611), .ZN(RoundOutput[109]) );
  NAND2_X1 U1158 ( .A1(MixColumnsOutput[10]), .A2(n577), .ZN(n614) );
  NAND2_X1 U1159 ( .A1(n579), .A2(MixColumnsInput[10]), .ZN(n613) );
  NAND2_X1 U1160 ( .A1(n614), .A2(n613), .ZN(RoundOutput[10]) );
  NAND2_X1 U1161 ( .A1(MixColumnsOutput[110]), .A2(n577), .ZN(n616) );
  NAND2_X1 U1162 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[15]), .ZN(n615) );
  NAND2_X1 U1163 ( .A1(n616), .A2(n615), .ZN(RoundOutput[110]) );
  NAND2_X1 U1164 ( .A1(MixColumnsOutput[111]), .A2(n577), .ZN(n618) );
  NAND2_X1 U1165 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]), .ZN(n617) );
  NAND2_X1 U1166 ( .A1(n618), .A2(n617), .ZN(RoundOutput[111]) );
  NAND2_X1 U1167 ( .A1(MixColumnsOutput[112]), .A2(n577), .ZN(n620) );
  NAND2_X1 U1168 ( .A1(n579), .A2(MixColumnsInput[112]), .ZN(n619) );
  NAND2_X1 U1169 ( .A1(n620), .A2(n619), .ZN(RoundOutput[112]) );
  NAND2_X1 U1170 ( .A1(MixColumnsOutput[113]), .A2(n577), .ZN(n622) );
  NAND2_X1 U1171 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[18]), .ZN(n621) );
  NAND2_X1 U1172 ( .A1(n622), .A2(n621), .ZN(RoundOutput[113]) );
  NAND2_X1 U1173 ( .A1(MixColumnsOutput[114]), .A2(n577), .ZN(n624) );
  NAND2_X1 U1174 ( .A1(n579), .A2(MixColumnsInput[114]), .ZN(n623) );
  NAND2_X1 U1175 ( .A1(n624), .A2(n623), .ZN(RoundOutput[114]) );
  NAND2_X1 U1176 ( .A1(MixColumnsOutput[115]), .A2(n577), .ZN(n626) );
  NAND2_X1 U1177 ( .A1(n579), .A2(MixColumnsInput[115]), .ZN(n625) );
  NAND2_X1 U1178 ( .A1(n626), .A2(n625), .ZN(RoundOutput[115]) );
  NAND2_X1 U1179 ( .A1(MixColumnsOutput[116]), .A2(n577), .ZN(n628) );
  NAND2_X1 U1180 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[21]), .ZN(n627) );
  NAND2_X1 U1181 ( .A1(n628), .A2(n627), .ZN(RoundOutput[116]) );
  NAND2_X1 U1182 ( .A1(MixColumnsOutput[117]), .A2(n577), .ZN(n630) );
  NAND2_X1 U1183 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[22]), .ZN(n629) );
  NAND2_X1 U1184 ( .A1(n630), .A2(n629), .ZN(RoundOutput[117]) );
  NAND2_X1 U1185 ( .A1(MixColumnsOutput[118]), .A2(n576), .ZN(n632) );
  NAND2_X1 U1186 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[23]), .ZN(n631) );
  NAND2_X1 U1187 ( .A1(n632), .A2(n631), .ZN(RoundOutput[118]) );
  NAND2_X1 U1188 ( .A1(MixColumnsOutput[119]), .A2(n576), .ZN(n634) );
  NAND2_X1 U1189 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]), .ZN(n633) );
  NAND2_X1 U1190 ( .A1(n634), .A2(n633), .ZN(RoundOutput[119]) );
  NAND2_X1 U1191 ( .A1(MixColumnsOutput[11]), .A2(n576), .ZN(n636) );
  NAND2_X1 U1192 ( .A1(n579), .A2(MixColumnsInput[11]), .ZN(n635) );
  NAND2_X1 U1193 ( .A1(n636), .A2(n635), .ZN(RoundOutput[11]) );
  NAND2_X1 U1194 ( .A1(MixColumnsOutput[120]), .A2(n576), .ZN(n638) );
  NAND2_X1 U1195 ( .A1(n579), .A2(MixColumnsInput[120]), .ZN(n637) );
  NAND2_X1 U1196 ( .A1(n638), .A2(n637), .ZN(RoundOutput[120]) );
  NAND2_X1 U1197 ( .A1(MixColumnsOutput[121]), .A2(n576), .ZN(n640) );
  NAND2_X1 U1198 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[26]), .ZN(n639) );
  NAND2_X1 U1199 ( .A1(n640), .A2(n639), .ZN(RoundOutput[121]) );
  NAND2_X1 U1200 ( .A1(MixColumnsOutput[122]), .A2(n576), .ZN(n642) );
  NAND2_X1 U1201 ( .A1(n579), .A2(MixColumnsInput[122]), .ZN(n641) );
  NAND2_X1 U1202 ( .A1(n642), .A2(n641), .ZN(RoundOutput[122]) );
  NAND2_X1 U1203 ( .A1(MixColumnsOutput[123]), .A2(n576), .ZN(n644) );
  NAND2_X1 U1204 ( .A1(n579), .A2(MixColumnsInput[123]), .ZN(n643) );
  NAND2_X1 U1205 ( .A1(n644), .A2(n643), .ZN(RoundOutput[123]) );
  NAND2_X1 U1206 ( .A1(MixColumnsOutput[124]), .A2(n576), .ZN(n646) );
  NAND2_X1 U1207 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[29]), .ZN(n645) );
  NAND2_X1 U1208 ( .A1(n646), .A2(n645), .ZN(RoundOutput[124]) );
  NAND2_X1 U1209 ( .A1(MixColumnsOutput[125]), .A2(n576), .ZN(n648) );
  NAND2_X1 U1210 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[30]), .ZN(n647) );
  NAND2_X1 U1211 ( .A1(n648), .A2(n647), .ZN(RoundOutput[125]) );
  NAND2_X1 U1212 ( .A1(MixColumnsOutput[126]), .A2(n576), .ZN(n650) );
  NAND2_X1 U1213 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[31]), .ZN(n649) );
  NAND2_X1 U1214 ( .A1(n650), .A2(n649), .ZN(RoundOutput[126]) );
  NAND2_X1 U1215 ( .A1(MixColumnsOutput[127]), .A2(n576), .ZN(n652) );
  NAND2_X1 U1216 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]), .ZN(n651) );
  NAND2_X1 U1217 ( .A1(n652), .A2(n651), .ZN(RoundOutput[127]) );
  NAND2_X1 U1218 ( .A1(MixColumnsOutput[12]), .A2(n576), .ZN(n654) );
  NAND2_X1 U1219 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[13]), .ZN(n653) );
  NAND2_X1 U1220 ( .A1(n654), .A2(n653), .ZN(RoundOutput[12]) );
  NAND2_X1 U1221 ( .A1(MixColumnsOutput[13]), .A2(n575), .ZN(n656) );
  NAND2_X1 U1222 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[14]), .ZN(n655) );
  NAND2_X1 U1223 ( .A1(n656), .A2(n655), .ZN(RoundOutput[13]) );
  NAND2_X1 U1224 ( .A1(MixColumnsOutput[14]), .A2(n575), .ZN(n658) );
  NAND2_X1 U1225 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[15]), .ZN(n657) );
  NAND2_X1 U1226 ( .A1(n658), .A2(n657), .ZN(RoundOutput[14]) );
  NAND2_X1 U1227 ( .A1(MixColumnsOutput[15]), .A2(n575), .ZN(n660) );
  NAND2_X1 U1228 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]), .ZN(n659) );
  NAND2_X1 U1229 ( .A1(n660), .A2(n659), .ZN(RoundOutput[15]) );
  NAND2_X1 U1230 ( .A1(MixColumnsOutput[16]), .A2(n575), .ZN(n662) );
  NAND2_X1 U1231 ( .A1(n579), .A2(MixColumnsInput[16]), .ZN(n661) );
  NAND2_X1 U1232 ( .A1(n662), .A2(n661), .ZN(RoundOutput[16]) );
  NAND2_X1 U1233 ( .A1(MixColumnsOutput[17]), .A2(n575), .ZN(n664) );
  NAND2_X1 U1234 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[18]), .ZN(n663) );
  NAND2_X1 U1235 ( .A1(n664), .A2(n663), .ZN(RoundOutput[17]) );
  NAND2_X1 U1236 ( .A1(MixColumnsOutput[18]), .A2(n575), .ZN(n666) );
  NAND2_X1 U1237 ( .A1(n579), .A2(MixColumnsInput[18]), .ZN(n665) );
  NAND2_X1 U1238 ( .A1(n666), .A2(n665), .ZN(RoundOutput[18]) );
  NAND2_X1 U1239 ( .A1(MixColumnsOutput[19]), .A2(n575), .ZN(n668) );
  NAND2_X1 U1240 ( .A1(n579), .A2(MixColumnsInput[19]), .ZN(n667) );
  NAND2_X1 U1241 ( .A1(n668), .A2(n667), .ZN(RoundOutput[19]) );
  NAND2_X1 U1242 ( .A1(MixColumnsOutput[1]), .A2(n575), .ZN(n670) );
  NAND2_X1 U1243 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[2]), .ZN(n669) );
  NAND2_X1 U1244 ( .A1(n670), .A2(n669), .ZN(RoundOutput[1]) );
  NAND2_X1 U1245 ( .A1(MixColumnsOutput[20]), .A2(n575), .ZN(n672) );
  NAND2_X1 U1246 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[21]), .ZN(n671) );
  NAND2_X1 U1247 ( .A1(n672), .A2(n671), .ZN(RoundOutput[20]) );
  NAND2_X1 U1248 ( .A1(MixColumnsOutput[21]), .A2(n575), .ZN(n674) );
  NAND2_X1 U1249 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[22]), .ZN(n673) );
  NAND2_X1 U1250 ( .A1(n674), .A2(n673), .ZN(RoundOutput[21]) );
  NAND2_X1 U1251 ( .A1(MixColumnsOutput[22]), .A2(n575), .ZN(n676) );
  NAND2_X1 U1252 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[23]), .ZN(n675) );
  NAND2_X1 U1253 ( .A1(n676), .A2(n675), .ZN(RoundOutput[22]) );
  NAND2_X1 U1254 ( .A1(MixColumnsOutput[23]), .A2(n575), .ZN(n678) );
  NAND2_X1 U1255 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]), .ZN(n677) );
  NAND2_X1 U1256 ( .A1(n678), .A2(n677), .ZN(RoundOutput[23]) );
  NAND2_X1 U1257 ( .A1(MixColumnsOutput[24]), .A2(n574), .ZN(n680) );
  NAND2_X1 U1258 ( .A1(n579), .A2(MixColumnsInput[24]), .ZN(n679) );
  NAND2_X1 U1259 ( .A1(n680), .A2(n679), .ZN(RoundOutput[24]) );
  NAND2_X1 U1260 ( .A1(MixColumnsOutput[25]), .A2(n574), .ZN(n682) );
  NAND2_X1 U1261 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[26]), .ZN(n681) );
  NAND2_X1 U1262 ( .A1(n682), .A2(n681), .ZN(RoundOutput[25]) );
  NAND2_X1 U1263 ( .A1(MixColumnsOutput[26]), .A2(n574), .ZN(n684) );
  NAND2_X1 U1264 ( .A1(n579), .A2(MixColumnsInput[26]), .ZN(n683) );
  NAND2_X1 U1265 ( .A1(n684), .A2(n683), .ZN(RoundOutput[26]) );
  NAND2_X1 U1266 ( .A1(MixColumnsOutput[27]), .A2(n574), .ZN(n686) );
  NAND2_X1 U1267 ( .A1(n579), .A2(MixColumnsInput[27]), .ZN(n685) );
  NAND2_X1 U1268 ( .A1(n686), .A2(n685), .ZN(RoundOutput[27]) );
  NAND2_X1 U1269 ( .A1(MixColumnsOutput[28]), .A2(n574), .ZN(n688) );
  NAND2_X1 U1270 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[29]), .ZN(n687) );
  NAND2_X1 U1271 ( .A1(n688), .A2(n687), .ZN(RoundOutput[28]) );
  NAND2_X1 U1272 ( .A1(MixColumnsOutput[29]), .A2(n574), .ZN(n690) );
  NAND2_X1 U1273 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[30]), .ZN(n689) );
  NAND2_X1 U1274 ( .A1(n690), .A2(n689), .ZN(RoundOutput[29]) );
  NAND2_X1 U1275 ( .A1(MixColumnsOutput[2]), .A2(n574), .ZN(n692) );
  NAND2_X1 U1276 ( .A1(n579), .A2(MixColumnsInput[2]), .ZN(n691) );
  NAND2_X1 U1277 ( .A1(n692), .A2(n691), .ZN(RoundOutput[2]) );
  NAND2_X1 U1278 ( .A1(MixColumnsOutput[30]), .A2(n574), .ZN(n694) );
  NAND2_X1 U1279 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[31]), .ZN(n693) );
  NAND2_X1 U1280 ( .A1(n694), .A2(n693), .ZN(RoundOutput[30]) );
  NAND2_X1 U1281 ( .A1(MixColumnsOutput[31]), .A2(n574), .ZN(n696) );
  NAND2_X1 U1282 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]), .ZN(n695) );
  NAND2_X1 U1283 ( .A1(n696), .A2(n695), .ZN(RoundOutput[31]) );
  NAND2_X1 U1284 ( .A1(MixColumnsOutput[32]), .A2(n574), .ZN(n698) );
  NAND2_X1 U1285 ( .A1(n579), .A2(MixColumnsInput[32]), .ZN(n697) );
  NAND2_X1 U1286 ( .A1(n698), .A2(n697), .ZN(RoundOutput[32]) );
  NAND2_X1 U1287 ( .A1(MixColumnsOutput[33]), .A2(n574), .ZN(n700) );
  NAND2_X1 U1288 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[2]), .ZN(n699) );
  NAND2_X1 U1289 ( .A1(n700), .A2(n699), .ZN(RoundOutput[33]) );
  NAND2_X1 U1290 ( .A1(MixColumnsOutput[34]), .A2(n574), .ZN(n702) );
  NAND2_X1 U1291 ( .A1(n579), .A2(MixColumnsInput[34]), .ZN(n701) );
  NAND2_X1 U1292 ( .A1(n702), .A2(n701), .ZN(RoundOutput[34]) );
  NAND2_X1 U1293 ( .A1(MixColumnsOutput[35]), .A2(n845), .ZN(n704) );
  NAND2_X1 U1294 ( .A1(n579), .A2(MixColumnsInput[35]), .ZN(n703) );
  NAND2_X1 U1295 ( .A1(n704), .A2(n703), .ZN(RoundOutput[35]) );
  NAND2_X1 U1296 ( .A1(MixColumnsOutput[36]), .A2(n578), .ZN(n706) );
  NAND2_X1 U1297 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[5]), .ZN(n705) );
  NAND2_X1 U1298 ( .A1(n706), .A2(n705), .ZN(RoundOutput[36]) );
  NAND2_X1 U1299 ( .A1(MixColumnsOutput[37]), .A2(n578), .ZN(n708) );
  NAND2_X1 U1300 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[6]), .ZN(n707) );
  NAND2_X1 U1301 ( .A1(n708), .A2(n707), .ZN(RoundOutput[37]) );
  NAND2_X1 U1302 ( .A1(MixColumnsOutput[38]), .A2(n845), .ZN(n710) );
  NAND2_X1 U1303 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[7]), .ZN(n709) );
  NAND2_X1 U1304 ( .A1(n710), .A2(n709), .ZN(RoundOutput[38]) );
  NAND2_X1 U1305 ( .A1(MixColumnsOutput[39]), .A2(n845), .ZN(n712) );
  NAND2_X1 U1306 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]), .ZN(n711) );
  NAND2_X1 U1307 ( .A1(n712), .A2(n711), .ZN(RoundOutput[39]) );
  NAND2_X1 U1308 ( .A1(MixColumnsOutput[3]), .A2(n578), .ZN(n714) );
  NAND2_X1 U1309 ( .A1(n579), .A2(MixColumnsInput[3]), .ZN(n713) );
  NAND2_X1 U1310 ( .A1(n714), .A2(n713), .ZN(RoundOutput[3]) );
  NAND2_X1 U1311 ( .A1(MixColumnsOutput[40]), .A2(n845), .ZN(n716) );
  NAND2_X1 U1312 ( .A1(n579), .A2(MixColumnsInput[40]), .ZN(n715) );
  NAND2_X1 U1313 ( .A1(n716), .A2(n715), .ZN(RoundOutput[40]) );
  NAND2_X1 U1314 ( .A1(MixColumnsOutput[41]), .A2(n845), .ZN(n718) );
  NAND2_X1 U1315 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[10]), .ZN(n717) );
  NAND2_X1 U1316 ( .A1(n718), .A2(n717), .ZN(RoundOutput[41]) );
  NAND2_X1 U1317 ( .A1(MixColumnsOutput[42]), .A2(n845), .ZN(n720) );
  NAND2_X1 U1318 ( .A1(n579), .A2(MixColumnsInput[42]), .ZN(n719) );
  NAND2_X1 U1319 ( .A1(n720), .A2(n719), .ZN(RoundOutput[42]) );
  NAND2_X1 U1320 ( .A1(MixColumnsOutput[43]), .A2(n845), .ZN(n722) );
  NAND2_X1 U1321 ( .A1(n579), .A2(MixColumnsInput[43]), .ZN(n721) );
  NAND2_X1 U1322 ( .A1(n722), .A2(n721), .ZN(RoundOutput[43]) );
  NAND2_X1 U1323 ( .A1(MixColumnsOutput[44]), .A2(n578), .ZN(n724) );
  NAND2_X1 U1324 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[13]), .ZN(n723) );
  NAND2_X1 U1325 ( .A1(n724), .A2(n723), .ZN(RoundOutput[44]) );
  NAND2_X1 U1326 ( .A1(MixColumnsOutput[45]), .A2(n578), .ZN(n726) );
  NAND2_X1 U1327 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[14]), .ZN(n725) );
  NAND2_X1 U1328 ( .A1(n726), .A2(n725), .ZN(RoundOutput[45]) );
  NAND2_X1 U1329 ( .A1(MixColumnsOutput[46]), .A2(n578), .ZN(n728) );
  NAND2_X1 U1330 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[15]), .ZN(n727) );
  NAND2_X1 U1331 ( .A1(n728), .A2(n727), .ZN(RoundOutput[46]) );
  NAND2_X1 U1332 ( .A1(MixColumnsOutput[47]), .A2(n578), .ZN(n730) );
  NAND2_X1 U1333 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]), .ZN(n729) );
  NAND2_X1 U1334 ( .A1(n730), .A2(n729), .ZN(RoundOutput[47]) );
  NAND2_X1 U1335 ( .A1(MixColumnsOutput[48]), .A2(n578), .ZN(n732) );
  NAND2_X1 U1336 ( .A1(n579), .A2(MixColumnsInput[48]), .ZN(n731) );
  NAND2_X1 U1337 ( .A1(n732), .A2(n731), .ZN(RoundOutput[48]) );
  NAND2_X1 U1338 ( .A1(MixColumnsOutput[49]), .A2(n574), .ZN(n734) );
  NAND2_X1 U1339 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[18]), .ZN(n733) );
  NAND2_X1 U1340 ( .A1(n734), .A2(n733), .ZN(RoundOutput[49]) );
  NAND2_X1 U1341 ( .A1(MixColumnsOutput[4]), .A2(n574), .ZN(n736) );
  NAND2_X1 U1342 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[5]), .ZN(n735) );
  NAND2_X1 U1343 ( .A1(n736), .A2(n735), .ZN(RoundOutput[4]) );
  NAND2_X1 U1344 ( .A1(MixColumnsOutput[50]), .A2(n576), .ZN(n738) );
  NAND2_X1 U1345 ( .A1(n579), .A2(MixColumnsInput[50]), .ZN(n737) );
  NAND2_X1 U1346 ( .A1(n738), .A2(n737), .ZN(RoundOutput[50]) );
  NAND2_X1 U1347 ( .A1(MixColumnsOutput[51]), .A2(n575), .ZN(n740) );
  NAND2_X1 U1348 ( .A1(n579), .A2(MixColumnsInput[51]), .ZN(n739) );
  NAND2_X1 U1349 ( .A1(n740), .A2(n739), .ZN(RoundOutput[51]) );
  NAND2_X1 U1350 ( .A1(MixColumnsOutput[52]), .A2(n576), .ZN(n742) );
  NAND2_X1 U1351 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[21]), .ZN(n741) );
  NAND2_X1 U1352 ( .A1(n742), .A2(n741), .ZN(RoundOutput[52]) );
  NAND2_X1 U1353 ( .A1(MixColumnsOutput[53]), .A2(n578), .ZN(n744) );
  NAND2_X1 U1354 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[22]), .ZN(n743) );
  NAND2_X1 U1355 ( .A1(n744), .A2(n743), .ZN(RoundOutput[53]) );
  NAND2_X1 U1356 ( .A1(MixColumnsOutput[54]), .A2(n845), .ZN(n746) );
  NAND2_X1 U1357 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[23]), .ZN(n745) );
  NAND2_X1 U1358 ( .A1(n746), .A2(n745), .ZN(RoundOutput[54]) );
  NAND2_X1 U1359 ( .A1(MixColumnsOutput[55]), .A2(n575), .ZN(n748) );
  NAND2_X1 U1360 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]), .ZN(n747) );
  NAND2_X1 U1361 ( .A1(n748), .A2(n747), .ZN(RoundOutput[55]) );
  NAND2_X1 U1362 ( .A1(MixColumnsOutput[56]), .A2(n845), .ZN(n750) );
  NAND2_X1 U1363 ( .A1(n579), .A2(MixColumnsInput[56]), .ZN(n749) );
  NAND2_X1 U1364 ( .A1(n750), .A2(n749), .ZN(RoundOutput[56]) );
  NAND2_X1 U1365 ( .A1(MixColumnsOutput[57]), .A2(n574), .ZN(n752) );
  NAND2_X1 U1366 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[26]), .ZN(n751) );
  NAND2_X1 U1367 ( .A1(n752), .A2(n751), .ZN(RoundOutput[57]) );
  NAND2_X1 U1368 ( .A1(MixColumnsOutput[58]), .A2(n576), .ZN(n754) );
  NAND2_X1 U1369 ( .A1(n579), .A2(MixColumnsInput[58]), .ZN(n753) );
  NAND2_X1 U1370 ( .A1(n754), .A2(n753), .ZN(RoundOutput[58]) );
  NAND2_X1 U1371 ( .A1(MixColumnsOutput[59]), .A2(n577), .ZN(n756) );
  NAND2_X1 U1372 ( .A1(n579), .A2(MixColumnsInput[59]), .ZN(n755) );
  NAND2_X1 U1373 ( .A1(n756), .A2(n755), .ZN(RoundOutput[59]) );
  NAND2_X1 U1374 ( .A1(MixColumnsOutput[5]), .A2(n575), .ZN(n758) );
  NAND2_X1 U1375 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[6]), .ZN(n757) );
  NAND2_X1 U1376 ( .A1(n758), .A2(n757), .ZN(RoundOutput[5]) );
  NAND2_X1 U1377 ( .A1(MixColumnsOutput[60]), .A2(n577), .ZN(n760) );
  NAND2_X1 U1378 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[29]), .ZN(n759) );
  NAND2_X1 U1379 ( .A1(n760), .A2(n759), .ZN(RoundOutput[60]) );
  NAND2_X1 U1380 ( .A1(MixColumnsOutput[61]), .A2(n845), .ZN(n762) );
  NAND2_X1 U1381 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[30]), .ZN(n761) );
  NAND2_X1 U1382 ( .A1(n762), .A2(n761), .ZN(RoundOutput[61]) );
  NAND2_X1 U1383 ( .A1(MixColumnsOutput[62]), .A2(n845), .ZN(n764) );
  NAND2_X1 U1384 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[31]), .ZN(n763) );
  NAND2_X1 U1385 ( .A1(n764), .A2(n763), .ZN(RoundOutput[62]) );
  NAND2_X1 U1386 ( .A1(MixColumnsOutput[63]), .A2(n574), .ZN(n766) );
  NAND2_X1 U1387 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]), .ZN(n765) );
  NAND2_X1 U1388 ( .A1(n766), .A2(n765), .ZN(RoundOutput[63]) );
  NAND2_X1 U1389 ( .A1(MixColumnsOutput[64]), .A2(n574), .ZN(n768) );
  NAND2_X1 U1390 ( .A1(n579), .A2(MixColumnsInput[64]), .ZN(n767) );
  NAND2_X1 U1391 ( .A1(n768), .A2(n767), .ZN(RoundOutput[64]) );
  NAND2_X1 U1392 ( .A1(MixColumnsOutput[65]), .A2(n576), .ZN(n770) );
  NAND2_X1 U1393 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[2]), .ZN(n769) );
  NAND2_X1 U1394 ( .A1(n770), .A2(n769), .ZN(RoundOutput[65]) );
  NAND2_X1 U1395 ( .A1(MixColumnsOutput[66]), .A2(n575), .ZN(n772) );
  NAND2_X1 U1396 ( .A1(n579), .A2(MixColumnsInput[66]), .ZN(n771) );
  NAND2_X1 U1397 ( .A1(n772), .A2(n771), .ZN(RoundOutput[66]) );
  NAND2_X1 U1398 ( .A1(MixColumnsOutput[67]), .A2(n577), .ZN(n774) );
  NAND2_X1 U1399 ( .A1(n579), .A2(MixColumnsInput[67]), .ZN(n773) );
  NAND2_X1 U1400 ( .A1(n774), .A2(n773), .ZN(RoundOutput[67]) );
  NAND2_X1 U1401 ( .A1(MixColumnsOutput[68]), .A2(n845), .ZN(n776) );
  NAND2_X1 U1402 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[5]), .ZN(n775) );
  NAND2_X1 U1403 ( .A1(n776), .A2(n775), .ZN(RoundOutput[68]) );
  NAND2_X1 U1404 ( .A1(MixColumnsOutput[69]), .A2(n845), .ZN(n778) );
  NAND2_X1 U1405 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[6]), .ZN(n777) );
  NAND2_X1 U1406 ( .A1(n778), .A2(n777), .ZN(RoundOutput[69]) );
  NAND2_X1 U1407 ( .A1(MixColumnsOutput[6]), .A2(n845), .ZN(n780) );
  NAND2_X1 U1408 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[7]), .ZN(n779) );
  NAND2_X1 U1409 ( .A1(n780), .A2(n779), .ZN(RoundOutput[6]) );
  NAND2_X1 U1410 ( .A1(MixColumnsOutput[70]), .A2(n574), .ZN(n782) );
  NAND2_X1 U1411 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[7]), .ZN(n781) );
  NAND2_X1 U1412 ( .A1(n782), .A2(n781), .ZN(RoundOutput[70]) );
  NAND2_X1 U1413 ( .A1(MixColumnsOutput[71]), .A2(n574), .ZN(n784) );
  NAND2_X1 U1414 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]), .ZN(n783) );
  NAND2_X1 U1415 ( .A1(n784), .A2(n783), .ZN(RoundOutput[71]) );
  NAND2_X1 U1416 ( .A1(MixColumnsOutput[72]), .A2(n574), .ZN(n786) );
  NAND2_X1 U1417 ( .A1(n579), .A2(MixColumnsInput[72]), .ZN(n785) );
  NAND2_X1 U1418 ( .A1(n786), .A2(n785), .ZN(RoundOutput[72]) );
  NAND2_X1 U1419 ( .A1(MixColumnsOutput[73]), .A2(n576), .ZN(n788) );
  NAND2_X1 U1420 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[10]), .ZN(n787) );
  NAND2_X1 U1421 ( .A1(n788), .A2(n787), .ZN(RoundOutput[73]) );
  NAND2_X1 U1422 ( .A1(MixColumnsOutput[74]), .A2(n575), .ZN(n790) );
  NAND2_X1 U1423 ( .A1(n579), .A2(MixColumnsInput[74]), .ZN(n789) );
  NAND2_X1 U1424 ( .A1(n790), .A2(n789), .ZN(RoundOutput[74]) );
  NAND2_X1 U1425 ( .A1(MixColumnsOutput[75]), .A2(n577), .ZN(n792) );
  NAND2_X1 U1426 ( .A1(n579), .A2(MixColumnsInput[75]), .ZN(n791) );
  NAND2_X1 U1427 ( .A1(n792), .A2(n791), .ZN(RoundOutput[75]) );
  NAND2_X1 U1428 ( .A1(MixColumnsOutput[76]), .A2(n576), .ZN(n794) );
  NAND2_X1 U1429 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[13]), .ZN(n793) );
  NAND2_X1 U1430 ( .A1(n794), .A2(n793), .ZN(RoundOutput[76]) );
  NAND2_X1 U1431 ( .A1(MixColumnsOutput[77]), .A2(n575), .ZN(n796) );
  NAND2_X1 U1432 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[14]), .ZN(n795) );
  NAND2_X1 U1433 ( .A1(n796), .A2(n795), .ZN(RoundOutput[77]) );
  NAND2_X1 U1434 ( .A1(MixColumnsOutput[78]), .A2(n845), .ZN(n798) );
  NAND2_X1 U1435 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[15]), .ZN(n797) );
  NAND2_X1 U1436 ( .A1(n798), .A2(n797), .ZN(RoundOutput[78]) );
  NAND2_X1 U1437 ( .A1(MixColumnsOutput[79]), .A2(n577), .ZN(n800) );
  NAND2_X1 U1438 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]), .ZN(n799) );
  NAND2_X1 U1439 ( .A1(n800), .A2(n799), .ZN(RoundOutput[79]) );
  NAND2_X1 U1440 ( .A1(MixColumnsOutput[7]), .A2(n576), .ZN(n802) );
  NAND2_X1 U1441 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]), .ZN(n801) );
  NAND2_X1 U1442 ( .A1(n802), .A2(n801), .ZN(RoundOutput[7]) );
  NAND2_X1 U1443 ( .A1(MixColumnsOutput[80]), .A2(n575), .ZN(n804) );
  NAND2_X1 U1444 ( .A1(n579), .A2(MixColumnsInput[80]), .ZN(n803) );
  NAND2_X1 U1445 ( .A1(n804), .A2(n803), .ZN(RoundOutput[80]) );
  NAND2_X1 U1446 ( .A1(MixColumnsOutput[81]), .A2(n577), .ZN(n806) );
  NAND2_X1 U1447 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[18]), .ZN(n805) );
  NAND2_X1 U1448 ( .A1(n806), .A2(n805), .ZN(RoundOutput[81]) );
  NAND2_X1 U1449 ( .A1(MixColumnsOutput[82]), .A2(n845), .ZN(n808) );
  NAND2_X1 U1450 ( .A1(n579), .A2(MixColumnsInput[82]), .ZN(n807) );
  NAND2_X1 U1451 ( .A1(n808), .A2(n807), .ZN(RoundOutput[82]) );
  NAND2_X1 U1452 ( .A1(MixColumnsOutput[83]), .A2(n576), .ZN(n810) );
  NAND2_X1 U1453 ( .A1(n579), .A2(MixColumnsInput[83]), .ZN(n809) );
  NAND2_X1 U1454 ( .A1(n810), .A2(n809), .ZN(RoundOutput[83]) );
  NAND2_X1 U1455 ( .A1(MixColumnsOutput[84]), .A2(n574), .ZN(n812) );
  NAND2_X1 U1456 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[21]), .ZN(n811) );
  NAND2_X1 U1457 ( .A1(n812), .A2(n811), .ZN(RoundOutput[84]) );
  NAND2_X1 U1458 ( .A1(MixColumnsOutput[85]), .A2(n576), .ZN(n814) );
  NAND2_X1 U1459 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[22]), .ZN(n813) );
  NAND2_X1 U1460 ( .A1(n814), .A2(n813), .ZN(RoundOutput[85]) );
  NAND2_X1 U1461 ( .A1(MixColumnsOutput[86]), .A2(n575), .ZN(n816) );
  NAND2_X1 U1462 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[23]), .ZN(n815) );
  NAND2_X1 U1463 ( .A1(n816), .A2(n815), .ZN(RoundOutput[86]) );
  NAND2_X1 U1464 ( .A1(MixColumnsOutput[87]), .A2(n577), .ZN(n818) );
  NAND2_X1 U1465 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]), .ZN(n817) );
  NAND2_X1 U1466 ( .A1(n818), .A2(n817), .ZN(RoundOutput[87]) );
  NAND2_X1 U1467 ( .A1(MixColumnsOutput[88]), .A2(n577), .ZN(n820) );
  NAND2_X1 U1468 ( .A1(n579), .A2(MixColumnsInput[88]), .ZN(n819) );
  NAND2_X1 U1469 ( .A1(n820), .A2(n819), .ZN(RoundOutput[88]) );
  NAND2_X1 U1470 ( .A1(MixColumnsOutput[89]), .A2(n845), .ZN(n822) );
  NAND2_X1 U1471 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[26]), .ZN(n821) );
  NAND2_X1 U1472 ( .A1(n822), .A2(n821), .ZN(RoundOutput[89]) );
  NAND2_X1 U1473 ( .A1(MixColumnsOutput[8]), .A2(n575), .ZN(n824) );
  NAND2_X1 U1474 ( .A1(n579), .A2(MixColumnsInput[8]), .ZN(n823) );
  NAND2_X1 U1475 ( .A1(n824), .A2(n823), .ZN(RoundOutput[8]) );
  NAND2_X1 U1476 ( .A1(MixColumnsOutput[90]), .A2(n574), .ZN(n826) );
  NAND2_X1 U1477 ( .A1(n579), .A2(MixColumnsInput[90]), .ZN(n825) );
  NAND2_X1 U1478 ( .A1(n826), .A2(n825), .ZN(RoundOutput[90]) );
  NAND2_X1 U1479 ( .A1(MixColumnsOutput[91]), .A2(n576), .ZN(n828) );
  NAND2_X1 U1480 ( .A1(n579), .A2(MixColumnsInput[91]), .ZN(n827) );
  NAND2_X1 U1481 ( .A1(n828), .A2(n827), .ZN(RoundOutput[91]) );
  NAND2_X1 U1482 ( .A1(MixColumnsOutput[92]), .A2(n575), .ZN(n830) );
  NAND2_X1 U1483 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[29]), .ZN(n829) );
  NAND2_X1 U1484 ( .A1(n830), .A2(n829), .ZN(RoundOutput[92]) );
  NAND2_X1 U1485 ( .A1(MixColumnsOutput[93]), .A2(n577), .ZN(n832) );
  NAND2_X1 U1486 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[30]), .ZN(n831) );
  NAND2_X1 U1487 ( .A1(n832), .A2(n831), .ZN(RoundOutput[93]) );
  NAND2_X1 U1488 ( .A1(MixColumnsOutput[94]), .A2(n575), .ZN(n834) );
  NAND2_X1 U1489 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[31]), .ZN(n833) );
  NAND2_X1 U1490 ( .A1(n834), .A2(n833), .ZN(RoundOutput[94]) );
  NAND2_X1 U1491 ( .A1(MixColumnsOutput[95]), .A2(n576), .ZN(n836) );
  NAND2_X1 U1492 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]), .ZN(n835) );
  NAND2_X1 U1493 ( .A1(n836), .A2(n835), .ZN(RoundOutput[95]) );
  NAND2_X1 U1494 ( .A1(MixColumnsOutput[96]), .A2(n577), .ZN(n838) );
  NAND2_X1 U1495 ( .A1(n579), .A2(MixColumnsInput[96]), .ZN(n837) );
  NAND2_X1 U1496 ( .A1(n838), .A2(n837), .ZN(RoundOutput[96]) );
  NAND2_X1 U1497 ( .A1(MixColumnsOutput[97]), .A2(n578), .ZN(n840) );
  NAND2_X1 U1498 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[2]), .ZN(n839) );
  NAND2_X1 U1499 ( .A1(n840), .A2(n839), .ZN(RoundOutput[97]) );
  NAND2_X1 U1500 ( .A1(MixColumnsOutput[98]), .A2(n577), .ZN(n842) );
  NAND2_X1 U1501 ( .A1(n579), .A2(MixColumnsInput[98]), .ZN(n841) );
  NAND2_X1 U1502 ( .A1(n842), .A2(n841), .ZN(RoundOutput[98]) );
  NAND2_X1 U1503 ( .A1(MixColumnsOutput[99]), .A2(n574), .ZN(n844) );
  NAND2_X1 U1504 ( .A1(n579), .A2(MixColumnsInput[99]), .ZN(n843) );
  NAND2_X1 U1505 ( .A1(n844), .A2(n843), .ZN(RoundOutput[99]) );
  NAND2_X1 U1506 ( .A1(MixColumnsOutput[9]), .A2(n578), .ZN(n847) );
  NAND2_X1 U1507 ( .A1(n579), .A2(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[10]), .ZN(n846) );
  NAND2_X1 U1508 ( .A1(n847), .A2(n846), .ZN(RoundOutput[9]) );
  XOR2_X1 U1509 ( .A(key_shifted[8]), .B(state_shifted[8]), .Z(
        SubBytesInput[0]) );
  XOR2_X1 U1510 ( .A(key_shifted[108]), .B(state_shifted[108]), .Z(
        SubBytesInput[100]) );
  XOR2_X1 U1511 ( .A(key_shifted[109]), .B(state_shifted[109]), .Z(
        SubBytesInput[101]) );
  XOR2_X1 U1512 ( .A(key_shifted[110]), .B(state_shifted[110]), .Z(
        SubBytesInput[102]) );
  XOR2_X1 U1513 ( .A(key_shifted[111]), .B(state_shifted[111]), .Z(
        SubBytesInput[103]) );
  XOR2_X1 U1514 ( .A(key_shifted[112]), .B(state_shifted[112]), .Z(
        SubBytesInput[104]) );
  XOR2_X1 U1515 ( .A(key_shifted[113]), .B(state_shifted[113]), .Z(
        SubBytesInput[105]) );
  XOR2_X1 U1516 ( .A(key_shifted[114]), .B(state_shifted[114]), .Z(
        SubBytesInput[106]) );
  XOR2_X1 U1517 ( .A(key_shifted[115]), .B(state_shifted[115]), .Z(
        SubBytesInput[107]) );
  XOR2_X1 U1518 ( .A(key_shifted[116]), .B(state_shifted[116]), .Z(
        SubBytesInput[108]) );
  XOR2_X1 U1519 ( .A(key_shifted[117]), .B(state_shifted[117]), .Z(
        SubBytesInput[109]) );
  XOR2_X1 U1520 ( .A(key_shifted[18]), .B(state_shifted[18]), .Z(
        SubBytesInput[10]) );
  XOR2_X1 U1521 ( .A(key_shifted[118]), .B(state_shifted[118]), .Z(
        SubBytesInput[110]) );
  XOR2_X1 U1522 ( .A(key_shifted[119]), .B(state_shifted[119]), .Z(
        SubBytesInput[111]) );
  XOR2_X1 U1523 ( .A(key_shifted[120]), .B(state_shifted[120]), .Z(
        SubBytesInput[112]) );
  XOR2_X1 U1524 ( .A(key_shifted[121]), .B(state_shifted[121]), .Z(
        SubBytesInput[113]) );
  XOR2_X1 U1525 ( .A(key_shifted[122]), .B(state_shifted[122]), .Z(
        SubBytesInput[114]) );
  XOR2_X1 U1526 ( .A(key_shifted[123]), .B(state_shifted[123]), .Z(
        SubBytesInput[115]) );
  XOR2_X1 U1527 ( .A(key_shifted[124]), .B(state_shifted[124]), .Z(
        SubBytesInput[116]) );
  XOR2_X1 U1528 ( .A(key_shifted[125]), .B(state_shifted[125]), .Z(
        SubBytesInput[117]) );
  XOR2_X1 U1529 ( .A(key_shifted[126]), .B(state_shifted[126]), .Z(
        SubBytesInput[118]) );
  XOR2_X1 U1530 ( .A(key_shifted[127]), .B(state_shifted[127]), .Z(
        SubBytesInput[119]) );
  XOR2_X1 U1531 ( .A(key_shifted[19]), .B(state_shifted[19]), .Z(
        SubBytesInput[11]) );
  XOR2_X1 U1532 ( .A(key_shifted[20]), .B(state_shifted[20]), .Z(
        SubBytesInput[12]) );
  XOR2_X1 U1533 ( .A(key_shifted[21]), .B(state_shifted[21]), .Z(
        SubBytesInput[13]) );
  XOR2_X1 U1534 ( .A(key_shifted[22]), .B(state_shifted[22]), .Z(
        SubBytesInput[14]) );
  XOR2_X1 U1535 ( .A(key_shifted[23]), .B(state_shifted[23]), .Z(
        SubBytesInput[15]) );
  XOR2_X1 U1536 ( .A(key_shifted[24]), .B(state_shifted[24]), .Z(
        SubBytesInput[16]) );
  XOR2_X1 U1537 ( .A(key_shifted[25]), .B(state_shifted[25]), .Z(
        SubBytesInput[17]) );
  XOR2_X1 U1538 ( .A(key_shifted[26]), .B(state_shifted[26]), .Z(
        SubBytesInput[18]) );
  XOR2_X1 U1539 ( .A(key_shifted[27]), .B(state_shifted[27]), .Z(
        SubBytesInput[19]) );
  XOR2_X1 U1540 ( .A(key_shifted[9]), .B(state_shifted[9]), .Z(
        SubBytesInput[1]) );
  XOR2_X1 U1541 ( .A(key_shifted[28]), .B(state_shifted[28]), .Z(
        SubBytesInput[20]) );
  XOR2_X1 U1542 ( .A(key_shifted[29]), .B(state_shifted[29]), .Z(
        SubBytesInput[21]) );
  XOR2_X1 U1543 ( .A(key_shifted[30]), .B(state_shifted[30]), .Z(
        SubBytesInput[22]) );
  XOR2_X1 U1544 ( .A(key_shifted[31]), .B(state_shifted[31]), .Z(
        SubBytesInput[23]) );
  XOR2_X1 U1545 ( .A(key_shifted[32]), .B(state_shifted[32]), .Z(
        SubBytesInput[24]) );
  XOR2_X1 U1546 ( .A(key_shifted[33]), .B(state_shifted[33]), .Z(
        SubBytesInput[25]) );
  XOR2_X1 U1547 ( .A(key_shifted[34]), .B(state_shifted[34]), .Z(
        SubBytesInput[26]) );
  XOR2_X1 U1548 ( .A(key_shifted[35]), .B(state_shifted[35]), .Z(
        SubBytesInput[27]) );
  XOR2_X1 U1549 ( .A(key_shifted[36]), .B(state_shifted[36]), .Z(
        SubBytesInput[28]) );
  XOR2_X1 U1550 ( .A(key_shifted[37]), .B(state_shifted[37]), .Z(
        SubBytesInput[29]) );
  XOR2_X1 U1551 ( .A(key_shifted[10]), .B(state_shifted[10]), .Z(
        SubBytesInput[2]) );
  XOR2_X1 U1552 ( .A(key_shifted[38]), .B(state_shifted[38]), .Z(
        SubBytesInput[30]) );
  XOR2_X1 U1553 ( .A(key_shifted[39]), .B(state_shifted[39]), .Z(
        SubBytesInput[31]) );
  XOR2_X1 U1554 ( .A(key_shifted[40]), .B(state_shifted[40]), .Z(
        SubBytesInput[32]) );
  XOR2_X1 U1555 ( .A(key_shifted[41]), .B(state_shifted[41]), .Z(
        SubBytesInput[33]) );
  XOR2_X1 U1556 ( .A(key_shifted[42]), .B(state_shifted[42]), .Z(
        SubBytesInput[34]) );
  XOR2_X1 U1557 ( .A(key_shifted[43]), .B(state_shifted[43]), .Z(
        SubBytesInput[35]) );
  XOR2_X1 U1558 ( .A(key_shifted[44]), .B(state_shifted[44]), .Z(
        SubBytesInput[36]) );
  XOR2_X1 U1559 ( .A(key_shifted[45]), .B(state_shifted[45]), .Z(
        SubBytesInput[37]) );
  XOR2_X1 U1560 ( .A(key_shifted[46]), .B(state_shifted[46]), .Z(
        SubBytesInput[38]) );
  XOR2_X1 U1561 ( .A(key_shifted[47]), .B(state_shifted[47]), .Z(
        SubBytesInput[39]) );
  XOR2_X1 U1562 ( .A(key_shifted[11]), .B(state_shifted[11]), .Z(
        SubBytesInput[3]) );
  XOR2_X1 U1563 ( .A(key_shifted[48]), .B(state_shifted[48]), .Z(
        SubBytesInput[40]) );
  XOR2_X1 U1564 ( .A(key_shifted[49]), .B(state_shifted[49]), .Z(
        SubBytesInput[41]) );
  XOR2_X1 U1565 ( .A(key_shifted[50]), .B(state_shifted[50]), .Z(
        SubBytesInput[42]) );
  XOR2_X1 U1566 ( .A(key_shifted[51]), .B(state_shifted[51]), .Z(
        SubBytesInput[43]) );
  XOR2_X1 U1567 ( .A(key_shifted[52]), .B(state_shifted[52]), .Z(
        SubBytesInput[44]) );
  XOR2_X1 U1568 ( .A(key_shifted[53]), .B(state_shifted[53]), .Z(
        SubBytesInput[45]) );
  XOR2_X1 U1569 ( .A(key_shifted[54]), .B(state_shifted[54]), .Z(
        SubBytesInput[46]) );
  XOR2_X1 U1570 ( .A(key_shifted[55]), .B(state_shifted[55]), .Z(
        SubBytesInput[47]) );
  XOR2_X1 U1571 ( .A(key_shifted[56]), .B(state_shifted[56]), .Z(
        SubBytesInput[48]) );
  XOR2_X1 U1572 ( .A(key_shifted[57]), .B(state_shifted[57]), .Z(
        SubBytesInput[49]) );
  XOR2_X1 U1573 ( .A(key_shifted[12]), .B(state_shifted[12]), .Z(
        SubBytesInput[4]) );
  XOR2_X1 U1574 ( .A(key_shifted[58]), .B(state_shifted[58]), .Z(
        SubBytesInput[50]) );
  XOR2_X1 U1575 ( .A(key_shifted[59]), .B(state_shifted[59]), .Z(
        SubBytesInput[51]) );
  XOR2_X1 U1576 ( .A(key_shifted[60]), .B(state_shifted[60]), .Z(
        SubBytesInput[52]) );
  XOR2_X1 U1577 ( .A(key_shifted[61]), .B(state_shifted[61]), .Z(
        SubBytesInput[53]) );
  XOR2_X1 U1578 ( .A(key_shifted[62]), .B(state_shifted[62]), .Z(
        SubBytesInput[54]) );
  XOR2_X1 U1579 ( .A(key_shifted[63]), .B(state_shifted[63]), .Z(
        SubBytesInput[55]) );
  XOR2_X1 U1580 ( .A(key_shifted[64]), .B(state_shifted[64]), .Z(
        SubBytesInput[56]) );
  XOR2_X1 U1581 ( .A(key_shifted[65]), .B(state_shifted[65]), .Z(
        SubBytesInput[57]) );
  XOR2_X1 U1582 ( .A(key_shifted[66]), .B(state_shifted[66]), .Z(
        SubBytesInput[58]) );
  XOR2_X1 U1583 ( .A(key_shifted[67]), .B(state_shifted[67]), .Z(
        SubBytesInput[59]) );
  XOR2_X1 U1584 ( .A(key_shifted[13]), .B(state_shifted[13]), .Z(
        SubBytesInput[5]) );
  XOR2_X1 U1585 ( .A(key_shifted[68]), .B(state_shifted[68]), .Z(
        SubBytesInput[60]) );
  XOR2_X1 U1586 ( .A(key_shifted[69]), .B(state_shifted[69]), .Z(
        SubBytesInput[61]) );
  XOR2_X1 U1587 ( .A(key_shifted[70]), .B(state_shifted[70]), .Z(
        SubBytesInput[62]) );
  XOR2_X1 U1588 ( .A(key_shifted[71]), .B(state_shifted[71]), .Z(
        SubBytesInput[63]) );
  XOR2_X1 U1589 ( .A(key_shifted[72]), .B(state_shifted[72]), .Z(
        SubBytesInput[64]) );
  XOR2_X1 U1590 ( .A(key_shifted[73]), .B(state_shifted[73]), .Z(
        SubBytesInput[65]) );
  XOR2_X1 U1591 ( .A(key_shifted[74]), .B(state_shifted[74]), .Z(
        SubBytesInput[66]) );
  XOR2_X1 U1592 ( .A(key_shifted[75]), .B(state_shifted[75]), .Z(
        SubBytesInput[67]) );
  XOR2_X1 U1593 ( .A(key_shifted[76]), .B(state_shifted[76]), .Z(
        SubBytesInput[68]) );
  XOR2_X1 U1594 ( .A(key_shifted[77]), .B(state_shifted[77]), .Z(
        SubBytesInput[69]) );
  XOR2_X1 U1595 ( .A(key_shifted[14]), .B(state_shifted[14]), .Z(
        SubBytesInput[6]) );
  XOR2_X1 U1596 ( .A(key_shifted[78]), .B(state_shifted[78]), .Z(
        SubBytesInput[70]) );
  XOR2_X1 U1597 ( .A(key_shifted[79]), .B(state_shifted[79]), .Z(
        SubBytesInput[71]) );
  XOR2_X1 U1598 ( .A(key_shifted[80]), .B(state_shifted[80]), .Z(
        SubBytesInput[72]) );
  XOR2_X1 U1599 ( .A(key_shifted[81]), .B(state_shifted[81]), .Z(
        SubBytesInput[73]) );
  XOR2_X1 U1600 ( .A(key_shifted[82]), .B(state_shifted[82]), .Z(
        SubBytesInput[74]) );
  XOR2_X1 U1601 ( .A(key_shifted[83]), .B(state_shifted[83]), .Z(
        SubBytesInput[75]) );
  XOR2_X1 U1602 ( .A(key_shifted[84]), .B(state_shifted[84]), .Z(
        SubBytesInput[76]) );
  XOR2_X1 U1603 ( .A(key_shifted[85]), .B(state_shifted[85]), .Z(
        SubBytesInput[77]) );
  XOR2_X1 U1604 ( .A(key_shifted[86]), .B(state_shifted[86]), .Z(
        SubBytesInput[78]) );
  XOR2_X1 U1605 ( .A(key_shifted[87]), .B(state_shifted[87]), .Z(
        SubBytesInput[79]) );
  XOR2_X1 U1606 ( .A(key_shifted[15]), .B(state_shifted[15]), .Z(
        SubBytesInput[7]) );
  XOR2_X1 U1607 ( .A(key_shifted[88]), .B(state_shifted[88]), .Z(
        SubBytesInput[80]) );
  XOR2_X1 U1608 ( .A(key_shifted[89]), .B(state_shifted[89]), .Z(
        SubBytesInput[81]) );
  XOR2_X1 U1609 ( .A(key_shifted[90]), .B(state_shifted[90]), .Z(
        SubBytesInput[82]) );
  XOR2_X1 U1610 ( .A(key_shifted[91]), .B(state_shifted[91]), .Z(
        SubBytesInput[83]) );
  XOR2_X1 U1611 ( .A(key_shifted[92]), .B(state_shifted[92]), .Z(
        SubBytesInput[84]) );
  XOR2_X1 U1612 ( .A(key_shifted[93]), .B(state_shifted[93]), .Z(
        SubBytesInput[85]) );
  XOR2_X1 U1613 ( .A(key_shifted[94]), .B(state_shifted[94]), .Z(
        SubBytesInput[86]) );
  XOR2_X1 U1614 ( .A(key_shifted[95]), .B(state_shifted[95]), .Z(
        SubBytesInput[87]) );
  XOR2_X1 U1615 ( .A(key_shifted[96]), .B(state_shifted[96]), .Z(
        SubBytesInput[88]) );
  XOR2_X1 U1616 ( .A(key_shifted[97]), .B(state_shifted[97]), .Z(
        SubBytesInput[89]) );
  XOR2_X1 U1617 ( .A(key_shifted[16]), .B(state_shifted[16]), .Z(
        SubBytesInput[8]) );
  XOR2_X1 U1618 ( .A(key_shifted[98]), .B(state_shifted[98]), .Z(
        SubBytesInput[90]) );
  XOR2_X1 U1619 ( .A(key_shifted[99]), .B(state_shifted[99]), .Z(
        SubBytesInput[91]) );
  XOR2_X1 U1620 ( .A(key_shifted[100]), .B(state_shifted[100]), .Z(
        SubBytesInput[92]) );
  XOR2_X1 U1621 ( .A(key_shifted[101]), .B(state_shifted[101]), .Z(
        SubBytesInput[93]) );
  XOR2_X1 U1622 ( .A(key_shifted[102]), .B(state_shifted[102]), .Z(
        SubBytesInput[94]) );
  XOR2_X1 U1623 ( .A(key_shifted[103]), .B(state_shifted[103]), .Z(
        SubBytesInput[95]) );
  XOR2_X1 U1624 ( .A(key_shifted[104]), .B(state_shifted[104]), .Z(
        SubBytesInput[96]) );
  XOR2_X1 U1625 ( .A(key_shifted[105]), .B(state_shifted[105]), .Z(
        SubBytesInput[97]) );
  XOR2_X1 U1626 ( .A(key_shifted[106]), .B(state_shifted[106]), .Z(
        SubBytesInput[98]) );
  XOR2_X1 U1627 ( .A(key_shifted[107]), .B(state_shifted[107]), .Z(
        SubBytesInput[99]) );
  XOR2_X1 U1628 ( .A(key_shifted[17]), .B(state_shifted[17]), .Z(
        SubBytesInput[9]) );
  AND2_X1 U1629 ( .A1(RoundCounter[2]), .A2(n848), .ZN(n286) );
  NAND2_X1 U1630 ( .A1(RoundCounter[1]), .A2(n849), .ZN(n850) );
  NOR2_X1 U1631 ( .A1(n851), .A2(n850), .ZN(n287) );
  XOR2_X1 U1632 ( .A(RoundInput[120]), .B(RoundKey[120]), .Z(port_out[0]) );
  XOR2_X1 U1633 ( .A(RoundInput[121]), .B(RoundKey[121]), .Z(port_out[1]) );
  XOR2_X1 U1634 ( .A(RoundInput[122]), .B(RoundKey[122]), .Z(port_out[2]) );
  XOR2_X1 U1635 ( .A(RoundInput[123]), .B(RoundKey[123]), .Z(port_out[3]) );
  XOR2_X1 U1636 ( .A(RoundInput[124]), .B(RoundKey[124]), .Z(port_out[4]) );
  XOR2_X1 U1637 ( .A(RoundInput[125]), .B(RoundKey[125]), .Z(port_out[5]) );
  XOR2_X1 U1638 ( .A(RoundInput[126]), .B(RoundKey[126]), .Z(port_out[6]) );
  XOR2_X1 U1639 ( .A(RoundInput[127]), .B(RoundKey[127]), .Z(port_out[7]) );
  INV_X1 RoundReg_U5 ( .A(start_done), .ZN(RoundReg_n10) );
  INV_X1 RoundReg_U4 ( .A(RoundReg_n10), .ZN(RoundReg_n9) );
  INV_X1 RoundReg_U3 ( .A(RoundReg_n10), .ZN(RoundReg_n8) );
  INV_X1 RoundReg_U2 ( .A(RoundReg_n10), .ZN(RoundReg_n7) );
  INV_X1 RoundReg_U1 ( .A(RoundReg_n10), .ZN(RoundReg_n6) );
  XOR2_X1 RoundReg_Inst_ff_SDE_0_MUX_inst_XOR1_U1 ( .A(RoundOutput[0]), .B(
        port_in[0]), .Z(RoundReg_Inst_ff_SDE_0_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_0_MUX_inst_AND1_U1 ( .A1(RoundReg_n6), .A2(
        RoundReg_Inst_ff_SDE_0_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_0_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_0_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_0_MUX_inst_Y), .B(RoundOutput[0]), .Z(
        RoundReg_Inst_ff_SDE_0_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_0_current_state_reg_U1 ( .A(state_shifted[8]), 
        .ZN(RoundReg_Inst_ff_SDE_0_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_0_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_0_next_state), .CK(clk), .Q(state_shifted[8]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_1_MUX_inst_XOR1_U1 ( .A(RoundOutput[1]), .B(
        port_in[1]), .Z(RoundReg_Inst_ff_SDE_1_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_1_MUX_inst_AND1_U1 ( .A1(RoundReg_n7), .A2(
        RoundReg_Inst_ff_SDE_1_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_1_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_1_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_1_MUX_inst_Y), .B(RoundOutput[1]), .Z(
        RoundReg_Inst_ff_SDE_1_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_1_current_state_reg_U1 ( .A(state_shifted[9]), 
        .ZN(RoundReg_Inst_ff_SDE_1_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_1_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_1_next_state), .CK(clk), .Q(state_shifted[9]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_2_MUX_inst_XOR1_U1 ( .A(RoundOutput[2]), .B(
        port_in[2]), .Z(RoundReg_Inst_ff_SDE_2_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_2_MUX_inst_AND1_U1 ( .A1(RoundReg_n8), .A2(
        RoundReg_Inst_ff_SDE_2_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_2_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_2_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_2_MUX_inst_Y), .B(RoundOutput[2]), .Z(
        RoundReg_Inst_ff_SDE_2_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_2_current_state_reg_U1 ( .A(state_shifted[10]), 
        .ZN(RoundReg_Inst_ff_SDE_2_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_2_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_2_next_state), .CK(clk), .Q(state_shifted[10]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_3_MUX_inst_XOR1_U1 ( .A(RoundOutput[3]), .B(
        port_in[3]), .Z(RoundReg_Inst_ff_SDE_3_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_3_MUX_inst_AND1_U1 ( .A1(RoundReg_n9), .A2(
        RoundReg_Inst_ff_SDE_3_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_3_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_3_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_3_MUX_inst_Y), .B(RoundOutput[3]), .Z(
        RoundReg_Inst_ff_SDE_3_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_3_current_state_reg_U1 ( .A(state_shifted[11]), 
        .ZN(RoundReg_Inst_ff_SDE_3_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_3_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_3_next_state), .CK(clk), .Q(state_shifted[11]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_4_MUX_inst_XOR1_U1 ( .A(RoundOutput[4]), .B(
        port_in[4]), .Z(RoundReg_Inst_ff_SDE_4_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_4_MUX_inst_AND1_U1 ( .A1(RoundReg_n7), .A2(
        RoundReg_Inst_ff_SDE_4_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_4_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_4_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_4_MUX_inst_Y), .B(RoundOutput[4]), .Z(
        RoundReg_Inst_ff_SDE_4_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_4_current_state_reg_U1 ( .A(state_shifted[12]), 
        .ZN(RoundReg_Inst_ff_SDE_4_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_4_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_4_next_state), .CK(clk), .Q(state_shifted[12]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_5_MUX_inst_XOR1_U1 ( .A(RoundOutput[5]), .B(
        port_in[5]), .Z(RoundReg_Inst_ff_SDE_5_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_5_MUX_inst_AND1_U1 ( .A1(RoundReg_n6), .A2(
        RoundReg_Inst_ff_SDE_5_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_5_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_5_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_5_MUX_inst_Y), .B(RoundOutput[5]), .Z(
        RoundReg_Inst_ff_SDE_5_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_5_current_state_reg_U1 ( .A(state_shifted[13]), 
        .ZN(RoundReg_Inst_ff_SDE_5_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_5_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_5_next_state), .CK(clk), .Q(state_shifted[13]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_6_MUX_inst_XOR1_U1 ( .A(RoundOutput[6]), .B(
        port_in[6]), .Z(RoundReg_Inst_ff_SDE_6_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_6_MUX_inst_AND1_U1 ( .A1(RoundReg_n7), .A2(
        RoundReg_Inst_ff_SDE_6_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_6_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_6_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_6_MUX_inst_Y), .B(RoundOutput[6]), .Z(
        RoundReg_Inst_ff_SDE_6_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_6_current_state_reg_U1 ( .A(state_shifted[14]), 
        .ZN(RoundReg_Inst_ff_SDE_6_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_6_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_6_next_state), .CK(clk), .Q(state_shifted[14]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_7_MUX_inst_XOR1_U1 ( .A(RoundOutput[7]), .B(
        port_in[7]), .Z(RoundReg_Inst_ff_SDE_7_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_7_MUX_inst_AND1_U1 ( .A1(start_done), .A2(
        RoundReg_Inst_ff_SDE_7_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_7_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_7_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_7_MUX_inst_Y), .B(RoundOutput[7]), .Z(
        RoundReg_Inst_ff_SDE_7_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_7_current_state_reg_U1 ( .A(state_shifted[15]), 
        .ZN(RoundReg_Inst_ff_SDE_7_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_7_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_7_next_state), .CK(clk), .Q(state_shifted[15]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_8_MUX_inst_XOR1_U1 ( .A(RoundOutput[8]), .B(
        state_shifted[8]), .Z(RoundReg_Inst_ff_SDE_8_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_8_MUX_inst_AND1_U1 ( .A1(RoundReg_n6), .A2(
        RoundReg_Inst_ff_SDE_8_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_8_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_8_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_8_MUX_inst_Y), .B(RoundOutput[8]), .Z(
        RoundReg_Inst_ff_SDE_8_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_8_current_state_reg_U1 ( .A(state_shifted[16]), 
        .ZN(RoundReg_Inst_ff_SDE_8_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_8_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_8_next_state), .CK(clk), .Q(state_shifted[16]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_9_MUX_inst_XOR1_U1 ( .A(RoundOutput[9]), .B(
        state_shifted[9]), .Z(RoundReg_Inst_ff_SDE_9_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_9_MUX_inst_AND1_U1 ( .A1(start_done), .A2(
        RoundReg_Inst_ff_SDE_9_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_9_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_9_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_9_MUX_inst_Y), .B(RoundOutput[9]), .Z(
        RoundReg_Inst_ff_SDE_9_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_9_current_state_reg_U1 ( .A(state_shifted[17]), 
        .ZN(RoundReg_Inst_ff_SDE_9_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_9_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_9_next_state), .CK(clk), .Q(state_shifted[17]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_10_MUX_inst_XOR1_U1 ( .A(RoundOutput[10]), .B(
        state_shifted[10]), .Z(RoundReg_Inst_ff_SDE_10_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_10_MUX_inst_AND1_U1 ( .A1(start_done), .A2(
        RoundReg_Inst_ff_SDE_10_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_10_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_10_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_10_MUX_inst_Y), .B(RoundOutput[10]), .Z(
        RoundReg_Inst_ff_SDE_10_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_10_current_state_reg_U1 ( .A(state_shifted[18]), 
        .ZN(RoundReg_Inst_ff_SDE_10_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_10_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_10_next_state), .CK(clk), .Q(state_shifted[18]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_11_MUX_inst_XOR1_U1 ( .A(RoundOutput[11]), .B(
        state_shifted[11]), .Z(RoundReg_Inst_ff_SDE_11_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_11_MUX_inst_AND1_U1 ( .A1(start_done), .A2(
        RoundReg_Inst_ff_SDE_11_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_11_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_11_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_11_MUX_inst_Y), .B(RoundOutput[11]), .Z(
        RoundReg_Inst_ff_SDE_11_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_11_current_state_reg_U1 ( .A(state_shifted[19]), 
        .ZN(RoundReg_Inst_ff_SDE_11_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_11_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_11_next_state), .CK(clk), .Q(state_shifted[19]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_12_MUX_inst_XOR1_U1 ( .A(RoundOutput[12]), .B(
        state_shifted[12]), .Z(RoundReg_Inst_ff_SDE_12_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_12_MUX_inst_AND1_U1 ( .A1(start_done), .A2(
        RoundReg_Inst_ff_SDE_12_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_12_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_12_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_12_MUX_inst_Y), .B(RoundOutput[12]), .Z(
        RoundReg_Inst_ff_SDE_12_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_12_current_state_reg_U1 ( .A(state_shifted[20]), 
        .ZN(RoundReg_Inst_ff_SDE_12_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_12_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_12_next_state), .CK(clk), .Q(state_shifted[20]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_13_MUX_inst_XOR1_U1 ( .A(RoundOutput[13]), .B(
        state_shifted[13]), .Z(RoundReg_Inst_ff_SDE_13_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_13_MUX_inst_AND1_U1 ( .A1(start_done), .A2(
        RoundReg_Inst_ff_SDE_13_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_13_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_13_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_13_MUX_inst_Y), .B(RoundOutput[13]), .Z(
        RoundReg_Inst_ff_SDE_13_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_13_current_state_reg_U1 ( .A(state_shifted[21]), 
        .ZN(RoundReg_Inst_ff_SDE_13_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_13_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_13_next_state), .CK(clk), .Q(state_shifted[21]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_14_MUX_inst_XOR1_U1 ( .A(RoundOutput[14]), .B(
        state_shifted[14]), .Z(RoundReg_Inst_ff_SDE_14_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_14_MUX_inst_AND1_U1 ( .A1(start_done), .A2(
        RoundReg_Inst_ff_SDE_14_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_14_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_14_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_14_MUX_inst_Y), .B(RoundOutput[14]), .Z(
        RoundReg_Inst_ff_SDE_14_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_14_current_state_reg_U1 ( .A(state_shifted[22]), 
        .ZN(RoundReg_Inst_ff_SDE_14_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_14_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_14_next_state), .CK(clk), .Q(state_shifted[22]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_15_MUX_inst_XOR1_U1 ( .A(RoundOutput[15]), .B(
        state_shifted[15]), .Z(RoundReg_Inst_ff_SDE_15_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_15_MUX_inst_AND1_U1 ( .A1(start_done), .A2(
        RoundReg_Inst_ff_SDE_15_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_15_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_15_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_15_MUX_inst_Y), .B(RoundOutput[15]), .Z(
        RoundReg_Inst_ff_SDE_15_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_15_current_state_reg_U1 ( .A(state_shifted[23]), 
        .ZN(RoundReg_Inst_ff_SDE_15_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_15_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_15_next_state), .CK(clk), .Q(state_shifted[23]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_16_MUX_inst_XOR1_U1 ( .A(RoundOutput[16]), .B(
        state_shifted[16]), .Z(RoundReg_Inst_ff_SDE_16_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_16_MUX_inst_AND1_U1 ( .A1(start_done), .A2(
        RoundReg_Inst_ff_SDE_16_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_16_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_16_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_16_MUX_inst_Y), .B(RoundOutput[16]), .Z(
        RoundReg_Inst_ff_SDE_16_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_16_current_state_reg_U1 ( .A(state_shifted[24]), 
        .ZN(RoundReg_Inst_ff_SDE_16_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_16_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_16_next_state), .CK(clk), .Q(state_shifted[24]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_17_MUX_inst_XOR1_U1 ( .A(RoundOutput[17]), .B(
        state_shifted[17]), .Z(RoundReg_Inst_ff_SDE_17_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_17_MUX_inst_AND1_U1 ( .A1(start_done), .A2(
        RoundReg_Inst_ff_SDE_17_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_17_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_17_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_17_MUX_inst_Y), .B(RoundOutput[17]), .Z(
        RoundReg_Inst_ff_SDE_17_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_17_current_state_reg_U1 ( .A(state_shifted[25]), 
        .ZN(RoundReg_Inst_ff_SDE_17_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_17_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_17_next_state), .CK(clk), .Q(state_shifted[25]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_18_MUX_inst_XOR1_U1 ( .A(RoundOutput[18]), .B(
        state_shifted[18]), .Z(RoundReg_Inst_ff_SDE_18_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_18_MUX_inst_AND1_U1 ( .A1(start_done), .A2(
        RoundReg_Inst_ff_SDE_18_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_18_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_18_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_18_MUX_inst_Y), .B(RoundOutput[18]), .Z(
        RoundReg_Inst_ff_SDE_18_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_18_current_state_reg_U1 ( .A(state_shifted[26]), 
        .ZN(RoundReg_Inst_ff_SDE_18_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_18_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_18_next_state), .CK(clk), .Q(state_shifted[26]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_19_MUX_inst_XOR1_U1 ( .A(RoundOutput[19]), .B(
        state_shifted[19]), .Z(RoundReg_Inst_ff_SDE_19_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_19_MUX_inst_AND1_U1 ( .A1(start_done), .A2(
        RoundReg_Inst_ff_SDE_19_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_19_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_19_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_19_MUX_inst_Y), .B(RoundOutput[19]), .Z(
        RoundReg_Inst_ff_SDE_19_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_19_current_state_reg_U1 ( .A(state_shifted[27]), 
        .ZN(RoundReg_Inst_ff_SDE_19_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_19_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_19_next_state), .CK(clk), .Q(state_shifted[27]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_20_MUX_inst_XOR1_U1 ( .A(RoundOutput[20]), .B(
        state_shifted[20]), .Z(RoundReg_Inst_ff_SDE_20_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_20_MUX_inst_AND1_U1 ( .A1(RoundReg_n7), .A2(
        RoundReg_Inst_ff_SDE_20_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_20_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_20_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_20_MUX_inst_Y), .B(RoundOutput[20]), .Z(
        RoundReg_Inst_ff_SDE_20_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_20_current_state_reg_U1 ( .A(state_shifted[28]), 
        .ZN(RoundReg_Inst_ff_SDE_20_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_20_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_20_next_state), .CK(clk), .Q(state_shifted[28]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_21_MUX_inst_XOR1_U1 ( .A(RoundOutput[21]), .B(
        state_shifted[21]), .Z(RoundReg_Inst_ff_SDE_21_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_21_MUX_inst_AND1_U1 ( .A1(RoundReg_n8), .A2(
        RoundReg_Inst_ff_SDE_21_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_21_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_21_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_21_MUX_inst_Y), .B(RoundOutput[21]), .Z(
        RoundReg_Inst_ff_SDE_21_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_21_current_state_reg_U1 ( .A(state_shifted[29]), 
        .ZN(RoundReg_Inst_ff_SDE_21_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_21_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_21_next_state), .CK(clk), .Q(state_shifted[29]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_22_MUX_inst_XOR1_U1 ( .A(RoundOutput[22]), .B(
        state_shifted[22]), .Z(RoundReg_Inst_ff_SDE_22_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_22_MUX_inst_AND1_U1 ( .A1(RoundReg_n9), .A2(
        RoundReg_Inst_ff_SDE_22_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_22_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_22_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_22_MUX_inst_Y), .B(RoundOutput[22]), .Z(
        RoundReg_Inst_ff_SDE_22_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_22_current_state_reg_U1 ( .A(state_shifted[30]), 
        .ZN(RoundReg_Inst_ff_SDE_22_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_22_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_22_next_state), .CK(clk), .Q(state_shifted[30]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_23_MUX_inst_XOR1_U1 ( .A(RoundOutput[23]), .B(
        state_shifted[23]), .Z(RoundReg_Inst_ff_SDE_23_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_23_MUX_inst_AND1_U1 ( .A1(RoundReg_n8), .A2(
        RoundReg_Inst_ff_SDE_23_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_23_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_23_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_23_MUX_inst_Y), .B(RoundOutput[23]), .Z(
        RoundReg_Inst_ff_SDE_23_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_23_current_state_reg_U1 ( .A(state_shifted[31]), 
        .ZN(RoundReg_Inst_ff_SDE_23_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_23_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_23_next_state), .CK(clk), .Q(state_shifted[31]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_24_MUX_inst_XOR1_U1 ( .A(RoundOutput[24]), .B(
        state_shifted[24]), .Z(RoundReg_Inst_ff_SDE_24_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_24_MUX_inst_AND1_U1 ( .A1(RoundReg_n6), .A2(
        RoundReg_Inst_ff_SDE_24_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_24_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_24_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_24_MUX_inst_Y), .B(RoundOutput[24]), .Z(
        RoundReg_Inst_ff_SDE_24_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_24_current_state_reg_U1 ( .A(state_shifted[32]), 
        .ZN(RoundReg_Inst_ff_SDE_24_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_24_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_24_next_state), .CK(clk), .Q(state_shifted[32]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_25_MUX_inst_XOR1_U1 ( .A(RoundOutput[25]), .B(
        state_shifted[25]), .Z(RoundReg_Inst_ff_SDE_25_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_25_MUX_inst_AND1_U1 ( .A1(RoundReg_n7), .A2(
        RoundReg_Inst_ff_SDE_25_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_25_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_25_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_25_MUX_inst_Y), .B(RoundOutput[25]), .Z(
        RoundReg_Inst_ff_SDE_25_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_25_current_state_reg_U1 ( .A(state_shifted[33]), 
        .ZN(RoundReg_Inst_ff_SDE_25_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_25_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_25_next_state), .CK(clk), .Q(state_shifted[33]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_26_MUX_inst_XOR1_U1 ( .A(RoundOutput[26]), .B(
        state_shifted[26]), .Z(RoundReg_Inst_ff_SDE_26_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_26_MUX_inst_AND1_U1 ( .A1(RoundReg_n7), .A2(
        RoundReg_Inst_ff_SDE_26_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_26_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_26_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_26_MUX_inst_Y), .B(RoundOutput[26]), .Z(
        RoundReg_Inst_ff_SDE_26_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_26_current_state_reg_U1 ( .A(state_shifted[34]), 
        .ZN(RoundReg_Inst_ff_SDE_26_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_26_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_26_next_state), .CK(clk), .Q(state_shifted[34]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_27_MUX_inst_XOR1_U1 ( .A(RoundOutput[27]), .B(
        state_shifted[27]), .Z(RoundReg_Inst_ff_SDE_27_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_27_MUX_inst_AND1_U1 ( .A1(start_done), .A2(
        RoundReg_Inst_ff_SDE_27_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_27_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_27_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_27_MUX_inst_Y), .B(RoundOutput[27]), .Z(
        RoundReg_Inst_ff_SDE_27_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_27_current_state_reg_U1 ( .A(state_shifted[35]), 
        .ZN(RoundReg_Inst_ff_SDE_27_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_27_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_27_next_state), .CK(clk), .Q(state_shifted[35]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_28_MUX_inst_XOR1_U1 ( .A(RoundOutput[28]), .B(
        state_shifted[28]), .Z(RoundReg_Inst_ff_SDE_28_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_28_MUX_inst_AND1_U1 ( .A1(start_done), .A2(
        RoundReg_Inst_ff_SDE_28_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_28_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_28_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_28_MUX_inst_Y), .B(RoundOutput[28]), .Z(
        RoundReg_Inst_ff_SDE_28_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_28_current_state_reg_U1 ( .A(state_shifted[36]), 
        .ZN(RoundReg_Inst_ff_SDE_28_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_28_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_28_next_state), .CK(clk), .Q(state_shifted[36]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_29_MUX_inst_XOR1_U1 ( .A(RoundOutput[29]), .B(
        state_shifted[29]), .Z(RoundReg_Inst_ff_SDE_29_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_29_MUX_inst_AND1_U1 ( .A1(start_done), .A2(
        RoundReg_Inst_ff_SDE_29_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_29_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_29_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_29_MUX_inst_Y), .B(RoundOutput[29]), .Z(
        RoundReg_Inst_ff_SDE_29_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_29_current_state_reg_U1 ( .A(state_shifted[37]), 
        .ZN(RoundReg_Inst_ff_SDE_29_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_29_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_29_next_state), .CK(clk), .Q(state_shifted[37]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_30_MUX_inst_XOR1_U1 ( .A(RoundOutput[30]), .B(
        state_shifted[30]), .Z(RoundReg_Inst_ff_SDE_30_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_30_MUX_inst_AND1_U1 ( .A1(start_done), .A2(
        RoundReg_Inst_ff_SDE_30_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_30_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_30_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_30_MUX_inst_Y), .B(RoundOutput[30]), .Z(
        RoundReg_Inst_ff_SDE_30_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_30_current_state_reg_U1 ( .A(state_shifted[38]), 
        .ZN(RoundReg_Inst_ff_SDE_30_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_30_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_30_next_state), .CK(clk), .Q(state_shifted[38]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_31_MUX_inst_XOR1_U1 ( .A(RoundOutput[31]), .B(
        state_shifted[31]), .Z(RoundReg_Inst_ff_SDE_31_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_31_MUX_inst_AND1_U1 ( .A1(start_done), .A2(
        RoundReg_Inst_ff_SDE_31_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_31_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_31_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_31_MUX_inst_Y), .B(RoundOutput[31]), .Z(
        RoundReg_Inst_ff_SDE_31_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_31_current_state_reg_U1 ( .A(state_shifted[39]), 
        .ZN(RoundReg_Inst_ff_SDE_31_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_31_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_31_next_state), .CK(clk), .Q(state_shifted[39]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_32_MUX_inst_XOR1_U1 ( .A(RoundOutput[32]), .B(
        state_shifted[32]), .Z(RoundReg_Inst_ff_SDE_32_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_32_MUX_inst_AND1_U1 ( .A1(RoundReg_n8), .A2(
        RoundReg_Inst_ff_SDE_32_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_32_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_32_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_32_MUX_inst_Y), .B(RoundOutput[32]), .Z(
        RoundReg_Inst_ff_SDE_32_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_32_current_state_reg_U1 ( .A(state_shifted[40]), 
        .ZN(RoundReg_Inst_ff_SDE_32_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_32_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_32_next_state), .CK(clk), .Q(state_shifted[40]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_33_MUX_inst_XOR1_U1 ( .A(RoundOutput[33]), .B(
        state_shifted[33]), .Z(RoundReg_Inst_ff_SDE_33_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_33_MUX_inst_AND1_U1 ( .A1(RoundReg_n9), .A2(
        RoundReg_Inst_ff_SDE_33_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_33_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_33_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_33_MUX_inst_Y), .B(RoundOutput[33]), .Z(
        RoundReg_Inst_ff_SDE_33_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_33_current_state_reg_U1 ( .A(state_shifted[41]), 
        .ZN(RoundReg_Inst_ff_SDE_33_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_33_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_33_next_state), .CK(clk), .Q(state_shifted[41]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_34_MUX_inst_XOR1_U1 ( .A(RoundOutput[34]), .B(
        state_shifted[34]), .Z(RoundReg_Inst_ff_SDE_34_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_34_MUX_inst_AND1_U1 ( .A1(RoundReg_n9), .A2(
        RoundReg_Inst_ff_SDE_34_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_34_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_34_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_34_MUX_inst_Y), .B(RoundOutput[34]), .Z(
        RoundReg_Inst_ff_SDE_34_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_34_current_state_reg_U1 ( .A(state_shifted[42]), 
        .ZN(RoundReg_Inst_ff_SDE_34_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_34_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_34_next_state), .CK(clk), .Q(state_shifted[42]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_35_MUX_inst_XOR1_U1 ( .A(RoundOutput[35]), .B(
        state_shifted[35]), .Z(RoundReg_Inst_ff_SDE_35_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_35_MUX_inst_AND1_U1 ( .A1(RoundReg_n7), .A2(
        RoundReg_Inst_ff_SDE_35_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_35_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_35_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_35_MUX_inst_Y), .B(RoundOutput[35]), .Z(
        RoundReg_Inst_ff_SDE_35_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_35_current_state_reg_U1 ( .A(state_shifted[43]), 
        .ZN(RoundReg_Inst_ff_SDE_35_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_35_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_35_next_state), .CK(clk), .Q(state_shifted[43]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_36_MUX_inst_XOR1_U1 ( .A(RoundOutput[36]), .B(
        state_shifted[36]), .Z(RoundReg_Inst_ff_SDE_36_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_36_MUX_inst_AND1_U1 ( .A1(RoundReg_n8), .A2(
        RoundReg_Inst_ff_SDE_36_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_36_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_36_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_36_MUX_inst_Y), .B(RoundOutput[36]), .Z(
        RoundReg_Inst_ff_SDE_36_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_36_current_state_reg_U1 ( .A(state_shifted[44]), 
        .ZN(RoundReg_Inst_ff_SDE_36_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_36_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_36_next_state), .CK(clk), .Q(state_shifted[44]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_37_MUX_inst_XOR1_U1 ( .A(RoundOutput[37]), .B(
        state_shifted[37]), .Z(RoundReg_Inst_ff_SDE_37_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_37_MUX_inst_AND1_U1 ( .A1(RoundReg_n6), .A2(
        RoundReg_Inst_ff_SDE_37_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_37_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_37_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_37_MUX_inst_Y), .B(RoundOutput[37]), .Z(
        RoundReg_Inst_ff_SDE_37_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_37_current_state_reg_U1 ( .A(state_shifted[45]), 
        .ZN(RoundReg_Inst_ff_SDE_37_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_37_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_37_next_state), .CK(clk), .Q(state_shifted[45]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_38_MUX_inst_XOR1_U1 ( .A(RoundOutput[38]), .B(
        state_shifted[38]), .Z(RoundReg_Inst_ff_SDE_38_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_38_MUX_inst_AND1_U1 ( .A1(start_done), .A2(
        RoundReg_Inst_ff_SDE_38_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_38_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_38_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_38_MUX_inst_Y), .B(RoundOutput[38]), .Z(
        RoundReg_Inst_ff_SDE_38_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_38_current_state_reg_U1 ( .A(state_shifted[46]), 
        .ZN(RoundReg_Inst_ff_SDE_38_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_38_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_38_next_state), .CK(clk), .Q(state_shifted[46]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_39_MUX_inst_XOR1_U1 ( .A(RoundOutput[39]), .B(
        state_shifted[39]), .Z(RoundReg_Inst_ff_SDE_39_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_39_MUX_inst_AND1_U1 ( .A1(start_done), .A2(
        RoundReg_Inst_ff_SDE_39_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_39_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_39_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_39_MUX_inst_Y), .B(RoundOutput[39]), .Z(
        RoundReg_Inst_ff_SDE_39_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_39_current_state_reg_U1 ( .A(state_shifted[47]), 
        .ZN(RoundReg_Inst_ff_SDE_39_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_39_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_39_next_state), .CK(clk), .Q(state_shifted[47]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_40_MUX_inst_XOR1_U1 ( .A(RoundOutput[40]), .B(
        state_shifted[40]), .Z(RoundReg_Inst_ff_SDE_40_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_40_MUX_inst_AND1_U1 ( .A1(start_done), .A2(
        RoundReg_Inst_ff_SDE_40_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_40_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_40_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_40_MUX_inst_Y), .B(RoundOutput[40]), .Z(
        RoundReg_Inst_ff_SDE_40_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_40_current_state_reg_U1 ( .A(state_shifted[48]), 
        .ZN(RoundReg_Inst_ff_SDE_40_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_40_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_40_next_state), .CK(clk), .Q(state_shifted[48]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_41_MUX_inst_XOR1_U1 ( .A(RoundOutput[41]), .B(
        state_shifted[41]), .Z(RoundReg_Inst_ff_SDE_41_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_41_MUX_inst_AND1_U1 ( .A1(start_done), .A2(
        RoundReg_Inst_ff_SDE_41_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_41_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_41_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_41_MUX_inst_Y), .B(RoundOutput[41]), .Z(
        RoundReg_Inst_ff_SDE_41_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_41_current_state_reg_U1 ( .A(state_shifted[49]), 
        .ZN(RoundReg_Inst_ff_SDE_41_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_41_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_41_next_state), .CK(clk), .Q(state_shifted[49]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_42_MUX_inst_XOR1_U1 ( .A(RoundOutput[42]), .B(
        state_shifted[42]), .Z(RoundReg_Inst_ff_SDE_42_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_42_MUX_inst_AND1_U1 ( .A1(start_done), .A2(
        RoundReg_Inst_ff_SDE_42_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_42_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_42_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_42_MUX_inst_Y), .B(RoundOutput[42]), .Z(
        RoundReg_Inst_ff_SDE_42_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_42_current_state_reg_U1 ( .A(state_shifted[50]), 
        .ZN(RoundReg_Inst_ff_SDE_42_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_42_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_42_next_state), .CK(clk), .Q(state_shifted[50]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_43_MUX_inst_XOR1_U1 ( .A(RoundOutput[43]), .B(
        state_shifted[43]), .Z(RoundReg_Inst_ff_SDE_43_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_43_MUX_inst_AND1_U1 ( .A1(start_done), .A2(
        RoundReg_Inst_ff_SDE_43_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_43_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_43_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_43_MUX_inst_Y), .B(RoundOutput[43]), .Z(
        RoundReg_Inst_ff_SDE_43_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_43_current_state_reg_U1 ( .A(state_shifted[51]), 
        .ZN(RoundReg_Inst_ff_SDE_43_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_43_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_43_next_state), .CK(clk), .Q(state_shifted[51]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_44_MUX_inst_XOR1_U1 ( .A(RoundOutput[44]), .B(
        state_shifted[44]), .Z(RoundReg_Inst_ff_SDE_44_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_44_MUX_inst_AND1_U1 ( .A1(RoundReg_n9), .A2(
        RoundReg_Inst_ff_SDE_44_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_44_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_44_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_44_MUX_inst_Y), .B(RoundOutput[44]), .Z(
        RoundReg_Inst_ff_SDE_44_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_44_current_state_reg_U1 ( .A(state_shifted[52]), 
        .ZN(RoundReg_Inst_ff_SDE_44_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_44_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_44_next_state), .CK(clk), .Q(state_shifted[52]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_45_MUX_inst_XOR1_U1 ( .A(RoundOutput[45]), .B(
        state_shifted[45]), .Z(RoundReg_Inst_ff_SDE_45_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_45_MUX_inst_AND1_U1 ( .A1(RoundReg_n6), .A2(
        RoundReg_Inst_ff_SDE_45_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_45_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_45_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_45_MUX_inst_Y), .B(RoundOutput[45]), .Z(
        RoundReg_Inst_ff_SDE_45_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_45_current_state_reg_U1 ( .A(state_shifted[53]), 
        .ZN(RoundReg_Inst_ff_SDE_45_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_45_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_45_next_state), .CK(clk), .Q(state_shifted[53]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_46_MUX_inst_XOR1_U1 ( .A(RoundOutput[46]), .B(
        state_shifted[46]), .Z(RoundReg_Inst_ff_SDE_46_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_46_MUX_inst_AND1_U1 ( .A1(RoundReg_n8), .A2(
        RoundReg_Inst_ff_SDE_46_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_46_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_46_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_46_MUX_inst_Y), .B(RoundOutput[46]), .Z(
        RoundReg_Inst_ff_SDE_46_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_46_current_state_reg_U1 ( .A(state_shifted[54]), 
        .ZN(RoundReg_Inst_ff_SDE_46_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_46_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_46_next_state), .CK(clk), .Q(state_shifted[54]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_47_MUX_inst_XOR1_U1 ( .A(RoundOutput[47]), .B(
        state_shifted[47]), .Z(RoundReg_Inst_ff_SDE_47_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_47_MUX_inst_AND1_U1 ( .A1(RoundReg_n6), .A2(
        RoundReg_Inst_ff_SDE_47_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_47_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_47_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_47_MUX_inst_Y), .B(RoundOutput[47]), .Z(
        RoundReg_Inst_ff_SDE_47_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_47_current_state_reg_U1 ( .A(state_shifted[55]), 
        .ZN(RoundReg_Inst_ff_SDE_47_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_47_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_47_next_state), .CK(clk), .Q(state_shifted[55]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_48_MUX_inst_XOR1_U1 ( .A(RoundOutput[48]), .B(
        state_shifted[48]), .Z(RoundReg_Inst_ff_SDE_48_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_48_MUX_inst_AND1_U1 ( .A1(start_done), .A2(
        RoundReg_Inst_ff_SDE_48_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_48_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_48_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_48_MUX_inst_Y), .B(RoundOutput[48]), .Z(
        RoundReg_Inst_ff_SDE_48_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_48_current_state_reg_U1 ( .A(state_shifted[56]), 
        .ZN(RoundReg_Inst_ff_SDE_48_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_48_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_48_next_state), .CK(clk), .Q(state_shifted[56]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_49_MUX_inst_XOR1_U1 ( .A(RoundOutput[49]), .B(
        state_shifted[49]), .Z(RoundReg_Inst_ff_SDE_49_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_49_MUX_inst_AND1_U1 ( .A1(start_done), .A2(
        RoundReg_Inst_ff_SDE_49_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_49_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_49_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_49_MUX_inst_Y), .B(RoundOutput[49]), .Z(
        RoundReg_Inst_ff_SDE_49_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_49_current_state_reg_U1 ( .A(state_shifted[57]), 
        .ZN(RoundReg_Inst_ff_SDE_49_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_49_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_49_next_state), .CK(clk), .Q(state_shifted[57]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_50_MUX_inst_XOR1_U1 ( .A(RoundOutput[50]), .B(
        state_shifted[50]), .Z(RoundReg_Inst_ff_SDE_50_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_50_MUX_inst_AND1_U1 ( .A1(start_done), .A2(
        RoundReg_Inst_ff_SDE_50_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_50_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_50_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_50_MUX_inst_Y), .B(RoundOutput[50]), .Z(
        RoundReg_Inst_ff_SDE_50_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_50_current_state_reg_U1 ( .A(state_shifted[58]), 
        .ZN(RoundReg_Inst_ff_SDE_50_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_50_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_50_next_state), .CK(clk), .Q(state_shifted[58]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_51_MUX_inst_XOR1_U1 ( .A(RoundOutput[51]), .B(
        state_shifted[51]), .Z(RoundReg_Inst_ff_SDE_51_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_51_MUX_inst_AND1_U1 ( .A1(start_done), .A2(
        RoundReg_Inst_ff_SDE_51_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_51_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_51_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_51_MUX_inst_Y), .B(RoundOutput[51]), .Z(
        RoundReg_Inst_ff_SDE_51_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_51_current_state_reg_U1 ( .A(state_shifted[59]), 
        .ZN(RoundReg_Inst_ff_SDE_51_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_51_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_51_next_state), .CK(clk), .Q(state_shifted[59]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_52_MUX_inst_XOR1_U1 ( .A(RoundOutput[52]), .B(
        state_shifted[52]), .Z(RoundReg_Inst_ff_SDE_52_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_52_MUX_inst_AND1_U1 ( .A1(RoundReg_n7), .A2(
        RoundReg_Inst_ff_SDE_52_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_52_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_52_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_52_MUX_inst_Y), .B(RoundOutput[52]), .Z(
        RoundReg_Inst_ff_SDE_52_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_52_current_state_reg_U1 ( .A(state_shifted[60]), 
        .ZN(RoundReg_Inst_ff_SDE_52_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_52_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_52_next_state), .CK(clk), .Q(state_shifted[60]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_53_MUX_inst_XOR1_U1 ( .A(RoundOutput[53]), .B(
        state_shifted[53]), .Z(RoundReg_Inst_ff_SDE_53_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_53_MUX_inst_AND1_U1 ( .A1(RoundReg_n8), .A2(
        RoundReg_Inst_ff_SDE_53_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_53_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_53_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_53_MUX_inst_Y), .B(RoundOutput[53]), .Z(
        RoundReg_Inst_ff_SDE_53_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_53_current_state_reg_U1 ( .A(state_shifted[61]), 
        .ZN(RoundReg_Inst_ff_SDE_53_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_53_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_53_next_state), .CK(clk), .Q(state_shifted[61]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_54_MUX_inst_XOR1_U1 ( .A(RoundOutput[54]), .B(
        state_shifted[54]), .Z(RoundReg_Inst_ff_SDE_54_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_54_MUX_inst_AND1_U1 ( .A1(RoundReg_n9), .A2(
        RoundReg_Inst_ff_SDE_54_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_54_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_54_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_54_MUX_inst_Y), .B(RoundOutput[54]), .Z(
        RoundReg_Inst_ff_SDE_54_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_54_current_state_reg_U1 ( .A(state_shifted[62]), 
        .ZN(RoundReg_Inst_ff_SDE_54_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_54_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_54_next_state), .CK(clk), .Q(state_shifted[62]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_55_MUX_inst_XOR1_U1 ( .A(RoundOutput[55]), .B(
        state_shifted[55]), .Z(RoundReg_Inst_ff_SDE_55_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_55_MUX_inst_AND1_U1 ( .A1(RoundReg_n7), .A2(
        RoundReg_Inst_ff_SDE_55_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_55_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_55_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_55_MUX_inst_Y), .B(RoundOutput[55]), .Z(
        RoundReg_Inst_ff_SDE_55_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_55_current_state_reg_U1 ( .A(state_shifted[63]), 
        .ZN(RoundReg_Inst_ff_SDE_55_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_55_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_55_next_state), .CK(clk), .Q(state_shifted[63]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_56_MUX_inst_XOR1_U1 ( .A(RoundOutput[56]), .B(
        state_shifted[56]), .Z(RoundReg_Inst_ff_SDE_56_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_56_MUX_inst_AND1_U1 ( .A1(RoundReg_n9), .A2(
        RoundReg_Inst_ff_SDE_56_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_56_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_56_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_56_MUX_inst_Y), .B(RoundOutput[56]), .Z(
        RoundReg_Inst_ff_SDE_56_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_56_current_state_reg_U1 ( .A(state_shifted[64]), 
        .ZN(RoundReg_Inst_ff_SDE_56_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_56_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_56_next_state), .CK(clk), .Q(state_shifted[64]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_57_MUX_inst_XOR1_U1 ( .A(RoundOutput[57]), .B(
        state_shifted[57]), .Z(RoundReg_Inst_ff_SDE_57_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_57_MUX_inst_AND1_U1 ( .A1(RoundReg_n8), .A2(
        RoundReg_Inst_ff_SDE_57_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_57_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_57_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_57_MUX_inst_Y), .B(RoundOutput[57]), .Z(
        RoundReg_Inst_ff_SDE_57_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_57_current_state_reg_U1 ( .A(state_shifted[65]), 
        .ZN(RoundReg_Inst_ff_SDE_57_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_57_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_57_next_state), .CK(clk), .Q(state_shifted[65]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_58_MUX_inst_XOR1_U1 ( .A(RoundOutput[58]), .B(
        state_shifted[58]), .Z(RoundReg_Inst_ff_SDE_58_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_58_MUX_inst_AND1_U1 ( .A1(RoundReg_n6), .A2(
        RoundReg_Inst_ff_SDE_58_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_58_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_58_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_58_MUX_inst_Y), .B(RoundOutput[58]), .Z(
        RoundReg_Inst_ff_SDE_58_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_58_current_state_reg_U1 ( .A(state_shifted[66]), 
        .ZN(RoundReg_Inst_ff_SDE_58_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_58_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_58_next_state), .CK(clk), .Q(state_shifted[66]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_59_MUX_inst_XOR1_U1 ( .A(RoundOutput[59]), .B(
        state_shifted[59]), .Z(RoundReg_Inst_ff_SDE_59_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_59_MUX_inst_AND1_U1 ( .A1(RoundReg_n7), .A2(
        RoundReg_Inst_ff_SDE_59_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_59_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_59_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_59_MUX_inst_Y), .B(RoundOutput[59]), .Z(
        RoundReg_Inst_ff_SDE_59_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_59_current_state_reg_U1 ( .A(state_shifted[67]), 
        .ZN(RoundReg_Inst_ff_SDE_59_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_59_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_59_next_state), .CK(clk), .Q(state_shifted[67]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_60_MUX_inst_XOR1_U1 ( .A(RoundOutput[60]), .B(
        state_shifted[60]), .Z(RoundReg_Inst_ff_SDE_60_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_60_MUX_inst_AND1_U1 ( .A1(RoundReg_n8), .A2(
        RoundReg_Inst_ff_SDE_60_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_60_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_60_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_60_MUX_inst_Y), .B(RoundOutput[60]), .Z(
        RoundReg_Inst_ff_SDE_60_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_60_current_state_reg_U1 ( .A(state_shifted[68]), 
        .ZN(RoundReg_Inst_ff_SDE_60_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_60_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_60_next_state), .CK(clk), .Q(state_shifted[68]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_61_MUX_inst_XOR1_U1 ( .A(RoundOutput[61]), .B(
        state_shifted[61]), .Z(RoundReg_Inst_ff_SDE_61_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_61_MUX_inst_AND1_U1 ( .A1(RoundReg_n9), .A2(
        RoundReg_Inst_ff_SDE_61_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_61_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_61_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_61_MUX_inst_Y), .B(RoundOutput[61]), .Z(
        RoundReg_Inst_ff_SDE_61_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_61_current_state_reg_U1 ( .A(state_shifted[69]), 
        .ZN(RoundReg_Inst_ff_SDE_61_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_61_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_61_next_state), .CK(clk), .Q(state_shifted[69]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_62_MUX_inst_XOR1_U1 ( .A(RoundOutput[62]), .B(
        state_shifted[62]), .Z(RoundReg_Inst_ff_SDE_62_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_62_MUX_inst_AND1_U1 ( .A1(RoundReg_n9), .A2(
        RoundReg_Inst_ff_SDE_62_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_62_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_62_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_62_MUX_inst_Y), .B(RoundOutput[62]), .Z(
        RoundReg_Inst_ff_SDE_62_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_62_current_state_reg_U1 ( .A(state_shifted[70]), 
        .ZN(RoundReg_Inst_ff_SDE_62_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_62_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_62_next_state), .CK(clk), .Q(state_shifted[70]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_63_MUX_inst_XOR1_U1 ( .A(RoundOutput[63]), .B(
        state_shifted[63]), .Z(RoundReg_Inst_ff_SDE_63_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_63_MUX_inst_AND1_U1 ( .A1(RoundReg_n6), .A2(
        RoundReg_Inst_ff_SDE_63_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_63_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_63_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_63_MUX_inst_Y), .B(RoundOutput[63]), .Z(
        RoundReg_Inst_ff_SDE_63_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_63_current_state_reg_U1 ( .A(state_shifted[71]), 
        .ZN(RoundReg_Inst_ff_SDE_63_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_63_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_63_next_state), .CK(clk), .Q(state_shifted[71]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_64_MUX_inst_XOR1_U1 ( .A(RoundOutput[64]), .B(
        state_shifted[64]), .Z(RoundReg_Inst_ff_SDE_64_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_64_MUX_inst_AND1_U1 ( .A1(RoundReg_n7), .A2(
        RoundReg_Inst_ff_SDE_64_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_64_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_64_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_64_MUX_inst_Y), .B(RoundOutput[64]), .Z(
        RoundReg_Inst_ff_SDE_64_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_64_current_state_reg_U1 ( .A(state_shifted[72]), 
        .ZN(RoundReg_Inst_ff_SDE_64_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_64_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_64_next_state), .CK(clk), .Q(state_shifted[72]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_65_MUX_inst_XOR1_U1 ( .A(RoundOutput[65]), .B(
        state_shifted[65]), .Z(RoundReg_Inst_ff_SDE_65_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_65_MUX_inst_AND1_U1 ( .A1(RoundReg_n8), .A2(
        RoundReg_Inst_ff_SDE_65_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_65_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_65_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_65_MUX_inst_Y), .B(RoundOutput[65]), .Z(
        RoundReg_Inst_ff_SDE_65_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_65_current_state_reg_U1 ( .A(state_shifted[73]), 
        .ZN(RoundReg_Inst_ff_SDE_65_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_65_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_65_next_state), .CK(clk), .Q(state_shifted[73]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_66_MUX_inst_XOR1_U1 ( .A(RoundOutput[66]), .B(
        state_shifted[66]), .Z(RoundReg_Inst_ff_SDE_66_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_66_MUX_inst_AND1_U1 ( .A1(RoundReg_n9), .A2(
        RoundReg_Inst_ff_SDE_66_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_66_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_66_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_66_MUX_inst_Y), .B(RoundOutput[66]), .Z(
        RoundReg_Inst_ff_SDE_66_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_66_current_state_reg_U1 ( .A(state_shifted[74]), 
        .ZN(RoundReg_Inst_ff_SDE_66_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_66_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_66_next_state), .CK(clk), .Q(state_shifted[74]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_67_MUX_inst_XOR1_U1 ( .A(RoundOutput[67]), .B(
        state_shifted[67]), .Z(RoundReg_Inst_ff_SDE_67_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_67_MUX_inst_AND1_U1 ( .A1(RoundReg_n6), .A2(
        RoundReg_Inst_ff_SDE_67_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_67_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_67_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_67_MUX_inst_Y), .B(RoundOutput[67]), .Z(
        RoundReg_Inst_ff_SDE_67_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_67_current_state_reg_U1 ( .A(state_shifted[75]), 
        .ZN(RoundReg_Inst_ff_SDE_67_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_67_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_67_next_state), .CK(clk), .Q(state_shifted[75]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_68_MUX_inst_XOR1_U1 ( .A(RoundOutput[68]), .B(
        state_shifted[68]), .Z(RoundReg_Inst_ff_SDE_68_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_68_MUX_inst_AND1_U1 ( .A1(RoundReg_n7), .A2(
        RoundReg_Inst_ff_SDE_68_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_68_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_68_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_68_MUX_inst_Y), .B(RoundOutput[68]), .Z(
        RoundReg_Inst_ff_SDE_68_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_68_current_state_reg_U1 ( .A(state_shifted[76]), 
        .ZN(RoundReg_Inst_ff_SDE_68_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_68_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_68_next_state), .CK(clk), .Q(state_shifted[76]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_69_MUX_inst_XOR1_U1 ( .A(RoundOutput[69]), .B(
        state_shifted[69]), .Z(RoundReg_Inst_ff_SDE_69_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_69_MUX_inst_AND1_U1 ( .A1(RoundReg_n8), .A2(
        RoundReg_Inst_ff_SDE_69_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_69_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_69_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_69_MUX_inst_Y), .B(RoundOutput[69]), .Z(
        RoundReg_Inst_ff_SDE_69_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_69_current_state_reg_U1 ( .A(state_shifted[77]), 
        .ZN(RoundReg_Inst_ff_SDE_69_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_69_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_69_next_state), .CK(clk), .Q(state_shifted[77]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_70_MUX_inst_XOR1_U1 ( .A(RoundOutput[70]), .B(
        state_shifted[70]), .Z(RoundReg_Inst_ff_SDE_70_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_70_MUX_inst_AND1_U1 ( .A1(RoundReg_n9), .A2(
        RoundReg_Inst_ff_SDE_70_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_70_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_70_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_70_MUX_inst_Y), .B(RoundOutput[70]), .Z(
        RoundReg_Inst_ff_SDE_70_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_70_current_state_reg_U1 ( .A(state_shifted[78]), 
        .ZN(RoundReg_Inst_ff_SDE_70_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_70_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_70_next_state), .CK(clk), .Q(state_shifted[78]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_71_MUX_inst_XOR1_U1 ( .A(RoundOutput[71]), .B(
        state_shifted[71]), .Z(RoundReg_Inst_ff_SDE_71_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_71_MUX_inst_AND1_U1 ( .A1(RoundReg_n6), .A2(
        RoundReg_Inst_ff_SDE_71_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_71_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_71_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_71_MUX_inst_Y), .B(RoundOutput[71]), .Z(
        RoundReg_Inst_ff_SDE_71_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_71_current_state_reg_U1 ( .A(state_shifted[79]), 
        .ZN(RoundReg_Inst_ff_SDE_71_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_71_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_71_next_state), .CK(clk), .Q(state_shifted[79]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_72_MUX_inst_XOR1_U1 ( .A(RoundOutput[72]), .B(
        state_shifted[72]), .Z(RoundReg_Inst_ff_SDE_72_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_72_MUX_inst_AND1_U1 ( .A1(RoundReg_n7), .A2(
        RoundReg_Inst_ff_SDE_72_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_72_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_72_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_72_MUX_inst_Y), .B(RoundOutput[72]), .Z(
        RoundReg_Inst_ff_SDE_72_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_72_current_state_reg_U1 ( .A(state_shifted[80]), 
        .ZN(RoundReg_Inst_ff_SDE_72_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_72_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_72_next_state), .CK(clk), .Q(state_shifted[80]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_73_MUX_inst_XOR1_U1 ( .A(RoundOutput[73]), .B(
        state_shifted[73]), .Z(RoundReg_Inst_ff_SDE_73_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_73_MUX_inst_AND1_U1 ( .A1(RoundReg_n8), .A2(
        RoundReg_Inst_ff_SDE_73_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_73_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_73_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_73_MUX_inst_Y), .B(RoundOutput[73]), .Z(
        RoundReg_Inst_ff_SDE_73_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_73_current_state_reg_U1 ( .A(state_shifted[81]), 
        .ZN(RoundReg_Inst_ff_SDE_73_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_73_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_73_next_state), .CK(clk), .Q(state_shifted[81]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_74_MUX_inst_XOR1_U1 ( .A(RoundOutput[74]), .B(
        state_shifted[74]), .Z(RoundReg_Inst_ff_SDE_74_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_74_MUX_inst_AND1_U1 ( .A1(RoundReg_n9), .A2(
        RoundReg_Inst_ff_SDE_74_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_74_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_74_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_74_MUX_inst_Y), .B(RoundOutput[74]), .Z(
        RoundReg_Inst_ff_SDE_74_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_74_current_state_reg_U1 ( .A(state_shifted[82]), 
        .ZN(RoundReg_Inst_ff_SDE_74_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_74_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_74_next_state), .CK(clk), .Q(state_shifted[82]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_75_MUX_inst_XOR1_U1 ( .A(RoundOutput[75]), .B(
        state_shifted[75]), .Z(RoundReg_Inst_ff_SDE_75_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_75_MUX_inst_AND1_U1 ( .A1(RoundReg_n6), .A2(
        RoundReg_Inst_ff_SDE_75_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_75_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_75_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_75_MUX_inst_Y), .B(RoundOutput[75]), .Z(
        RoundReg_Inst_ff_SDE_75_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_75_current_state_reg_U1 ( .A(state_shifted[83]), 
        .ZN(RoundReg_Inst_ff_SDE_75_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_75_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_75_next_state), .CK(clk), .Q(state_shifted[83]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_76_MUX_inst_XOR1_U1 ( .A(RoundOutput[76]), .B(
        state_shifted[76]), .Z(RoundReg_Inst_ff_SDE_76_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_76_MUX_inst_AND1_U1 ( .A1(RoundReg_n7), .A2(
        RoundReg_Inst_ff_SDE_76_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_76_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_76_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_76_MUX_inst_Y), .B(RoundOutput[76]), .Z(
        RoundReg_Inst_ff_SDE_76_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_76_current_state_reg_U1 ( .A(state_shifted[84]), 
        .ZN(RoundReg_Inst_ff_SDE_76_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_76_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_76_next_state), .CK(clk), .Q(state_shifted[84]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_77_MUX_inst_XOR1_U1 ( .A(RoundOutput[77]), .B(
        state_shifted[77]), .Z(RoundReg_Inst_ff_SDE_77_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_77_MUX_inst_AND1_U1 ( .A1(RoundReg_n8), .A2(
        RoundReg_Inst_ff_SDE_77_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_77_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_77_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_77_MUX_inst_Y), .B(RoundOutput[77]), .Z(
        RoundReg_Inst_ff_SDE_77_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_77_current_state_reg_U1 ( .A(state_shifted[85]), 
        .ZN(RoundReg_Inst_ff_SDE_77_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_77_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_77_next_state), .CK(clk), .Q(state_shifted[85]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_78_MUX_inst_XOR1_U1 ( .A(RoundOutput[78]), .B(
        state_shifted[78]), .Z(RoundReg_Inst_ff_SDE_78_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_78_MUX_inst_AND1_U1 ( .A1(RoundReg_n9), .A2(
        RoundReg_Inst_ff_SDE_78_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_78_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_78_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_78_MUX_inst_Y), .B(RoundOutput[78]), .Z(
        RoundReg_Inst_ff_SDE_78_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_78_current_state_reg_U1 ( .A(state_shifted[86]), 
        .ZN(RoundReg_Inst_ff_SDE_78_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_78_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_78_next_state), .CK(clk), .Q(state_shifted[86]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_79_MUX_inst_XOR1_U1 ( .A(RoundOutput[79]), .B(
        state_shifted[79]), .Z(RoundReg_Inst_ff_SDE_79_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_79_MUX_inst_AND1_U1 ( .A1(RoundReg_n6), .A2(
        RoundReg_Inst_ff_SDE_79_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_79_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_79_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_79_MUX_inst_Y), .B(RoundOutput[79]), .Z(
        RoundReg_Inst_ff_SDE_79_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_79_current_state_reg_U1 ( .A(state_shifted[87]), 
        .ZN(RoundReg_Inst_ff_SDE_79_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_79_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_79_next_state), .CK(clk), .Q(state_shifted[87]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_80_MUX_inst_XOR1_U1 ( .A(RoundOutput[80]), .B(
        state_shifted[80]), .Z(RoundReg_Inst_ff_SDE_80_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_80_MUX_inst_AND1_U1 ( .A1(RoundReg_n9), .A2(
        RoundReg_Inst_ff_SDE_80_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_80_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_80_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_80_MUX_inst_Y), .B(RoundOutput[80]), .Z(
        RoundReg_Inst_ff_SDE_80_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_80_current_state_reg_U1 ( .A(state_shifted[88]), 
        .ZN(RoundReg_Inst_ff_SDE_80_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_80_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_80_next_state), .CK(clk), .Q(state_shifted[88]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_81_MUX_inst_XOR1_U1 ( .A(RoundOutput[81]), .B(
        state_shifted[81]), .Z(RoundReg_Inst_ff_SDE_81_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_81_MUX_inst_AND1_U1 ( .A1(RoundReg_n9), .A2(
        RoundReg_Inst_ff_SDE_81_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_81_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_81_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_81_MUX_inst_Y), .B(RoundOutput[81]), .Z(
        RoundReg_Inst_ff_SDE_81_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_81_current_state_reg_U1 ( .A(state_shifted[89]), 
        .ZN(RoundReg_Inst_ff_SDE_81_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_81_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_81_next_state), .CK(clk), .Q(state_shifted[89]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_82_MUX_inst_XOR1_U1 ( .A(RoundOutput[82]), .B(
        state_shifted[82]), .Z(RoundReg_Inst_ff_SDE_82_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_82_MUX_inst_AND1_U1 ( .A1(RoundReg_n9), .A2(
        RoundReg_Inst_ff_SDE_82_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_82_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_82_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_82_MUX_inst_Y), .B(RoundOutput[82]), .Z(
        RoundReg_Inst_ff_SDE_82_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_82_current_state_reg_U1 ( .A(state_shifted[90]), 
        .ZN(RoundReg_Inst_ff_SDE_82_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_82_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_82_next_state), .CK(clk), .Q(state_shifted[90]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_83_MUX_inst_XOR1_U1 ( .A(RoundOutput[83]), .B(
        state_shifted[83]), .Z(RoundReg_Inst_ff_SDE_83_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_83_MUX_inst_AND1_U1 ( .A1(RoundReg_n9), .A2(
        RoundReg_Inst_ff_SDE_83_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_83_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_83_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_83_MUX_inst_Y), .B(RoundOutput[83]), .Z(
        RoundReg_Inst_ff_SDE_83_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_83_current_state_reg_U1 ( .A(state_shifted[91]), 
        .ZN(RoundReg_Inst_ff_SDE_83_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_83_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_83_next_state), .CK(clk), .Q(state_shifted[91]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_84_MUX_inst_XOR1_U1 ( .A(RoundOutput[84]), .B(
        state_shifted[84]), .Z(RoundReg_Inst_ff_SDE_84_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_84_MUX_inst_AND1_U1 ( .A1(RoundReg_n9), .A2(
        RoundReg_Inst_ff_SDE_84_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_84_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_84_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_84_MUX_inst_Y), .B(RoundOutput[84]), .Z(
        RoundReg_Inst_ff_SDE_84_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_84_current_state_reg_U1 ( .A(state_shifted[92]), 
        .ZN(RoundReg_Inst_ff_SDE_84_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_84_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_84_next_state), .CK(clk), .Q(state_shifted[92]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_85_MUX_inst_XOR1_U1 ( .A(RoundOutput[85]), .B(
        state_shifted[85]), .Z(RoundReg_Inst_ff_SDE_85_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_85_MUX_inst_AND1_U1 ( .A1(RoundReg_n9), .A2(
        RoundReg_Inst_ff_SDE_85_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_85_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_85_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_85_MUX_inst_Y), .B(RoundOutput[85]), .Z(
        RoundReg_Inst_ff_SDE_85_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_85_current_state_reg_U1 ( .A(state_shifted[93]), 
        .ZN(RoundReg_Inst_ff_SDE_85_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_85_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_85_next_state), .CK(clk), .Q(state_shifted[93]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_86_MUX_inst_XOR1_U1 ( .A(RoundOutput[86]), .B(
        state_shifted[86]), .Z(RoundReg_Inst_ff_SDE_86_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_86_MUX_inst_AND1_U1 ( .A1(RoundReg_n9), .A2(
        RoundReg_Inst_ff_SDE_86_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_86_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_86_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_86_MUX_inst_Y), .B(RoundOutput[86]), .Z(
        RoundReg_Inst_ff_SDE_86_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_86_current_state_reg_U1 ( .A(state_shifted[94]), 
        .ZN(RoundReg_Inst_ff_SDE_86_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_86_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_86_next_state), .CK(clk), .Q(state_shifted[94]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_87_MUX_inst_XOR1_U1 ( .A(RoundOutput[87]), .B(
        state_shifted[87]), .Z(RoundReg_Inst_ff_SDE_87_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_87_MUX_inst_AND1_U1 ( .A1(RoundReg_n9), .A2(
        RoundReg_Inst_ff_SDE_87_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_87_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_87_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_87_MUX_inst_Y), .B(RoundOutput[87]), .Z(
        RoundReg_Inst_ff_SDE_87_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_87_current_state_reg_U1 ( .A(state_shifted[95]), 
        .ZN(RoundReg_Inst_ff_SDE_87_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_87_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_87_next_state), .CK(clk), .Q(state_shifted[95]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_88_MUX_inst_XOR1_U1 ( .A(RoundOutput[88]), .B(
        state_shifted[88]), .Z(RoundReg_Inst_ff_SDE_88_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_88_MUX_inst_AND1_U1 ( .A1(RoundReg_n9), .A2(
        RoundReg_Inst_ff_SDE_88_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_88_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_88_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_88_MUX_inst_Y), .B(RoundOutput[88]), .Z(
        RoundReg_Inst_ff_SDE_88_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_88_current_state_reg_U1 ( .A(state_shifted[96]), 
        .ZN(RoundReg_Inst_ff_SDE_88_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_88_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_88_next_state), .CK(clk), .Q(state_shifted[96]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_89_MUX_inst_XOR1_U1 ( .A(RoundOutput[89]), .B(
        state_shifted[89]), .Z(RoundReg_Inst_ff_SDE_89_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_89_MUX_inst_AND1_U1 ( .A1(RoundReg_n9), .A2(
        RoundReg_Inst_ff_SDE_89_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_89_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_89_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_89_MUX_inst_Y), .B(RoundOutput[89]), .Z(
        RoundReg_Inst_ff_SDE_89_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_89_current_state_reg_U1 ( .A(state_shifted[97]), 
        .ZN(RoundReg_Inst_ff_SDE_89_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_89_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_89_next_state), .CK(clk), .Q(state_shifted[97]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_90_MUX_inst_XOR1_U1 ( .A(RoundOutput[90]), .B(
        state_shifted[90]), .Z(RoundReg_Inst_ff_SDE_90_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_90_MUX_inst_AND1_U1 ( .A1(RoundReg_n9), .A2(
        RoundReg_Inst_ff_SDE_90_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_90_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_90_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_90_MUX_inst_Y), .B(RoundOutput[90]), .Z(
        RoundReg_Inst_ff_SDE_90_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_90_current_state_reg_U1 ( .A(state_shifted[98]), 
        .ZN(RoundReg_Inst_ff_SDE_90_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_90_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_90_next_state), .CK(clk), .Q(state_shifted[98]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_91_MUX_inst_XOR1_U1 ( .A(RoundOutput[91]), .B(
        state_shifted[91]), .Z(RoundReg_Inst_ff_SDE_91_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_91_MUX_inst_AND1_U1 ( .A1(RoundReg_n9), .A2(
        RoundReg_Inst_ff_SDE_91_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_91_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_91_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_91_MUX_inst_Y), .B(RoundOutput[91]), .Z(
        RoundReg_Inst_ff_SDE_91_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_91_current_state_reg_U1 ( .A(state_shifted[99]), 
        .ZN(RoundReg_Inst_ff_SDE_91_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_91_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_91_next_state), .CK(clk), .Q(state_shifted[99]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_92_MUX_inst_XOR1_U1 ( .A(RoundOutput[92]), .B(
        state_shifted[92]), .Z(RoundReg_Inst_ff_SDE_92_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_92_MUX_inst_AND1_U1 ( .A1(RoundReg_n8), .A2(
        RoundReg_Inst_ff_SDE_92_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_92_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_92_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_92_MUX_inst_Y), .B(RoundOutput[92]), .Z(
        RoundReg_Inst_ff_SDE_92_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_92_current_state_reg_U1 ( .A(state_shifted[100]), 
        .ZN(RoundReg_Inst_ff_SDE_92_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_92_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_92_next_state), .CK(clk), .Q(state_shifted[100]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_93_MUX_inst_XOR1_U1 ( .A(RoundOutput[93]), .B(
        state_shifted[93]), .Z(RoundReg_Inst_ff_SDE_93_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_93_MUX_inst_AND1_U1 ( .A1(RoundReg_n8), .A2(
        RoundReg_Inst_ff_SDE_93_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_93_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_93_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_93_MUX_inst_Y), .B(RoundOutput[93]), .Z(
        RoundReg_Inst_ff_SDE_93_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_93_current_state_reg_U1 ( .A(state_shifted[101]), 
        .ZN(RoundReg_Inst_ff_SDE_93_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_93_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_93_next_state), .CK(clk), .Q(state_shifted[101]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_94_MUX_inst_XOR1_U1 ( .A(RoundOutput[94]), .B(
        state_shifted[94]), .Z(RoundReg_Inst_ff_SDE_94_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_94_MUX_inst_AND1_U1 ( .A1(RoundReg_n8), .A2(
        RoundReg_Inst_ff_SDE_94_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_94_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_94_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_94_MUX_inst_Y), .B(RoundOutput[94]), .Z(
        RoundReg_Inst_ff_SDE_94_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_94_current_state_reg_U1 ( .A(state_shifted[102]), 
        .ZN(RoundReg_Inst_ff_SDE_94_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_94_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_94_next_state), .CK(clk), .Q(state_shifted[102]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_95_MUX_inst_XOR1_U1 ( .A(RoundOutput[95]), .B(
        state_shifted[95]), .Z(RoundReg_Inst_ff_SDE_95_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_95_MUX_inst_AND1_U1 ( .A1(RoundReg_n8), .A2(
        RoundReg_Inst_ff_SDE_95_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_95_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_95_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_95_MUX_inst_Y), .B(RoundOutput[95]), .Z(
        RoundReg_Inst_ff_SDE_95_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_95_current_state_reg_U1 ( .A(state_shifted[103]), 
        .ZN(RoundReg_Inst_ff_SDE_95_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_95_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_95_next_state), .CK(clk), .Q(state_shifted[103]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_96_MUX_inst_XOR1_U1 ( .A(RoundOutput[96]), .B(
        state_shifted[96]), .Z(RoundReg_Inst_ff_SDE_96_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_96_MUX_inst_AND1_U1 ( .A1(RoundReg_n8), .A2(
        RoundReg_Inst_ff_SDE_96_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_96_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_96_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_96_MUX_inst_Y), .B(RoundOutput[96]), .Z(
        RoundReg_Inst_ff_SDE_96_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_96_current_state_reg_U1 ( .A(state_shifted[104]), 
        .ZN(RoundReg_Inst_ff_SDE_96_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_96_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_96_next_state), .CK(clk), .Q(state_shifted[104]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_97_MUX_inst_XOR1_U1 ( .A(RoundOutput[97]), .B(
        state_shifted[97]), .Z(RoundReg_Inst_ff_SDE_97_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_97_MUX_inst_AND1_U1 ( .A1(RoundReg_n8), .A2(
        RoundReg_Inst_ff_SDE_97_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_97_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_97_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_97_MUX_inst_Y), .B(RoundOutput[97]), .Z(
        RoundReg_Inst_ff_SDE_97_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_97_current_state_reg_U1 ( .A(state_shifted[105]), 
        .ZN(RoundReg_Inst_ff_SDE_97_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_97_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_97_next_state), .CK(clk), .Q(state_shifted[105]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_98_MUX_inst_XOR1_U1 ( .A(RoundOutput[98]), .B(
        state_shifted[98]), .Z(RoundReg_Inst_ff_SDE_98_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_98_MUX_inst_AND1_U1 ( .A1(RoundReg_n8), .A2(
        RoundReg_Inst_ff_SDE_98_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_98_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_98_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_98_MUX_inst_Y), .B(RoundOutput[98]), .Z(
        RoundReg_Inst_ff_SDE_98_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_98_current_state_reg_U1 ( .A(state_shifted[106]), 
        .ZN(RoundReg_Inst_ff_SDE_98_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_98_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_98_next_state), .CK(clk), .Q(state_shifted[106]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_99_MUX_inst_XOR1_U1 ( .A(RoundOutput[99]), .B(
        state_shifted[99]), .Z(RoundReg_Inst_ff_SDE_99_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_99_MUX_inst_AND1_U1 ( .A1(RoundReg_n8), .A2(
        RoundReg_Inst_ff_SDE_99_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_99_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_99_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_99_MUX_inst_Y), .B(RoundOutput[99]), .Z(
        RoundReg_Inst_ff_SDE_99_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_99_current_state_reg_U1 ( .A(state_shifted[107]), 
        .ZN(RoundReg_Inst_ff_SDE_99_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_99_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_99_next_state), .CK(clk), .Q(state_shifted[107]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_100_MUX_inst_XOR1_U1 ( .A(RoundOutput[100]), 
        .B(state_shifted[100]), .Z(RoundReg_Inst_ff_SDE_100_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_100_MUX_inst_AND1_U1 ( .A1(RoundReg_n8), .A2(
        RoundReg_Inst_ff_SDE_100_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_100_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_100_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_100_MUX_inst_Y), .B(RoundOutput[100]), .Z(
        RoundReg_Inst_ff_SDE_100_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_100_current_state_reg_U1 ( .A(state_shifted[108]), .ZN(RoundReg_Inst_ff_SDE_100_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_100_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_100_next_state), .CK(clk), .Q(state_shifted[108]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_101_MUX_inst_XOR1_U1 ( .A(RoundOutput[101]), 
        .B(state_shifted[101]), .Z(RoundReg_Inst_ff_SDE_101_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_101_MUX_inst_AND1_U1 ( .A1(RoundReg_n8), .A2(
        RoundReg_Inst_ff_SDE_101_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_101_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_101_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_101_MUX_inst_Y), .B(RoundOutput[101]), .Z(
        RoundReg_Inst_ff_SDE_101_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_101_current_state_reg_U1 ( .A(state_shifted[109]), .ZN(RoundReg_Inst_ff_SDE_101_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_101_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_101_next_state), .CK(clk), .Q(state_shifted[109]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_102_MUX_inst_XOR1_U1 ( .A(RoundOutput[102]), 
        .B(state_shifted[102]), .Z(RoundReg_Inst_ff_SDE_102_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_102_MUX_inst_AND1_U1 ( .A1(RoundReg_n8), .A2(
        RoundReg_Inst_ff_SDE_102_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_102_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_102_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_102_MUX_inst_Y), .B(RoundOutput[102]), .Z(
        RoundReg_Inst_ff_SDE_102_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_102_current_state_reg_U1 ( .A(state_shifted[110]), .ZN(RoundReg_Inst_ff_SDE_102_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_102_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_102_next_state), .CK(clk), .Q(state_shifted[110]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_103_MUX_inst_XOR1_U1 ( .A(RoundOutput[103]), 
        .B(state_shifted[103]), .Z(RoundReg_Inst_ff_SDE_103_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_103_MUX_inst_AND1_U1 ( .A1(RoundReg_n8), .A2(
        RoundReg_Inst_ff_SDE_103_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_103_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_103_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_103_MUX_inst_Y), .B(RoundOutput[103]), .Z(
        RoundReg_Inst_ff_SDE_103_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_103_current_state_reg_U1 ( .A(state_shifted[111]), .ZN(RoundReg_Inst_ff_SDE_103_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_103_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_103_next_state), .CK(clk), .Q(state_shifted[111]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_104_MUX_inst_XOR1_U1 ( .A(RoundOutput[104]), 
        .B(state_shifted[104]), .Z(RoundReg_Inst_ff_SDE_104_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_104_MUX_inst_AND1_U1 ( .A1(RoundReg_n7), .A2(
        RoundReg_Inst_ff_SDE_104_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_104_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_104_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_104_MUX_inst_Y), .B(RoundOutput[104]), .Z(
        RoundReg_Inst_ff_SDE_104_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_104_current_state_reg_U1 ( .A(state_shifted[112]), .ZN(RoundReg_Inst_ff_SDE_104_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_104_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_104_next_state), .CK(clk), .Q(state_shifted[112]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_105_MUX_inst_XOR1_U1 ( .A(RoundOutput[105]), 
        .B(state_shifted[105]), .Z(RoundReg_Inst_ff_SDE_105_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_105_MUX_inst_AND1_U1 ( .A1(RoundReg_n7), .A2(
        RoundReg_Inst_ff_SDE_105_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_105_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_105_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_105_MUX_inst_Y), .B(RoundOutput[105]), .Z(
        RoundReg_Inst_ff_SDE_105_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_105_current_state_reg_U1 ( .A(state_shifted[113]), .ZN(RoundReg_Inst_ff_SDE_105_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_105_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_105_next_state), .CK(clk), .Q(state_shifted[113]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_106_MUX_inst_XOR1_U1 ( .A(RoundOutput[106]), 
        .B(state_shifted[106]), .Z(RoundReg_Inst_ff_SDE_106_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_106_MUX_inst_AND1_U1 ( .A1(RoundReg_n7), .A2(
        RoundReg_Inst_ff_SDE_106_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_106_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_106_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_106_MUX_inst_Y), .B(RoundOutput[106]), .Z(
        RoundReg_Inst_ff_SDE_106_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_106_current_state_reg_U1 ( .A(state_shifted[114]), .ZN(RoundReg_Inst_ff_SDE_106_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_106_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_106_next_state), .CK(clk), .Q(state_shifted[114]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_107_MUX_inst_XOR1_U1 ( .A(RoundOutput[107]), 
        .B(state_shifted[107]), .Z(RoundReg_Inst_ff_SDE_107_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_107_MUX_inst_AND1_U1 ( .A1(RoundReg_n7), .A2(
        RoundReg_Inst_ff_SDE_107_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_107_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_107_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_107_MUX_inst_Y), .B(RoundOutput[107]), .Z(
        RoundReg_Inst_ff_SDE_107_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_107_current_state_reg_U1 ( .A(state_shifted[115]), .ZN(RoundReg_Inst_ff_SDE_107_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_107_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_107_next_state), .CK(clk), .Q(state_shifted[115]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_108_MUX_inst_XOR1_U1 ( .A(RoundOutput[108]), 
        .B(state_shifted[108]), .Z(RoundReg_Inst_ff_SDE_108_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_108_MUX_inst_AND1_U1 ( .A1(RoundReg_n7), .A2(
        RoundReg_Inst_ff_SDE_108_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_108_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_108_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_108_MUX_inst_Y), .B(RoundOutput[108]), .Z(
        RoundReg_Inst_ff_SDE_108_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_108_current_state_reg_U1 ( .A(state_shifted[116]), .ZN(RoundReg_Inst_ff_SDE_108_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_108_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_108_next_state), .CK(clk), .Q(state_shifted[116]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_109_MUX_inst_XOR1_U1 ( .A(RoundOutput[109]), 
        .B(state_shifted[109]), .Z(RoundReg_Inst_ff_SDE_109_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_109_MUX_inst_AND1_U1 ( .A1(RoundReg_n7), .A2(
        RoundReg_Inst_ff_SDE_109_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_109_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_109_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_109_MUX_inst_Y), .B(RoundOutput[109]), .Z(
        RoundReg_Inst_ff_SDE_109_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_109_current_state_reg_U1 ( .A(state_shifted[117]), .ZN(RoundReg_Inst_ff_SDE_109_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_109_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_109_next_state), .CK(clk), .Q(state_shifted[117]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_110_MUX_inst_XOR1_U1 ( .A(RoundOutput[110]), 
        .B(state_shifted[110]), .Z(RoundReg_Inst_ff_SDE_110_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_110_MUX_inst_AND1_U1 ( .A1(RoundReg_n7), .A2(
        RoundReg_Inst_ff_SDE_110_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_110_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_110_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_110_MUX_inst_Y), .B(RoundOutput[110]), .Z(
        RoundReg_Inst_ff_SDE_110_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_110_current_state_reg_U1 ( .A(state_shifted[118]), .ZN(RoundReg_Inst_ff_SDE_110_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_110_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_110_next_state), .CK(clk), .Q(state_shifted[118]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_111_MUX_inst_XOR1_U1 ( .A(RoundOutput[111]), 
        .B(state_shifted[111]), .Z(RoundReg_Inst_ff_SDE_111_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_111_MUX_inst_AND1_U1 ( .A1(RoundReg_n7), .A2(
        RoundReg_Inst_ff_SDE_111_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_111_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_111_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_111_MUX_inst_Y), .B(RoundOutput[111]), .Z(
        RoundReg_Inst_ff_SDE_111_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_111_current_state_reg_U1 ( .A(state_shifted[119]), .ZN(RoundReg_Inst_ff_SDE_111_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_111_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_111_next_state), .CK(clk), .Q(state_shifted[119]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_112_MUX_inst_XOR1_U1 ( .A(RoundOutput[112]), 
        .B(state_shifted[112]), .Z(RoundReg_Inst_ff_SDE_112_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_112_MUX_inst_AND1_U1 ( .A1(RoundReg_n7), .A2(
        RoundReg_Inst_ff_SDE_112_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_112_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_112_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_112_MUX_inst_Y), .B(RoundOutput[112]), .Z(
        RoundReg_Inst_ff_SDE_112_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_112_current_state_reg_U1 ( .A(state_shifted[120]), .ZN(RoundReg_Inst_ff_SDE_112_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_112_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_112_next_state), .CK(clk), .Q(state_shifted[120]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_113_MUX_inst_XOR1_U1 ( .A(RoundOutput[113]), 
        .B(state_shifted[113]), .Z(RoundReg_Inst_ff_SDE_113_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_113_MUX_inst_AND1_U1 ( .A1(RoundReg_n7), .A2(
        RoundReg_Inst_ff_SDE_113_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_113_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_113_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_113_MUX_inst_Y), .B(RoundOutput[113]), .Z(
        RoundReg_Inst_ff_SDE_113_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_113_current_state_reg_U1 ( .A(state_shifted[121]), .ZN(RoundReg_Inst_ff_SDE_113_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_113_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_113_next_state), .CK(clk), .Q(state_shifted[121]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_114_MUX_inst_XOR1_U1 ( .A(RoundOutput[114]), 
        .B(state_shifted[114]), .Z(RoundReg_Inst_ff_SDE_114_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_114_MUX_inst_AND1_U1 ( .A1(RoundReg_n7), .A2(
        RoundReg_Inst_ff_SDE_114_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_114_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_114_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_114_MUX_inst_Y), .B(RoundOutput[114]), .Z(
        RoundReg_Inst_ff_SDE_114_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_114_current_state_reg_U1 ( .A(state_shifted[122]), .ZN(RoundReg_Inst_ff_SDE_114_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_114_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_114_next_state), .CK(clk), .Q(state_shifted[122]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_115_MUX_inst_XOR1_U1 ( .A(RoundOutput[115]), 
        .B(state_shifted[115]), .Z(RoundReg_Inst_ff_SDE_115_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_115_MUX_inst_AND1_U1 ( .A1(RoundReg_n7), .A2(
        RoundReg_Inst_ff_SDE_115_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_115_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_115_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_115_MUX_inst_Y), .B(RoundOutput[115]), .Z(
        RoundReg_Inst_ff_SDE_115_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_115_current_state_reg_U1 ( .A(state_shifted[123]), .ZN(RoundReg_Inst_ff_SDE_115_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_115_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_115_next_state), .CK(clk), .Q(state_shifted[123]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_116_MUX_inst_XOR1_U1 ( .A(RoundOutput[116]), 
        .B(state_shifted[116]), .Z(RoundReg_Inst_ff_SDE_116_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_116_MUX_inst_AND1_U1 ( .A1(RoundReg_n6), .A2(
        RoundReg_Inst_ff_SDE_116_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_116_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_116_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_116_MUX_inst_Y), .B(RoundOutput[116]), .Z(
        RoundReg_Inst_ff_SDE_116_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_116_current_state_reg_U1 ( .A(state_shifted[124]), .ZN(RoundReg_Inst_ff_SDE_116_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_116_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_116_next_state), .CK(clk), .Q(state_shifted[124]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_117_MUX_inst_XOR1_U1 ( .A(RoundOutput[117]), 
        .B(state_shifted[117]), .Z(RoundReg_Inst_ff_SDE_117_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_117_MUX_inst_AND1_U1 ( .A1(RoundReg_n6), .A2(
        RoundReg_Inst_ff_SDE_117_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_117_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_117_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_117_MUX_inst_Y), .B(RoundOutput[117]), .Z(
        RoundReg_Inst_ff_SDE_117_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_117_current_state_reg_U1 ( .A(state_shifted[125]), .ZN(RoundReg_Inst_ff_SDE_117_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_117_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_117_next_state), .CK(clk), .Q(state_shifted[125]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_118_MUX_inst_XOR1_U1 ( .A(RoundOutput[118]), 
        .B(state_shifted[118]), .Z(RoundReg_Inst_ff_SDE_118_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_118_MUX_inst_AND1_U1 ( .A1(RoundReg_n6), .A2(
        RoundReg_Inst_ff_SDE_118_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_118_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_118_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_118_MUX_inst_Y), .B(RoundOutput[118]), .Z(
        RoundReg_Inst_ff_SDE_118_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_118_current_state_reg_U1 ( .A(state_shifted[126]), .ZN(RoundReg_Inst_ff_SDE_118_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_118_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_118_next_state), .CK(clk), .Q(state_shifted[126]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_119_MUX_inst_XOR1_U1 ( .A(RoundOutput[119]), 
        .B(state_shifted[119]), .Z(RoundReg_Inst_ff_SDE_119_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_119_MUX_inst_AND1_U1 ( .A1(RoundReg_n6), .A2(
        RoundReg_Inst_ff_SDE_119_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_119_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_119_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_119_MUX_inst_Y), .B(RoundOutput[119]), .Z(
        RoundReg_Inst_ff_SDE_119_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_119_current_state_reg_U1 ( .A(state_shifted[127]), .ZN(RoundReg_Inst_ff_SDE_119_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_119_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_119_next_state), .CK(clk), .Q(state_shifted[127]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_120_MUX_inst_XOR1_U1 ( .A(RoundOutput[120]), 
        .B(state_shifted[120]), .Z(RoundReg_Inst_ff_SDE_120_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_120_MUX_inst_AND1_U1 ( .A1(RoundReg_n6), .A2(
        RoundReg_Inst_ff_SDE_120_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_120_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_120_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_120_MUX_inst_Y), .B(RoundOutput[120]), .Z(
        RoundReg_Inst_ff_SDE_120_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_120_current_state_reg_U1 ( .A(RoundInput[120]), 
        .ZN(RoundReg_Inst_ff_SDE_120_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_120_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_120_next_state), .CK(clk), .Q(RoundInput[120]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_121_MUX_inst_XOR1_U1 ( .A(RoundOutput[121]), 
        .B(state_shifted[121]), .Z(RoundReg_Inst_ff_SDE_121_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_121_MUX_inst_AND1_U1 ( .A1(RoundReg_n6), .A2(
        RoundReg_Inst_ff_SDE_121_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_121_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_121_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_121_MUX_inst_Y), .B(RoundOutput[121]), .Z(
        RoundReg_Inst_ff_SDE_121_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_121_current_state_reg_U1 ( .A(RoundInput[121]), 
        .ZN(RoundReg_Inst_ff_SDE_121_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_121_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_121_next_state), .CK(clk), .Q(RoundInput[121]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_122_MUX_inst_XOR1_U1 ( .A(RoundOutput[122]), 
        .B(state_shifted[122]), .Z(RoundReg_Inst_ff_SDE_122_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_122_MUX_inst_AND1_U1 ( .A1(RoundReg_n6), .A2(
        RoundReg_Inst_ff_SDE_122_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_122_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_122_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_122_MUX_inst_Y), .B(RoundOutput[122]), .Z(
        RoundReg_Inst_ff_SDE_122_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_122_current_state_reg_U1 ( .A(RoundInput[122]), 
        .ZN(RoundReg_Inst_ff_SDE_122_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_122_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_122_next_state), .CK(clk), .Q(RoundInput[122]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_123_MUX_inst_XOR1_U1 ( .A(RoundOutput[123]), 
        .B(state_shifted[123]), .Z(RoundReg_Inst_ff_SDE_123_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_123_MUX_inst_AND1_U1 ( .A1(RoundReg_n6), .A2(
        RoundReg_Inst_ff_SDE_123_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_123_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_123_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_123_MUX_inst_Y), .B(RoundOutput[123]), .Z(
        RoundReg_Inst_ff_SDE_123_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_123_current_state_reg_U1 ( .A(RoundInput[123]), 
        .ZN(RoundReg_Inst_ff_SDE_123_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_123_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_123_next_state), .CK(clk), .Q(RoundInput[123]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_124_MUX_inst_XOR1_U1 ( .A(RoundOutput[124]), 
        .B(state_shifted[124]), .Z(RoundReg_Inst_ff_SDE_124_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_124_MUX_inst_AND1_U1 ( .A1(RoundReg_n6), .A2(
        RoundReg_Inst_ff_SDE_124_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_124_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_124_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_124_MUX_inst_Y), .B(RoundOutput[124]), .Z(
        RoundReg_Inst_ff_SDE_124_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_124_current_state_reg_U1 ( .A(RoundInput[124]), 
        .ZN(RoundReg_Inst_ff_SDE_124_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_124_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_124_next_state), .CK(clk), .Q(RoundInput[124]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_125_MUX_inst_XOR1_U1 ( .A(RoundOutput[125]), 
        .B(state_shifted[125]), .Z(RoundReg_Inst_ff_SDE_125_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_125_MUX_inst_AND1_U1 ( .A1(RoundReg_n6), .A2(
        RoundReg_Inst_ff_SDE_125_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_125_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_125_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_125_MUX_inst_Y), .B(RoundOutput[125]), .Z(
        RoundReg_Inst_ff_SDE_125_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_125_current_state_reg_U1 ( .A(RoundInput[125]), 
        .ZN(RoundReg_Inst_ff_SDE_125_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_125_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_125_next_state), .CK(clk), .Q(RoundInput[125]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_126_MUX_inst_XOR1_U1 ( .A(RoundOutput[126]), 
        .B(state_shifted[126]), .Z(RoundReg_Inst_ff_SDE_126_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_126_MUX_inst_AND1_U1 ( .A1(RoundReg_n6), .A2(
        RoundReg_Inst_ff_SDE_126_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_126_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_126_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_126_MUX_inst_Y), .B(RoundOutput[126]), .Z(
        RoundReg_Inst_ff_SDE_126_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_126_current_state_reg_U1 ( .A(RoundInput[126]), 
        .ZN(RoundReg_Inst_ff_SDE_126_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_126_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_126_next_state), .CK(clk), .Q(RoundInput[126]), 
        .QN() );
  XOR2_X1 RoundReg_Inst_ff_SDE_127_MUX_inst_XOR1_U1 ( .A(RoundOutput[127]), 
        .B(state_shifted[127]), .Z(RoundReg_Inst_ff_SDE_127_MUX_inst_X) );
  AND2_X1 RoundReg_Inst_ff_SDE_127_MUX_inst_AND1_U1 ( .A1(RoundReg_n6), .A2(
        RoundReg_Inst_ff_SDE_127_MUX_inst_X), .ZN(
        RoundReg_Inst_ff_SDE_127_MUX_inst_Y) );
  XOR2_X1 RoundReg_Inst_ff_SDE_127_MUX_inst_XOR2_U1 ( .A(
        RoundReg_Inst_ff_SDE_127_MUX_inst_Y), .B(RoundOutput[127]), .Z(
        RoundReg_Inst_ff_SDE_127_next_state) );
  INV_X1 RoundReg_Inst_ff_SDE_127_current_state_reg_U1 ( .A(RoundInput[127]), 
        .ZN(RoundReg_Inst_ff_SDE_127_current_state_reg_QN) );
  DFF_X1 RoundReg_Inst_ff_SDE_127_current_state_reg_FF_FF ( .D(
        RoundReg_Inst_ff_SDE_127_next_state), .CK(clk), .Q(RoundInput[127]), 
        .QN() );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T1_U1 ( .A(SubBytesInput[7]), .B(
        SubBytesInput[4]), .Z(SubBytesIns_Inst_Sbox_0_T1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T2_U1 ( .A(SubBytesInput[7]), .B(
        SubBytesInput[2]), .Z(SubBytesIns_Inst_Sbox_0_T2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T3_U1 ( .A(SubBytesInput[7]), .B(
        SubBytesInput[1]), .Z(SubBytesIns_Inst_Sbox_0_T3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T4_U1 ( .A(SubBytesInput[4]), .B(
        SubBytesInput[2]), .Z(SubBytesIns_Inst_Sbox_0_T4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T5_U1 ( .A(SubBytesInput[3]), .B(
        SubBytesInput[1]), .Z(SubBytesIns_Inst_Sbox_0_T5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T6_U1 ( .A(SubBytesIns_Inst_Sbox_0_T1), 
        .B(SubBytesIns_Inst_Sbox_0_T5), .Z(SubBytesIns_Inst_Sbox_0_T6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T7_U1 ( .A(SubBytesInput[6]), .B(
        SubBytesInput[5]), .Z(SubBytesIns_Inst_Sbox_0_T7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T8_U1 ( .A(SubBytesInput[0]), .B(
        SubBytesIns_Inst_Sbox_0_T6), .Z(SubBytesIns_Inst_Sbox_0_T8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T9_U1 ( .A(SubBytesInput[0]), .B(
        SubBytesIns_Inst_Sbox_0_T7), .Z(SubBytesIns_Inst_Sbox_0_T9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T10_U1 ( .A(SubBytesIns_Inst_Sbox_0_T6), 
        .B(SubBytesIns_Inst_Sbox_0_T7), .Z(SubBytesIns_Inst_Sbox_0_T10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T11_U1 ( .A(SubBytesInput[6]), .B(
        SubBytesInput[2]), .Z(SubBytesIns_Inst_Sbox_0_T11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T12_U1 ( .A(SubBytesInput[5]), .B(
        SubBytesInput[2]), .Z(SubBytesIns_Inst_Sbox_0_T12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T13_U1 ( .A(SubBytesIns_Inst_Sbox_0_T3), 
        .B(SubBytesIns_Inst_Sbox_0_T4), .Z(SubBytesIns_Inst_Sbox_0_T13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T14_U1 ( .A(SubBytesIns_Inst_Sbox_0_T6), 
        .B(SubBytesIns_Inst_Sbox_0_T11), .Z(SubBytesIns_Inst_Sbox_0_T14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T15_U1 ( .A(SubBytesIns_Inst_Sbox_0_T5), 
        .B(SubBytesIns_Inst_Sbox_0_T11), .Z(SubBytesIns_Inst_Sbox_0_T15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T16_U1 ( .A(SubBytesIns_Inst_Sbox_0_T5), 
        .B(SubBytesIns_Inst_Sbox_0_T12), .Z(SubBytesIns_Inst_Sbox_0_T16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T17_U1 ( .A(SubBytesIns_Inst_Sbox_0_T9), 
        .B(SubBytesIns_Inst_Sbox_0_T16), .Z(SubBytesIns_Inst_Sbox_0_T17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T18_U1 ( .A(SubBytesInput[4]), .B(
        SubBytesInput[0]), .Z(SubBytesIns_Inst_Sbox_0_T18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T19_U1 ( .A(SubBytesIns_Inst_Sbox_0_T7), 
        .B(SubBytesIns_Inst_Sbox_0_T18), .Z(SubBytesIns_Inst_Sbox_0_T19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T20_U1 ( .A(SubBytesIns_Inst_Sbox_0_T1), 
        .B(SubBytesIns_Inst_Sbox_0_T19), .Z(SubBytesIns_Inst_Sbox_0_T20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T21_U1 ( .A(SubBytesInput[1]), .B(
        SubBytesInput[0]), .Z(SubBytesIns_Inst_Sbox_0_T21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T22_U1 ( .A(SubBytesIns_Inst_Sbox_0_T7), 
        .B(SubBytesIns_Inst_Sbox_0_T21), .Z(SubBytesIns_Inst_Sbox_0_T22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T23_U1 ( .A(SubBytesIns_Inst_Sbox_0_T2), 
        .B(SubBytesIns_Inst_Sbox_0_T22), .Z(SubBytesIns_Inst_Sbox_0_T23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T24_U1 ( .A(SubBytesIns_Inst_Sbox_0_T2), 
        .B(SubBytesIns_Inst_Sbox_0_T10), .Z(SubBytesIns_Inst_Sbox_0_T24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T25_U1 ( .A(SubBytesIns_Inst_Sbox_0_T20), 
        .B(SubBytesIns_Inst_Sbox_0_T17), .Z(SubBytesIns_Inst_Sbox_0_T25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T26_U1 ( .A(SubBytesIns_Inst_Sbox_0_T3), 
        .B(SubBytesIns_Inst_Sbox_0_T16), .Z(SubBytesIns_Inst_Sbox_0_T26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_T27_U1 ( .A(SubBytesIns_Inst_Sbox_0_T1), 
        .B(SubBytesIns_Inst_Sbox_0_T12), .Z(SubBytesIns_Inst_Sbox_0_T27) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M1_U1 ( .A1(SubBytesIns_Inst_Sbox_0_T13), 
        .A2(SubBytesIns_Inst_Sbox_0_T6), .ZN(SubBytesIns_Inst_Sbox_0_M1) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M2_U1 ( .A1(SubBytesIns_Inst_Sbox_0_T23), 
        .A2(SubBytesIns_Inst_Sbox_0_T8), .ZN(SubBytesIns_Inst_Sbox_0_M2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M3_U1 ( .A(SubBytesIns_Inst_Sbox_0_T14), 
        .B(SubBytesIns_Inst_Sbox_0_M1), .Z(SubBytesIns_Inst_Sbox_0_M3) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M4_U1 ( .A1(SubBytesIns_Inst_Sbox_0_T19), 
        .A2(SubBytesInput[0]), .ZN(SubBytesIns_Inst_Sbox_0_M4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M5_U1 ( .A(SubBytesIns_Inst_Sbox_0_M4), 
        .B(SubBytesIns_Inst_Sbox_0_M1), .Z(SubBytesIns_Inst_Sbox_0_M5) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M6_U1 ( .A1(SubBytesIns_Inst_Sbox_0_T3), 
        .A2(SubBytesIns_Inst_Sbox_0_T16), .ZN(SubBytesIns_Inst_Sbox_0_M6) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M7_U1 ( .A1(SubBytesIns_Inst_Sbox_0_T22), 
        .A2(SubBytesIns_Inst_Sbox_0_T9), .ZN(SubBytesIns_Inst_Sbox_0_M7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M8_U1 ( .A(SubBytesIns_Inst_Sbox_0_T26), 
        .B(SubBytesIns_Inst_Sbox_0_M6), .Z(SubBytesIns_Inst_Sbox_0_M8) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M9_U1 ( .A1(SubBytesIns_Inst_Sbox_0_T20), 
        .A2(SubBytesIns_Inst_Sbox_0_T17), .ZN(SubBytesIns_Inst_Sbox_0_M9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M10_U1 ( .A(SubBytesIns_Inst_Sbox_0_M9), 
        .B(SubBytesIns_Inst_Sbox_0_M6), .Z(SubBytesIns_Inst_Sbox_0_M10) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M11_U1 ( .A1(SubBytesIns_Inst_Sbox_0_T1), 
        .A2(SubBytesIns_Inst_Sbox_0_T15), .ZN(SubBytesIns_Inst_Sbox_0_M11) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M12_U1 ( .A1(SubBytesIns_Inst_Sbox_0_T4), 
        .A2(SubBytesIns_Inst_Sbox_0_T27), .ZN(SubBytesIns_Inst_Sbox_0_M12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M13_U1 ( .A(SubBytesIns_Inst_Sbox_0_M12), 
        .B(SubBytesIns_Inst_Sbox_0_M11), .Z(SubBytesIns_Inst_Sbox_0_M13) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M14_U1 ( .A1(SubBytesIns_Inst_Sbox_0_T2), 
        .A2(SubBytesIns_Inst_Sbox_0_T10), .ZN(SubBytesIns_Inst_Sbox_0_M14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M15_U1 ( .A(SubBytesIns_Inst_Sbox_0_M14), 
        .B(SubBytesIns_Inst_Sbox_0_M11), .Z(SubBytesIns_Inst_Sbox_0_M15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M16_U1 ( .A(SubBytesIns_Inst_Sbox_0_M3), 
        .B(SubBytesIns_Inst_Sbox_0_M2), .Z(SubBytesIns_Inst_Sbox_0_M16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M17_U1 ( .A(SubBytesIns_Inst_Sbox_0_M5), 
        .B(SubBytesIns_Inst_Sbox_0_T24), .Z(SubBytesIns_Inst_Sbox_0_M17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M18_U1 ( .A(SubBytesIns_Inst_Sbox_0_M8), 
        .B(SubBytesIns_Inst_Sbox_0_M7), .Z(SubBytesIns_Inst_Sbox_0_M18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M19_U1 ( .A(SubBytesIns_Inst_Sbox_0_M10), 
        .B(SubBytesIns_Inst_Sbox_0_M15), .Z(SubBytesIns_Inst_Sbox_0_M19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M20_U1 ( .A(SubBytesIns_Inst_Sbox_0_M16), 
        .B(SubBytesIns_Inst_Sbox_0_M13), .Z(SubBytesIns_Inst_Sbox_0_M20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M21_U1 ( .A(SubBytesIns_Inst_Sbox_0_M17), 
        .B(SubBytesIns_Inst_Sbox_0_M15), .Z(SubBytesIns_Inst_Sbox_0_M21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M22_U1 ( .A(SubBytesIns_Inst_Sbox_0_M18), 
        .B(SubBytesIns_Inst_Sbox_0_M13), .Z(SubBytesIns_Inst_Sbox_0_M22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M23_U1 ( .A(SubBytesIns_Inst_Sbox_0_M19), 
        .B(SubBytesIns_Inst_Sbox_0_T25), .Z(SubBytesIns_Inst_Sbox_0_M23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M24_U1 ( .A(SubBytesIns_Inst_Sbox_0_M22), 
        .B(SubBytesIns_Inst_Sbox_0_M23), .Z(SubBytesIns_Inst_Sbox_0_M24) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M25_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M22), .A2(SubBytesIns_Inst_Sbox_0_M20), .ZN(SubBytesIns_Inst_Sbox_0_M25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M26_U1 ( .A(SubBytesIns_Inst_Sbox_0_M21), 
        .B(SubBytesIns_Inst_Sbox_0_M25), .Z(SubBytesIns_Inst_Sbox_0_M26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M27_U1 ( .A(SubBytesIns_Inst_Sbox_0_M20), 
        .B(SubBytesIns_Inst_Sbox_0_M21), .Z(SubBytesIns_Inst_Sbox_0_M27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M28_U1 ( .A(SubBytesIns_Inst_Sbox_0_M23), 
        .B(SubBytesIns_Inst_Sbox_0_M25), .Z(SubBytesIns_Inst_Sbox_0_M28) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M29_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M28), .A2(SubBytesIns_Inst_Sbox_0_M27), .ZN(SubBytesIns_Inst_Sbox_0_M29) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M30_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M26), .A2(SubBytesIns_Inst_Sbox_0_M24), .ZN(SubBytesIns_Inst_Sbox_0_M30) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M31_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M20), .A2(SubBytesIns_Inst_Sbox_0_M23), .ZN(SubBytesIns_Inst_Sbox_0_M31) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M32_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M27), .A2(SubBytesIns_Inst_Sbox_0_M31), .ZN(SubBytesIns_Inst_Sbox_0_M32) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M33_U1 ( .A(SubBytesIns_Inst_Sbox_0_M27), 
        .B(SubBytesIns_Inst_Sbox_0_M25), .Z(SubBytesIns_Inst_Sbox_0_M33) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M34_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M21), .A2(SubBytesIns_Inst_Sbox_0_M22), .ZN(SubBytesIns_Inst_Sbox_0_M34) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M35_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M24), .A2(SubBytesIns_Inst_Sbox_0_M34), .ZN(SubBytesIns_Inst_Sbox_0_M35) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M36_U1 ( .A(SubBytesIns_Inst_Sbox_0_M24), 
        .B(SubBytesIns_Inst_Sbox_0_M25), .Z(SubBytesIns_Inst_Sbox_0_M36) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M37_U1 ( .A(SubBytesIns_Inst_Sbox_0_M21), 
        .B(SubBytesIns_Inst_Sbox_0_M29), .Z(SubBytesIns_Inst_Sbox_0_M37) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M38_U1 ( .A(SubBytesIns_Inst_Sbox_0_M32), 
        .B(SubBytesIns_Inst_Sbox_0_M33), .Z(SubBytesIns_Inst_Sbox_0_M38) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M39_U1 ( .A(SubBytesIns_Inst_Sbox_0_M23), 
        .B(SubBytesIns_Inst_Sbox_0_M30), .Z(SubBytesIns_Inst_Sbox_0_M39) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M40_U1 ( .A(SubBytesIns_Inst_Sbox_0_M35), 
        .B(SubBytesIns_Inst_Sbox_0_M36), .Z(SubBytesIns_Inst_Sbox_0_M40) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M41_U1 ( .A(SubBytesIns_Inst_Sbox_0_M38), 
        .B(SubBytesIns_Inst_Sbox_0_M40), .Z(SubBytesIns_Inst_Sbox_0_M41) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M42_U1 ( .A(SubBytesIns_Inst_Sbox_0_M37), 
        .B(SubBytesIns_Inst_Sbox_0_M39), .Z(SubBytesIns_Inst_Sbox_0_M42) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M43_U1 ( .A(SubBytesIns_Inst_Sbox_0_M37), 
        .B(SubBytesIns_Inst_Sbox_0_M38), .Z(SubBytesIns_Inst_Sbox_0_M43) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M44_U1 ( .A(SubBytesIns_Inst_Sbox_0_M39), 
        .B(SubBytesIns_Inst_Sbox_0_M40), .Z(SubBytesIns_Inst_Sbox_0_M44) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_M45_U1 ( .A(SubBytesIns_Inst_Sbox_0_M42), 
        .B(SubBytesIns_Inst_Sbox_0_M41), .Z(SubBytesIns_Inst_Sbox_0_M45) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M46_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M44), .A2(SubBytesIns_Inst_Sbox_0_T6), .ZN(SubBytesIns_Inst_Sbox_0_M46) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M47_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M40), .A2(SubBytesIns_Inst_Sbox_0_T8), .ZN(SubBytesIns_Inst_Sbox_0_M47) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M48_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M39), .A2(SubBytesInput[0]), .ZN(SubBytesIns_Inst_Sbox_0_M48) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M49_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M43), .A2(SubBytesIns_Inst_Sbox_0_T16), .ZN(SubBytesIns_Inst_Sbox_0_M49) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M50_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M38), .A2(SubBytesIns_Inst_Sbox_0_T9), .ZN(SubBytesIns_Inst_Sbox_0_M50) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M51_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M37), .A2(SubBytesIns_Inst_Sbox_0_T17), .ZN(SubBytesIns_Inst_Sbox_0_M51) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M52_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M42), .A2(SubBytesIns_Inst_Sbox_0_T15), .ZN(SubBytesIns_Inst_Sbox_0_M52) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M53_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M45), .A2(SubBytesIns_Inst_Sbox_0_T27), .ZN(SubBytesIns_Inst_Sbox_0_M53) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M54_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M41), .A2(SubBytesIns_Inst_Sbox_0_T10), .ZN(SubBytesIns_Inst_Sbox_0_M54) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M55_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M44), .A2(SubBytesIns_Inst_Sbox_0_T13), .ZN(SubBytesIns_Inst_Sbox_0_M55) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M56_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M40), .A2(SubBytesIns_Inst_Sbox_0_T23), .ZN(SubBytesIns_Inst_Sbox_0_M56) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M57_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M39), .A2(SubBytesIns_Inst_Sbox_0_T19), .ZN(SubBytesIns_Inst_Sbox_0_M57) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M58_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M43), .A2(SubBytesIns_Inst_Sbox_0_T3), .ZN(SubBytesIns_Inst_Sbox_0_M58) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M59_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M38), .A2(SubBytesIns_Inst_Sbox_0_T22), .ZN(SubBytesIns_Inst_Sbox_0_M59) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M60_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M37), .A2(SubBytesIns_Inst_Sbox_0_T20), .ZN(SubBytesIns_Inst_Sbox_0_M60) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M61_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M42), .A2(SubBytesIns_Inst_Sbox_0_T1), .ZN(SubBytesIns_Inst_Sbox_0_M61) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M62_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M45), .A2(SubBytesIns_Inst_Sbox_0_T4), .ZN(SubBytesIns_Inst_Sbox_0_M62) );
  AND2_X1 SubBytesIns_Inst_Sbox_0_AND_M63_U1 ( .A1(SubBytesIns_Inst_Sbox_0_M41), .A2(SubBytesIns_Inst_Sbox_0_T2), .ZN(SubBytesIns_Inst_Sbox_0_M63) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L0_U1 ( .A(SubBytesIns_Inst_Sbox_0_M61), 
        .B(SubBytesIns_Inst_Sbox_0_M62), .Z(SubBytesIns_Inst_Sbox_0_L0) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L1_U1 ( .A(SubBytesIns_Inst_Sbox_0_M50), 
        .B(SubBytesIns_Inst_Sbox_0_M56), .Z(SubBytesIns_Inst_Sbox_0_L1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L2_U1 ( .A(SubBytesIns_Inst_Sbox_0_M46), 
        .B(SubBytesIns_Inst_Sbox_0_M48), .Z(SubBytesIns_Inst_Sbox_0_L2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L3_U1 ( .A(SubBytesIns_Inst_Sbox_0_M47), 
        .B(SubBytesIns_Inst_Sbox_0_M55), .Z(SubBytesIns_Inst_Sbox_0_L3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L4_U1 ( .A(SubBytesIns_Inst_Sbox_0_M54), 
        .B(SubBytesIns_Inst_Sbox_0_M58), .Z(SubBytesIns_Inst_Sbox_0_L4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L5_U1 ( .A(SubBytesIns_Inst_Sbox_0_M49), 
        .B(SubBytesIns_Inst_Sbox_0_M61), .Z(SubBytesIns_Inst_Sbox_0_L5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L6_U1 ( .A(SubBytesIns_Inst_Sbox_0_M62), 
        .B(SubBytesIns_Inst_Sbox_0_L5), .Z(SubBytesIns_Inst_Sbox_0_L6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L7_U1 ( .A(SubBytesIns_Inst_Sbox_0_M46), 
        .B(SubBytesIns_Inst_Sbox_0_L3), .Z(SubBytesIns_Inst_Sbox_0_L7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L8_U1 ( .A(SubBytesIns_Inst_Sbox_0_M51), 
        .B(SubBytesIns_Inst_Sbox_0_M59), .Z(SubBytesIns_Inst_Sbox_0_L8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L9_U1 ( .A(SubBytesIns_Inst_Sbox_0_M52), 
        .B(SubBytesIns_Inst_Sbox_0_M53), .Z(SubBytesIns_Inst_Sbox_0_L9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L10_U1 ( .A(SubBytesIns_Inst_Sbox_0_M53), 
        .B(SubBytesIns_Inst_Sbox_0_L4), .Z(SubBytesIns_Inst_Sbox_0_L10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L11_U1 ( .A(SubBytesIns_Inst_Sbox_0_M60), 
        .B(SubBytesIns_Inst_Sbox_0_L2), .Z(SubBytesIns_Inst_Sbox_0_L11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L12_U1 ( .A(SubBytesIns_Inst_Sbox_0_M48), 
        .B(SubBytesIns_Inst_Sbox_0_M51), .Z(SubBytesIns_Inst_Sbox_0_L12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L13_U1 ( .A(SubBytesIns_Inst_Sbox_0_M50), 
        .B(SubBytesIns_Inst_Sbox_0_L0), .Z(SubBytesIns_Inst_Sbox_0_L13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L14_U1 ( .A(SubBytesIns_Inst_Sbox_0_M52), 
        .B(SubBytesIns_Inst_Sbox_0_M61), .Z(SubBytesIns_Inst_Sbox_0_L14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L15_U1 ( .A(SubBytesIns_Inst_Sbox_0_M55), 
        .B(SubBytesIns_Inst_Sbox_0_L1), .Z(SubBytesIns_Inst_Sbox_0_L15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L16_U1 ( .A(SubBytesIns_Inst_Sbox_0_M56), 
        .B(SubBytesIns_Inst_Sbox_0_L0), .Z(SubBytesIns_Inst_Sbox_0_L16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L17_U1 ( .A(SubBytesIns_Inst_Sbox_0_M57), 
        .B(SubBytesIns_Inst_Sbox_0_L1), .Z(SubBytesIns_Inst_Sbox_0_L17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L18_U1 ( .A(SubBytesIns_Inst_Sbox_0_M58), 
        .B(SubBytesIns_Inst_Sbox_0_L8), .Z(SubBytesIns_Inst_Sbox_0_L18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L19_U1 ( .A(SubBytesIns_Inst_Sbox_0_M63), 
        .B(SubBytesIns_Inst_Sbox_0_L4), .Z(SubBytesIns_Inst_Sbox_0_L19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L20_U1 ( .A(SubBytesIns_Inst_Sbox_0_L0), 
        .B(SubBytesIns_Inst_Sbox_0_L1), .Z(SubBytesIns_Inst_Sbox_0_L20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L21_U1 ( .A(SubBytesIns_Inst_Sbox_0_L1), 
        .B(SubBytesIns_Inst_Sbox_0_L7), .Z(SubBytesIns_Inst_Sbox_0_L21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L22_U1 ( .A(SubBytesIns_Inst_Sbox_0_L3), 
        .B(SubBytesIns_Inst_Sbox_0_L12), .Z(SubBytesIns_Inst_Sbox_0_L22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L23_U1 ( .A(SubBytesIns_Inst_Sbox_0_L18), 
        .B(SubBytesIns_Inst_Sbox_0_L2), .Z(SubBytesIns_Inst_Sbox_0_L23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L24_U1 ( .A(SubBytesIns_Inst_Sbox_0_L15), 
        .B(SubBytesIns_Inst_Sbox_0_L9), .Z(SubBytesIns_Inst_Sbox_0_L24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L25_U1 ( .A(SubBytesIns_Inst_Sbox_0_L6), 
        .B(SubBytesIns_Inst_Sbox_0_L10), .Z(SubBytesIns_Inst_Sbox_0_L25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L26_U1 ( .A(SubBytesIns_Inst_Sbox_0_L7), 
        .B(SubBytesIns_Inst_Sbox_0_L9), .Z(SubBytesIns_Inst_Sbox_0_L26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L27_U1 ( .A(SubBytesIns_Inst_Sbox_0_L8), 
        .B(SubBytesIns_Inst_Sbox_0_L10), .Z(SubBytesIns_Inst_Sbox_0_L27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L28_U1 ( .A(SubBytesIns_Inst_Sbox_0_L11), 
        .B(SubBytesIns_Inst_Sbox_0_L14), .Z(SubBytesIns_Inst_Sbox_0_L28) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_L29_U1 ( .A(SubBytesIns_Inst_Sbox_0_L11), 
        .B(SubBytesIns_Inst_Sbox_0_L17), .Z(SubBytesIns_Inst_Sbox_0_L29) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_S0_U1 ( .A(SubBytesIns_Inst_Sbox_0_L6), 
        .B(SubBytesIns_Inst_Sbox_0_L24), .Z(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_S1_U1 ( .A(SubBytesIns_Inst_Sbox_0_L16), 
        .B(SubBytesIns_Inst_Sbox_0_L26), .ZN(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[7]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_S2_U1 ( .A(SubBytesIns_Inst_Sbox_0_L19), 
        .B(SubBytesIns_Inst_Sbox_0_L28), .ZN(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[6]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_S3_U1 ( .A(SubBytesIns_Inst_Sbox_0_L6), 
        .B(SubBytesIns_Inst_Sbox_0_L21), .Z(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[5]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_S4_U1 ( .A(SubBytesIns_Inst_Sbox_0_L20), 
        .B(SubBytesIns_Inst_Sbox_0_L22), .Z(MixColumnsInput[99]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_S5_U1 ( .A(SubBytesIns_Inst_Sbox_0_L25), 
        .B(SubBytesIns_Inst_Sbox_0_L29), .Z(MixColumnsInput[98]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_S6_U1 ( .A(SubBytesIns_Inst_Sbox_0_L13), 
        .B(SubBytesIns_Inst_Sbox_0_L27), .ZN(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[2]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_0_XOR_S7_U1 ( .A(SubBytesIns_Inst_Sbox_0_L6), 
        .B(SubBytesIns_Inst_Sbox_0_L23), .ZN(MixColumnsInput[96]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T1_U1 ( .A(SubBytesInput[15]), .B(
        SubBytesInput[12]), .Z(SubBytesIns_Inst_Sbox_1_T1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T2_U1 ( .A(SubBytesInput[15]), .B(
        SubBytesInput[10]), .Z(SubBytesIns_Inst_Sbox_1_T2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T3_U1 ( .A(SubBytesInput[15]), .B(
        SubBytesInput[9]), .Z(SubBytesIns_Inst_Sbox_1_T3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T4_U1 ( .A(SubBytesInput[12]), .B(
        SubBytesInput[10]), .Z(SubBytesIns_Inst_Sbox_1_T4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T5_U1 ( .A(SubBytesInput[11]), .B(
        SubBytesInput[9]), .Z(SubBytesIns_Inst_Sbox_1_T5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T6_U1 ( .A(SubBytesIns_Inst_Sbox_1_T1), 
        .B(SubBytesIns_Inst_Sbox_1_T5), .Z(SubBytesIns_Inst_Sbox_1_T6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T7_U1 ( .A(SubBytesInput[14]), .B(
        SubBytesInput[13]), .Z(SubBytesIns_Inst_Sbox_1_T7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T8_U1 ( .A(SubBytesInput[8]), .B(
        SubBytesIns_Inst_Sbox_1_T6), .Z(SubBytesIns_Inst_Sbox_1_T8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T9_U1 ( .A(SubBytesInput[8]), .B(
        SubBytesIns_Inst_Sbox_1_T7), .Z(SubBytesIns_Inst_Sbox_1_T9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T10_U1 ( .A(SubBytesIns_Inst_Sbox_1_T6), 
        .B(SubBytesIns_Inst_Sbox_1_T7), .Z(SubBytesIns_Inst_Sbox_1_T10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T11_U1 ( .A(SubBytesInput[14]), .B(
        SubBytesInput[10]), .Z(SubBytesIns_Inst_Sbox_1_T11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T12_U1 ( .A(SubBytesInput[13]), .B(
        SubBytesInput[10]), .Z(SubBytesIns_Inst_Sbox_1_T12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T13_U1 ( .A(SubBytesIns_Inst_Sbox_1_T3), 
        .B(SubBytesIns_Inst_Sbox_1_T4), .Z(SubBytesIns_Inst_Sbox_1_T13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T14_U1 ( .A(SubBytesIns_Inst_Sbox_1_T6), 
        .B(SubBytesIns_Inst_Sbox_1_T11), .Z(SubBytesIns_Inst_Sbox_1_T14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T15_U1 ( .A(SubBytesIns_Inst_Sbox_1_T5), 
        .B(SubBytesIns_Inst_Sbox_1_T11), .Z(SubBytesIns_Inst_Sbox_1_T15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T16_U1 ( .A(SubBytesIns_Inst_Sbox_1_T5), 
        .B(SubBytesIns_Inst_Sbox_1_T12), .Z(SubBytesIns_Inst_Sbox_1_T16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T17_U1 ( .A(SubBytesIns_Inst_Sbox_1_T9), 
        .B(SubBytesIns_Inst_Sbox_1_T16), .Z(SubBytesIns_Inst_Sbox_1_T17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T18_U1 ( .A(SubBytesInput[12]), .B(
        SubBytesInput[8]), .Z(SubBytesIns_Inst_Sbox_1_T18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T19_U1 ( .A(SubBytesIns_Inst_Sbox_1_T7), 
        .B(SubBytesIns_Inst_Sbox_1_T18), .Z(SubBytesIns_Inst_Sbox_1_T19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T20_U1 ( .A(SubBytesIns_Inst_Sbox_1_T1), 
        .B(SubBytesIns_Inst_Sbox_1_T19), .Z(SubBytesIns_Inst_Sbox_1_T20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T21_U1 ( .A(SubBytesInput[9]), .B(
        SubBytesInput[8]), .Z(SubBytesIns_Inst_Sbox_1_T21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T22_U1 ( .A(SubBytesIns_Inst_Sbox_1_T7), 
        .B(SubBytesIns_Inst_Sbox_1_T21), .Z(SubBytesIns_Inst_Sbox_1_T22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T23_U1 ( .A(SubBytesIns_Inst_Sbox_1_T2), 
        .B(SubBytesIns_Inst_Sbox_1_T22), .Z(SubBytesIns_Inst_Sbox_1_T23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T24_U1 ( .A(SubBytesIns_Inst_Sbox_1_T2), 
        .B(SubBytesIns_Inst_Sbox_1_T10), .Z(SubBytesIns_Inst_Sbox_1_T24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T25_U1 ( .A(SubBytesIns_Inst_Sbox_1_T20), 
        .B(SubBytesIns_Inst_Sbox_1_T17), .Z(SubBytesIns_Inst_Sbox_1_T25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T26_U1 ( .A(SubBytesIns_Inst_Sbox_1_T3), 
        .B(SubBytesIns_Inst_Sbox_1_T16), .Z(SubBytesIns_Inst_Sbox_1_T26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_T27_U1 ( .A(SubBytesIns_Inst_Sbox_1_T1), 
        .B(SubBytesIns_Inst_Sbox_1_T12), .Z(SubBytesIns_Inst_Sbox_1_T27) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M1_U1 ( .A1(SubBytesIns_Inst_Sbox_1_T13), 
        .A2(SubBytesIns_Inst_Sbox_1_T6), .ZN(SubBytesIns_Inst_Sbox_1_M1) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M2_U1 ( .A1(SubBytesIns_Inst_Sbox_1_T23), 
        .A2(SubBytesIns_Inst_Sbox_1_T8), .ZN(SubBytesIns_Inst_Sbox_1_M2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M3_U1 ( .A(SubBytesIns_Inst_Sbox_1_T14), 
        .B(SubBytesIns_Inst_Sbox_1_M1), .Z(SubBytesIns_Inst_Sbox_1_M3) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M4_U1 ( .A1(SubBytesIns_Inst_Sbox_1_T19), 
        .A2(SubBytesInput[8]), .ZN(SubBytesIns_Inst_Sbox_1_M4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M5_U1 ( .A(SubBytesIns_Inst_Sbox_1_M4), 
        .B(SubBytesIns_Inst_Sbox_1_M1), .Z(SubBytesIns_Inst_Sbox_1_M5) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M6_U1 ( .A1(SubBytesIns_Inst_Sbox_1_T3), 
        .A2(SubBytesIns_Inst_Sbox_1_T16), .ZN(SubBytesIns_Inst_Sbox_1_M6) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M7_U1 ( .A1(SubBytesIns_Inst_Sbox_1_T22), 
        .A2(SubBytesIns_Inst_Sbox_1_T9), .ZN(SubBytesIns_Inst_Sbox_1_M7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M8_U1 ( .A(SubBytesIns_Inst_Sbox_1_T26), 
        .B(SubBytesIns_Inst_Sbox_1_M6), .Z(SubBytesIns_Inst_Sbox_1_M8) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M9_U1 ( .A1(SubBytesIns_Inst_Sbox_1_T20), 
        .A2(SubBytesIns_Inst_Sbox_1_T17), .ZN(SubBytesIns_Inst_Sbox_1_M9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M10_U1 ( .A(SubBytesIns_Inst_Sbox_1_M9), 
        .B(SubBytesIns_Inst_Sbox_1_M6), .Z(SubBytesIns_Inst_Sbox_1_M10) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M11_U1 ( .A1(SubBytesIns_Inst_Sbox_1_T1), 
        .A2(SubBytesIns_Inst_Sbox_1_T15), .ZN(SubBytesIns_Inst_Sbox_1_M11) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M12_U1 ( .A1(SubBytesIns_Inst_Sbox_1_T4), 
        .A2(SubBytesIns_Inst_Sbox_1_T27), .ZN(SubBytesIns_Inst_Sbox_1_M12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M13_U1 ( .A(SubBytesIns_Inst_Sbox_1_M12), 
        .B(SubBytesIns_Inst_Sbox_1_M11), .Z(SubBytesIns_Inst_Sbox_1_M13) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M14_U1 ( .A1(SubBytesIns_Inst_Sbox_1_T2), 
        .A2(SubBytesIns_Inst_Sbox_1_T10), .ZN(SubBytesIns_Inst_Sbox_1_M14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M15_U1 ( .A(SubBytesIns_Inst_Sbox_1_M14), 
        .B(SubBytesIns_Inst_Sbox_1_M11), .Z(SubBytesIns_Inst_Sbox_1_M15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M16_U1 ( .A(SubBytesIns_Inst_Sbox_1_M3), 
        .B(SubBytesIns_Inst_Sbox_1_M2), .Z(SubBytesIns_Inst_Sbox_1_M16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M17_U1 ( .A(SubBytesIns_Inst_Sbox_1_M5), 
        .B(SubBytesIns_Inst_Sbox_1_T24), .Z(SubBytesIns_Inst_Sbox_1_M17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M18_U1 ( .A(SubBytesIns_Inst_Sbox_1_M8), 
        .B(SubBytesIns_Inst_Sbox_1_M7), .Z(SubBytesIns_Inst_Sbox_1_M18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M19_U1 ( .A(SubBytesIns_Inst_Sbox_1_M10), 
        .B(SubBytesIns_Inst_Sbox_1_M15), .Z(SubBytesIns_Inst_Sbox_1_M19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M20_U1 ( .A(SubBytesIns_Inst_Sbox_1_M16), 
        .B(SubBytesIns_Inst_Sbox_1_M13), .Z(SubBytesIns_Inst_Sbox_1_M20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M21_U1 ( .A(SubBytesIns_Inst_Sbox_1_M17), 
        .B(SubBytesIns_Inst_Sbox_1_M15), .Z(SubBytesIns_Inst_Sbox_1_M21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M22_U1 ( .A(SubBytesIns_Inst_Sbox_1_M18), 
        .B(SubBytesIns_Inst_Sbox_1_M13), .Z(SubBytesIns_Inst_Sbox_1_M22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M23_U1 ( .A(SubBytesIns_Inst_Sbox_1_M19), 
        .B(SubBytesIns_Inst_Sbox_1_T25), .Z(SubBytesIns_Inst_Sbox_1_M23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M24_U1 ( .A(SubBytesIns_Inst_Sbox_1_M22), 
        .B(SubBytesIns_Inst_Sbox_1_M23), .Z(SubBytesIns_Inst_Sbox_1_M24) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M25_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M22), .A2(SubBytesIns_Inst_Sbox_1_M20), .ZN(SubBytesIns_Inst_Sbox_1_M25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M26_U1 ( .A(SubBytesIns_Inst_Sbox_1_M21), 
        .B(SubBytesIns_Inst_Sbox_1_M25), .Z(SubBytesIns_Inst_Sbox_1_M26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M27_U1 ( .A(SubBytesIns_Inst_Sbox_1_M20), 
        .B(SubBytesIns_Inst_Sbox_1_M21), .Z(SubBytesIns_Inst_Sbox_1_M27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M28_U1 ( .A(SubBytesIns_Inst_Sbox_1_M23), 
        .B(SubBytesIns_Inst_Sbox_1_M25), .Z(SubBytesIns_Inst_Sbox_1_M28) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M29_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M28), .A2(SubBytesIns_Inst_Sbox_1_M27), .ZN(SubBytesIns_Inst_Sbox_1_M29) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M30_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M26), .A2(SubBytesIns_Inst_Sbox_1_M24), .ZN(SubBytesIns_Inst_Sbox_1_M30) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M31_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M20), .A2(SubBytesIns_Inst_Sbox_1_M23), .ZN(SubBytesIns_Inst_Sbox_1_M31) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M32_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M27), .A2(SubBytesIns_Inst_Sbox_1_M31), .ZN(SubBytesIns_Inst_Sbox_1_M32) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M33_U1 ( .A(SubBytesIns_Inst_Sbox_1_M27), 
        .B(SubBytesIns_Inst_Sbox_1_M25), .Z(SubBytesIns_Inst_Sbox_1_M33) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M34_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M21), .A2(SubBytesIns_Inst_Sbox_1_M22), .ZN(SubBytesIns_Inst_Sbox_1_M34) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M35_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M24), .A2(SubBytesIns_Inst_Sbox_1_M34), .ZN(SubBytesIns_Inst_Sbox_1_M35) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M36_U1 ( .A(SubBytesIns_Inst_Sbox_1_M24), 
        .B(SubBytesIns_Inst_Sbox_1_M25), .Z(SubBytesIns_Inst_Sbox_1_M36) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M37_U1 ( .A(SubBytesIns_Inst_Sbox_1_M21), 
        .B(SubBytesIns_Inst_Sbox_1_M29), .Z(SubBytesIns_Inst_Sbox_1_M37) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M38_U1 ( .A(SubBytesIns_Inst_Sbox_1_M32), 
        .B(SubBytesIns_Inst_Sbox_1_M33), .Z(SubBytesIns_Inst_Sbox_1_M38) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M39_U1 ( .A(SubBytesIns_Inst_Sbox_1_M23), 
        .B(SubBytesIns_Inst_Sbox_1_M30), .Z(SubBytesIns_Inst_Sbox_1_M39) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M40_U1 ( .A(SubBytesIns_Inst_Sbox_1_M35), 
        .B(SubBytesIns_Inst_Sbox_1_M36), .Z(SubBytesIns_Inst_Sbox_1_M40) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M41_U1 ( .A(SubBytesIns_Inst_Sbox_1_M38), 
        .B(SubBytesIns_Inst_Sbox_1_M40), .Z(SubBytesIns_Inst_Sbox_1_M41) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M42_U1 ( .A(SubBytesIns_Inst_Sbox_1_M37), 
        .B(SubBytesIns_Inst_Sbox_1_M39), .Z(SubBytesIns_Inst_Sbox_1_M42) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M43_U1 ( .A(SubBytesIns_Inst_Sbox_1_M37), 
        .B(SubBytesIns_Inst_Sbox_1_M38), .Z(SubBytesIns_Inst_Sbox_1_M43) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M44_U1 ( .A(SubBytesIns_Inst_Sbox_1_M39), 
        .B(SubBytesIns_Inst_Sbox_1_M40), .Z(SubBytesIns_Inst_Sbox_1_M44) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_M45_U1 ( .A(SubBytesIns_Inst_Sbox_1_M42), 
        .B(SubBytesIns_Inst_Sbox_1_M41), .Z(SubBytesIns_Inst_Sbox_1_M45) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M46_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M44), .A2(SubBytesIns_Inst_Sbox_1_T6), .ZN(SubBytesIns_Inst_Sbox_1_M46) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M47_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M40), .A2(SubBytesIns_Inst_Sbox_1_T8), .ZN(SubBytesIns_Inst_Sbox_1_M47) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M48_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M39), .A2(SubBytesInput[8]), .ZN(SubBytesIns_Inst_Sbox_1_M48) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M49_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M43), .A2(SubBytesIns_Inst_Sbox_1_T16), .ZN(SubBytesIns_Inst_Sbox_1_M49) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M50_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M38), .A2(SubBytesIns_Inst_Sbox_1_T9), .ZN(SubBytesIns_Inst_Sbox_1_M50) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M51_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M37), .A2(SubBytesIns_Inst_Sbox_1_T17), .ZN(SubBytesIns_Inst_Sbox_1_M51) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M52_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M42), .A2(SubBytesIns_Inst_Sbox_1_T15), .ZN(SubBytesIns_Inst_Sbox_1_M52) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M53_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M45), .A2(SubBytesIns_Inst_Sbox_1_T27), .ZN(SubBytesIns_Inst_Sbox_1_M53) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M54_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M41), .A2(SubBytesIns_Inst_Sbox_1_T10), .ZN(SubBytesIns_Inst_Sbox_1_M54) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M55_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M44), .A2(SubBytesIns_Inst_Sbox_1_T13), .ZN(SubBytesIns_Inst_Sbox_1_M55) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M56_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M40), .A2(SubBytesIns_Inst_Sbox_1_T23), .ZN(SubBytesIns_Inst_Sbox_1_M56) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M57_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M39), .A2(SubBytesIns_Inst_Sbox_1_T19), .ZN(SubBytesIns_Inst_Sbox_1_M57) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M58_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M43), .A2(SubBytesIns_Inst_Sbox_1_T3), .ZN(SubBytesIns_Inst_Sbox_1_M58) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M59_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M38), .A2(SubBytesIns_Inst_Sbox_1_T22), .ZN(SubBytesIns_Inst_Sbox_1_M59) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M60_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M37), .A2(SubBytesIns_Inst_Sbox_1_T20), .ZN(SubBytesIns_Inst_Sbox_1_M60) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M61_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M42), .A2(SubBytesIns_Inst_Sbox_1_T1), .ZN(SubBytesIns_Inst_Sbox_1_M61) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M62_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M45), .A2(SubBytesIns_Inst_Sbox_1_T4), .ZN(SubBytesIns_Inst_Sbox_1_M62) );
  AND2_X1 SubBytesIns_Inst_Sbox_1_AND_M63_U1 ( .A1(SubBytesIns_Inst_Sbox_1_M41), .A2(SubBytesIns_Inst_Sbox_1_T2), .ZN(SubBytesIns_Inst_Sbox_1_M63) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L0_U1 ( .A(SubBytesIns_Inst_Sbox_1_M61), 
        .B(SubBytesIns_Inst_Sbox_1_M62), .Z(SubBytesIns_Inst_Sbox_1_L0) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L1_U1 ( .A(SubBytesIns_Inst_Sbox_1_M50), 
        .B(SubBytesIns_Inst_Sbox_1_M56), .Z(SubBytesIns_Inst_Sbox_1_L1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L2_U1 ( .A(SubBytesIns_Inst_Sbox_1_M46), 
        .B(SubBytesIns_Inst_Sbox_1_M48), .Z(SubBytesIns_Inst_Sbox_1_L2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L3_U1 ( .A(SubBytesIns_Inst_Sbox_1_M47), 
        .B(SubBytesIns_Inst_Sbox_1_M55), .Z(SubBytesIns_Inst_Sbox_1_L3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L4_U1 ( .A(SubBytesIns_Inst_Sbox_1_M54), 
        .B(SubBytesIns_Inst_Sbox_1_M58), .Z(SubBytesIns_Inst_Sbox_1_L4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L5_U1 ( .A(SubBytesIns_Inst_Sbox_1_M49), 
        .B(SubBytesIns_Inst_Sbox_1_M61), .Z(SubBytesIns_Inst_Sbox_1_L5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L6_U1 ( .A(SubBytesIns_Inst_Sbox_1_M62), 
        .B(SubBytesIns_Inst_Sbox_1_L5), .Z(SubBytesIns_Inst_Sbox_1_L6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L7_U1 ( .A(SubBytesIns_Inst_Sbox_1_M46), 
        .B(SubBytesIns_Inst_Sbox_1_L3), .Z(SubBytesIns_Inst_Sbox_1_L7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L8_U1 ( .A(SubBytesIns_Inst_Sbox_1_M51), 
        .B(SubBytesIns_Inst_Sbox_1_M59), .Z(SubBytesIns_Inst_Sbox_1_L8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L9_U1 ( .A(SubBytesIns_Inst_Sbox_1_M52), 
        .B(SubBytesIns_Inst_Sbox_1_M53), .Z(SubBytesIns_Inst_Sbox_1_L9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L10_U1 ( .A(SubBytesIns_Inst_Sbox_1_M53), 
        .B(SubBytesIns_Inst_Sbox_1_L4), .Z(SubBytesIns_Inst_Sbox_1_L10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L11_U1 ( .A(SubBytesIns_Inst_Sbox_1_M60), 
        .B(SubBytesIns_Inst_Sbox_1_L2), .Z(SubBytesIns_Inst_Sbox_1_L11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L12_U1 ( .A(SubBytesIns_Inst_Sbox_1_M48), 
        .B(SubBytesIns_Inst_Sbox_1_M51), .Z(SubBytesIns_Inst_Sbox_1_L12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L13_U1 ( .A(SubBytesIns_Inst_Sbox_1_M50), 
        .B(SubBytesIns_Inst_Sbox_1_L0), .Z(SubBytesIns_Inst_Sbox_1_L13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L14_U1 ( .A(SubBytesIns_Inst_Sbox_1_M52), 
        .B(SubBytesIns_Inst_Sbox_1_M61), .Z(SubBytesIns_Inst_Sbox_1_L14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L15_U1 ( .A(SubBytesIns_Inst_Sbox_1_M55), 
        .B(SubBytesIns_Inst_Sbox_1_L1), .Z(SubBytesIns_Inst_Sbox_1_L15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L16_U1 ( .A(SubBytesIns_Inst_Sbox_1_M56), 
        .B(SubBytesIns_Inst_Sbox_1_L0), .Z(SubBytesIns_Inst_Sbox_1_L16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L17_U1 ( .A(SubBytesIns_Inst_Sbox_1_M57), 
        .B(SubBytesIns_Inst_Sbox_1_L1), .Z(SubBytesIns_Inst_Sbox_1_L17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L18_U1 ( .A(SubBytesIns_Inst_Sbox_1_M58), 
        .B(SubBytesIns_Inst_Sbox_1_L8), .Z(SubBytesIns_Inst_Sbox_1_L18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L19_U1 ( .A(SubBytesIns_Inst_Sbox_1_M63), 
        .B(SubBytesIns_Inst_Sbox_1_L4), .Z(SubBytesIns_Inst_Sbox_1_L19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L20_U1 ( .A(SubBytesIns_Inst_Sbox_1_L0), 
        .B(SubBytesIns_Inst_Sbox_1_L1), .Z(SubBytesIns_Inst_Sbox_1_L20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L21_U1 ( .A(SubBytesIns_Inst_Sbox_1_L1), 
        .B(SubBytesIns_Inst_Sbox_1_L7), .Z(SubBytesIns_Inst_Sbox_1_L21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L22_U1 ( .A(SubBytesIns_Inst_Sbox_1_L3), 
        .B(SubBytesIns_Inst_Sbox_1_L12), .Z(SubBytesIns_Inst_Sbox_1_L22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L23_U1 ( .A(SubBytesIns_Inst_Sbox_1_L18), 
        .B(SubBytesIns_Inst_Sbox_1_L2), .Z(SubBytesIns_Inst_Sbox_1_L23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L24_U1 ( .A(SubBytesIns_Inst_Sbox_1_L15), 
        .B(SubBytesIns_Inst_Sbox_1_L9), .Z(SubBytesIns_Inst_Sbox_1_L24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L25_U1 ( .A(SubBytesIns_Inst_Sbox_1_L6), 
        .B(SubBytesIns_Inst_Sbox_1_L10), .Z(SubBytesIns_Inst_Sbox_1_L25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L26_U1 ( .A(SubBytesIns_Inst_Sbox_1_L7), 
        .B(SubBytesIns_Inst_Sbox_1_L9), .Z(SubBytesIns_Inst_Sbox_1_L26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L27_U1 ( .A(SubBytesIns_Inst_Sbox_1_L8), 
        .B(SubBytesIns_Inst_Sbox_1_L10), .Z(SubBytesIns_Inst_Sbox_1_L27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L28_U1 ( .A(SubBytesIns_Inst_Sbox_1_L11), 
        .B(SubBytesIns_Inst_Sbox_1_L14), .Z(SubBytesIns_Inst_Sbox_1_L28) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_L29_U1 ( .A(SubBytesIns_Inst_Sbox_1_L11), 
        .B(SubBytesIns_Inst_Sbox_1_L17), .Z(SubBytesIns_Inst_Sbox_1_L29) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_S0_U1 ( .A(SubBytesIns_Inst_Sbox_1_L6), 
        .B(SubBytesIns_Inst_Sbox_1_L24), .Z(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_S1_U1 ( .A(SubBytesIns_Inst_Sbox_1_L16), 
        .B(SubBytesIns_Inst_Sbox_1_L26), .ZN(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[15]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_S2_U1 ( .A(SubBytesIns_Inst_Sbox_1_L19), 
        .B(SubBytesIns_Inst_Sbox_1_L28), .ZN(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[14]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_S3_U1 ( .A(SubBytesIns_Inst_Sbox_1_L6), 
        .B(SubBytesIns_Inst_Sbox_1_L21), .Z(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[13]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_S4_U1 ( .A(SubBytesIns_Inst_Sbox_1_L20), 
        .B(SubBytesIns_Inst_Sbox_1_L22), .Z(MixColumnsInput[75]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_S5_U1 ( .A(SubBytesIns_Inst_Sbox_1_L25), 
        .B(SubBytesIns_Inst_Sbox_1_L29), .Z(MixColumnsInput[74]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_S6_U1 ( .A(SubBytesIns_Inst_Sbox_1_L13), 
        .B(SubBytesIns_Inst_Sbox_1_L27), .ZN(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[10]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_1_XOR_S7_U1 ( .A(SubBytesIns_Inst_Sbox_1_L6), 
        .B(SubBytesIns_Inst_Sbox_1_L23), .ZN(MixColumnsInput[72]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T1_U1 ( .A(SubBytesInput[23]), .B(
        SubBytesInput[20]), .Z(SubBytesIns_Inst_Sbox_2_T1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T2_U1 ( .A(SubBytesInput[23]), .B(
        SubBytesInput[18]), .Z(SubBytesIns_Inst_Sbox_2_T2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T3_U1 ( .A(SubBytesInput[23]), .B(
        SubBytesInput[17]), .Z(SubBytesIns_Inst_Sbox_2_T3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T4_U1 ( .A(SubBytesInput[20]), .B(
        SubBytesInput[18]), .Z(SubBytesIns_Inst_Sbox_2_T4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T5_U1 ( .A(SubBytesInput[19]), .B(
        SubBytesInput[17]), .Z(SubBytesIns_Inst_Sbox_2_T5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T6_U1 ( .A(SubBytesIns_Inst_Sbox_2_T1), 
        .B(SubBytesIns_Inst_Sbox_2_T5), .Z(SubBytesIns_Inst_Sbox_2_T6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T7_U1 ( .A(SubBytesInput[22]), .B(
        SubBytesInput[21]), .Z(SubBytesIns_Inst_Sbox_2_T7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T8_U1 ( .A(SubBytesInput[16]), .B(
        SubBytesIns_Inst_Sbox_2_T6), .Z(SubBytesIns_Inst_Sbox_2_T8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T9_U1 ( .A(SubBytesInput[16]), .B(
        SubBytesIns_Inst_Sbox_2_T7), .Z(SubBytesIns_Inst_Sbox_2_T9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T10_U1 ( .A(SubBytesIns_Inst_Sbox_2_T6), 
        .B(SubBytesIns_Inst_Sbox_2_T7), .Z(SubBytesIns_Inst_Sbox_2_T10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T11_U1 ( .A(SubBytesInput[22]), .B(
        SubBytesInput[18]), .Z(SubBytesIns_Inst_Sbox_2_T11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T12_U1 ( .A(SubBytesInput[21]), .B(
        SubBytesInput[18]), .Z(SubBytesIns_Inst_Sbox_2_T12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T13_U1 ( .A(SubBytesIns_Inst_Sbox_2_T3), 
        .B(SubBytesIns_Inst_Sbox_2_T4), .Z(SubBytesIns_Inst_Sbox_2_T13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T14_U1 ( .A(SubBytesIns_Inst_Sbox_2_T6), 
        .B(SubBytesIns_Inst_Sbox_2_T11), .Z(SubBytesIns_Inst_Sbox_2_T14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T15_U1 ( .A(SubBytesIns_Inst_Sbox_2_T5), 
        .B(SubBytesIns_Inst_Sbox_2_T11), .Z(SubBytesIns_Inst_Sbox_2_T15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T16_U1 ( .A(SubBytesIns_Inst_Sbox_2_T5), 
        .B(SubBytesIns_Inst_Sbox_2_T12), .Z(SubBytesIns_Inst_Sbox_2_T16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T17_U1 ( .A(SubBytesIns_Inst_Sbox_2_T9), 
        .B(SubBytesIns_Inst_Sbox_2_T16), .Z(SubBytesIns_Inst_Sbox_2_T17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T18_U1 ( .A(SubBytesInput[20]), .B(
        SubBytesInput[16]), .Z(SubBytesIns_Inst_Sbox_2_T18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T19_U1 ( .A(SubBytesIns_Inst_Sbox_2_T7), 
        .B(SubBytesIns_Inst_Sbox_2_T18), .Z(SubBytesIns_Inst_Sbox_2_T19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T20_U1 ( .A(SubBytesIns_Inst_Sbox_2_T1), 
        .B(SubBytesIns_Inst_Sbox_2_T19), .Z(SubBytesIns_Inst_Sbox_2_T20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T21_U1 ( .A(SubBytesInput[17]), .B(
        SubBytesInput[16]), .Z(SubBytesIns_Inst_Sbox_2_T21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T22_U1 ( .A(SubBytesIns_Inst_Sbox_2_T7), 
        .B(SubBytesIns_Inst_Sbox_2_T21), .Z(SubBytesIns_Inst_Sbox_2_T22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T23_U1 ( .A(SubBytesIns_Inst_Sbox_2_T2), 
        .B(SubBytesIns_Inst_Sbox_2_T22), .Z(SubBytesIns_Inst_Sbox_2_T23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T24_U1 ( .A(SubBytesIns_Inst_Sbox_2_T2), 
        .B(SubBytesIns_Inst_Sbox_2_T10), .Z(SubBytesIns_Inst_Sbox_2_T24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T25_U1 ( .A(SubBytesIns_Inst_Sbox_2_T20), 
        .B(SubBytesIns_Inst_Sbox_2_T17), .Z(SubBytesIns_Inst_Sbox_2_T25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T26_U1 ( .A(SubBytesIns_Inst_Sbox_2_T3), 
        .B(SubBytesIns_Inst_Sbox_2_T16), .Z(SubBytesIns_Inst_Sbox_2_T26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_T27_U1 ( .A(SubBytesIns_Inst_Sbox_2_T1), 
        .B(SubBytesIns_Inst_Sbox_2_T12), .Z(SubBytesIns_Inst_Sbox_2_T27) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M1_U1 ( .A1(SubBytesIns_Inst_Sbox_2_T13), 
        .A2(SubBytesIns_Inst_Sbox_2_T6), .ZN(SubBytesIns_Inst_Sbox_2_M1) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M2_U1 ( .A1(SubBytesIns_Inst_Sbox_2_T23), 
        .A2(SubBytesIns_Inst_Sbox_2_T8), .ZN(SubBytesIns_Inst_Sbox_2_M2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M3_U1 ( .A(SubBytesIns_Inst_Sbox_2_T14), 
        .B(SubBytesIns_Inst_Sbox_2_M1), .Z(SubBytesIns_Inst_Sbox_2_M3) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M4_U1 ( .A1(SubBytesIns_Inst_Sbox_2_T19), 
        .A2(SubBytesInput[16]), .ZN(SubBytesIns_Inst_Sbox_2_M4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M5_U1 ( .A(SubBytesIns_Inst_Sbox_2_M4), 
        .B(SubBytesIns_Inst_Sbox_2_M1), .Z(SubBytesIns_Inst_Sbox_2_M5) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M6_U1 ( .A1(SubBytesIns_Inst_Sbox_2_T3), 
        .A2(SubBytesIns_Inst_Sbox_2_T16), .ZN(SubBytesIns_Inst_Sbox_2_M6) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M7_U1 ( .A1(SubBytesIns_Inst_Sbox_2_T22), 
        .A2(SubBytesIns_Inst_Sbox_2_T9), .ZN(SubBytesIns_Inst_Sbox_2_M7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M8_U1 ( .A(SubBytesIns_Inst_Sbox_2_T26), 
        .B(SubBytesIns_Inst_Sbox_2_M6), .Z(SubBytesIns_Inst_Sbox_2_M8) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M9_U1 ( .A1(SubBytesIns_Inst_Sbox_2_T20), 
        .A2(SubBytesIns_Inst_Sbox_2_T17), .ZN(SubBytesIns_Inst_Sbox_2_M9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M10_U1 ( .A(SubBytesIns_Inst_Sbox_2_M9), 
        .B(SubBytesIns_Inst_Sbox_2_M6), .Z(SubBytesIns_Inst_Sbox_2_M10) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M11_U1 ( .A1(SubBytesIns_Inst_Sbox_2_T1), 
        .A2(SubBytesIns_Inst_Sbox_2_T15), .ZN(SubBytesIns_Inst_Sbox_2_M11) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M12_U1 ( .A1(SubBytesIns_Inst_Sbox_2_T4), 
        .A2(SubBytesIns_Inst_Sbox_2_T27), .ZN(SubBytesIns_Inst_Sbox_2_M12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M13_U1 ( .A(SubBytesIns_Inst_Sbox_2_M12), 
        .B(SubBytesIns_Inst_Sbox_2_M11), .Z(SubBytesIns_Inst_Sbox_2_M13) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M14_U1 ( .A1(SubBytesIns_Inst_Sbox_2_T2), 
        .A2(SubBytesIns_Inst_Sbox_2_T10), .ZN(SubBytesIns_Inst_Sbox_2_M14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M15_U1 ( .A(SubBytesIns_Inst_Sbox_2_M14), 
        .B(SubBytesIns_Inst_Sbox_2_M11), .Z(SubBytesIns_Inst_Sbox_2_M15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M16_U1 ( .A(SubBytesIns_Inst_Sbox_2_M3), 
        .B(SubBytesIns_Inst_Sbox_2_M2), .Z(SubBytesIns_Inst_Sbox_2_M16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M17_U1 ( .A(SubBytesIns_Inst_Sbox_2_M5), 
        .B(SubBytesIns_Inst_Sbox_2_T24), .Z(SubBytesIns_Inst_Sbox_2_M17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M18_U1 ( .A(SubBytesIns_Inst_Sbox_2_M8), 
        .B(SubBytesIns_Inst_Sbox_2_M7), .Z(SubBytesIns_Inst_Sbox_2_M18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M19_U1 ( .A(SubBytesIns_Inst_Sbox_2_M10), 
        .B(SubBytesIns_Inst_Sbox_2_M15), .Z(SubBytesIns_Inst_Sbox_2_M19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M20_U1 ( .A(SubBytesIns_Inst_Sbox_2_M16), 
        .B(SubBytesIns_Inst_Sbox_2_M13), .Z(SubBytesIns_Inst_Sbox_2_M20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M21_U1 ( .A(SubBytesIns_Inst_Sbox_2_M17), 
        .B(SubBytesIns_Inst_Sbox_2_M15), .Z(SubBytesIns_Inst_Sbox_2_M21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M22_U1 ( .A(SubBytesIns_Inst_Sbox_2_M18), 
        .B(SubBytesIns_Inst_Sbox_2_M13), .Z(SubBytesIns_Inst_Sbox_2_M22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M23_U1 ( .A(SubBytesIns_Inst_Sbox_2_M19), 
        .B(SubBytesIns_Inst_Sbox_2_T25), .Z(SubBytesIns_Inst_Sbox_2_M23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M24_U1 ( .A(SubBytesIns_Inst_Sbox_2_M22), 
        .B(SubBytesIns_Inst_Sbox_2_M23), .Z(SubBytesIns_Inst_Sbox_2_M24) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M25_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M22), .A2(SubBytesIns_Inst_Sbox_2_M20), .ZN(SubBytesIns_Inst_Sbox_2_M25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M26_U1 ( .A(SubBytesIns_Inst_Sbox_2_M21), 
        .B(SubBytesIns_Inst_Sbox_2_M25), .Z(SubBytesIns_Inst_Sbox_2_M26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M27_U1 ( .A(SubBytesIns_Inst_Sbox_2_M20), 
        .B(SubBytesIns_Inst_Sbox_2_M21), .Z(SubBytesIns_Inst_Sbox_2_M27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M28_U1 ( .A(SubBytesIns_Inst_Sbox_2_M23), 
        .B(SubBytesIns_Inst_Sbox_2_M25), .Z(SubBytesIns_Inst_Sbox_2_M28) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M29_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M28), .A2(SubBytesIns_Inst_Sbox_2_M27), .ZN(SubBytesIns_Inst_Sbox_2_M29) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M30_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M26), .A2(SubBytesIns_Inst_Sbox_2_M24), .ZN(SubBytesIns_Inst_Sbox_2_M30) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M31_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M20), .A2(SubBytesIns_Inst_Sbox_2_M23), .ZN(SubBytesIns_Inst_Sbox_2_M31) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M32_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M27), .A2(SubBytesIns_Inst_Sbox_2_M31), .ZN(SubBytesIns_Inst_Sbox_2_M32) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M33_U1 ( .A(SubBytesIns_Inst_Sbox_2_M27), 
        .B(SubBytesIns_Inst_Sbox_2_M25), .Z(SubBytesIns_Inst_Sbox_2_M33) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M34_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M21), .A2(SubBytesIns_Inst_Sbox_2_M22), .ZN(SubBytesIns_Inst_Sbox_2_M34) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M35_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M24), .A2(SubBytesIns_Inst_Sbox_2_M34), .ZN(SubBytesIns_Inst_Sbox_2_M35) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M36_U1 ( .A(SubBytesIns_Inst_Sbox_2_M24), 
        .B(SubBytesIns_Inst_Sbox_2_M25), .Z(SubBytesIns_Inst_Sbox_2_M36) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M37_U1 ( .A(SubBytesIns_Inst_Sbox_2_M21), 
        .B(SubBytesIns_Inst_Sbox_2_M29), .Z(SubBytesIns_Inst_Sbox_2_M37) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M38_U1 ( .A(SubBytesIns_Inst_Sbox_2_M32), 
        .B(SubBytesIns_Inst_Sbox_2_M33), .Z(SubBytesIns_Inst_Sbox_2_M38) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M39_U1 ( .A(SubBytesIns_Inst_Sbox_2_M23), 
        .B(SubBytesIns_Inst_Sbox_2_M30), .Z(SubBytesIns_Inst_Sbox_2_M39) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M40_U1 ( .A(SubBytesIns_Inst_Sbox_2_M35), 
        .B(SubBytesIns_Inst_Sbox_2_M36), .Z(SubBytesIns_Inst_Sbox_2_M40) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M41_U1 ( .A(SubBytesIns_Inst_Sbox_2_M38), 
        .B(SubBytesIns_Inst_Sbox_2_M40), .Z(SubBytesIns_Inst_Sbox_2_M41) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M42_U1 ( .A(SubBytesIns_Inst_Sbox_2_M37), 
        .B(SubBytesIns_Inst_Sbox_2_M39), .Z(SubBytesIns_Inst_Sbox_2_M42) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M43_U1 ( .A(SubBytesIns_Inst_Sbox_2_M37), 
        .B(SubBytesIns_Inst_Sbox_2_M38), .Z(SubBytesIns_Inst_Sbox_2_M43) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M44_U1 ( .A(SubBytesIns_Inst_Sbox_2_M39), 
        .B(SubBytesIns_Inst_Sbox_2_M40), .Z(SubBytesIns_Inst_Sbox_2_M44) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_M45_U1 ( .A(SubBytesIns_Inst_Sbox_2_M42), 
        .B(SubBytesIns_Inst_Sbox_2_M41), .Z(SubBytesIns_Inst_Sbox_2_M45) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M46_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M44), .A2(SubBytesIns_Inst_Sbox_2_T6), .ZN(SubBytesIns_Inst_Sbox_2_M46) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M47_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M40), .A2(SubBytesIns_Inst_Sbox_2_T8), .ZN(SubBytesIns_Inst_Sbox_2_M47) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M48_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M39), .A2(SubBytesInput[16]), .ZN(SubBytesIns_Inst_Sbox_2_M48) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M49_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M43), .A2(SubBytesIns_Inst_Sbox_2_T16), .ZN(SubBytesIns_Inst_Sbox_2_M49) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M50_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M38), .A2(SubBytesIns_Inst_Sbox_2_T9), .ZN(SubBytesIns_Inst_Sbox_2_M50) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M51_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M37), .A2(SubBytesIns_Inst_Sbox_2_T17), .ZN(SubBytesIns_Inst_Sbox_2_M51) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M52_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M42), .A2(SubBytesIns_Inst_Sbox_2_T15), .ZN(SubBytesIns_Inst_Sbox_2_M52) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M53_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M45), .A2(SubBytesIns_Inst_Sbox_2_T27), .ZN(SubBytesIns_Inst_Sbox_2_M53) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M54_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M41), .A2(SubBytesIns_Inst_Sbox_2_T10), .ZN(SubBytesIns_Inst_Sbox_2_M54) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M55_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M44), .A2(SubBytesIns_Inst_Sbox_2_T13), .ZN(SubBytesIns_Inst_Sbox_2_M55) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M56_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M40), .A2(SubBytesIns_Inst_Sbox_2_T23), .ZN(SubBytesIns_Inst_Sbox_2_M56) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M57_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M39), .A2(SubBytesIns_Inst_Sbox_2_T19), .ZN(SubBytesIns_Inst_Sbox_2_M57) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M58_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M43), .A2(SubBytesIns_Inst_Sbox_2_T3), .ZN(SubBytesIns_Inst_Sbox_2_M58) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M59_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M38), .A2(SubBytesIns_Inst_Sbox_2_T22), .ZN(SubBytesIns_Inst_Sbox_2_M59) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M60_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M37), .A2(SubBytesIns_Inst_Sbox_2_T20), .ZN(SubBytesIns_Inst_Sbox_2_M60) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M61_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M42), .A2(SubBytesIns_Inst_Sbox_2_T1), .ZN(SubBytesIns_Inst_Sbox_2_M61) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M62_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M45), .A2(SubBytesIns_Inst_Sbox_2_T4), .ZN(SubBytesIns_Inst_Sbox_2_M62) );
  AND2_X1 SubBytesIns_Inst_Sbox_2_AND_M63_U1 ( .A1(SubBytesIns_Inst_Sbox_2_M41), .A2(SubBytesIns_Inst_Sbox_2_T2), .ZN(SubBytesIns_Inst_Sbox_2_M63) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L0_U1 ( .A(SubBytesIns_Inst_Sbox_2_M61), 
        .B(SubBytesIns_Inst_Sbox_2_M62), .Z(SubBytesIns_Inst_Sbox_2_L0) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L1_U1 ( .A(SubBytesIns_Inst_Sbox_2_M50), 
        .B(SubBytesIns_Inst_Sbox_2_M56), .Z(SubBytesIns_Inst_Sbox_2_L1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L2_U1 ( .A(SubBytesIns_Inst_Sbox_2_M46), 
        .B(SubBytesIns_Inst_Sbox_2_M48), .Z(SubBytesIns_Inst_Sbox_2_L2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L3_U1 ( .A(SubBytesIns_Inst_Sbox_2_M47), 
        .B(SubBytesIns_Inst_Sbox_2_M55), .Z(SubBytesIns_Inst_Sbox_2_L3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L4_U1 ( .A(SubBytesIns_Inst_Sbox_2_M54), 
        .B(SubBytesIns_Inst_Sbox_2_M58), .Z(SubBytesIns_Inst_Sbox_2_L4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L5_U1 ( .A(SubBytesIns_Inst_Sbox_2_M49), 
        .B(SubBytesIns_Inst_Sbox_2_M61), .Z(SubBytesIns_Inst_Sbox_2_L5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L6_U1 ( .A(SubBytesIns_Inst_Sbox_2_M62), 
        .B(SubBytesIns_Inst_Sbox_2_L5), .Z(SubBytesIns_Inst_Sbox_2_L6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L7_U1 ( .A(SubBytesIns_Inst_Sbox_2_M46), 
        .B(SubBytesIns_Inst_Sbox_2_L3), .Z(SubBytesIns_Inst_Sbox_2_L7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L8_U1 ( .A(SubBytesIns_Inst_Sbox_2_M51), 
        .B(SubBytesIns_Inst_Sbox_2_M59), .Z(SubBytesIns_Inst_Sbox_2_L8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L9_U1 ( .A(SubBytesIns_Inst_Sbox_2_M52), 
        .B(SubBytesIns_Inst_Sbox_2_M53), .Z(SubBytesIns_Inst_Sbox_2_L9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L10_U1 ( .A(SubBytesIns_Inst_Sbox_2_M53), 
        .B(SubBytesIns_Inst_Sbox_2_L4), .Z(SubBytesIns_Inst_Sbox_2_L10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L11_U1 ( .A(SubBytesIns_Inst_Sbox_2_M60), 
        .B(SubBytesIns_Inst_Sbox_2_L2), .Z(SubBytesIns_Inst_Sbox_2_L11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L12_U1 ( .A(SubBytesIns_Inst_Sbox_2_M48), 
        .B(SubBytesIns_Inst_Sbox_2_M51), .Z(SubBytesIns_Inst_Sbox_2_L12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L13_U1 ( .A(SubBytesIns_Inst_Sbox_2_M50), 
        .B(SubBytesIns_Inst_Sbox_2_L0), .Z(SubBytesIns_Inst_Sbox_2_L13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L14_U1 ( .A(SubBytesIns_Inst_Sbox_2_M52), 
        .B(SubBytesIns_Inst_Sbox_2_M61), .Z(SubBytesIns_Inst_Sbox_2_L14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L15_U1 ( .A(SubBytesIns_Inst_Sbox_2_M55), 
        .B(SubBytesIns_Inst_Sbox_2_L1), .Z(SubBytesIns_Inst_Sbox_2_L15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L16_U1 ( .A(SubBytesIns_Inst_Sbox_2_M56), 
        .B(SubBytesIns_Inst_Sbox_2_L0), .Z(SubBytesIns_Inst_Sbox_2_L16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L17_U1 ( .A(SubBytesIns_Inst_Sbox_2_M57), 
        .B(SubBytesIns_Inst_Sbox_2_L1), .Z(SubBytesIns_Inst_Sbox_2_L17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L18_U1 ( .A(SubBytesIns_Inst_Sbox_2_M58), 
        .B(SubBytesIns_Inst_Sbox_2_L8), .Z(SubBytesIns_Inst_Sbox_2_L18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L19_U1 ( .A(SubBytesIns_Inst_Sbox_2_M63), 
        .B(SubBytesIns_Inst_Sbox_2_L4), .Z(SubBytesIns_Inst_Sbox_2_L19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L20_U1 ( .A(SubBytesIns_Inst_Sbox_2_L0), 
        .B(SubBytesIns_Inst_Sbox_2_L1), .Z(SubBytesIns_Inst_Sbox_2_L20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L21_U1 ( .A(SubBytesIns_Inst_Sbox_2_L1), 
        .B(SubBytesIns_Inst_Sbox_2_L7), .Z(SubBytesIns_Inst_Sbox_2_L21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L22_U1 ( .A(SubBytesIns_Inst_Sbox_2_L3), 
        .B(SubBytesIns_Inst_Sbox_2_L12), .Z(SubBytesIns_Inst_Sbox_2_L22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L23_U1 ( .A(SubBytesIns_Inst_Sbox_2_L18), 
        .B(SubBytesIns_Inst_Sbox_2_L2), .Z(SubBytesIns_Inst_Sbox_2_L23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L24_U1 ( .A(SubBytesIns_Inst_Sbox_2_L15), 
        .B(SubBytesIns_Inst_Sbox_2_L9), .Z(SubBytesIns_Inst_Sbox_2_L24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L25_U1 ( .A(SubBytesIns_Inst_Sbox_2_L6), 
        .B(SubBytesIns_Inst_Sbox_2_L10), .Z(SubBytesIns_Inst_Sbox_2_L25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L26_U1 ( .A(SubBytesIns_Inst_Sbox_2_L7), 
        .B(SubBytesIns_Inst_Sbox_2_L9), .Z(SubBytesIns_Inst_Sbox_2_L26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L27_U1 ( .A(SubBytesIns_Inst_Sbox_2_L8), 
        .B(SubBytesIns_Inst_Sbox_2_L10), .Z(SubBytesIns_Inst_Sbox_2_L27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L28_U1 ( .A(SubBytesIns_Inst_Sbox_2_L11), 
        .B(SubBytesIns_Inst_Sbox_2_L14), .Z(SubBytesIns_Inst_Sbox_2_L28) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_L29_U1 ( .A(SubBytesIns_Inst_Sbox_2_L11), 
        .B(SubBytesIns_Inst_Sbox_2_L17), .Z(SubBytesIns_Inst_Sbox_2_L29) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_S0_U1 ( .A(SubBytesIns_Inst_Sbox_2_L6), 
        .B(SubBytesIns_Inst_Sbox_2_L24), .Z(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_S1_U1 ( .A(SubBytesIns_Inst_Sbox_2_L16), 
        .B(SubBytesIns_Inst_Sbox_2_L26), .ZN(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[23]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_S2_U1 ( .A(SubBytesIns_Inst_Sbox_2_L19), 
        .B(SubBytesIns_Inst_Sbox_2_L28), .ZN(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[22]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_S3_U1 ( .A(SubBytesIns_Inst_Sbox_2_L6), 
        .B(SubBytesIns_Inst_Sbox_2_L21), .Z(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[21]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_S4_U1 ( .A(SubBytesIns_Inst_Sbox_2_L20), 
        .B(SubBytesIns_Inst_Sbox_2_L22), .Z(MixColumnsInput[51]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_S5_U1 ( .A(SubBytesIns_Inst_Sbox_2_L25), 
        .B(SubBytesIns_Inst_Sbox_2_L29), .Z(MixColumnsInput[50]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_S6_U1 ( .A(SubBytesIns_Inst_Sbox_2_L13), 
        .B(SubBytesIns_Inst_Sbox_2_L27), .ZN(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[18]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_2_XOR_S7_U1 ( .A(SubBytesIns_Inst_Sbox_2_L6), 
        .B(SubBytesIns_Inst_Sbox_2_L23), .ZN(MixColumnsInput[48]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T1_U1 ( .A(SubBytesInput[31]), .B(
        SubBytesInput[28]), .Z(SubBytesIns_Inst_Sbox_3_T1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T2_U1 ( .A(SubBytesInput[31]), .B(
        SubBytesInput[26]), .Z(SubBytesIns_Inst_Sbox_3_T2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T3_U1 ( .A(SubBytesInput[31]), .B(
        SubBytesInput[25]), .Z(SubBytesIns_Inst_Sbox_3_T3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T4_U1 ( .A(SubBytesInput[28]), .B(
        SubBytesInput[26]), .Z(SubBytesIns_Inst_Sbox_3_T4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T5_U1 ( .A(SubBytesInput[27]), .B(
        SubBytesInput[25]), .Z(SubBytesIns_Inst_Sbox_3_T5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T6_U1 ( .A(SubBytesIns_Inst_Sbox_3_T1), 
        .B(SubBytesIns_Inst_Sbox_3_T5), .Z(SubBytesIns_Inst_Sbox_3_T6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T7_U1 ( .A(SubBytesInput[30]), .B(
        SubBytesInput[29]), .Z(SubBytesIns_Inst_Sbox_3_T7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T8_U1 ( .A(SubBytesInput[24]), .B(
        SubBytesIns_Inst_Sbox_3_T6), .Z(SubBytesIns_Inst_Sbox_3_T8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T9_U1 ( .A(SubBytesInput[24]), .B(
        SubBytesIns_Inst_Sbox_3_T7), .Z(SubBytesIns_Inst_Sbox_3_T9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T10_U1 ( .A(SubBytesIns_Inst_Sbox_3_T6), 
        .B(SubBytesIns_Inst_Sbox_3_T7), .Z(SubBytesIns_Inst_Sbox_3_T10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T11_U1 ( .A(SubBytesInput[30]), .B(
        SubBytesInput[26]), .Z(SubBytesIns_Inst_Sbox_3_T11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T12_U1 ( .A(SubBytesInput[29]), .B(
        SubBytesInput[26]), .Z(SubBytesIns_Inst_Sbox_3_T12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T13_U1 ( .A(SubBytesIns_Inst_Sbox_3_T3), 
        .B(SubBytesIns_Inst_Sbox_3_T4), .Z(SubBytesIns_Inst_Sbox_3_T13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T14_U1 ( .A(SubBytesIns_Inst_Sbox_3_T6), 
        .B(SubBytesIns_Inst_Sbox_3_T11), .Z(SubBytesIns_Inst_Sbox_3_T14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T15_U1 ( .A(SubBytesIns_Inst_Sbox_3_T5), 
        .B(SubBytesIns_Inst_Sbox_3_T11), .Z(SubBytesIns_Inst_Sbox_3_T15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T16_U1 ( .A(SubBytesIns_Inst_Sbox_3_T5), 
        .B(SubBytesIns_Inst_Sbox_3_T12), .Z(SubBytesIns_Inst_Sbox_3_T16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T17_U1 ( .A(SubBytesIns_Inst_Sbox_3_T9), 
        .B(SubBytesIns_Inst_Sbox_3_T16), .Z(SubBytesIns_Inst_Sbox_3_T17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T18_U1 ( .A(SubBytesInput[28]), .B(
        SubBytesInput[24]), .Z(SubBytesIns_Inst_Sbox_3_T18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T19_U1 ( .A(SubBytesIns_Inst_Sbox_3_T7), 
        .B(SubBytesIns_Inst_Sbox_3_T18), .Z(SubBytesIns_Inst_Sbox_3_T19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T20_U1 ( .A(SubBytesIns_Inst_Sbox_3_T1), 
        .B(SubBytesIns_Inst_Sbox_3_T19), .Z(SubBytesIns_Inst_Sbox_3_T20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T21_U1 ( .A(SubBytesInput[25]), .B(
        SubBytesInput[24]), .Z(SubBytesIns_Inst_Sbox_3_T21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T22_U1 ( .A(SubBytesIns_Inst_Sbox_3_T7), 
        .B(SubBytesIns_Inst_Sbox_3_T21), .Z(SubBytesIns_Inst_Sbox_3_T22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T23_U1 ( .A(SubBytesIns_Inst_Sbox_3_T2), 
        .B(SubBytesIns_Inst_Sbox_3_T22), .Z(SubBytesIns_Inst_Sbox_3_T23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T24_U1 ( .A(SubBytesIns_Inst_Sbox_3_T2), 
        .B(SubBytesIns_Inst_Sbox_3_T10), .Z(SubBytesIns_Inst_Sbox_3_T24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T25_U1 ( .A(SubBytesIns_Inst_Sbox_3_T20), 
        .B(SubBytesIns_Inst_Sbox_3_T17), .Z(SubBytesIns_Inst_Sbox_3_T25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T26_U1 ( .A(SubBytesIns_Inst_Sbox_3_T3), 
        .B(SubBytesIns_Inst_Sbox_3_T16), .Z(SubBytesIns_Inst_Sbox_3_T26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_T27_U1 ( .A(SubBytesIns_Inst_Sbox_3_T1), 
        .B(SubBytesIns_Inst_Sbox_3_T12), .Z(SubBytesIns_Inst_Sbox_3_T27) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M1_U1 ( .A1(SubBytesIns_Inst_Sbox_3_T13), 
        .A2(SubBytesIns_Inst_Sbox_3_T6), .ZN(SubBytesIns_Inst_Sbox_3_M1) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M2_U1 ( .A1(SubBytesIns_Inst_Sbox_3_T23), 
        .A2(SubBytesIns_Inst_Sbox_3_T8), .ZN(SubBytesIns_Inst_Sbox_3_M2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M3_U1 ( .A(SubBytesIns_Inst_Sbox_3_T14), 
        .B(SubBytesIns_Inst_Sbox_3_M1), .Z(SubBytesIns_Inst_Sbox_3_M3) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M4_U1 ( .A1(SubBytesIns_Inst_Sbox_3_T19), 
        .A2(SubBytesInput[24]), .ZN(SubBytesIns_Inst_Sbox_3_M4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M5_U1 ( .A(SubBytesIns_Inst_Sbox_3_M4), 
        .B(SubBytesIns_Inst_Sbox_3_M1), .Z(SubBytesIns_Inst_Sbox_3_M5) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M6_U1 ( .A1(SubBytesIns_Inst_Sbox_3_T3), 
        .A2(SubBytesIns_Inst_Sbox_3_T16), .ZN(SubBytesIns_Inst_Sbox_3_M6) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M7_U1 ( .A1(SubBytesIns_Inst_Sbox_3_T22), 
        .A2(SubBytesIns_Inst_Sbox_3_T9), .ZN(SubBytesIns_Inst_Sbox_3_M7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M8_U1 ( .A(SubBytesIns_Inst_Sbox_3_T26), 
        .B(SubBytesIns_Inst_Sbox_3_M6), .Z(SubBytesIns_Inst_Sbox_3_M8) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M9_U1 ( .A1(SubBytesIns_Inst_Sbox_3_T20), 
        .A2(SubBytesIns_Inst_Sbox_3_T17), .ZN(SubBytesIns_Inst_Sbox_3_M9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M10_U1 ( .A(SubBytesIns_Inst_Sbox_3_M9), 
        .B(SubBytesIns_Inst_Sbox_3_M6), .Z(SubBytesIns_Inst_Sbox_3_M10) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M11_U1 ( .A1(SubBytesIns_Inst_Sbox_3_T1), 
        .A2(SubBytesIns_Inst_Sbox_3_T15), .ZN(SubBytesIns_Inst_Sbox_3_M11) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M12_U1 ( .A1(SubBytesIns_Inst_Sbox_3_T4), 
        .A2(SubBytesIns_Inst_Sbox_3_T27), .ZN(SubBytesIns_Inst_Sbox_3_M12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M13_U1 ( .A(SubBytesIns_Inst_Sbox_3_M12), 
        .B(SubBytesIns_Inst_Sbox_3_M11), .Z(SubBytesIns_Inst_Sbox_3_M13) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M14_U1 ( .A1(SubBytesIns_Inst_Sbox_3_T2), 
        .A2(SubBytesIns_Inst_Sbox_3_T10), .ZN(SubBytesIns_Inst_Sbox_3_M14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M15_U1 ( .A(SubBytesIns_Inst_Sbox_3_M14), 
        .B(SubBytesIns_Inst_Sbox_3_M11), .Z(SubBytesIns_Inst_Sbox_3_M15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M16_U1 ( .A(SubBytesIns_Inst_Sbox_3_M3), 
        .B(SubBytesIns_Inst_Sbox_3_M2), .Z(SubBytesIns_Inst_Sbox_3_M16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M17_U1 ( .A(SubBytesIns_Inst_Sbox_3_M5), 
        .B(SubBytesIns_Inst_Sbox_3_T24), .Z(SubBytesIns_Inst_Sbox_3_M17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M18_U1 ( .A(SubBytesIns_Inst_Sbox_3_M8), 
        .B(SubBytesIns_Inst_Sbox_3_M7), .Z(SubBytesIns_Inst_Sbox_3_M18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M19_U1 ( .A(SubBytesIns_Inst_Sbox_3_M10), 
        .B(SubBytesIns_Inst_Sbox_3_M15), .Z(SubBytesIns_Inst_Sbox_3_M19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M20_U1 ( .A(SubBytesIns_Inst_Sbox_3_M16), 
        .B(SubBytesIns_Inst_Sbox_3_M13), .Z(SubBytesIns_Inst_Sbox_3_M20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M21_U1 ( .A(SubBytesIns_Inst_Sbox_3_M17), 
        .B(SubBytesIns_Inst_Sbox_3_M15), .Z(SubBytesIns_Inst_Sbox_3_M21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M22_U1 ( .A(SubBytesIns_Inst_Sbox_3_M18), 
        .B(SubBytesIns_Inst_Sbox_3_M13), .Z(SubBytesIns_Inst_Sbox_3_M22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M23_U1 ( .A(SubBytesIns_Inst_Sbox_3_M19), 
        .B(SubBytesIns_Inst_Sbox_3_T25), .Z(SubBytesIns_Inst_Sbox_3_M23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M24_U1 ( .A(SubBytesIns_Inst_Sbox_3_M22), 
        .B(SubBytesIns_Inst_Sbox_3_M23), .Z(SubBytesIns_Inst_Sbox_3_M24) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M25_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M22), .A2(SubBytesIns_Inst_Sbox_3_M20), .ZN(SubBytesIns_Inst_Sbox_3_M25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M26_U1 ( .A(SubBytesIns_Inst_Sbox_3_M21), 
        .B(SubBytesIns_Inst_Sbox_3_M25), .Z(SubBytesIns_Inst_Sbox_3_M26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M27_U1 ( .A(SubBytesIns_Inst_Sbox_3_M20), 
        .B(SubBytesIns_Inst_Sbox_3_M21), .Z(SubBytesIns_Inst_Sbox_3_M27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M28_U1 ( .A(SubBytesIns_Inst_Sbox_3_M23), 
        .B(SubBytesIns_Inst_Sbox_3_M25), .Z(SubBytesIns_Inst_Sbox_3_M28) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M29_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M28), .A2(SubBytesIns_Inst_Sbox_3_M27), .ZN(SubBytesIns_Inst_Sbox_3_M29) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M30_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M26), .A2(SubBytesIns_Inst_Sbox_3_M24), .ZN(SubBytesIns_Inst_Sbox_3_M30) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M31_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M20), .A2(SubBytesIns_Inst_Sbox_3_M23), .ZN(SubBytesIns_Inst_Sbox_3_M31) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M32_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M27), .A2(SubBytesIns_Inst_Sbox_3_M31), .ZN(SubBytesIns_Inst_Sbox_3_M32) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M33_U1 ( .A(SubBytesIns_Inst_Sbox_3_M27), 
        .B(SubBytesIns_Inst_Sbox_3_M25), .Z(SubBytesIns_Inst_Sbox_3_M33) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M34_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M21), .A2(SubBytesIns_Inst_Sbox_3_M22), .ZN(SubBytesIns_Inst_Sbox_3_M34) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M35_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M24), .A2(SubBytesIns_Inst_Sbox_3_M34), .ZN(SubBytesIns_Inst_Sbox_3_M35) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M36_U1 ( .A(SubBytesIns_Inst_Sbox_3_M24), 
        .B(SubBytesIns_Inst_Sbox_3_M25), .Z(SubBytesIns_Inst_Sbox_3_M36) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M37_U1 ( .A(SubBytesIns_Inst_Sbox_3_M21), 
        .B(SubBytesIns_Inst_Sbox_3_M29), .Z(SubBytesIns_Inst_Sbox_3_M37) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M38_U1 ( .A(SubBytesIns_Inst_Sbox_3_M32), 
        .B(SubBytesIns_Inst_Sbox_3_M33), .Z(SubBytesIns_Inst_Sbox_3_M38) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M39_U1 ( .A(SubBytesIns_Inst_Sbox_3_M23), 
        .B(SubBytesIns_Inst_Sbox_3_M30), .Z(SubBytesIns_Inst_Sbox_3_M39) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M40_U1 ( .A(SubBytesIns_Inst_Sbox_3_M35), 
        .B(SubBytesIns_Inst_Sbox_3_M36), .Z(SubBytesIns_Inst_Sbox_3_M40) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M41_U1 ( .A(SubBytesIns_Inst_Sbox_3_M38), 
        .B(SubBytesIns_Inst_Sbox_3_M40), .Z(SubBytesIns_Inst_Sbox_3_M41) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M42_U1 ( .A(SubBytesIns_Inst_Sbox_3_M37), 
        .B(SubBytesIns_Inst_Sbox_3_M39), .Z(SubBytesIns_Inst_Sbox_3_M42) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M43_U1 ( .A(SubBytesIns_Inst_Sbox_3_M37), 
        .B(SubBytesIns_Inst_Sbox_3_M38), .Z(SubBytesIns_Inst_Sbox_3_M43) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M44_U1 ( .A(SubBytesIns_Inst_Sbox_3_M39), 
        .B(SubBytesIns_Inst_Sbox_3_M40), .Z(SubBytesIns_Inst_Sbox_3_M44) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_M45_U1 ( .A(SubBytesIns_Inst_Sbox_3_M42), 
        .B(SubBytesIns_Inst_Sbox_3_M41), .Z(SubBytesIns_Inst_Sbox_3_M45) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M46_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M44), .A2(SubBytesIns_Inst_Sbox_3_T6), .ZN(SubBytesIns_Inst_Sbox_3_M46) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M47_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M40), .A2(SubBytesIns_Inst_Sbox_3_T8), .ZN(SubBytesIns_Inst_Sbox_3_M47) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M48_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M39), .A2(SubBytesInput[24]), .ZN(SubBytesIns_Inst_Sbox_3_M48) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M49_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M43), .A2(SubBytesIns_Inst_Sbox_3_T16), .ZN(SubBytesIns_Inst_Sbox_3_M49) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M50_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M38), .A2(SubBytesIns_Inst_Sbox_3_T9), .ZN(SubBytesIns_Inst_Sbox_3_M50) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M51_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M37), .A2(SubBytesIns_Inst_Sbox_3_T17), .ZN(SubBytesIns_Inst_Sbox_3_M51) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M52_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M42), .A2(SubBytesIns_Inst_Sbox_3_T15), .ZN(SubBytesIns_Inst_Sbox_3_M52) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M53_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M45), .A2(SubBytesIns_Inst_Sbox_3_T27), .ZN(SubBytesIns_Inst_Sbox_3_M53) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M54_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M41), .A2(SubBytesIns_Inst_Sbox_3_T10), .ZN(SubBytesIns_Inst_Sbox_3_M54) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M55_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M44), .A2(SubBytesIns_Inst_Sbox_3_T13), .ZN(SubBytesIns_Inst_Sbox_3_M55) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M56_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M40), .A2(SubBytesIns_Inst_Sbox_3_T23), .ZN(SubBytesIns_Inst_Sbox_3_M56) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M57_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M39), .A2(SubBytesIns_Inst_Sbox_3_T19), .ZN(SubBytesIns_Inst_Sbox_3_M57) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M58_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M43), .A2(SubBytesIns_Inst_Sbox_3_T3), .ZN(SubBytesIns_Inst_Sbox_3_M58) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M59_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M38), .A2(SubBytesIns_Inst_Sbox_3_T22), .ZN(SubBytesIns_Inst_Sbox_3_M59) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M60_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M37), .A2(SubBytesIns_Inst_Sbox_3_T20), .ZN(SubBytesIns_Inst_Sbox_3_M60) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M61_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M42), .A2(SubBytesIns_Inst_Sbox_3_T1), .ZN(SubBytesIns_Inst_Sbox_3_M61) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M62_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M45), .A2(SubBytesIns_Inst_Sbox_3_T4), .ZN(SubBytesIns_Inst_Sbox_3_M62) );
  AND2_X1 SubBytesIns_Inst_Sbox_3_AND_M63_U1 ( .A1(SubBytesIns_Inst_Sbox_3_M41), .A2(SubBytesIns_Inst_Sbox_3_T2), .ZN(SubBytesIns_Inst_Sbox_3_M63) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L0_U1 ( .A(SubBytesIns_Inst_Sbox_3_M61), 
        .B(SubBytesIns_Inst_Sbox_3_M62), .Z(SubBytesIns_Inst_Sbox_3_L0) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L1_U1 ( .A(SubBytesIns_Inst_Sbox_3_M50), 
        .B(SubBytesIns_Inst_Sbox_3_M56), .Z(SubBytesIns_Inst_Sbox_3_L1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L2_U1 ( .A(SubBytesIns_Inst_Sbox_3_M46), 
        .B(SubBytesIns_Inst_Sbox_3_M48), .Z(SubBytesIns_Inst_Sbox_3_L2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L3_U1 ( .A(SubBytesIns_Inst_Sbox_3_M47), 
        .B(SubBytesIns_Inst_Sbox_3_M55), .Z(SubBytesIns_Inst_Sbox_3_L3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L4_U1 ( .A(SubBytesIns_Inst_Sbox_3_M54), 
        .B(SubBytesIns_Inst_Sbox_3_M58), .Z(SubBytesIns_Inst_Sbox_3_L4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L5_U1 ( .A(SubBytesIns_Inst_Sbox_3_M49), 
        .B(SubBytesIns_Inst_Sbox_3_M61), .Z(SubBytesIns_Inst_Sbox_3_L5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L6_U1 ( .A(SubBytesIns_Inst_Sbox_3_M62), 
        .B(SubBytesIns_Inst_Sbox_3_L5), .Z(SubBytesIns_Inst_Sbox_3_L6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L7_U1 ( .A(SubBytesIns_Inst_Sbox_3_M46), 
        .B(SubBytesIns_Inst_Sbox_3_L3), .Z(SubBytesIns_Inst_Sbox_3_L7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L8_U1 ( .A(SubBytesIns_Inst_Sbox_3_M51), 
        .B(SubBytesIns_Inst_Sbox_3_M59), .Z(SubBytesIns_Inst_Sbox_3_L8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L9_U1 ( .A(SubBytesIns_Inst_Sbox_3_M52), 
        .B(SubBytesIns_Inst_Sbox_3_M53), .Z(SubBytesIns_Inst_Sbox_3_L9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L10_U1 ( .A(SubBytesIns_Inst_Sbox_3_M53), 
        .B(SubBytesIns_Inst_Sbox_3_L4), .Z(SubBytesIns_Inst_Sbox_3_L10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L11_U1 ( .A(SubBytesIns_Inst_Sbox_3_M60), 
        .B(SubBytesIns_Inst_Sbox_3_L2), .Z(SubBytesIns_Inst_Sbox_3_L11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L12_U1 ( .A(SubBytesIns_Inst_Sbox_3_M48), 
        .B(SubBytesIns_Inst_Sbox_3_M51), .Z(SubBytesIns_Inst_Sbox_3_L12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L13_U1 ( .A(SubBytesIns_Inst_Sbox_3_M50), 
        .B(SubBytesIns_Inst_Sbox_3_L0), .Z(SubBytesIns_Inst_Sbox_3_L13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L14_U1 ( .A(SubBytesIns_Inst_Sbox_3_M52), 
        .B(SubBytesIns_Inst_Sbox_3_M61), .Z(SubBytesIns_Inst_Sbox_3_L14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L15_U1 ( .A(SubBytesIns_Inst_Sbox_3_M55), 
        .B(SubBytesIns_Inst_Sbox_3_L1), .Z(SubBytesIns_Inst_Sbox_3_L15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L16_U1 ( .A(SubBytesIns_Inst_Sbox_3_M56), 
        .B(SubBytesIns_Inst_Sbox_3_L0), .Z(SubBytesIns_Inst_Sbox_3_L16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L17_U1 ( .A(SubBytesIns_Inst_Sbox_3_M57), 
        .B(SubBytesIns_Inst_Sbox_3_L1), .Z(SubBytesIns_Inst_Sbox_3_L17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L18_U1 ( .A(SubBytesIns_Inst_Sbox_3_M58), 
        .B(SubBytesIns_Inst_Sbox_3_L8), .Z(SubBytesIns_Inst_Sbox_3_L18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L19_U1 ( .A(SubBytesIns_Inst_Sbox_3_M63), 
        .B(SubBytesIns_Inst_Sbox_3_L4), .Z(SubBytesIns_Inst_Sbox_3_L19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L20_U1 ( .A(SubBytesIns_Inst_Sbox_3_L0), 
        .B(SubBytesIns_Inst_Sbox_3_L1), .Z(SubBytesIns_Inst_Sbox_3_L20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L21_U1 ( .A(SubBytesIns_Inst_Sbox_3_L1), 
        .B(SubBytesIns_Inst_Sbox_3_L7), .Z(SubBytesIns_Inst_Sbox_3_L21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L22_U1 ( .A(SubBytesIns_Inst_Sbox_3_L3), 
        .B(SubBytesIns_Inst_Sbox_3_L12), .Z(SubBytesIns_Inst_Sbox_3_L22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L23_U1 ( .A(SubBytesIns_Inst_Sbox_3_L18), 
        .B(SubBytesIns_Inst_Sbox_3_L2), .Z(SubBytesIns_Inst_Sbox_3_L23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L24_U1 ( .A(SubBytesIns_Inst_Sbox_3_L15), 
        .B(SubBytesIns_Inst_Sbox_3_L9), .Z(SubBytesIns_Inst_Sbox_3_L24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L25_U1 ( .A(SubBytesIns_Inst_Sbox_3_L6), 
        .B(SubBytesIns_Inst_Sbox_3_L10), .Z(SubBytesIns_Inst_Sbox_3_L25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L26_U1 ( .A(SubBytesIns_Inst_Sbox_3_L7), 
        .B(SubBytesIns_Inst_Sbox_3_L9), .Z(SubBytesIns_Inst_Sbox_3_L26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L27_U1 ( .A(SubBytesIns_Inst_Sbox_3_L8), 
        .B(SubBytesIns_Inst_Sbox_3_L10), .Z(SubBytesIns_Inst_Sbox_3_L27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L28_U1 ( .A(SubBytesIns_Inst_Sbox_3_L11), 
        .B(SubBytesIns_Inst_Sbox_3_L14), .Z(SubBytesIns_Inst_Sbox_3_L28) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_L29_U1 ( .A(SubBytesIns_Inst_Sbox_3_L11), 
        .B(SubBytesIns_Inst_Sbox_3_L17), .Z(SubBytesIns_Inst_Sbox_3_L29) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_S0_U1 ( .A(SubBytesIns_Inst_Sbox_3_L6), 
        .B(SubBytesIns_Inst_Sbox_3_L24), .Z(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_S1_U1 ( .A(SubBytesIns_Inst_Sbox_3_L16), 
        .B(SubBytesIns_Inst_Sbox_3_L26), .ZN(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[31]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_S2_U1 ( .A(SubBytesIns_Inst_Sbox_3_L19), 
        .B(SubBytesIns_Inst_Sbox_3_L28), .ZN(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[30]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_S3_U1 ( .A(SubBytesIns_Inst_Sbox_3_L6), 
        .B(SubBytesIns_Inst_Sbox_3_L21), .Z(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[29]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_S4_U1 ( .A(SubBytesIns_Inst_Sbox_3_L20), 
        .B(SubBytesIns_Inst_Sbox_3_L22), .Z(MixColumnsInput[27]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_S5_U1 ( .A(SubBytesIns_Inst_Sbox_3_L25), 
        .B(SubBytesIns_Inst_Sbox_3_L29), .Z(MixColumnsInput[26]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_S6_U1 ( .A(SubBytesIns_Inst_Sbox_3_L13), 
        .B(SubBytesIns_Inst_Sbox_3_L27), .ZN(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[26]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_3_XOR_S7_U1 ( .A(SubBytesIns_Inst_Sbox_3_L6), 
        .B(SubBytesIns_Inst_Sbox_3_L23), .ZN(MixColumnsInput[24]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_T1_U1 ( .A(SubBytesInput[39]), .B(
        SubBytesInput[36]), .Z(SubBytesIns_Inst_Sbox_4_T1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_T2_U1 ( .A(SubBytesInput[39]), .B(
        SubBytesInput[34]), .Z(SubBytesIns_Inst_Sbox_4_T2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_T3_U1 ( .A(SubBytesInput[39]), .B(
        SubBytesInput[33]), .Z(SubBytesIns_Inst_Sbox_4_T3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_T4_U1 ( .A(SubBytesInput[36]), .B(
        SubBytesInput[34]), .Z(SubBytesIns_Inst_Sbox_4_T4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_T5_U1 ( .A(SubBytesInput[35]), .B(
        SubBytesInput[33]), .Z(SubBytesIns_Inst_Sbox_4_T5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_T6_U1 ( .A(SubBytesIns_Inst_Sbox_4_T1), 
        .B(SubBytesIns_Inst_Sbox_4_T5), .Z(SubBytesIns_Inst_Sbox_4_T6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_T7_U1 ( .A(SubBytesInput[38]), .B(
        SubBytesInput[37]), .Z(SubBytesIns_Inst_Sbox_4_T7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_T8_U1 ( .A(SubBytesInput[32]), .B(
        SubBytesIns_Inst_Sbox_4_T6), .Z(SubBytesIns_Inst_Sbox_4_T8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_T9_U1 ( .A(SubBytesInput[32]), .B(
        SubBytesIns_Inst_Sbox_4_T7), .Z(SubBytesIns_Inst_Sbox_4_T9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_T10_U1 ( .A(SubBytesIns_Inst_Sbox_4_T6), 
        .B(SubBytesIns_Inst_Sbox_4_T7), .Z(SubBytesIns_Inst_Sbox_4_T10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_T11_U1 ( .A(SubBytesInput[38]), .B(
        SubBytesInput[34]), .Z(SubBytesIns_Inst_Sbox_4_T11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_T12_U1 ( .A(SubBytesInput[37]), .B(
        SubBytesInput[34]), .Z(SubBytesIns_Inst_Sbox_4_T12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_T13_U1 ( .A(SubBytesIns_Inst_Sbox_4_T3), 
        .B(SubBytesIns_Inst_Sbox_4_T4), .Z(SubBytesIns_Inst_Sbox_4_T13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_T14_U1 ( .A(SubBytesIns_Inst_Sbox_4_T6), 
        .B(SubBytesIns_Inst_Sbox_4_T11), .Z(SubBytesIns_Inst_Sbox_4_T14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_T15_U1 ( .A(SubBytesIns_Inst_Sbox_4_T5), 
        .B(SubBytesIns_Inst_Sbox_4_T11), .Z(SubBytesIns_Inst_Sbox_4_T15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_T16_U1 ( .A(SubBytesIns_Inst_Sbox_4_T5), 
        .B(SubBytesIns_Inst_Sbox_4_T12), .Z(SubBytesIns_Inst_Sbox_4_T16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_T17_U1 ( .A(SubBytesIns_Inst_Sbox_4_T9), 
        .B(SubBytesIns_Inst_Sbox_4_T16), .Z(SubBytesIns_Inst_Sbox_4_T17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_T18_U1 ( .A(SubBytesInput[36]), .B(
        SubBytesInput[32]), .Z(SubBytesIns_Inst_Sbox_4_T18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_T19_U1 ( .A(SubBytesIns_Inst_Sbox_4_T7), 
        .B(SubBytesIns_Inst_Sbox_4_T18), .Z(SubBytesIns_Inst_Sbox_4_T19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_T20_U1 ( .A(SubBytesIns_Inst_Sbox_4_T1), 
        .B(SubBytesIns_Inst_Sbox_4_T19), .Z(SubBytesIns_Inst_Sbox_4_T20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_T21_U1 ( .A(SubBytesInput[33]), .B(
        SubBytesInput[32]), .Z(SubBytesIns_Inst_Sbox_4_T21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_T22_U1 ( .A(SubBytesIns_Inst_Sbox_4_T7), 
        .B(SubBytesIns_Inst_Sbox_4_T21), .Z(SubBytesIns_Inst_Sbox_4_T22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_T23_U1 ( .A(SubBytesIns_Inst_Sbox_4_T2), 
        .B(SubBytesIns_Inst_Sbox_4_T22), .Z(SubBytesIns_Inst_Sbox_4_T23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_T24_U1 ( .A(SubBytesIns_Inst_Sbox_4_T2), 
        .B(SubBytesIns_Inst_Sbox_4_T10), .Z(SubBytesIns_Inst_Sbox_4_T24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_T25_U1 ( .A(SubBytesIns_Inst_Sbox_4_T20), 
        .B(SubBytesIns_Inst_Sbox_4_T17), .Z(SubBytesIns_Inst_Sbox_4_T25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_T26_U1 ( .A(SubBytesIns_Inst_Sbox_4_T3), 
        .B(SubBytesIns_Inst_Sbox_4_T16), .Z(SubBytesIns_Inst_Sbox_4_T26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_T27_U1 ( .A(SubBytesIns_Inst_Sbox_4_T1), 
        .B(SubBytesIns_Inst_Sbox_4_T12), .Z(SubBytesIns_Inst_Sbox_4_T27) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M1_U1 ( .A1(SubBytesIns_Inst_Sbox_4_T13), 
        .A2(SubBytesIns_Inst_Sbox_4_T6), .ZN(SubBytesIns_Inst_Sbox_4_M1) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M2_U1 ( .A1(SubBytesIns_Inst_Sbox_4_T23), 
        .A2(SubBytesIns_Inst_Sbox_4_T8), .ZN(SubBytesIns_Inst_Sbox_4_M2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_M3_U1 ( .A(SubBytesIns_Inst_Sbox_4_T14), 
        .B(SubBytesIns_Inst_Sbox_4_M1), .Z(SubBytesIns_Inst_Sbox_4_M3) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M4_U1 ( .A1(SubBytesIns_Inst_Sbox_4_T19), 
        .A2(SubBytesInput[32]), .ZN(SubBytesIns_Inst_Sbox_4_M4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_M5_U1 ( .A(SubBytesIns_Inst_Sbox_4_M4), 
        .B(SubBytesIns_Inst_Sbox_4_M1), .Z(SubBytesIns_Inst_Sbox_4_M5) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M6_U1 ( .A1(SubBytesIns_Inst_Sbox_4_T3), 
        .A2(SubBytesIns_Inst_Sbox_4_T16), .ZN(SubBytesIns_Inst_Sbox_4_M6) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M7_U1 ( .A1(SubBytesIns_Inst_Sbox_4_T22), 
        .A2(SubBytesIns_Inst_Sbox_4_T9), .ZN(SubBytesIns_Inst_Sbox_4_M7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_M8_U1 ( .A(SubBytesIns_Inst_Sbox_4_T26), 
        .B(SubBytesIns_Inst_Sbox_4_M6), .Z(SubBytesIns_Inst_Sbox_4_M8) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M9_U1 ( .A1(SubBytesIns_Inst_Sbox_4_T20), 
        .A2(SubBytesIns_Inst_Sbox_4_T17), .ZN(SubBytesIns_Inst_Sbox_4_M9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_M10_U1 ( .A(SubBytesIns_Inst_Sbox_4_M9), 
        .B(SubBytesIns_Inst_Sbox_4_M6), .Z(SubBytesIns_Inst_Sbox_4_M10) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M11_U1 ( .A1(SubBytesIns_Inst_Sbox_4_T1), 
        .A2(SubBytesIns_Inst_Sbox_4_T15), .ZN(SubBytesIns_Inst_Sbox_4_M11) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M12_U1 ( .A1(SubBytesIns_Inst_Sbox_4_T4), 
        .A2(SubBytesIns_Inst_Sbox_4_T27), .ZN(SubBytesIns_Inst_Sbox_4_M12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_M13_U1 ( .A(SubBytesIns_Inst_Sbox_4_M12), 
        .B(SubBytesIns_Inst_Sbox_4_M11), .Z(SubBytesIns_Inst_Sbox_4_M13) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M14_U1 ( .A1(SubBytesIns_Inst_Sbox_4_T2), 
        .A2(SubBytesIns_Inst_Sbox_4_T10), .ZN(SubBytesIns_Inst_Sbox_4_M14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_M15_U1 ( .A(SubBytesIns_Inst_Sbox_4_M14), 
        .B(SubBytesIns_Inst_Sbox_4_M11), .Z(SubBytesIns_Inst_Sbox_4_M15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_M16_U1 ( .A(SubBytesIns_Inst_Sbox_4_M3), 
        .B(SubBytesIns_Inst_Sbox_4_M2), .Z(SubBytesIns_Inst_Sbox_4_M16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_M17_U1 ( .A(SubBytesIns_Inst_Sbox_4_M5), 
        .B(SubBytesIns_Inst_Sbox_4_T24), .Z(SubBytesIns_Inst_Sbox_4_M17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_M18_U1 ( .A(SubBytesIns_Inst_Sbox_4_M8), 
        .B(SubBytesIns_Inst_Sbox_4_M7), .Z(SubBytesIns_Inst_Sbox_4_M18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_M19_U1 ( .A(SubBytesIns_Inst_Sbox_4_M10), 
        .B(SubBytesIns_Inst_Sbox_4_M15), .Z(SubBytesIns_Inst_Sbox_4_M19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_M20_U1 ( .A(SubBytesIns_Inst_Sbox_4_M16), 
        .B(SubBytesIns_Inst_Sbox_4_M13), .Z(SubBytesIns_Inst_Sbox_4_M20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_M21_U1 ( .A(SubBytesIns_Inst_Sbox_4_M17), 
        .B(SubBytesIns_Inst_Sbox_4_M15), .Z(SubBytesIns_Inst_Sbox_4_M21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_M22_U1 ( .A(SubBytesIns_Inst_Sbox_4_M18), 
        .B(SubBytesIns_Inst_Sbox_4_M13), .Z(SubBytesIns_Inst_Sbox_4_M22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_M23_U1 ( .A(SubBytesIns_Inst_Sbox_4_M19), 
        .B(SubBytesIns_Inst_Sbox_4_T25), .Z(SubBytesIns_Inst_Sbox_4_M23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_M24_U1 ( .A(SubBytesIns_Inst_Sbox_4_M22), 
        .B(SubBytesIns_Inst_Sbox_4_M23), .Z(SubBytesIns_Inst_Sbox_4_M24) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M25_U1 ( .A1(SubBytesIns_Inst_Sbox_4_M22), .A2(SubBytesIns_Inst_Sbox_4_M20), .ZN(SubBytesIns_Inst_Sbox_4_M25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_M26_U1 ( .A(SubBytesIns_Inst_Sbox_4_M21), 
        .B(SubBytesIns_Inst_Sbox_4_M25), .Z(SubBytesIns_Inst_Sbox_4_M26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_M27_U1 ( .A(SubBytesIns_Inst_Sbox_4_M20), 
        .B(SubBytesIns_Inst_Sbox_4_M21), .Z(SubBytesIns_Inst_Sbox_4_M27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_M28_U1 ( .A(SubBytesIns_Inst_Sbox_4_M23), 
        .B(SubBytesIns_Inst_Sbox_4_M25), .Z(SubBytesIns_Inst_Sbox_4_M28) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M29_U1 ( .A1(SubBytesIns_Inst_Sbox_4_M28), .A2(SubBytesIns_Inst_Sbox_4_M27), .ZN(SubBytesIns_Inst_Sbox_4_M29) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M30_U1 ( .A1(SubBytesIns_Inst_Sbox_4_M26), .A2(SubBytesIns_Inst_Sbox_4_M24), .ZN(SubBytesIns_Inst_Sbox_4_M30) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M31_U1 ( .A1(SubBytesIns_Inst_Sbox_4_M20), .A2(SubBytesIns_Inst_Sbox_4_M23), .ZN(SubBytesIns_Inst_Sbox_4_M31) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M32_U1 ( .A1(SubBytesIns_Inst_Sbox_4_M27), .A2(SubBytesIns_Inst_Sbox_4_M31), .ZN(SubBytesIns_Inst_Sbox_4_M32) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_M33_U1 ( .A(SubBytesIns_Inst_Sbox_4_M27), 
        .B(SubBytesIns_Inst_Sbox_4_M25), .Z(SubBytesIns_Inst_Sbox_4_M33) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M34_U1 ( .A1(SubBytesIns_Inst_Sbox_4_M21), .A2(SubBytesIns_Inst_Sbox_4_M22), .ZN(SubBytesIns_Inst_Sbox_4_M34) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M35_U1 ( .A1(SubBytesIns_Inst_Sbox_4_M24), .A2(SubBytesIns_Inst_Sbox_4_M34), .ZN(SubBytesIns_Inst_Sbox_4_M35) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_M36_U1 ( .A(SubBytesIns_Inst_Sbox_4_M24), 
        .B(SubBytesIns_Inst_Sbox_4_M25), .Z(SubBytesIns_Inst_Sbox_4_M36) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_M37_U1 ( .A(SubBytesIns_Inst_Sbox_4_M21), 
        .B(SubBytesIns_Inst_Sbox_4_M29), .Z(SubBytesIns_Inst_Sbox_4_M37) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_M38_U1 ( .A(SubBytesIns_Inst_Sbox_4_M32), 
        .B(SubBytesIns_Inst_Sbox_4_M33), .Z(SubBytesIns_Inst_Sbox_4_M38) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_M39_U1 ( .A(SubBytesIns_Inst_Sbox_4_M23), 
        .B(SubBytesIns_Inst_Sbox_4_M30), .Z(SubBytesIns_Inst_Sbox_4_M39) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_M40_U1 ( .A(SubBytesIns_Inst_Sbox_4_M35), 
        .B(SubBytesIns_Inst_Sbox_4_M36), .Z(SubBytesIns_Inst_Sbox_4_M40) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_M41_U1 ( .A(SubBytesIns_Inst_Sbox_4_M38), 
        .B(SubBytesIns_Inst_Sbox_4_M40), .Z(SubBytesIns_Inst_Sbox_4_M41) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_M42_U1 ( .A(SubBytesIns_Inst_Sbox_4_M37), 
        .B(SubBytesIns_Inst_Sbox_4_M39), .Z(SubBytesIns_Inst_Sbox_4_M42) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_M43_U1 ( .A(SubBytesIns_Inst_Sbox_4_M37), 
        .B(SubBytesIns_Inst_Sbox_4_M38), .Z(SubBytesIns_Inst_Sbox_4_M43) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_M44_U1 ( .A(SubBytesIns_Inst_Sbox_4_M39), 
        .B(SubBytesIns_Inst_Sbox_4_M40), .Z(SubBytesIns_Inst_Sbox_4_M44) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_M45_U1 ( .A(SubBytesIns_Inst_Sbox_4_M42), 
        .B(SubBytesIns_Inst_Sbox_4_M41), .Z(SubBytesIns_Inst_Sbox_4_M45) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M46_U1 ( .A1(SubBytesIns_Inst_Sbox_4_M44), .A2(SubBytesIns_Inst_Sbox_4_T6), .ZN(SubBytesIns_Inst_Sbox_4_M46) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M47_U1 ( .A1(SubBytesIns_Inst_Sbox_4_M40), .A2(SubBytesIns_Inst_Sbox_4_T8), .ZN(SubBytesIns_Inst_Sbox_4_M47) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M48_U1 ( .A1(SubBytesIns_Inst_Sbox_4_M39), .A2(SubBytesInput[32]), .ZN(SubBytesIns_Inst_Sbox_4_M48) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M49_U1 ( .A1(SubBytesIns_Inst_Sbox_4_M43), .A2(SubBytesIns_Inst_Sbox_4_T16), .ZN(SubBytesIns_Inst_Sbox_4_M49) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M50_U1 ( .A1(SubBytesIns_Inst_Sbox_4_M38), .A2(SubBytesIns_Inst_Sbox_4_T9), .ZN(SubBytesIns_Inst_Sbox_4_M50) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M51_U1 ( .A1(SubBytesIns_Inst_Sbox_4_M37), .A2(SubBytesIns_Inst_Sbox_4_T17), .ZN(SubBytesIns_Inst_Sbox_4_M51) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M52_U1 ( .A1(SubBytesIns_Inst_Sbox_4_M42), .A2(SubBytesIns_Inst_Sbox_4_T15), .ZN(SubBytesIns_Inst_Sbox_4_M52) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M53_U1 ( .A1(SubBytesIns_Inst_Sbox_4_M45), .A2(SubBytesIns_Inst_Sbox_4_T27), .ZN(SubBytesIns_Inst_Sbox_4_M53) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M54_U1 ( .A1(SubBytesIns_Inst_Sbox_4_M41), .A2(SubBytesIns_Inst_Sbox_4_T10), .ZN(SubBytesIns_Inst_Sbox_4_M54) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M55_U1 ( .A1(SubBytesIns_Inst_Sbox_4_M44), .A2(SubBytesIns_Inst_Sbox_4_T13), .ZN(SubBytesIns_Inst_Sbox_4_M55) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M56_U1 ( .A1(SubBytesIns_Inst_Sbox_4_M40), .A2(SubBytesIns_Inst_Sbox_4_T23), .ZN(SubBytesIns_Inst_Sbox_4_M56) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M57_U1 ( .A1(SubBytesIns_Inst_Sbox_4_M39), .A2(SubBytesIns_Inst_Sbox_4_T19), .ZN(SubBytesIns_Inst_Sbox_4_M57) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M58_U1 ( .A1(SubBytesIns_Inst_Sbox_4_M43), .A2(SubBytesIns_Inst_Sbox_4_T3), .ZN(SubBytesIns_Inst_Sbox_4_M58) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M59_U1 ( .A1(SubBytesIns_Inst_Sbox_4_M38), .A2(SubBytesIns_Inst_Sbox_4_T22), .ZN(SubBytesIns_Inst_Sbox_4_M59) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M60_U1 ( .A1(SubBytesIns_Inst_Sbox_4_M37), .A2(SubBytesIns_Inst_Sbox_4_T20), .ZN(SubBytesIns_Inst_Sbox_4_M60) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M61_U1 ( .A1(SubBytesIns_Inst_Sbox_4_M42), .A2(SubBytesIns_Inst_Sbox_4_T1), .ZN(SubBytesIns_Inst_Sbox_4_M61) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M62_U1 ( .A1(SubBytesIns_Inst_Sbox_4_M45), .A2(SubBytesIns_Inst_Sbox_4_T4), .ZN(SubBytesIns_Inst_Sbox_4_M62) );
  AND2_X1 SubBytesIns_Inst_Sbox_4_AND_M63_U1 ( .A1(SubBytesIns_Inst_Sbox_4_M41), .A2(SubBytesIns_Inst_Sbox_4_T2), .ZN(SubBytesIns_Inst_Sbox_4_M63) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_L0_U1 ( .A(SubBytesIns_Inst_Sbox_4_M61), 
        .B(SubBytesIns_Inst_Sbox_4_M62), .Z(SubBytesIns_Inst_Sbox_4_L0) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_L1_U1 ( .A(SubBytesIns_Inst_Sbox_4_M50), 
        .B(SubBytesIns_Inst_Sbox_4_M56), .Z(SubBytesIns_Inst_Sbox_4_L1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_L2_U1 ( .A(SubBytesIns_Inst_Sbox_4_M46), 
        .B(SubBytesIns_Inst_Sbox_4_M48), .Z(SubBytesIns_Inst_Sbox_4_L2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_L3_U1 ( .A(SubBytesIns_Inst_Sbox_4_M47), 
        .B(SubBytesIns_Inst_Sbox_4_M55), .Z(SubBytesIns_Inst_Sbox_4_L3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_L4_U1 ( .A(SubBytesIns_Inst_Sbox_4_M54), 
        .B(SubBytesIns_Inst_Sbox_4_M58), .Z(SubBytesIns_Inst_Sbox_4_L4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_L5_U1 ( .A(SubBytesIns_Inst_Sbox_4_M49), 
        .B(SubBytesIns_Inst_Sbox_4_M61), .Z(SubBytesIns_Inst_Sbox_4_L5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_L6_U1 ( .A(SubBytesIns_Inst_Sbox_4_M62), 
        .B(SubBytesIns_Inst_Sbox_4_L5), .Z(SubBytesIns_Inst_Sbox_4_L6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_L7_U1 ( .A(SubBytesIns_Inst_Sbox_4_M46), 
        .B(SubBytesIns_Inst_Sbox_4_L3), .Z(SubBytesIns_Inst_Sbox_4_L7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_L8_U1 ( .A(SubBytesIns_Inst_Sbox_4_M51), 
        .B(SubBytesIns_Inst_Sbox_4_M59), .Z(SubBytesIns_Inst_Sbox_4_L8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_L9_U1 ( .A(SubBytesIns_Inst_Sbox_4_M52), 
        .B(SubBytesIns_Inst_Sbox_4_M53), .Z(SubBytesIns_Inst_Sbox_4_L9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_L10_U1 ( .A(SubBytesIns_Inst_Sbox_4_M53), 
        .B(SubBytesIns_Inst_Sbox_4_L4), .Z(SubBytesIns_Inst_Sbox_4_L10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_L11_U1 ( .A(SubBytesIns_Inst_Sbox_4_M60), 
        .B(SubBytesIns_Inst_Sbox_4_L2), .Z(SubBytesIns_Inst_Sbox_4_L11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_L12_U1 ( .A(SubBytesIns_Inst_Sbox_4_M48), 
        .B(SubBytesIns_Inst_Sbox_4_M51), .Z(SubBytesIns_Inst_Sbox_4_L12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_L13_U1 ( .A(SubBytesIns_Inst_Sbox_4_M50), 
        .B(SubBytesIns_Inst_Sbox_4_L0), .Z(SubBytesIns_Inst_Sbox_4_L13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_L14_U1 ( .A(SubBytesIns_Inst_Sbox_4_M52), 
        .B(SubBytesIns_Inst_Sbox_4_M61), .Z(SubBytesIns_Inst_Sbox_4_L14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_L15_U1 ( .A(SubBytesIns_Inst_Sbox_4_M55), 
        .B(SubBytesIns_Inst_Sbox_4_L1), .Z(SubBytesIns_Inst_Sbox_4_L15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_L16_U1 ( .A(SubBytesIns_Inst_Sbox_4_M56), 
        .B(SubBytesIns_Inst_Sbox_4_L0), .Z(SubBytesIns_Inst_Sbox_4_L16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_L17_U1 ( .A(SubBytesIns_Inst_Sbox_4_M57), 
        .B(SubBytesIns_Inst_Sbox_4_L1), .Z(SubBytesIns_Inst_Sbox_4_L17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_L18_U1 ( .A(SubBytesIns_Inst_Sbox_4_M58), 
        .B(SubBytesIns_Inst_Sbox_4_L8), .Z(SubBytesIns_Inst_Sbox_4_L18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_L19_U1 ( .A(SubBytesIns_Inst_Sbox_4_M63), 
        .B(SubBytesIns_Inst_Sbox_4_L4), .Z(SubBytesIns_Inst_Sbox_4_L19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_L20_U1 ( .A(SubBytesIns_Inst_Sbox_4_L0), 
        .B(SubBytesIns_Inst_Sbox_4_L1), .Z(SubBytesIns_Inst_Sbox_4_L20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_L21_U1 ( .A(SubBytesIns_Inst_Sbox_4_L1), 
        .B(SubBytesIns_Inst_Sbox_4_L7), .Z(SubBytesIns_Inst_Sbox_4_L21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_L22_U1 ( .A(SubBytesIns_Inst_Sbox_4_L3), 
        .B(SubBytesIns_Inst_Sbox_4_L12), .Z(SubBytesIns_Inst_Sbox_4_L22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_L23_U1 ( .A(SubBytesIns_Inst_Sbox_4_L18), 
        .B(SubBytesIns_Inst_Sbox_4_L2), .Z(SubBytesIns_Inst_Sbox_4_L23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_L24_U1 ( .A(SubBytesIns_Inst_Sbox_4_L15), 
        .B(SubBytesIns_Inst_Sbox_4_L9), .Z(SubBytesIns_Inst_Sbox_4_L24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_L25_U1 ( .A(SubBytesIns_Inst_Sbox_4_L6), 
        .B(SubBytesIns_Inst_Sbox_4_L10), .Z(SubBytesIns_Inst_Sbox_4_L25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_L26_U1 ( .A(SubBytesIns_Inst_Sbox_4_L7), 
        .B(SubBytesIns_Inst_Sbox_4_L9), .Z(SubBytesIns_Inst_Sbox_4_L26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_L27_U1 ( .A(SubBytesIns_Inst_Sbox_4_L8), 
        .B(SubBytesIns_Inst_Sbox_4_L10), .Z(SubBytesIns_Inst_Sbox_4_L27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_L28_U1 ( .A(SubBytesIns_Inst_Sbox_4_L11), 
        .B(SubBytesIns_Inst_Sbox_4_L14), .Z(SubBytesIns_Inst_Sbox_4_L28) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_L29_U1 ( .A(SubBytesIns_Inst_Sbox_4_L11), 
        .B(SubBytesIns_Inst_Sbox_4_L17), .Z(SubBytesIns_Inst_Sbox_4_L29) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_S0_U1 ( .A(SubBytesIns_Inst_Sbox_4_L6), 
        .B(SubBytesIns_Inst_Sbox_4_L24), .Z(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_S1_U1 ( .A(SubBytesIns_Inst_Sbox_4_L16), 
        .B(SubBytesIns_Inst_Sbox_4_L26), .ZN(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[7]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_S2_U1 ( .A(SubBytesIns_Inst_Sbox_4_L19), 
        .B(SubBytesIns_Inst_Sbox_4_L28), .ZN(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[6]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_S3_U1 ( .A(SubBytesIns_Inst_Sbox_4_L6), 
        .B(SubBytesIns_Inst_Sbox_4_L21), .Z(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[5]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_S4_U1 ( .A(SubBytesIns_Inst_Sbox_4_L20), 
        .B(SubBytesIns_Inst_Sbox_4_L22), .Z(MixColumnsInput[3]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_S5_U1 ( .A(SubBytesIns_Inst_Sbox_4_L25), 
        .B(SubBytesIns_Inst_Sbox_4_L29), .Z(MixColumnsInput[2]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_S6_U1 ( .A(SubBytesIns_Inst_Sbox_4_L13), 
        .B(SubBytesIns_Inst_Sbox_4_L27), .ZN(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[2]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_4_XOR_S7_U1 ( .A(SubBytesIns_Inst_Sbox_4_L6), 
        .B(SubBytesIns_Inst_Sbox_4_L23), .ZN(MixColumnsInput[0]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_T1_U1 ( .A(SubBytesInput[47]), .B(
        SubBytesInput[44]), .Z(SubBytesIns_Inst_Sbox_5_T1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_T2_U1 ( .A(SubBytesInput[47]), .B(
        SubBytesInput[42]), .Z(SubBytesIns_Inst_Sbox_5_T2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_T3_U1 ( .A(SubBytesInput[47]), .B(
        SubBytesInput[41]), .Z(SubBytesIns_Inst_Sbox_5_T3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_T4_U1 ( .A(SubBytesInput[44]), .B(
        SubBytesInput[42]), .Z(SubBytesIns_Inst_Sbox_5_T4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_T5_U1 ( .A(SubBytesInput[43]), .B(
        SubBytesInput[41]), .Z(SubBytesIns_Inst_Sbox_5_T5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_T6_U1 ( .A(SubBytesIns_Inst_Sbox_5_T1), 
        .B(SubBytesIns_Inst_Sbox_5_T5), .Z(SubBytesIns_Inst_Sbox_5_T6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_T7_U1 ( .A(SubBytesInput[46]), .B(
        SubBytesInput[45]), .Z(SubBytesIns_Inst_Sbox_5_T7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_T8_U1 ( .A(SubBytesInput[40]), .B(
        SubBytesIns_Inst_Sbox_5_T6), .Z(SubBytesIns_Inst_Sbox_5_T8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_T9_U1 ( .A(SubBytesInput[40]), .B(
        SubBytesIns_Inst_Sbox_5_T7), .Z(SubBytesIns_Inst_Sbox_5_T9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_T10_U1 ( .A(SubBytesIns_Inst_Sbox_5_T6), 
        .B(SubBytesIns_Inst_Sbox_5_T7), .Z(SubBytesIns_Inst_Sbox_5_T10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_T11_U1 ( .A(SubBytesInput[46]), .B(
        SubBytesInput[42]), .Z(SubBytesIns_Inst_Sbox_5_T11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_T12_U1 ( .A(SubBytesInput[45]), .B(
        SubBytesInput[42]), .Z(SubBytesIns_Inst_Sbox_5_T12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_T13_U1 ( .A(SubBytesIns_Inst_Sbox_5_T3), 
        .B(SubBytesIns_Inst_Sbox_5_T4), .Z(SubBytesIns_Inst_Sbox_5_T13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_T14_U1 ( .A(SubBytesIns_Inst_Sbox_5_T6), 
        .B(SubBytesIns_Inst_Sbox_5_T11), .Z(SubBytesIns_Inst_Sbox_5_T14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_T15_U1 ( .A(SubBytesIns_Inst_Sbox_5_T5), 
        .B(SubBytesIns_Inst_Sbox_5_T11), .Z(SubBytesIns_Inst_Sbox_5_T15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_T16_U1 ( .A(SubBytesIns_Inst_Sbox_5_T5), 
        .B(SubBytesIns_Inst_Sbox_5_T12), .Z(SubBytesIns_Inst_Sbox_5_T16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_T17_U1 ( .A(SubBytesIns_Inst_Sbox_5_T9), 
        .B(SubBytesIns_Inst_Sbox_5_T16), .Z(SubBytesIns_Inst_Sbox_5_T17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_T18_U1 ( .A(SubBytesInput[44]), .B(
        SubBytesInput[40]), .Z(SubBytesIns_Inst_Sbox_5_T18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_T19_U1 ( .A(SubBytesIns_Inst_Sbox_5_T7), 
        .B(SubBytesIns_Inst_Sbox_5_T18), .Z(SubBytesIns_Inst_Sbox_5_T19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_T20_U1 ( .A(SubBytesIns_Inst_Sbox_5_T1), 
        .B(SubBytesIns_Inst_Sbox_5_T19), .Z(SubBytesIns_Inst_Sbox_5_T20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_T21_U1 ( .A(SubBytesInput[41]), .B(
        SubBytesInput[40]), .Z(SubBytesIns_Inst_Sbox_5_T21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_T22_U1 ( .A(SubBytesIns_Inst_Sbox_5_T7), 
        .B(SubBytesIns_Inst_Sbox_5_T21), .Z(SubBytesIns_Inst_Sbox_5_T22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_T23_U1 ( .A(SubBytesIns_Inst_Sbox_5_T2), 
        .B(SubBytesIns_Inst_Sbox_5_T22), .Z(SubBytesIns_Inst_Sbox_5_T23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_T24_U1 ( .A(SubBytesIns_Inst_Sbox_5_T2), 
        .B(SubBytesIns_Inst_Sbox_5_T10), .Z(SubBytesIns_Inst_Sbox_5_T24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_T25_U1 ( .A(SubBytesIns_Inst_Sbox_5_T20), 
        .B(SubBytesIns_Inst_Sbox_5_T17), .Z(SubBytesIns_Inst_Sbox_5_T25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_T26_U1 ( .A(SubBytesIns_Inst_Sbox_5_T3), 
        .B(SubBytesIns_Inst_Sbox_5_T16), .Z(SubBytesIns_Inst_Sbox_5_T26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_T27_U1 ( .A(SubBytesIns_Inst_Sbox_5_T1), 
        .B(SubBytesIns_Inst_Sbox_5_T12), .Z(SubBytesIns_Inst_Sbox_5_T27) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M1_U1 ( .A1(SubBytesIns_Inst_Sbox_5_T13), 
        .A2(SubBytesIns_Inst_Sbox_5_T6), .ZN(SubBytesIns_Inst_Sbox_5_M1) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M2_U1 ( .A1(SubBytesIns_Inst_Sbox_5_T23), 
        .A2(SubBytesIns_Inst_Sbox_5_T8), .ZN(SubBytesIns_Inst_Sbox_5_M2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_M3_U1 ( .A(SubBytesIns_Inst_Sbox_5_T14), 
        .B(SubBytesIns_Inst_Sbox_5_M1), .Z(SubBytesIns_Inst_Sbox_5_M3) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M4_U1 ( .A1(SubBytesIns_Inst_Sbox_5_T19), 
        .A2(SubBytesInput[40]), .ZN(SubBytesIns_Inst_Sbox_5_M4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_M5_U1 ( .A(SubBytesIns_Inst_Sbox_5_M4), 
        .B(SubBytesIns_Inst_Sbox_5_M1), .Z(SubBytesIns_Inst_Sbox_5_M5) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M6_U1 ( .A1(SubBytesIns_Inst_Sbox_5_T3), 
        .A2(SubBytesIns_Inst_Sbox_5_T16), .ZN(SubBytesIns_Inst_Sbox_5_M6) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M7_U1 ( .A1(SubBytesIns_Inst_Sbox_5_T22), 
        .A2(SubBytesIns_Inst_Sbox_5_T9), .ZN(SubBytesIns_Inst_Sbox_5_M7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_M8_U1 ( .A(SubBytesIns_Inst_Sbox_5_T26), 
        .B(SubBytesIns_Inst_Sbox_5_M6), .Z(SubBytesIns_Inst_Sbox_5_M8) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M9_U1 ( .A1(SubBytesIns_Inst_Sbox_5_T20), 
        .A2(SubBytesIns_Inst_Sbox_5_T17), .ZN(SubBytesIns_Inst_Sbox_5_M9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_M10_U1 ( .A(SubBytesIns_Inst_Sbox_5_M9), 
        .B(SubBytesIns_Inst_Sbox_5_M6), .Z(SubBytesIns_Inst_Sbox_5_M10) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M11_U1 ( .A1(SubBytesIns_Inst_Sbox_5_T1), 
        .A2(SubBytesIns_Inst_Sbox_5_T15), .ZN(SubBytesIns_Inst_Sbox_5_M11) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M12_U1 ( .A1(SubBytesIns_Inst_Sbox_5_T4), 
        .A2(SubBytesIns_Inst_Sbox_5_T27), .ZN(SubBytesIns_Inst_Sbox_5_M12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_M13_U1 ( .A(SubBytesIns_Inst_Sbox_5_M12), 
        .B(SubBytesIns_Inst_Sbox_5_M11), .Z(SubBytesIns_Inst_Sbox_5_M13) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M14_U1 ( .A1(SubBytesIns_Inst_Sbox_5_T2), 
        .A2(SubBytesIns_Inst_Sbox_5_T10), .ZN(SubBytesIns_Inst_Sbox_5_M14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_M15_U1 ( .A(SubBytesIns_Inst_Sbox_5_M14), 
        .B(SubBytesIns_Inst_Sbox_5_M11), .Z(SubBytesIns_Inst_Sbox_5_M15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_M16_U1 ( .A(SubBytesIns_Inst_Sbox_5_M3), 
        .B(SubBytesIns_Inst_Sbox_5_M2), .Z(SubBytesIns_Inst_Sbox_5_M16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_M17_U1 ( .A(SubBytesIns_Inst_Sbox_5_M5), 
        .B(SubBytesIns_Inst_Sbox_5_T24), .Z(SubBytesIns_Inst_Sbox_5_M17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_M18_U1 ( .A(SubBytesIns_Inst_Sbox_5_M8), 
        .B(SubBytesIns_Inst_Sbox_5_M7), .Z(SubBytesIns_Inst_Sbox_5_M18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_M19_U1 ( .A(SubBytesIns_Inst_Sbox_5_M10), 
        .B(SubBytesIns_Inst_Sbox_5_M15), .Z(SubBytesIns_Inst_Sbox_5_M19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_M20_U1 ( .A(SubBytesIns_Inst_Sbox_5_M16), 
        .B(SubBytesIns_Inst_Sbox_5_M13), .Z(SubBytesIns_Inst_Sbox_5_M20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_M21_U1 ( .A(SubBytesIns_Inst_Sbox_5_M17), 
        .B(SubBytesIns_Inst_Sbox_5_M15), .Z(SubBytesIns_Inst_Sbox_5_M21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_M22_U1 ( .A(SubBytesIns_Inst_Sbox_5_M18), 
        .B(SubBytesIns_Inst_Sbox_5_M13), .Z(SubBytesIns_Inst_Sbox_5_M22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_M23_U1 ( .A(SubBytesIns_Inst_Sbox_5_M19), 
        .B(SubBytesIns_Inst_Sbox_5_T25), .Z(SubBytesIns_Inst_Sbox_5_M23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_M24_U1 ( .A(SubBytesIns_Inst_Sbox_5_M22), 
        .B(SubBytesIns_Inst_Sbox_5_M23), .Z(SubBytesIns_Inst_Sbox_5_M24) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M25_U1 ( .A1(SubBytesIns_Inst_Sbox_5_M22), .A2(SubBytesIns_Inst_Sbox_5_M20), .ZN(SubBytesIns_Inst_Sbox_5_M25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_M26_U1 ( .A(SubBytesIns_Inst_Sbox_5_M21), 
        .B(SubBytesIns_Inst_Sbox_5_M25), .Z(SubBytesIns_Inst_Sbox_5_M26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_M27_U1 ( .A(SubBytesIns_Inst_Sbox_5_M20), 
        .B(SubBytesIns_Inst_Sbox_5_M21), .Z(SubBytesIns_Inst_Sbox_5_M27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_M28_U1 ( .A(SubBytesIns_Inst_Sbox_5_M23), 
        .B(SubBytesIns_Inst_Sbox_5_M25), .Z(SubBytesIns_Inst_Sbox_5_M28) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M29_U1 ( .A1(SubBytesIns_Inst_Sbox_5_M28), .A2(SubBytesIns_Inst_Sbox_5_M27), .ZN(SubBytesIns_Inst_Sbox_5_M29) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M30_U1 ( .A1(SubBytesIns_Inst_Sbox_5_M26), .A2(SubBytesIns_Inst_Sbox_5_M24), .ZN(SubBytesIns_Inst_Sbox_5_M30) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M31_U1 ( .A1(SubBytesIns_Inst_Sbox_5_M20), .A2(SubBytesIns_Inst_Sbox_5_M23), .ZN(SubBytesIns_Inst_Sbox_5_M31) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M32_U1 ( .A1(SubBytesIns_Inst_Sbox_5_M27), .A2(SubBytesIns_Inst_Sbox_5_M31), .ZN(SubBytesIns_Inst_Sbox_5_M32) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_M33_U1 ( .A(SubBytesIns_Inst_Sbox_5_M27), 
        .B(SubBytesIns_Inst_Sbox_5_M25), .Z(SubBytesIns_Inst_Sbox_5_M33) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M34_U1 ( .A1(SubBytesIns_Inst_Sbox_5_M21), .A2(SubBytesIns_Inst_Sbox_5_M22), .ZN(SubBytesIns_Inst_Sbox_5_M34) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M35_U1 ( .A1(SubBytesIns_Inst_Sbox_5_M24), .A2(SubBytesIns_Inst_Sbox_5_M34), .ZN(SubBytesIns_Inst_Sbox_5_M35) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_M36_U1 ( .A(SubBytesIns_Inst_Sbox_5_M24), 
        .B(SubBytesIns_Inst_Sbox_5_M25), .Z(SubBytesIns_Inst_Sbox_5_M36) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_M37_U1 ( .A(SubBytesIns_Inst_Sbox_5_M21), 
        .B(SubBytesIns_Inst_Sbox_5_M29), .Z(SubBytesIns_Inst_Sbox_5_M37) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_M38_U1 ( .A(SubBytesIns_Inst_Sbox_5_M32), 
        .B(SubBytesIns_Inst_Sbox_5_M33), .Z(SubBytesIns_Inst_Sbox_5_M38) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_M39_U1 ( .A(SubBytesIns_Inst_Sbox_5_M23), 
        .B(SubBytesIns_Inst_Sbox_5_M30), .Z(SubBytesIns_Inst_Sbox_5_M39) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_M40_U1 ( .A(SubBytesIns_Inst_Sbox_5_M35), 
        .B(SubBytesIns_Inst_Sbox_5_M36), .Z(SubBytesIns_Inst_Sbox_5_M40) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_M41_U1 ( .A(SubBytesIns_Inst_Sbox_5_M38), 
        .B(SubBytesIns_Inst_Sbox_5_M40), .Z(SubBytesIns_Inst_Sbox_5_M41) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_M42_U1 ( .A(SubBytesIns_Inst_Sbox_5_M37), 
        .B(SubBytesIns_Inst_Sbox_5_M39), .Z(SubBytesIns_Inst_Sbox_5_M42) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_M43_U1 ( .A(SubBytesIns_Inst_Sbox_5_M37), 
        .B(SubBytesIns_Inst_Sbox_5_M38), .Z(SubBytesIns_Inst_Sbox_5_M43) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_M44_U1 ( .A(SubBytesIns_Inst_Sbox_5_M39), 
        .B(SubBytesIns_Inst_Sbox_5_M40), .Z(SubBytesIns_Inst_Sbox_5_M44) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_M45_U1 ( .A(SubBytesIns_Inst_Sbox_5_M42), 
        .B(SubBytesIns_Inst_Sbox_5_M41), .Z(SubBytesIns_Inst_Sbox_5_M45) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M46_U1 ( .A1(SubBytesIns_Inst_Sbox_5_M44), .A2(SubBytesIns_Inst_Sbox_5_T6), .ZN(SubBytesIns_Inst_Sbox_5_M46) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M47_U1 ( .A1(SubBytesIns_Inst_Sbox_5_M40), .A2(SubBytesIns_Inst_Sbox_5_T8), .ZN(SubBytesIns_Inst_Sbox_5_M47) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M48_U1 ( .A1(SubBytesIns_Inst_Sbox_5_M39), .A2(SubBytesInput[40]), .ZN(SubBytesIns_Inst_Sbox_5_M48) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M49_U1 ( .A1(SubBytesIns_Inst_Sbox_5_M43), .A2(SubBytesIns_Inst_Sbox_5_T16), .ZN(SubBytesIns_Inst_Sbox_5_M49) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M50_U1 ( .A1(SubBytesIns_Inst_Sbox_5_M38), .A2(SubBytesIns_Inst_Sbox_5_T9), .ZN(SubBytesIns_Inst_Sbox_5_M50) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M51_U1 ( .A1(SubBytesIns_Inst_Sbox_5_M37), .A2(SubBytesIns_Inst_Sbox_5_T17), .ZN(SubBytesIns_Inst_Sbox_5_M51) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M52_U1 ( .A1(SubBytesIns_Inst_Sbox_5_M42), .A2(SubBytesIns_Inst_Sbox_5_T15), .ZN(SubBytesIns_Inst_Sbox_5_M52) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M53_U1 ( .A1(SubBytesIns_Inst_Sbox_5_M45), .A2(SubBytesIns_Inst_Sbox_5_T27), .ZN(SubBytesIns_Inst_Sbox_5_M53) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M54_U1 ( .A1(SubBytesIns_Inst_Sbox_5_M41), .A2(SubBytesIns_Inst_Sbox_5_T10), .ZN(SubBytesIns_Inst_Sbox_5_M54) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M55_U1 ( .A1(SubBytesIns_Inst_Sbox_5_M44), .A2(SubBytesIns_Inst_Sbox_5_T13), .ZN(SubBytesIns_Inst_Sbox_5_M55) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M56_U1 ( .A1(SubBytesIns_Inst_Sbox_5_M40), .A2(SubBytesIns_Inst_Sbox_5_T23), .ZN(SubBytesIns_Inst_Sbox_5_M56) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M57_U1 ( .A1(SubBytesIns_Inst_Sbox_5_M39), .A2(SubBytesIns_Inst_Sbox_5_T19), .ZN(SubBytesIns_Inst_Sbox_5_M57) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M58_U1 ( .A1(SubBytesIns_Inst_Sbox_5_M43), .A2(SubBytesIns_Inst_Sbox_5_T3), .ZN(SubBytesIns_Inst_Sbox_5_M58) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M59_U1 ( .A1(SubBytesIns_Inst_Sbox_5_M38), .A2(SubBytesIns_Inst_Sbox_5_T22), .ZN(SubBytesIns_Inst_Sbox_5_M59) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M60_U1 ( .A1(SubBytesIns_Inst_Sbox_5_M37), .A2(SubBytesIns_Inst_Sbox_5_T20), .ZN(SubBytesIns_Inst_Sbox_5_M60) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M61_U1 ( .A1(SubBytesIns_Inst_Sbox_5_M42), .A2(SubBytesIns_Inst_Sbox_5_T1), .ZN(SubBytesIns_Inst_Sbox_5_M61) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M62_U1 ( .A1(SubBytesIns_Inst_Sbox_5_M45), .A2(SubBytesIns_Inst_Sbox_5_T4), .ZN(SubBytesIns_Inst_Sbox_5_M62) );
  AND2_X1 SubBytesIns_Inst_Sbox_5_AND_M63_U1 ( .A1(SubBytesIns_Inst_Sbox_5_M41), .A2(SubBytesIns_Inst_Sbox_5_T2), .ZN(SubBytesIns_Inst_Sbox_5_M63) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_L0_U1 ( .A(SubBytesIns_Inst_Sbox_5_M61), 
        .B(SubBytesIns_Inst_Sbox_5_M62), .Z(SubBytesIns_Inst_Sbox_5_L0) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_L1_U1 ( .A(SubBytesIns_Inst_Sbox_5_M50), 
        .B(SubBytesIns_Inst_Sbox_5_M56), .Z(SubBytesIns_Inst_Sbox_5_L1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_L2_U1 ( .A(SubBytesIns_Inst_Sbox_5_M46), 
        .B(SubBytesIns_Inst_Sbox_5_M48), .Z(SubBytesIns_Inst_Sbox_5_L2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_L3_U1 ( .A(SubBytesIns_Inst_Sbox_5_M47), 
        .B(SubBytesIns_Inst_Sbox_5_M55), .Z(SubBytesIns_Inst_Sbox_5_L3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_L4_U1 ( .A(SubBytesIns_Inst_Sbox_5_M54), 
        .B(SubBytesIns_Inst_Sbox_5_M58), .Z(SubBytesIns_Inst_Sbox_5_L4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_L5_U1 ( .A(SubBytesIns_Inst_Sbox_5_M49), 
        .B(SubBytesIns_Inst_Sbox_5_M61), .Z(SubBytesIns_Inst_Sbox_5_L5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_L6_U1 ( .A(SubBytesIns_Inst_Sbox_5_M62), 
        .B(SubBytesIns_Inst_Sbox_5_L5), .Z(SubBytesIns_Inst_Sbox_5_L6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_L7_U1 ( .A(SubBytesIns_Inst_Sbox_5_M46), 
        .B(SubBytesIns_Inst_Sbox_5_L3), .Z(SubBytesIns_Inst_Sbox_5_L7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_L8_U1 ( .A(SubBytesIns_Inst_Sbox_5_M51), 
        .B(SubBytesIns_Inst_Sbox_5_M59), .Z(SubBytesIns_Inst_Sbox_5_L8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_L9_U1 ( .A(SubBytesIns_Inst_Sbox_5_M52), 
        .B(SubBytesIns_Inst_Sbox_5_M53), .Z(SubBytesIns_Inst_Sbox_5_L9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_L10_U1 ( .A(SubBytesIns_Inst_Sbox_5_M53), 
        .B(SubBytesIns_Inst_Sbox_5_L4), .Z(SubBytesIns_Inst_Sbox_5_L10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_L11_U1 ( .A(SubBytesIns_Inst_Sbox_5_M60), 
        .B(SubBytesIns_Inst_Sbox_5_L2), .Z(SubBytesIns_Inst_Sbox_5_L11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_L12_U1 ( .A(SubBytesIns_Inst_Sbox_5_M48), 
        .B(SubBytesIns_Inst_Sbox_5_M51), .Z(SubBytesIns_Inst_Sbox_5_L12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_L13_U1 ( .A(SubBytesIns_Inst_Sbox_5_M50), 
        .B(SubBytesIns_Inst_Sbox_5_L0), .Z(SubBytesIns_Inst_Sbox_5_L13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_L14_U1 ( .A(SubBytesIns_Inst_Sbox_5_M52), 
        .B(SubBytesIns_Inst_Sbox_5_M61), .Z(SubBytesIns_Inst_Sbox_5_L14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_L15_U1 ( .A(SubBytesIns_Inst_Sbox_5_M55), 
        .B(SubBytesIns_Inst_Sbox_5_L1), .Z(SubBytesIns_Inst_Sbox_5_L15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_L16_U1 ( .A(SubBytesIns_Inst_Sbox_5_M56), 
        .B(SubBytesIns_Inst_Sbox_5_L0), .Z(SubBytesIns_Inst_Sbox_5_L16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_L17_U1 ( .A(SubBytesIns_Inst_Sbox_5_M57), 
        .B(SubBytesIns_Inst_Sbox_5_L1), .Z(SubBytesIns_Inst_Sbox_5_L17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_L18_U1 ( .A(SubBytesIns_Inst_Sbox_5_M58), 
        .B(SubBytesIns_Inst_Sbox_5_L8), .Z(SubBytesIns_Inst_Sbox_5_L18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_L19_U1 ( .A(SubBytesIns_Inst_Sbox_5_M63), 
        .B(SubBytesIns_Inst_Sbox_5_L4), .Z(SubBytesIns_Inst_Sbox_5_L19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_L20_U1 ( .A(SubBytesIns_Inst_Sbox_5_L0), 
        .B(SubBytesIns_Inst_Sbox_5_L1), .Z(SubBytesIns_Inst_Sbox_5_L20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_L21_U1 ( .A(SubBytesIns_Inst_Sbox_5_L1), 
        .B(SubBytesIns_Inst_Sbox_5_L7), .Z(SubBytesIns_Inst_Sbox_5_L21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_L22_U1 ( .A(SubBytesIns_Inst_Sbox_5_L3), 
        .B(SubBytesIns_Inst_Sbox_5_L12), .Z(SubBytesIns_Inst_Sbox_5_L22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_L23_U1 ( .A(SubBytesIns_Inst_Sbox_5_L18), 
        .B(SubBytesIns_Inst_Sbox_5_L2), .Z(SubBytesIns_Inst_Sbox_5_L23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_L24_U1 ( .A(SubBytesIns_Inst_Sbox_5_L15), 
        .B(SubBytesIns_Inst_Sbox_5_L9), .Z(SubBytesIns_Inst_Sbox_5_L24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_L25_U1 ( .A(SubBytesIns_Inst_Sbox_5_L6), 
        .B(SubBytesIns_Inst_Sbox_5_L10), .Z(SubBytesIns_Inst_Sbox_5_L25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_L26_U1 ( .A(SubBytesIns_Inst_Sbox_5_L7), 
        .B(SubBytesIns_Inst_Sbox_5_L9), .Z(SubBytesIns_Inst_Sbox_5_L26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_L27_U1 ( .A(SubBytesIns_Inst_Sbox_5_L8), 
        .B(SubBytesIns_Inst_Sbox_5_L10), .Z(SubBytesIns_Inst_Sbox_5_L27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_L28_U1 ( .A(SubBytesIns_Inst_Sbox_5_L11), 
        .B(SubBytesIns_Inst_Sbox_5_L14), .Z(SubBytesIns_Inst_Sbox_5_L28) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_L29_U1 ( .A(SubBytesIns_Inst_Sbox_5_L11), 
        .B(SubBytesIns_Inst_Sbox_5_L17), .Z(SubBytesIns_Inst_Sbox_5_L29) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_S0_U1 ( .A(SubBytesIns_Inst_Sbox_5_L6), 
        .B(SubBytesIns_Inst_Sbox_5_L24), .Z(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_S1_U1 ( .A(SubBytesIns_Inst_Sbox_5_L16), 
        .B(SubBytesIns_Inst_Sbox_5_L26), .ZN(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[15]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_S2_U1 ( .A(SubBytesIns_Inst_Sbox_5_L19), 
        .B(SubBytesIns_Inst_Sbox_5_L28), .ZN(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[14]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_S3_U1 ( .A(SubBytesIns_Inst_Sbox_5_L6), 
        .B(SubBytesIns_Inst_Sbox_5_L21), .Z(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[13]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_S4_U1 ( .A(SubBytesIns_Inst_Sbox_5_L20), 
        .B(SubBytesIns_Inst_Sbox_5_L22), .Z(MixColumnsInput[107]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_S5_U1 ( .A(SubBytesIns_Inst_Sbox_5_L25), 
        .B(SubBytesIns_Inst_Sbox_5_L29), .Z(MixColumnsInput[106]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_S6_U1 ( .A(SubBytesIns_Inst_Sbox_5_L13), 
        .B(SubBytesIns_Inst_Sbox_5_L27), .ZN(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[10]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_5_XOR_S7_U1 ( .A(SubBytesIns_Inst_Sbox_5_L6), 
        .B(SubBytesIns_Inst_Sbox_5_L23), .ZN(MixColumnsInput[104]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_T1_U1 ( .A(SubBytesInput[55]), .B(
        SubBytesInput[52]), .Z(SubBytesIns_Inst_Sbox_6_T1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_T2_U1 ( .A(SubBytesInput[55]), .B(
        SubBytesInput[50]), .Z(SubBytesIns_Inst_Sbox_6_T2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_T3_U1 ( .A(SubBytesInput[55]), .B(
        SubBytesInput[49]), .Z(SubBytesIns_Inst_Sbox_6_T3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_T4_U1 ( .A(SubBytesInput[52]), .B(
        SubBytesInput[50]), .Z(SubBytesIns_Inst_Sbox_6_T4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_T5_U1 ( .A(SubBytesInput[51]), .B(
        SubBytesInput[49]), .Z(SubBytesIns_Inst_Sbox_6_T5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_T6_U1 ( .A(SubBytesIns_Inst_Sbox_6_T1), 
        .B(SubBytesIns_Inst_Sbox_6_T5), .Z(SubBytesIns_Inst_Sbox_6_T6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_T7_U1 ( .A(SubBytesInput[54]), .B(
        SubBytesInput[53]), .Z(SubBytesIns_Inst_Sbox_6_T7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_T8_U1 ( .A(SubBytesInput[48]), .B(
        SubBytesIns_Inst_Sbox_6_T6), .Z(SubBytesIns_Inst_Sbox_6_T8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_T9_U1 ( .A(SubBytesInput[48]), .B(
        SubBytesIns_Inst_Sbox_6_T7), .Z(SubBytesIns_Inst_Sbox_6_T9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_T10_U1 ( .A(SubBytesIns_Inst_Sbox_6_T6), 
        .B(SubBytesIns_Inst_Sbox_6_T7), .Z(SubBytesIns_Inst_Sbox_6_T10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_T11_U1 ( .A(SubBytesInput[54]), .B(
        SubBytesInput[50]), .Z(SubBytesIns_Inst_Sbox_6_T11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_T12_U1 ( .A(SubBytesInput[53]), .B(
        SubBytesInput[50]), .Z(SubBytesIns_Inst_Sbox_6_T12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_T13_U1 ( .A(SubBytesIns_Inst_Sbox_6_T3), 
        .B(SubBytesIns_Inst_Sbox_6_T4), .Z(SubBytesIns_Inst_Sbox_6_T13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_T14_U1 ( .A(SubBytesIns_Inst_Sbox_6_T6), 
        .B(SubBytesIns_Inst_Sbox_6_T11), .Z(SubBytesIns_Inst_Sbox_6_T14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_T15_U1 ( .A(SubBytesIns_Inst_Sbox_6_T5), 
        .B(SubBytesIns_Inst_Sbox_6_T11), .Z(SubBytesIns_Inst_Sbox_6_T15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_T16_U1 ( .A(SubBytesIns_Inst_Sbox_6_T5), 
        .B(SubBytesIns_Inst_Sbox_6_T12), .Z(SubBytesIns_Inst_Sbox_6_T16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_T17_U1 ( .A(SubBytesIns_Inst_Sbox_6_T9), 
        .B(SubBytesIns_Inst_Sbox_6_T16), .Z(SubBytesIns_Inst_Sbox_6_T17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_T18_U1 ( .A(SubBytesInput[52]), .B(
        SubBytesInput[48]), .Z(SubBytesIns_Inst_Sbox_6_T18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_T19_U1 ( .A(SubBytesIns_Inst_Sbox_6_T7), 
        .B(SubBytesIns_Inst_Sbox_6_T18), .Z(SubBytesIns_Inst_Sbox_6_T19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_T20_U1 ( .A(SubBytesIns_Inst_Sbox_6_T1), 
        .B(SubBytesIns_Inst_Sbox_6_T19), .Z(SubBytesIns_Inst_Sbox_6_T20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_T21_U1 ( .A(SubBytesInput[49]), .B(
        SubBytesInput[48]), .Z(SubBytesIns_Inst_Sbox_6_T21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_T22_U1 ( .A(SubBytesIns_Inst_Sbox_6_T7), 
        .B(SubBytesIns_Inst_Sbox_6_T21), .Z(SubBytesIns_Inst_Sbox_6_T22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_T23_U1 ( .A(SubBytesIns_Inst_Sbox_6_T2), 
        .B(SubBytesIns_Inst_Sbox_6_T22), .Z(SubBytesIns_Inst_Sbox_6_T23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_T24_U1 ( .A(SubBytesIns_Inst_Sbox_6_T2), 
        .B(SubBytesIns_Inst_Sbox_6_T10), .Z(SubBytesIns_Inst_Sbox_6_T24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_T25_U1 ( .A(SubBytesIns_Inst_Sbox_6_T20), 
        .B(SubBytesIns_Inst_Sbox_6_T17), .Z(SubBytesIns_Inst_Sbox_6_T25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_T26_U1 ( .A(SubBytesIns_Inst_Sbox_6_T3), 
        .B(SubBytesIns_Inst_Sbox_6_T16), .Z(SubBytesIns_Inst_Sbox_6_T26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_T27_U1 ( .A(SubBytesIns_Inst_Sbox_6_T1), 
        .B(SubBytesIns_Inst_Sbox_6_T12), .Z(SubBytesIns_Inst_Sbox_6_T27) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M1_U1 ( .A1(SubBytesIns_Inst_Sbox_6_T13), 
        .A2(SubBytesIns_Inst_Sbox_6_T6), .ZN(SubBytesIns_Inst_Sbox_6_M1) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M2_U1 ( .A1(SubBytesIns_Inst_Sbox_6_T23), 
        .A2(SubBytesIns_Inst_Sbox_6_T8), .ZN(SubBytesIns_Inst_Sbox_6_M2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_M3_U1 ( .A(SubBytesIns_Inst_Sbox_6_T14), 
        .B(SubBytesIns_Inst_Sbox_6_M1), .Z(SubBytesIns_Inst_Sbox_6_M3) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M4_U1 ( .A1(SubBytesIns_Inst_Sbox_6_T19), 
        .A2(SubBytesInput[48]), .ZN(SubBytesIns_Inst_Sbox_6_M4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_M5_U1 ( .A(SubBytesIns_Inst_Sbox_6_M4), 
        .B(SubBytesIns_Inst_Sbox_6_M1), .Z(SubBytesIns_Inst_Sbox_6_M5) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M6_U1 ( .A1(SubBytesIns_Inst_Sbox_6_T3), 
        .A2(SubBytesIns_Inst_Sbox_6_T16), .ZN(SubBytesIns_Inst_Sbox_6_M6) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M7_U1 ( .A1(SubBytesIns_Inst_Sbox_6_T22), 
        .A2(SubBytesIns_Inst_Sbox_6_T9), .ZN(SubBytesIns_Inst_Sbox_6_M7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_M8_U1 ( .A(SubBytesIns_Inst_Sbox_6_T26), 
        .B(SubBytesIns_Inst_Sbox_6_M6), .Z(SubBytesIns_Inst_Sbox_6_M8) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M9_U1 ( .A1(SubBytesIns_Inst_Sbox_6_T20), 
        .A2(SubBytesIns_Inst_Sbox_6_T17), .ZN(SubBytesIns_Inst_Sbox_6_M9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_M10_U1 ( .A(SubBytesIns_Inst_Sbox_6_M9), 
        .B(SubBytesIns_Inst_Sbox_6_M6), .Z(SubBytesIns_Inst_Sbox_6_M10) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M11_U1 ( .A1(SubBytesIns_Inst_Sbox_6_T1), 
        .A2(SubBytesIns_Inst_Sbox_6_T15), .ZN(SubBytesIns_Inst_Sbox_6_M11) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M12_U1 ( .A1(SubBytesIns_Inst_Sbox_6_T4), 
        .A2(SubBytesIns_Inst_Sbox_6_T27), .ZN(SubBytesIns_Inst_Sbox_6_M12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_M13_U1 ( .A(SubBytesIns_Inst_Sbox_6_M12), 
        .B(SubBytesIns_Inst_Sbox_6_M11), .Z(SubBytesIns_Inst_Sbox_6_M13) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M14_U1 ( .A1(SubBytesIns_Inst_Sbox_6_T2), 
        .A2(SubBytesIns_Inst_Sbox_6_T10), .ZN(SubBytesIns_Inst_Sbox_6_M14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_M15_U1 ( .A(SubBytesIns_Inst_Sbox_6_M14), 
        .B(SubBytesIns_Inst_Sbox_6_M11), .Z(SubBytesIns_Inst_Sbox_6_M15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_M16_U1 ( .A(SubBytesIns_Inst_Sbox_6_M3), 
        .B(SubBytesIns_Inst_Sbox_6_M2), .Z(SubBytesIns_Inst_Sbox_6_M16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_M17_U1 ( .A(SubBytesIns_Inst_Sbox_6_M5), 
        .B(SubBytesIns_Inst_Sbox_6_T24), .Z(SubBytesIns_Inst_Sbox_6_M17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_M18_U1 ( .A(SubBytesIns_Inst_Sbox_6_M8), 
        .B(SubBytesIns_Inst_Sbox_6_M7), .Z(SubBytesIns_Inst_Sbox_6_M18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_M19_U1 ( .A(SubBytesIns_Inst_Sbox_6_M10), 
        .B(SubBytesIns_Inst_Sbox_6_M15), .Z(SubBytesIns_Inst_Sbox_6_M19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_M20_U1 ( .A(SubBytesIns_Inst_Sbox_6_M16), 
        .B(SubBytesIns_Inst_Sbox_6_M13), .Z(SubBytesIns_Inst_Sbox_6_M20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_M21_U1 ( .A(SubBytesIns_Inst_Sbox_6_M17), 
        .B(SubBytesIns_Inst_Sbox_6_M15), .Z(SubBytesIns_Inst_Sbox_6_M21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_M22_U1 ( .A(SubBytesIns_Inst_Sbox_6_M18), 
        .B(SubBytesIns_Inst_Sbox_6_M13), .Z(SubBytesIns_Inst_Sbox_6_M22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_M23_U1 ( .A(SubBytesIns_Inst_Sbox_6_M19), 
        .B(SubBytesIns_Inst_Sbox_6_T25), .Z(SubBytesIns_Inst_Sbox_6_M23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_M24_U1 ( .A(SubBytesIns_Inst_Sbox_6_M22), 
        .B(SubBytesIns_Inst_Sbox_6_M23), .Z(SubBytesIns_Inst_Sbox_6_M24) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M25_U1 ( .A1(SubBytesIns_Inst_Sbox_6_M22), .A2(SubBytesIns_Inst_Sbox_6_M20), .ZN(SubBytesIns_Inst_Sbox_6_M25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_M26_U1 ( .A(SubBytesIns_Inst_Sbox_6_M21), 
        .B(SubBytesIns_Inst_Sbox_6_M25), .Z(SubBytesIns_Inst_Sbox_6_M26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_M27_U1 ( .A(SubBytesIns_Inst_Sbox_6_M20), 
        .B(SubBytesIns_Inst_Sbox_6_M21), .Z(SubBytesIns_Inst_Sbox_6_M27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_M28_U1 ( .A(SubBytesIns_Inst_Sbox_6_M23), 
        .B(SubBytesIns_Inst_Sbox_6_M25), .Z(SubBytesIns_Inst_Sbox_6_M28) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M29_U1 ( .A1(SubBytesIns_Inst_Sbox_6_M28), .A2(SubBytesIns_Inst_Sbox_6_M27), .ZN(SubBytesIns_Inst_Sbox_6_M29) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M30_U1 ( .A1(SubBytesIns_Inst_Sbox_6_M26), .A2(SubBytesIns_Inst_Sbox_6_M24), .ZN(SubBytesIns_Inst_Sbox_6_M30) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M31_U1 ( .A1(SubBytesIns_Inst_Sbox_6_M20), .A2(SubBytesIns_Inst_Sbox_6_M23), .ZN(SubBytesIns_Inst_Sbox_6_M31) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M32_U1 ( .A1(SubBytesIns_Inst_Sbox_6_M27), .A2(SubBytesIns_Inst_Sbox_6_M31), .ZN(SubBytesIns_Inst_Sbox_6_M32) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_M33_U1 ( .A(SubBytesIns_Inst_Sbox_6_M27), 
        .B(SubBytesIns_Inst_Sbox_6_M25), .Z(SubBytesIns_Inst_Sbox_6_M33) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M34_U1 ( .A1(SubBytesIns_Inst_Sbox_6_M21), .A2(SubBytesIns_Inst_Sbox_6_M22), .ZN(SubBytesIns_Inst_Sbox_6_M34) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M35_U1 ( .A1(SubBytesIns_Inst_Sbox_6_M24), .A2(SubBytesIns_Inst_Sbox_6_M34), .ZN(SubBytesIns_Inst_Sbox_6_M35) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_M36_U1 ( .A(SubBytesIns_Inst_Sbox_6_M24), 
        .B(SubBytesIns_Inst_Sbox_6_M25), .Z(SubBytesIns_Inst_Sbox_6_M36) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_M37_U1 ( .A(SubBytesIns_Inst_Sbox_6_M21), 
        .B(SubBytesIns_Inst_Sbox_6_M29), .Z(SubBytesIns_Inst_Sbox_6_M37) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_M38_U1 ( .A(SubBytesIns_Inst_Sbox_6_M32), 
        .B(SubBytesIns_Inst_Sbox_6_M33), .Z(SubBytesIns_Inst_Sbox_6_M38) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_M39_U1 ( .A(SubBytesIns_Inst_Sbox_6_M23), 
        .B(SubBytesIns_Inst_Sbox_6_M30), .Z(SubBytesIns_Inst_Sbox_6_M39) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_M40_U1 ( .A(SubBytesIns_Inst_Sbox_6_M35), 
        .B(SubBytesIns_Inst_Sbox_6_M36), .Z(SubBytesIns_Inst_Sbox_6_M40) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_M41_U1 ( .A(SubBytesIns_Inst_Sbox_6_M38), 
        .B(SubBytesIns_Inst_Sbox_6_M40), .Z(SubBytesIns_Inst_Sbox_6_M41) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_M42_U1 ( .A(SubBytesIns_Inst_Sbox_6_M37), 
        .B(SubBytesIns_Inst_Sbox_6_M39), .Z(SubBytesIns_Inst_Sbox_6_M42) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_M43_U1 ( .A(SubBytesIns_Inst_Sbox_6_M37), 
        .B(SubBytesIns_Inst_Sbox_6_M38), .Z(SubBytesIns_Inst_Sbox_6_M43) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_M44_U1 ( .A(SubBytesIns_Inst_Sbox_6_M39), 
        .B(SubBytesIns_Inst_Sbox_6_M40), .Z(SubBytesIns_Inst_Sbox_6_M44) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_M45_U1 ( .A(SubBytesIns_Inst_Sbox_6_M42), 
        .B(SubBytesIns_Inst_Sbox_6_M41), .Z(SubBytesIns_Inst_Sbox_6_M45) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M46_U1 ( .A1(SubBytesIns_Inst_Sbox_6_M44), .A2(SubBytesIns_Inst_Sbox_6_T6), .ZN(SubBytesIns_Inst_Sbox_6_M46) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M47_U1 ( .A1(SubBytesIns_Inst_Sbox_6_M40), .A2(SubBytesIns_Inst_Sbox_6_T8), .ZN(SubBytesIns_Inst_Sbox_6_M47) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M48_U1 ( .A1(SubBytesIns_Inst_Sbox_6_M39), .A2(SubBytesInput[48]), .ZN(SubBytesIns_Inst_Sbox_6_M48) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M49_U1 ( .A1(SubBytesIns_Inst_Sbox_6_M43), .A2(SubBytesIns_Inst_Sbox_6_T16), .ZN(SubBytesIns_Inst_Sbox_6_M49) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M50_U1 ( .A1(SubBytesIns_Inst_Sbox_6_M38), .A2(SubBytesIns_Inst_Sbox_6_T9), .ZN(SubBytesIns_Inst_Sbox_6_M50) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M51_U1 ( .A1(SubBytesIns_Inst_Sbox_6_M37), .A2(SubBytesIns_Inst_Sbox_6_T17), .ZN(SubBytesIns_Inst_Sbox_6_M51) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M52_U1 ( .A1(SubBytesIns_Inst_Sbox_6_M42), .A2(SubBytesIns_Inst_Sbox_6_T15), .ZN(SubBytesIns_Inst_Sbox_6_M52) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M53_U1 ( .A1(SubBytesIns_Inst_Sbox_6_M45), .A2(SubBytesIns_Inst_Sbox_6_T27), .ZN(SubBytesIns_Inst_Sbox_6_M53) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M54_U1 ( .A1(SubBytesIns_Inst_Sbox_6_M41), .A2(SubBytesIns_Inst_Sbox_6_T10), .ZN(SubBytesIns_Inst_Sbox_6_M54) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M55_U1 ( .A1(SubBytesIns_Inst_Sbox_6_M44), .A2(SubBytesIns_Inst_Sbox_6_T13), .ZN(SubBytesIns_Inst_Sbox_6_M55) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M56_U1 ( .A1(SubBytesIns_Inst_Sbox_6_M40), .A2(SubBytesIns_Inst_Sbox_6_T23), .ZN(SubBytesIns_Inst_Sbox_6_M56) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M57_U1 ( .A1(SubBytesIns_Inst_Sbox_6_M39), .A2(SubBytesIns_Inst_Sbox_6_T19), .ZN(SubBytesIns_Inst_Sbox_6_M57) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M58_U1 ( .A1(SubBytesIns_Inst_Sbox_6_M43), .A2(SubBytesIns_Inst_Sbox_6_T3), .ZN(SubBytesIns_Inst_Sbox_6_M58) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M59_U1 ( .A1(SubBytesIns_Inst_Sbox_6_M38), .A2(SubBytesIns_Inst_Sbox_6_T22), .ZN(SubBytesIns_Inst_Sbox_6_M59) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M60_U1 ( .A1(SubBytesIns_Inst_Sbox_6_M37), .A2(SubBytesIns_Inst_Sbox_6_T20), .ZN(SubBytesIns_Inst_Sbox_6_M60) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M61_U1 ( .A1(SubBytesIns_Inst_Sbox_6_M42), .A2(SubBytesIns_Inst_Sbox_6_T1), .ZN(SubBytesIns_Inst_Sbox_6_M61) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M62_U1 ( .A1(SubBytesIns_Inst_Sbox_6_M45), .A2(SubBytesIns_Inst_Sbox_6_T4), .ZN(SubBytesIns_Inst_Sbox_6_M62) );
  AND2_X1 SubBytesIns_Inst_Sbox_6_AND_M63_U1 ( .A1(SubBytesIns_Inst_Sbox_6_M41), .A2(SubBytesIns_Inst_Sbox_6_T2), .ZN(SubBytesIns_Inst_Sbox_6_M63) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_L0_U1 ( .A(SubBytesIns_Inst_Sbox_6_M61), 
        .B(SubBytesIns_Inst_Sbox_6_M62), .Z(SubBytesIns_Inst_Sbox_6_L0) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_L1_U1 ( .A(SubBytesIns_Inst_Sbox_6_M50), 
        .B(SubBytesIns_Inst_Sbox_6_M56), .Z(SubBytesIns_Inst_Sbox_6_L1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_L2_U1 ( .A(SubBytesIns_Inst_Sbox_6_M46), 
        .B(SubBytesIns_Inst_Sbox_6_M48), .Z(SubBytesIns_Inst_Sbox_6_L2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_L3_U1 ( .A(SubBytesIns_Inst_Sbox_6_M47), 
        .B(SubBytesIns_Inst_Sbox_6_M55), .Z(SubBytesIns_Inst_Sbox_6_L3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_L4_U1 ( .A(SubBytesIns_Inst_Sbox_6_M54), 
        .B(SubBytesIns_Inst_Sbox_6_M58), .Z(SubBytesIns_Inst_Sbox_6_L4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_L5_U1 ( .A(SubBytesIns_Inst_Sbox_6_M49), 
        .B(SubBytesIns_Inst_Sbox_6_M61), .Z(SubBytesIns_Inst_Sbox_6_L5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_L6_U1 ( .A(SubBytesIns_Inst_Sbox_6_M62), 
        .B(SubBytesIns_Inst_Sbox_6_L5), .Z(SubBytesIns_Inst_Sbox_6_L6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_L7_U1 ( .A(SubBytesIns_Inst_Sbox_6_M46), 
        .B(SubBytesIns_Inst_Sbox_6_L3), .Z(SubBytesIns_Inst_Sbox_6_L7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_L8_U1 ( .A(SubBytesIns_Inst_Sbox_6_M51), 
        .B(SubBytesIns_Inst_Sbox_6_M59), .Z(SubBytesIns_Inst_Sbox_6_L8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_L9_U1 ( .A(SubBytesIns_Inst_Sbox_6_M52), 
        .B(SubBytesIns_Inst_Sbox_6_M53), .Z(SubBytesIns_Inst_Sbox_6_L9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_L10_U1 ( .A(SubBytesIns_Inst_Sbox_6_M53), 
        .B(SubBytesIns_Inst_Sbox_6_L4), .Z(SubBytesIns_Inst_Sbox_6_L10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_L11_U1 ( .A(SubBytesIns_Inst_Sbox_6_M60), 
        .B(SubBytesIns_Inst_Sbox_6_L2), .Z(SubBytesIns_Inst_Sbox_6_L11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_L12_U1 ( .A(SubBytesIns_Inst_Sbox_6_M48), 
        .B(SubBytesIns_Inst_Sbox_6_M51), .Z(SubBytesIns_Inst_Sbox_6_L12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_L13_U1 ( .A(SubBytesIns_Inst_Sbox_6_M50), 
        .B(SubBytesIns_Inst_Sbox_6_L0), .Z(SubBytesIns_Inst_Sbox_6_L13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_L14_U1 ( .A(SubBytesIns_Inst_Sbox_6_M52), 
        .B(SubBytesIns_Inst_Sbox_6_M61), .Z(SubBytesIns_Inst_Sbox_6_L14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_L15_U1 ( .A(SubBytesIns_Inst_Sbox_6_M55), 
        .B(SubBytesIns_Inst_Sbox_6_L1), .Z(SubBytesIns_Inst_Sbox_6_L15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_L16_U1 ( .A(SubBytesIns_Inst_Sbox_6_M56), 
        .B(SubBytesIns_Inst_Sbox_6_L0), .Z(SubBytesIns_Inst_Sbox_6_L16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_L17_U1 ( .A(SubBytesIns_Inst_Sbox_6_M57), 
        .B(SubBytesIns_Inst_Sbox_6_L1), .Z(SubBytesIns_Inst_Sbox_6_L17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_L18_U1 ( .A(SubBytesIns_Inst_Sbox_6_M58), 
        .B(SubBytesIns_Inst_Sbox_6_L8), .Z(SubBytesIns_Inst_Sbox_6_L18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_L19_U1 ( .A(SubBytesIns_Inst_Sbox_6_M63), 
        .B(SubBytesIns_Inst_Sbox_6_L4), .Z(SubBytesIns_Inst_Sbox_6_L19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_L20_U1 ( .A(SubBytesIns_Inst_Sbox_6_L0), 
        .B(SubBytesIns_Inst_Sbox_6_L1), .Z(SubBytesIns_Inst_Sbox_6_L20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_L21_U1 ( .A(SubBytesIns_Inst_Sbox_6_L1), 
        .B(SubBytesIns_Inst_Sbox_6_L7), .Z(SubBytesIns_Inst_Sbox_6_L21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_L22_U1 ( .A(SubBytesIns_Inst_Sbox_6_L3), 
        .B(SubBytesIns_Inst_Sbox_6_L12), .Z(SubBytesIns_Inst_Sbox_6_L22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_L23_U1 ( .A(SubBytesIns_Inst_Sbox_6_L18), 
        .B(SubBytesIns_Inst_Sbox_6_L2), .Z(SubBytesIns_Inst_Sbox_6_L23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_L24_U1 ( .A(SubBytesIns_Inst_Sbox_6_L15), 
        .B(SubBytesIns_Inst_Sbox_6_L9), .Z(SubBytesIns_Inst_Sbox_6_L24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_L25_U1 ( .A(SubBytesIns_Inst_Sbox_6_L6), 
        .B(SubBytesIns_Inst_Sbox_6_L10), .Z(SubBytesIns_Inst_Sbox_6_L25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_L26_U1 ( .A(SubBytesIns_Inst_Sbox_6_L7), 
        .B(SubBytesIns_Inst_Sbox_6_L9), .Z(SubBytesIns_Inst_Sbox_6_L26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_L27_U1 ( .A(SubBytesIns_Inst_Sbox_6_L8), 
        .B(SubBytesIns_Inst_Sbox_6_L10), .Z(SubBytesIns_Inst_Sbox_6_L27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_L28_U1 ( .A(SubBytesIns_Inst_Sbox_6_L11), 
        .B(SubBytesIns_Inst_Sbox_6_L14), .Z(SubBytesIns_Inst_Sbox_6_L28) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_L29_U1 ( .A(SubBytesIns_Inst_Sbox_6_L11), 
        .B(SubBytesIns_Inst_Sbox_6_L17), .Z(SubBytesIns_Inst_Sbox_6_L29) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_S0_U1 ( .A(SubBytesIns_Inst_Sbox_6_L6), 
        .B(SubBytesIns_Inst_Sbox_6_L24), .Z(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_S1_U1 ( .A(SubBytesIns_Inst_Sbox_6_L16), 
        .B(SubBytesIns_Inst_Sbox_6_L26), .ZN(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[23]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_S2_U1 ( .A(SubBytesIns_Inst_Sbox_6_L19), 
        .B(SubBytesIns_Inst_Sbox_6_L28), .ZN(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[22]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_S3_U1 ( .A(SubBytesIns_Inst_Sbox_6_L6), 
        .B(SubBytesIns_Inst_Sbox_6_L21), .Z(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[21]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_S4_U1 ( .A(SubBytesIns_Inst_Sbox_6_L20), 
        .B(SubBytesIns_Inst_Sbox_6_L22), .Z(MixColumnsInput[83]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_S5_U1 ( .A(SubBytesIns_Inst_Sbox_6_L25), 
        .B(SubBytesIns_Inst_Sbox_6_L29), .Z(MixColumnsInput[82]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_S6_U1 ( .A(SubBytesIns_Inst_Sbox_6_L13), 
        .B(SubBytesIns_Inst_Sbox_6_L27), .ZN(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[18]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_6_XOR_S7_U1 ( .A(SubBytesIns_Inst_Sbox_6_L6), 
        .B(SubBytesIns_Inst_Sbox_6_L23), .ZN(MixColumnsInput[80]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_T1_U1 ( .A(SubBytesInput[63]), .B(
        SubBytesInput[60]), .Z(SubBytesIns_Inst_Sbox_7_T1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_T2_U1 ( .A(SubBytesInput[63]), .B(
        SubBytesInput[58]), .Z(SubBytesIns_Inst_Sbox_7_T2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_T3_U1 ( .A(SubBytesInput[63]), .B(
        SubBytesInput[57]), .Z(SubBytesIns_Inst_Sbox_7_T3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_T4_U1 ( .A(SubBytesInput[60]), .B(
        SubBytesInput[58]), .Z(SubBytesIns_Inst_Sbox_7_T4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_T5_U1 ( .A(SubBytesInput[59]), .B(
        SubBytesInput[57]), .Z(SubBytesIns_Inst_Sbox_7_T5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_T6_U1 ( .A(SubBytesIns_Inst_Sbox_7_T1), 
        .B(SubBytesIns_Inst_Sbox_7_T5), .Z(SubBytesIns_Inst_Sbox_7_T6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_T7_U1 ( .A(SubBytesInput[62]), .B(
        SubBytesInput[61]), .Z(SubBytesIns_Inst_Sbox_7_T7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_T8_U1 ( .A(SubBytesInput[56]), .B(
        SubBytesIns_Inst_Sbox_7_T6), .Z(SubBytesIns_Inst_Sbox_7_T8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_T9_U1 ( .A(SubBytesInput[56]), .B(
        SubBytesIns_Inst_Sbox_7_T7), .Z(SubBytesIns_Inst_Sbox_7_T9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_T10_U1 ( .A(SubBytesIns_Inst_Sbox_7_T6), 
        .B(SubBytesIns_Inst_Sbox_7_T7), .Z(SubBytesIns_Inst_Sbox_7_T10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_T11_U1 ( .A(SubBytesInput[62]), .B(
        SubBytesInput[58]), .Z(SubBytesIns_Inst_Sbox_7_T11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_T12_U1 ( .A(SubBytesInput[61]), .B(
        SubBytesInput[58]), .Z(SubBytesIns_Inst_Sbox_7_T12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_T13_U1 ( .A(SubBytesIns_Inst_Sbox_7_T3), 
        .B(SubBytesIns_Inst_Sbox_7_T4), .Z(SubBytesIns_Inst_Sbox_7_T13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_T14_U1 ( .A(SubBytesIns_Inst_Sbox_7_T6), 
        .B(SubBytesIns_Inst_Sbox_7_T11), .Z(SubBytesIns_Inst_Sbox_7_T14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_T15_U1 ( .A(SubBytesIns_Inst_Sbox_7_T5), 
        .B(SubBytesIns_Inst_Sbox_7_T11), .Z(SubBytesIns_Inst_Sbox_7_T15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_T16_U1 ( .A(SubBytesIns_Inst_Sbox_7_T5), 
        .B(SubBytesIns_Inst_Sbox_7_T12), .Z(SubBytesIns_Inst_Sbox_7_T16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_T17_U1 ( .A(SubBytesIns_Inst_Sbox_7_T9), 
        .B(SubBytesIns_Inst_Sbox_7_T16), .Z(SubBytesIns_Inst_Sbox_7_T17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_T18_U1 ( .A(SubBytesInput[60]), .B(
        SubBytesInput[56]), .Z(SubBytesIns_Inst_Sbox_7_T18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_T19_U1 ( .A(SubBytesIns_Inst_Sbox_7_T7), 
        .B(SubBytesIns_Inst_Sbox_7_T18), .Z(SubBytesIns_Inst_Sbox_7_T19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_T20_U1 ( .A(SubBytesIns_Inst_Sbox_7_T1), 
        .B(SubBytesIns_Inst_Sbox_7_T19), .Z(SubBytesIns_Inst_Sbox_7_T20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_T21_U1 ( .A(SubBytesInput[57]), .B(
        SubBytesInput[56]), .Z(SubBytesIns_Inst_Sbox_7_T21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_T22_U1 ( .A(SubBytesIns_Inst_Sbox_7_T7), 
        .B(SubBytesIns_Inst_Sbox_7_T21), .Z(SubBytesIns_Inst_Sbox_7_T22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_T23_U1 ( .A(SubBytesIns_Inst_Sbox_7_T2), 
        .B(SubBytesIns_Inst_Sbox_7_T22), .Z(SubBytesIns_Inst_Sbox_7_T23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_T24_U1 ( .A(SubBytesIns_Inst_Sbox_7_T2), 
        .B(SubBytesIns_Inst_Sbox_7_T10), .Z(SubBytesIns_Inst_Sbox_7_T24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_T25_U1 ( .A(SubBytesIns_Inst_Sbox_7_T20), 
        .B(SubBytesIns_Inst_Sbox_7_T17), .Z(SubBytesIns_Inst_Sbox_7_T25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_T26_U1 ( .A(SubBytesIns_Inst_Sbox_7_T3), 
        .B(SubBytesIns_Inst_Sbox_7_T16), .Z(SubBytesIns_Inst_Sbox_7_T26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_T27_U1 ( .A(SubBytesIns_Inst_Sbox_7_T1), 
        .B(SubBytesIns_Inst_Sbox_7_T12), .Z(SubBytesIns_Inst_Sbox_7_T27) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M1_U1 ( .A1(SubBytesIns_Inst_Sbox_7_T13), 
        .A2(SubBytesIns_Inst_Sbox_7_T6), .ZN(SubBytesIns_Inst_Sbox_7_M1) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M2_U1 ( .A1(SubBytesIns_Inst_Sbox_7_T23), 
        .A2(SubBytesIns_Inst_Sbox_7_T8), .ZN(SubBytesIns_Inst_Sbox_7_M2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_M3_U1 ( .A(SubBytesIns_Inst_Sbox_7_T14), 
        .B(SubBytesIns_Inst_Sbox_7_M1), .Z(SubBytesIns_Inst_Sbox_7_M3) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M4_U1 ( .A1(SubBytesIns_Inst_Sbox_7_T19), 
        .A2(SubBytesInput[56]), .ZN(SubBytesIns_Inst_Sbox_7_M4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_M5_U1 ( .A(SubBytesIns_Inst_Sbox_7_M4), 
        .B(SubBytesIns_Inst_Sbox_7_M1), .Z(SubBytesIns_Inst_Sbox_7_M5) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M6_U1 ( .A1(SubBytesIns_Inst_Sbox_7_T3), 
        .A2(SubBytesIns_Inst_Sbox_7_T16), .ZN(SubBytesIns_Inst_Sbox_7_M6) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M7_U1 ( .A1(SubBytesIns_Inst_Sbox_7_T22), 
        .A2(SubBytesIns_Inst_Sbox_7_T9), .ZN(SubBytesIns_Inst_Sbox_7_M7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_M8_U1 ( .A(SubBytesIns_Inst_Sbox_7_T26), 
        .B(SubBytesIns_Inst_Sbox_7_M6), .Z(SubBytesIns_Inst_Sbox_7_M8) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M9_U1 ( .A1(SubBytesIns_Inst_Sbox_7_T20), 
        .A2(SubBytesIns_Inst_Sbox_7_T17), .ZN(SubBytesIns_Inst_Sbox_7_M9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_M10_U1 ( .A(SubBytesIns_Inst_Sbox_7_M9), 
        .B(SubBytesIns_Inst_Sbox_7_M6), .Z(SubBytesIns_Inst_Sbox_7_M10) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M11_U1 ( .A1(SubBytesIns_Inst_Sbox_7_T1), 
        .A2(SubBytesIns_Inst_Sbox_7_T15), .ZN(SubBytesIns_Inst_Sbox_7_M11) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M12_U1 ( .A1(SubBytesIns_Inst_Sbox_7_T4), 
        .A2(SubBytesIns_Inst_Sbox_7_T27), .ZN(SubBytesIns_Inst_Sbox_7_M12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_M13_U1 ( .A(SubBytesIns_Inst_Sbox_7_M12), 
        .B(SubBytesIns_Inst_Sbox_7_M11), .Z(SubBytesIns_Inst_Sbox_7_M13) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M14_U1 ( .A1(SubBytesIns_Inst_Sbox_7_T2), 
        .A2(SubBytesIns_Inst_Sbox_7_T10), .ZN(SubBytesIns_Inst_Sbox_7_M14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_M15_U1 ( .A(SubBytesIns_Inst_Sbox_7_M14), 
        .B(SubBytesIns_Inst_Sbox_7_M11), .Z(SubBytesIns_Inst_Sbox_7_M15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_M16_U1 ( .A(SubBytesIns_Inst_Sbox_7_M3), 
        .B(SubBytesIns_Inst_Sbox_7_M2), .Z(SubBytesIns_Inst_Sbox_7_M16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_M17_U1 ( .A(SubBytesIns_Inst_Sbox_7_M5), 
        .B(SubBytesIns_Inst_Sbox_7_T24), .Z(SubBytesIns_Inst_Sbox_7_M17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_M18_U1 ( .A(SubBytesIns_Inst_Sbox_7_M8), 
        .B(SubBytesIns_Inst_Sbox_7_M7), .Z(SubBytesIns_Inst_Sbox_7_M18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_M19_U1 ( .A(SubBytesIns_Inst_Sbox_7_M10), 
        .B(SubBytesIns_Inst_Sbox_7_M15), .Z(SubBytesIns_Inst_Sbox_7_M19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_M20_U1 ( .A(SubBytesIns_Inst_Sbox_7_M16), 
        .B(SubBytesIns_Inst_Sbox_7_M13), .Z(SubBytesIns_Inst_Sbox_7_M20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_M21_U1 ( .A(SubBytesIns_Inst_Sbox_7_M17), 
        .B(SubBytesIns_Inst_Sbox_7_M15), .Z(SubBytesIns_Inst_Sbox_7_M21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_M22_U1 ( .A(SubBytesIns_Inst_Sbox_7_M18), 
        .B(SubBytesIns_Inst_Sbox_7_M13), .Z(SubBytesIns_Inst_Sbox_7_M22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_M23_U1 ( .A(SubBytesIns_Inst_Sbox_7_M19), 
        .B(SubBytesIns_Inst_Sbox_7_T25), .Z(SubBytesIns_Inst_Sbox_7_M23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_M24_U1 ( .A(SubBytesIns_Inst_Sbox_7_M22), 
        .B(SubBytesIns_Inst_Sbox_7_M23), .Z(SubBytesIns_Inst_Sbox_7_M24) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M25_U1 ( .A1(SubBytesIns_Inst_Sbox_7_M22), .A2(SubBytesIns_Inst_Sbox_7_M20), .ZN(SubBytesIns_Inst_Sbox_7_M25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_M26_U1 ( .A(SubBytesIns_Inst_Sbox_7_M21), 
        .B(SubBytesIns_Inst_Sbox_7_M25), .Z(SubBytesIns_Inst_Sbox_7_M26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_M27_U1 ( .A(SubBytesIns_Inst_Sbox_7_M20), 
        .B(SubBytesIns_Inst_Sbox_7_M21), .Z(SubBytesIns_Inst_Sbox_7_M27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_M28_U1 ( .A(SubBytesIns_Inst_Sbox_7_M23), 
        .B(SubBytesIns_Inst_Sbox_7_M25), .Z(SubBytesIns_Inst_Sbox_7_M28) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M29_U1 ( .A1(SubBytesIns_Inst_Sbox_7_M28), .A2(SubBytesIns_Inst_Sbox_7_M27), .ZN(SubBytesIns_Inst_Sbox_7_M29) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M30_U1 ( .A1(SubBytesIns_Inst_Sbox_7_M26), .A2(SubBytesIns_Inst_Sbox_7_M24), .ZN(SubBytesIns_Inst_Sbox_7_M30) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M31_U1 ( .A1(SubBytesIns_Inst_Sbox_7_M20), .A2(SubBytesIns_Inst_Sbox_7_M23), .ZN(SubBytesIns_Inst_Sbox_7_M31) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M32_U1 ( .A1(SubBytesIns_Inst_Sbox_7_M27), .A2(SubBytesIns_Inst_Sbox_7_M31), .ZN(SubBytesIns_Inst_Sbox_7_M32) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_M33_U1 ( .A(SubBytesIns_Inst_Sbox_7_M27), 
        .B(SubBytesIns_Inst_Sbox_7_M25), .Z(SubBytesIns_Inst_Sbox_7_M33) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M34_U1 ( .A1(SubBytesIns_Inst_Sbox_7_M21), .A2(SubBytesIns_Inst_Sbox_7_M22), .ZN(SubBytesIns_Inst_Sbox_7_M34) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M35_U1 ( .A1(SubBytesIns_Inst_Sbox_7_M24), .A2(SubBytesIns_Inst_Sbox_7_M34), .ZN(SubBytesIns_Inst_Sbox_7_M35) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_M36_U1 ( .A(SubBytesIns_Inst_Sbox_7_M24), 
        .B(SubBytesIns_Inst_Sbox_7_M25), .Z(SubBytesIns_Inst_Sbox_7_M36) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_M37_U1 ( .A(SubBytesIns_Inst_Sbox_7_M21), 
        .B(SubBytesIns_Inst_Sbox_7_M29), .Z(SubBytesIns_Inst_Sbox_7_M37) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_M38_U1 ( .A(SubBytesIns_Inst_Sbox_7_M32), 
        .B(SubBytesIns_Inst_Sbox_7_M33), .Z(SubBytesIns_Inst_Sbox_7_M38) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_M39_U1 ( .A(SubBytesIns_Inst_Sbox_7_M23), 
        .B(SubBytesIns_Inst_Sbox_7_M30), .Z(SubBytesIns_Inst_Sbox_7_M39) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_M40_U1 ( .A(SubBytesIns_Inst_Sbox_7_M35), 
        .B(SubBytesIns_Inst_Sbox_7_M36), .Z(SubBytesIns_Inst_Sbox_7_M40) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_M41_U1 ( .A(SubBytesIns_Inst_Sbox_7_M38), 
        .B(SubBytesIns_Inst_Sbox_7_M40), .Z(SubBytesIns_Inst_Sbox_7_M41) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_M42_U1 ( .A(SubBytesIns_Inst_Sbox_7_M37), 
        .B(SubBytesIns_Inst_Sbox_7_M39), .Z(SubBytesIns_Inst_Sbox_7_M42) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_M43_U1 ( .A(SubBytesIns_Inst_Sbox_7_M37), 
        .B(SubBytesIns_Inst_Sbox_7_M38), .Z(SubBytesIns_Inst_Sbox_7_M43) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_M44_U1 ( .A(SubBytesIns_Inst_Sbox_7_M39), 
        .B(SubBytesIns_Inst_Sbox_7_M40), .Z(SubBytesIns_Inst_Sbox_7_M44) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_M45_U1 ( .A(SubBytesIns_Inst_Sbox_7_M42), 
        .B(SubBytesIns_Inst_Sbox_7_M41), .Z(SubBytesIns_Inst_Sbox_7_M45) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M46_U1 ( .A1(SubBytesIns_Inst_Sbox_7_M44), .A2(SubBytesIns_Inst_Sbox_7_T6), .ZN(SubBytesIns_Inst_Sbox_7_M46) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M47_U1 ( .A1(SubBytesIns_Inst_Sbox_7_M40), .A2(SubBytesIns_Inst_Sbox_7_T8), .ZN(SubBytesIns_Inst_Sbox_7_M47) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M48_U1 ( .A1(SubBytesIns_Inst_Sbox_7_M39), .A2(SubBytesInput[56]), .ZN(SubBytesIns_Inst_Sbox_7_M48) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M49_U1 ( .A1(SubBytesIns_Inst_Sbox_7_M43), .A2(SubBytesIns_Inst_Sbox_7_T16), .ZN(SubBytesIns_Inst_Sbox_7_M49) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M50_U1 ( .A1(SubBytesIns_Inst_Sbox_7_M38), .A2(SubBytesIns_Inst_Sbox_7_T9), .ZN(SubBytesIns_Inst_Sbox_7_M50) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M51_U1 ( .A1(SubBytesIns_Inst_Sbox_7_M37), .A2(SubBytesIns_Inst_Sbox_7_T17), .ZN(SubBytesIns_Inst_Sbox_7_M51) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M52_U1 ( .A1(SubBytesIns_Inst_Sbox_7_M42), .A2(SubBytesIns_Inst_Sbox_7_T15), .ZN(SubBytesIns_Inst_Sbox_7_M52) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M53_U1 ( .A1(SubBytesIns_Inst_Sbox_7_M45), .A2(SubBytesIns_Inst_Sbox_7_T27), .ZN(SubBytesIns_Inst_Sbox_7_M53) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M54_U1 ( .A1(SubBytesIns_Inst_Sbox_7_M41), .A2(SubBytesIns_Inst_Sbox_7_T10), .ZN(SubBytesIns_Inst_Sbox_7_M54) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M55_U1 ( .A1(SubBytesIns_Inst_Sbox_7_M44), .A2(SubBytesIns_Inst_Sbox_7_T13), .ZN(SubBytesIns_Inst_Sbox_7_M55) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M56_U1 ( .A1(SubBytesIns_Inst_Sbox_7_M40), .A2(SubBytesIns_Inst_Sbox_7_T23), .ZN(SubBytesIns_Inst_Sbox_7_M56) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M57_U1 ( .A1(SubBytesIns_Inst_Sbox_7_M39), .A2(SubBytesIns_Inst_Sbox_7_T19), .ZN(SubBytesIns_Inst_Sbox_7_M57) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M58_U1 ( .A1(SubBytesIns_Inst_Sbox_7_M43), .A2(SubBytesIns_Inst_Sbox_7_T3), .ZN(SubBytesIns_Inst_Sbox_7_M58) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M59_U1 ( .A1(SubBytesIns_Inst_Sbox_7_M38), .A2(SubBytesIns_Inst_Sbox_7_T22), .ZN(SubBytesIns_Inst_Sbox_7_M59) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M60_U1 ( .A1(SubBytesIns_Inst_Sbox_7_M37), .A2(SubBytesIns_Inst_Sbox_7_T20), .ZN(SubBytesIns_Inst_Sbox_7_M60) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M61_U1 ( .A1(SubBytesIns_Inst_Sbox_7_M42), .A2(SubBytesIns_Inst_Sbox_7_T1), .ZN(SubBytesIns_Inst_Sbox_7_M61) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M62_U1 ( .A1(SubBytesIns_Inst_Sbox_7_M45), .A2(SubBytesIns_Inst_Sbox_7_T4), .ZN(SubBytesIns_Inst_Sbox_7_M62) );
  AND2_X1 SubBytesIns_Inst_Sbox_7_AND_M63_U1 ( .A1(SubBytesIns_Inst_Sbox_7_M41), .A2(SubBytesIns_Inst_Sbox_7_T2), .ZN(SubBytesIns_Inst_Sbox_7_M63) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_L0_U1 ( .A(SubBytesIns_Inst_Sbox_7_M61), 
        .B(SubBytesIns_Inst_Sbox_7_M62), .Z(SubBytesIns_Inst_Sbox_7_L0) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_L1_U1 ( .A(SubBytesIns_Inst_Sbox_7_M50), 
        .B(SubBytesIns_Inst_Sbox_7_M56), .Z(SubBytesIns_Inst_Sbox_7_L1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_L2_U1 ( .A(SubBytesIns_Inst_Sbox_7_M46), 
        .B(SubBytesIns_Inst_Sbox_7_M48), .Z(SubBytesIns_Inst_Sbox_7_L2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_L3_U1 ( .A(SubBytesIns_Inst_Sbox_7_M47), 
        .B(SubBytesIns_Inst_Sbox_7_M55), .Z(SubBytesIns_Inst_Sbox_7_L3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_L4_U1 ( .A(SubBytesIns_Inst_Sbox_7_M54), 
        .B(SubBytesIns_Inst_Sbox_7_M58), .Z(SubBytesIns_Inst_Sbox_7_L4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_L5_U1 ( .A(SubBytesIns_Inst_Sbox_7_M49), 
        .B(SubBytesIns_Inst_Sbox_7_M61), .Z(SubBytesIns_Inst_Sbox_7_L5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_L6_U1 ( .A(SubBytesIns_Inst_Sbox_7_M62), 
        .B(SubBytesIns_Inst_Sbox_7_L5), .Z(SubBytesIns_Inst_Sbox_7_L6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_L7_U1 ( .A(SubBytesIns_Inst_Sbox_7_M46), 
        .B(SubBytesIns_Inst_Sbox_7_L3), .Z(SubBytesIns_Inst_Sbox_7_L7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_L8_U1 ( .A(SubBytesIns_Inst_Sbox_7_M51), 
        .B(SubBytesIns_Inst_Sbox_7_M59), .Z(SubBytesIns_Inst_Sbox_7_L8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_L9_U1 ( .A(SubBytesIns_Inst_Sbox_7_M52), 
        .B(SubBytesIns_Inst_Sbox_7_M53), .Z(SubBytesIns_Inst_Sbox_7_L9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_L10_U1 ( .A(SubBytesIns_Inst_Sbox_7_M53), 
        .B(SubBytesIns_Inst_Sbox_7_L4), .Z(SubBytesIns_Inst_Sbox_7_L10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_L11_U1 ( .A(SubBytesIns_Inst_Sbox_7_M60), 
        .B(SubBytesIns_Inst_Sbox_7_L2), .Z(SubBytesIns_Inst_Sbox_7_L11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_L12_U1 ( .A(SubBytesIns_Inst_Sbox_7_M48), 
        .B(SubBytesIns_Inst_Sbox_7_M51), .Z(SubBytesIns_Inst_Sbox_7_L12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_L13_U1 ( .A(SubBytesIns_Inst_Sbox_7_M50), 
        .B(SubBytesIns_Inst_Sbox_7_L0), .Z(SubBytesIns_Inst_Sbox_7_L13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_L14_U1 ( .A(SubBytesIns_Inst_Sbox_7_M52), 
        .B(SubBytesIns_Inst_Sbox_7_M61), .Z(SubBytesIns_Inst_Sbox_7_L14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_L15_U1 ( .A(SubBytesIns_Inst_Sbox_7_M55), 
        .B(SubBytesIns_Inst_Sbox_7_L1), .Z(SubBytesIns_Inst_Sbox_7_L15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_L16_U1 ( .A(SubBytesIns_Inst_Sbox_7_M56), 
        .B(SubBytesIns_Inst_Sbox_7_L0), .Z(SubBytesIns_Inst_Sbox_7_L16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_L17_U1 ( .A(SubBytesIns_Inst_Sbox_7_M57), 
        .B(SubBytesIns_Inst_Sbox_7_L1), .Z(SubBytesIns_Inst_Sbox_7_L17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_L18_U1 ( .A(SubBytesIns_Inst_Sbox_7_M58), 
        .B(SubBytesIns_Inst_Sbox_7_L8), .Z(SubBytesIns_Inst_Sbox_7_L18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_L19_U1 ( .A(SubBytesIns_Inst_Sbox_7_M63), 
        .B(SubBytesIns_Inst_Sbox_7_L4), .Z(SubBytesIns_Inst_Sbox_7_L19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_L20_U1 ( .A(SubBytesIns_Inst_Sbox_7_L0), 
        .B(SubBytesIns_Inst_Sbox_7_L1), .Z(SubBytesIns_Inst_Sbox_7_L20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_L21_U1 ( .A(SubBytesIns_Inst_Sbox_7_L1), 
        .B(SubBytesIns_Inst_Sbox_7_L7), .Z(SubBytesIns_Inst_Sbox_7_L21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_L22_U1 ( .A(SubBytesIns_Inst_Sbox_7_L3), 
        .B(SubBytesIns_Inst_Sbox_7_L12), .Z(SubBytesIns_Inst_Sbox_7_L22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_L23_U1 ( .A(SubBytesIns_Inst_Sbox_7_L18), 
        .B(SubBytesIns_Inst_Sbox_7_L2), .Z(SubBytesIns_Inst_Sbox_7_L23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_L24_U1 ( .A(SubBytesIns_Inst_Sbox_7_L15), 
        .B(SubBytesIns_Inst_Sbox_7_L9), .Z(SubBytesIns_Inst_Sbox_7_L24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_L25_U1 ( .A(SubBytesIns_Inst_Sbox_7_L6), 
        .B(SubBytesIns_Inst_Sbox_7_L10), .Z(SubBytesIns_Inst_Sbox_7_L25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_L26_U1 ( .A(SubBytesIns_Inst_Sbox_7_L7), 
        .B(SubBytesIns_Inst_Sbox_7_L9), .Z(SubBytesIns_Inst_Sbox_7_L26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_L27_U1 ( .A(SubBytesIns_Inst_Sbox_7_L8), 
        .B(SubBytesIns_Inst_Sbox_7_L10), .Z(SubBytesIns_Inst_Sbox_7_L27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_L28_U1 ( .A(SubBytesIns_Inst_Sbox_7_L11), 
        .B(SubBytesIns_Inst_Sbox_7_L14), .Z(SubBytesIns_Inst_Sbox_7_L28) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_L29_U1 ( .A(SubBytesIns_Inst_Sbox_7_L11), 
        .B(SubBytesIns_Inst_Sbox_7_L17), .Z(SubBytesIns_Inst_Sbox_7_L29) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_S0_U1 ( .A(SubBytesIns_Inst_Sbox_7_L6), 
        .B(SubBytesIns_Inst_Sbox_7_L24), .Z(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_S1_U1 ( .A(SubBytesIns_Inst_Sbox_7_L16), 
        .B(SubBytesIns_Inst_Sbox_7_L26), .ZN(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[31]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_S2_U1 ( .A(SubBytesIns_Inst_Sbox_7_L19), 
        .B(SubBytesIns_Inst_Sbox_7_L28), .ZN(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[30]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_S3_U1 ( .A(SubBytesIns_Inst_Sbox_7_L6), 
        .B(SubBytesIns_Inst_Sbox_7_L21), .Z(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[29]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_S4_U1 ( .A(SubBytesIns_Inst_Sbox_7_L20), 
        .B(SubBytesIns_Inst_Sbox_7_L22), .Z(MixColumnsInput[59]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_S5_U1 ( .A(SubBytesIns_Inst_Sbox_7_L25), 
        .B(SubBytesIns_Inst_Sbox_7_L29), .Z(MixColumnsInput[58]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_S6_U1 ( .A(SubBytesIns_Inst_Sbox_7_L13), 
        .B(SubBytesIns_Inst_Sbox_7_L27), .ZN(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[26]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_7_XOR_S7_U1 ( .A(SubBytesIns_Inst_Sbox_7_L6), 
        .B(SubBytesIns_Inst_Sbox_7_L23), .ZN(MixColumnsInput[56]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_T1_U1 ( .A(SubBytesInput[71]), .B(
        SubBytesInput[68]), .Z(SubBytesIns_Inst_Sbox_8_T1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_T2_U1 ( .A(SubBytesInput[71]), .B(
        SubBytesInput[66]), .Z(SubBytesIns_Inst_Sbox_8_T2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_T3_U1 ( .A(SubBytesInput[71]), .B(
        SubBytesInput[65]), .Z(SubBytesIns_Inst_Sbox_8_T3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_T4_U1 ( .A(SubBytesInput[68]), .B(
        SubBytesInput[66]), .Z(SubBytesIns_Inst_Sbox_8_T4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_T5_U1 ( .A(SubBytesInput[67]), .B(
        SubBytesInput[65]), .Z(SubBytesIns_Inst_Sbox_8_T5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_T6_U1 ( .A(SubBytesIns_Inst_Sbox_8_T1), 
        .B(SubBytesIns_Inst_Sbox_8_T5), .Z(SubBytesIns_Inst_Sbox_8_T6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_T7_U1 ( .A(SubBytesInput[70]), .B(
        SubBytesInput[69]), .Z(SubBytesIns_Inst_Sbox_8_T7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_T8_U1 ( .A(SubBytesInput[64]), .B(
        SubBytesIns_Inst_Sbox_8_T6), .Z(SubBytesIns_Inst_Sbox_8_T8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_T9_U1 ( .A(SubBytesInput[64]), .B(
        SubBytesIns_Inst_Sbox_8_T7), .Z(SubBytesIns_Inst_Sbox_8_T9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_T10_U1 ( .A(SubBytesIns_Inst_Sbox_8_T6), 
        .B(SubBytesIns_Inst_Sbox_8_T7), .Z(SubBytesIns_Inst_Sbox_8_T10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_T11_U1 ( .A(SubBytesInput[70]), .B(
        SubBytesInput[66]), .Z(SubBytesIns_Inst_Sbox_8_T11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_T12_U1 ( .A(SubBytesInput[69]), .B(
        SubBytesInput[66]), .Z(SubBytesIns_Inst_Sbox_8_T12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_T13_U1 ( .A(SubBytesIns_Inst_Sbox_8_T3), 
        .B(SubBytesIns_Inst_Sbox_8_T4), .Z(SubBytesIns_Inst_Sbox_8_T13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_T14_U1 ( .A(SubBytesIns_Inst_Sbox_8_T6), 
        .B(SubBytesIns_Inst_Sbox_8_T11), .Z(SubBytesIns_Inst_Sbox_8_T14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_T15_U1 ( .A(SubBytesIns_Inst_Sbox_8_T5), 
        .B(SubBytesIns_Inst_Sbox_8_T11), .Z(SubBytesIns_Inst_Sbox_8_T15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_T16_U1 ( .A(SubBytesIns_Inst_Sbox_8_T5), 
        .B(SubBytesIns_Inst_Sbox_8_T12), .Z(SubBytesIns_Inst_Sbox_8_T16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_T17_U1 ( .A(SubBytesIns_Inst_Sbox_8_T9), 
        .B(SubBytesIns_Inst_Sbox_8_T16), .Z(SubBytesIns_Inst_Sbox_8_T17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_T18_U1 ( .A(SubBytesInput[68]), .B(
        SubBytesInput[64]), .Z(SubBytesIns_Inst_Sbox_8_T18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_T19_U1 ( .A(SubBytesIns_Inst_Sbox_8_T7), 
        .B(SubBytesIns_Inst_Sbox_8_T18), .Z(SubBytesIns_Inst_Sbox_8_T19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_T20_U1 ( .A(SubBytesIns_Inst_Sbox_8_T1), 
        .B(SubBytesIns_Inst_Sbox_8_T19), .Z(SubBytesIns_Inst_Sbox_8_T20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_T21_U1 ( .A(SubBytesInput[65]), .B(
        SubBytesInput[64]), .Z(SubBytesIns_Inst_Sbox_8_T21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_T22_U1 ( .A(SubBytesIns_Inst_Sbox_8_T7), 
        .B(SubBytesIns_Inst_Sbox_8_T21), .Z(SubBytesIns_Inst_Sbox_8_T22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_T23_U1 ( .A(SubBytesIns_Inst_Sbox_8_T2), 
        .B(SubBytesIns_Inst_Sbox_8_T22), .Z(SubBytesIns_Inst_Sbox_8_T23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_T24_U1 ( .A(SubBytesIns_Inst_Sbox_8_T2), 
        .B(SubBytesIns_Inst_Sbox_8_T10), .Z(SubBytesIns_Inst_Sbox_8_T24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_T25_U1 ( .A(SubBytesIns_Inst_Sbox_8_T20), 
        .B(SubBytesIns_Inst_Sbox_8_T17), .Z(SubBytesIns_Inst_Sbox_8_T25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_T26_U1 ( .A(SubBytesIns_Inst_Sbox_8_T3), 
        .B(SubBytesIns_Inst_Sbox_8_T16), .Z(SubBytesIns_Inst_Sbox_8_T26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_T27_U1 ( .A(SubBytesIns_Inst_Sbox_8_T1), 
        .B(SubBytesIns_Inst_Sbox_8_T12), .Z(SubBytesIns_Inst_Sbox_8_T27) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M1_U1 ( .A1(SubBytesIns_Inst_Sbox_8_T13), 
        .A2(SubBytesIns_Inst_Sbox_8_T6), .ZN(SubBytesIns_Inst_Sbox_8_M1) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M2_U1 ( .A1(SubBytesIns_Inst_Sbox_8_T23), 
        .A2(SubBytesIns_Inst_Sbox_8_T8), .ZN(SubBytesIns_Inst_Sbox_8_M2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_M3_U1 ( .A(SubBytesIns_Inst_Sbox_8_T14), 
        .B(SubBytesIns_Inst_Sbox_8_M1), .Z(SubBytesIns_Inst_Sbox_8_M3) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M4_U1 ( .A1(SubBytesIns_Inst_Sbox_8_T19), 
        .A2(SubBytesInput[64]), .ZN(SubBytesIns_Inst_Sbox_8_M4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_M5_U1 ( .A(SubBytesIns_Inst_Sbox_8_M4), 
        .B(SubBytesIns_Inst_Sbox_8_M1), .Z(SubBytesIns_Inst_Sbox_8_M5) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M6_U1 ( .A1(SubBytesIns_Inst_Sbox_8_T3), 
        .A2(SubBytesIns_Inst_Sbox_8_T16), .ZN(SubBytesIns_Inst_Sbox_8_M6) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M7_U1 ( .A1(SubBytesIns_Inst_Sbox_8_T22), 
        .A2(SubBytesIns_Inst_Sbox_8_T9), .ZN(SubBytesIns_Inst_Sbox_8_M7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_M8_U1 ( .A(SubBytesIns_Inst_Sbox_8_T26), 
        .B(SubBytesIns_Inst_Sbox_8_M6), .Z(SubBytesIns_Inst_Sbox_8_M8) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M9_U1 ( .A1(SubBytesIns_Inst_Sbox_8_T20), 
        .A2(SubBytesIns_Inst_Sbox_8_T17), .ZN(SubBytesIns_Inst_Sbox_8_M9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_M10_U1 ( .A(SubBytesIns_Inst_Sbox_8_M9), 
        .B(SubBytesIns_Inst_Sbox_8_M6), .Z(SubBytesIns_Inst_Sbox_8_M10) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M11_U1 ( .A1(SubBytesIns_Inst_Sbox_8_T1), 
        .A2(SubBytesIns_Inst_Sbox_8_T15), .ZN(SubBytesIns_Inst_Sbox_8_M11) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M12_U1 ( .A1(SubBytesIns_Inst_Sbox_8_T4), 
        .A2(SubBytesIns_Inst_Sbox_8_T27), .ZN(SubBytesIns_Inst_Sbox_8_M12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_M13_U1 ( .A(SubBytesIns_Inst_Sbox_8_M12), 
        .B(SubBytesIns_Inst_Sbox_8_M11), .Z(SubBytesIns_Inst_Sbox_8_M13) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M14_U1 ( .A1(SubBytesIns_Inst_Sbox_8_T2), 
        .A2(SubBytesIns_Inst_Sbox_8_T10), .ZN(SubBytesIns_Inst_Sbox_8_M14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_M15_U1 ( .A(SubBytesIns_Inst_Sbox_8_M14), 
        .B(SubBytesIns_Inst_Sbox_8_M11), .Z(SubBytesIns_Inst_Sbox_8_M15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_M16_U1 ( .A(SubBytesIns_Inst_Sbox_8_M3), 
        .B(SubBytesIns_Inst_Sbox_8_M2), .Z(SubBytesIns_Inst_Sbox_8_M16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_M17_U1 ( .A(SubBytesIns_Inst_Sbox_8_M5), 
        .B(SubBytesIns_Inst_Sbox_8_T24), .Z(SubBytesIns_Inst_Sbox_8_M17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_M18_U1 ( .A(SubBytesIns_Inst_Sbox_8_M8), 
        .B(SubBytesIns_Inst_Sbox_8_M7), .Z(SubBytesIns_Inst_Sbox_8_M18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_M19_U1 ( .A(SubBytesIns_Inst_Sbox_8_M10), 
        .B(SubBytesIns_Inst_Sbox_8_M15), .Z(SubBytesIns_Inst_Sbox_8_M19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_M20_U1 ( .A(SubBytesIns_Inst_Sbox_8_M16), 
        .B(SubBytesIns_Inst_Sbox_8_M13), .Z(SubBytesIns_Inst_Sbox_8_M20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_M21_U1 ( .A(SubBytesIns_Inst_Sbox_8_M17), 
        .B(SubBytesIns_Inst_Sbox_8_M15), .Z(SubBytesIns_Inst_Sbox_8_M21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_M22_U1 ( .A(SubBytesIns_Inst_Sbox_8_M18), 
        .B(SubBytesIns_Inst_Sbox_8_M13), .Z(SubBytesIns_Inst_Sbox_8_M22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_M23_U1 ( .A(SubBytesIns_Inst_Sbox_8_M19), 
        .B(SubBytesIns_Inst_Sbox_8_T25), .Z(SubBytesIns_Inst_Sbox_8_M23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_M24_U1 ( .A(SubBytesIns_Inst_Sbox_8_M22), 
        .B(SubBytesIns_Inst_Sbox_8_M23), .Z(SubBytesIns_Inst_Sbox_8_M24) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M25_U1 ( .A1(SubBytesIns_Inst_Sbox_8_M22), .A2(SubBytesIns_Inst_Sbox_8_M20), .ZN(SubBytesIns_Inst_Sbox_8_M25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_M26_U1 ( .A(SubBytesIns_Inst_Sbox_8_M21), 
        .B(SubBytesIns_Inst_Sbox_8_M25), .Z(SubBytesIns_Inst_Sbox_8_M26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_M27_U1 ( .A(SubBytesIns_Inst_Sbox_8_M20), 
        .B(SubBytesIns_Inst_Sbox_8_M21), .Z(SubBytesIns_Inst_Sbox_8_M27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_M28_U1 ( .A(SubBytesIns_Inst_Sbox_8_M23), 
        .B(SubBytesIns_Inst_Sbox_8_M25), .Z(SubBytesIns_Inst_Sbox_8_M28) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M29_U1 ( .A1(SubBytesIns_Inst_Sbox_8_M28), .A2(SubBytesIns_Inst_Sbox_8_M27), .ZN(SubBytesIns_Inst_Sbox_8_M29) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M30_U1 ( .A1(SubBytesIns_Inst_Sbox_8_M26), .A2(SubBytesIns_Inst_Sbox_8_M24), .ZN(SubBytesIns_Inst_Sbox_8_M30) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M31_U1 ( .A1(SubBytesIns_Inst_Sbox_8_M20), .A2(SubBytesIns_Inst_Sbox_8_M23), .ZN(SubBytesIns_Inst_Sbox_8_M31) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M32_U1 ( .A1(SubBytesIns_Inst_Sbox_8_M27), .A2(SubBytesIns_Inst_Sbox_8_M31), .ZN(SubBytesIns_Inst_Sbox_8_M32) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_M33_U1 ( .A(SubBytesIns_Inst_Sbox_8_M27), 
        .B(SubBytesIns_Inst_Sbox_8_M25), .Z(SubBytesIns_Inst_Sbox_8_M33) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M34_U1 ( .A1(SubBytesIns_Inst_Sbox_8_M21), .A2(SubBytesIns_Inst_Sbox_8_M22), .ZN(SubBytesIns_Inst_Sbox_8_M34) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M35_U1 ( .A1(SubBytesIns_Inst_Sbox_8_M24), .A2(SubBytesIns_Inst_Sbox_8_M34), .ZN(SubBytesIns_Inst_Sbox_8_M35) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_M36_U1 ( .A(SubBytesIns_Inst_Sbox_8_M24), 
        .B(SubBytesIns_Inst_Sbox_8_M25), .Z(SubBytesIns_Inst_Sbox_8_M36) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_M37_U1 ( .A(SubBytesIns_Inst_Sbox_8_M21), 
        .B(SubBytesIns_Inst_Sbox_8_M29), .Z(SubBytesIns_Inst_Sbox_8_M37) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_M38_U1 ( .A(SubBytesIns_Inst_Sbox_8_M32), 
        .B(SubBytesIns_Inst_Sbox_8_M33), .Z(SubBytesIns_Inst_Sbox_8_M38) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_M39_U1 ( .A(SubBytesIns_Inst_Sbox_8_M23), 
        .B(SubBytesIns_Inst_Sbox_8_M30), .Z(SubBytesIns_Inst_Sbox_8_M39) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_M40_U1 ( .A(SubBytesIns_Inst_Sbox_8_M35), 
        .B(SubBytesIns_Inst_Sbox_8_M36), .Z(SubBytesIns_Inst_Sbox_8_M40) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_M41_U1 ( .A(SubBytesIns_Inst_Sbox_8_M38), 
        .B(SubBytesIns_Inst_Sbox_8_M40), .Z(SubBytesIns_Inst_Sbox_8_M41) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_M42_U1 ( .A(SubBytesIns_Inst_Sbox_8_M37), 
        .B(SubBytesIns_Inst_Sbox_8_M39), .Z(SubBytesIns_Inst_Sbox_8_M42) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_M43_U1 ( .A(SubBytesIns_Inst_Sbox_8_M37), 
        .B(SubBytesIns_Inst_Sbox_8_M38), .Z(SubBytesIns_Inst_Sbox_8_M43) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_M44_U1 ( .A(SubBytesIns_Inst_Sbox_8_M39), 
        .B(SubBytesIns_Inst_Sbox_8_M40), .Z(SubBytesIns_Inst_Sbox_8_M44) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_M45_U1 ( .A(SubBytesIns_Inst_Sbox_8_M42), 
        .B(SubBytesIns_Inst_Sbox_8_M41), .Z(SubBytesIns_Inst_Sbox_8_M45) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M46_U1 ( .A1(SubBytesIns_Inst_Sbox_8_M44), .A2(SubBytesIns_Inst_Sbox_8_T6), .ZN(SubBytesIns_Inst_Sbox_8_M46) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M47_U1 ( .A1(SubBytesIns_Inst_Sbox_8_M40), .A2(SubBytesIns_Inst_Sbox_8_T8), .ZN(SubBytesIns_Inst_Sbox_8_M47) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M48_U1 ( .A1(SubBytesIns_Inst_Sbox_8_M39), .A2(SubBytesInput[64]), .ZN(SubBytesIns_Inst_Sbox_8_M48) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M49_U1 ( .A1(SubBytesIns_Inst_Sbox_8_M43), .A2(SubBytesIns_Inst_Sbox_8_T16), .ZN(SubBytesIns_Inst_Sbox_8_M49) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M50_U1 ( .A1(SubBytesIns_Inst_Sbox_8_M38), .A2(SubBytesIns_Inst_Sbox_8_T9), .ZN(SubBytesIns_Inst_Sbox_8_M50) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M51_U1 ( .A1(SubBytesIns_Inst_Sbox_8_M37), .A2(SubBytesIns_Inst_Sbox_8_T17), .ZN(SubBytesIns_Inst_Sbox_8_M51) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M52_U1 ( .A1(SubBytesIns_Inst_Sbox_8_M42), .A2(SubBytesIns_Inst_Sbox_8_T15), .ZN(SubBytesIns_Inst_Sbox_8_M52) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M53_U1 ( .A1(SubBytesIns_Inst_Sbox_8_M45), .A2(SubBytesIns_Inst_Sbox_8_T27), .ZN(SubBytesIns_Inst_Sbox_8_M53) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M54_U1 ( .A1(SubBytesIns_Inst_Sbox_8_M41), .A2(SubBytesIns_Inst_Sbox_8_T10), .ZN(SubBytesIns_Inst_Sbox_8_M54) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M55_U1 ( .A1(SubBytesIns_Inst_Sbox_8_M44), .A2(SubBytesIns_Inst_Sbox_8_T13), .ZN(SubBytesIns_Inst_Sbox_8_M55) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M56_U1 ( .A1(SubBytesIns_Inst_Sbox_8_M40), .A2(SubBytesIns_Inst_Sbox_8_T23), .ZN(SubBytesIns_Inst_Sbox_8_M56) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M57_U1 ( .A1(SubBytesIns_Inst_Sbox_8_M39), .A2(SubBytesIns_Inst_Sbox_8_T19), .ZN(SubBytesIns_Inst_Sbox_8_M57) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M58_U1 ( .A1(SubBytesIns_Inst_Sbox_8_M43), .A2(SubBytesIns_Inst_Sbox_8_T3), .ZN(SubBytesIns_Inst_Sbox_8_M58) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M59_U1 ( .A1(SubBytesIns_Inst_Sbox_8_M38), .A2(SubBytesIns_Inst_Sbox_8_T22), .ZN(SubBytesIns_Inst_Sbox_8_M59) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M60_U1 ( .A1(SubBytesIns_Inst_Sbox_8_M37), .A2(SubBytesIns_Inst_Sbox_8_T20), .ZN(SubBytesIns_Inst_Sbox_8_M60) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M61_U1 ( .A1(SubBytesIns_Inst_Sbox_8_M42), .A2(SubBytesIns_Inst_Sbox_8_T1), .ZN(SubBytesIns_Inst_Sbox_8_M61) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M62_U1 ( .A1(SubBytesIns_Inst_Sbox_8_M45), .A2(SubBytesIns_Inst_Sbox_8_T4), .ZN(SubBytesIns_Inst_Sbox_8_M62) );
  AND2_X1 SubBytesIns_Inst_Sbox_8_AND_M63_U1 ( .A1(SubBytesIns_Inst_Sbox_8_M41), .A2(SubBytesIns_Inst_Sbox_8_T2), .ZN(SubBytesIns_Inst_Sbox_8_M63) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_L0_U1 ( .A(SubBytesIns_Inst_Sbox_8_M61), 
        .B(SubBytesIns_Inst_Sbox_8_M62), .Z(SubBytesIns_Inst_Sbox_8_L0) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_L1_U1 ( .A(SubBytesIns_Inst_Sbox_8_M50), 
        .B(SubBytesIns_Inst_Sbox_8_M56), .Z(SubBytesIns_Inst_Sbox_8_L1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_L2_U1 ( .A(SubBytesIns_Inst_Sbox_8_M46), 
        .B(SubBytesIns_Inst_Sbox_8_M48), .Z(SubBytesIns_Inst_Sbox_8_L2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_L3_U1 ( .A(SubBytesIns_Inst_Sbox_8_M47), 
        .B(SubBytesIns_Inst_Sbox_8_M55), .Z(SubBytesIns_Inst_Sbox_8_L3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_L4_U1 ( .A(SubBytesIns_Inst_Sbox_8_M54), 
        .B(SubBytesIns_Inst_Sbox_8_M58), .Z(SubBytesIns_Inst_Sbox_8_L4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_L5_U1 ( .A(SubBytesIns_Inst_Sbox_8_M49), 
        .B(SubBytesIns_Inst_Sbox_8_M61), .Z(SubBytesIns_Inst_Sbox_8_L5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_L6_U1 ( .A(SubBytesIns_Inst_Sbox_8_M62), 
        .B(SubBytesIns_Inst_Sbox_8_L5), .Z(SubBytesIns_Inst_Sbox_8_L6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_L7_U1 ( .A(SubBytesIns_Inst_Sbox_8_M46), 
        .B(SubBytesIns_Inst_Sbox_8_L3), .Z(SubBytesIns_Inst_Sbox_8_L7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_L8_U1 ( .A(SubBytesIns_Inst_Sbox_8_M51), 
        .B(SubBytesIns_Inst_Sbox_8_M59), .Z(SubBytesIns_Inst_Sbox_8_L8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_L9_U1 ( .A(SubBytesIns_Inst_Sbox_8_M52), 
        .B(SubBytesIns_Inst_Sbox_8_M53), .Z(SubBytesIns_Inst_Sbox_8_L9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_L10_U1 ( .A(SubBytesIns_Inst_Sbox_8_M53), 
        .B(SubBytesIns_Inst_Sbox_8_L4), .Z(SubBytesIns_Inst_Sbox_8_L10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_L11_U1 ( .A(SubBytesIns_Inst_Sbox_8_M60), 
        .B(SubBytesIns_Inst_Sbox_8_L2), .Z(SubBytesIns_Inst_Sbox_8_L11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_L12_U1 ( .A(SubBytesIns_Inst_Sbox_8_M48), 
        .B(SubBytesIns_Inst_Sbox_8_M51), .Z(SubBytesIns_Inst_Sbox_8_L12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_L13_U1 ( .A(SubBytesIns_Inst_Sbox_8_M50), 
        .B(SubBytesIns_Inst_Sbox_8_L0), .Z(SubBytesIns_Inst_Sbox_8_L13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_L14_U1 ( .A(SubBytesIns_Inst_Sbox_8_M52), 
        .B(SubBytesIns_Inst_Sbox_8_M61), .Z(SubBytesIns_Inst_Sbox_8_L14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_L15_U1 ( .A(SubBytesIns_Inst_Sbox_8_M55), 
        .B(SubBytesIns_Inst_Sbox_8_L1), .Z(SubBytesIns_Inst_Sbox_8_L15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_L16_U1 ( .A(SubBytesIns_Inst_Sbox_8_M56), 
        .B(SubBytesIns_Inst_Sbox_8_L0), .Z(SubBytesIns_Inst_Sbox_8_L16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_L17_U1 ( .A(SubBytesIns_Inst_Sbox_8_M57), 
        .B(SubBytesIns_Inst_Sbox_8_L1), .Z(SubBytesIns_Inst_Sbox_8_L17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_L18_U1 ( .A(SubBytesIns_Inst_Sbox_8_M58), 
        .B(SubBytesIns_Inst_Sbox_8_L8), .Z(SubBytesIns_Inst_Sbox_8_L18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_L19_U1 ( .A(SubBytesIns_Inst_Sbox_8_M63), 
        .B(SubBytesIns_Inst_Sbox_8_L4), .Z(SubBytesIns_Inst_Sbox_8_L19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_L20_U1 ( .A(SubBytesIns_Inst_Sbox_8_L0), 
        .B(SubBytesIns_Inst_Sbox_8_L1), .Z(SubBytesIns_Inst_Sbox_8_L20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_L21_U1 ( .A(SubBytesIns_Inst_Sbox_8_L1), 
        .B(SubBytesIns_Inst_Sbox_8_L7), .Z(SubBytesIns_Inst_Sbox_8_L21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_L22_U1 ( .A(SubBytesIns_Inst_Sbox_8_L3), 
        .B(SubBytesIns_Inst_Sbox_8_L12), .Z(SubBytesIns_Inst_Sbox_8_L22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_L23_U1 ( .A(SubBytesIns_Inst_Sbox_8_L18), 
        .B(SubBytesIns_Inst_Sbox_8_L2), .Z(SubBytesIns_Inst_Sbox_8_L23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_L24_U1 ( .A(SubBytesIns_Inst_Sbox_8_L15), 
        .B(SubBytesIns_Inst_Sbox_8_L9), .Z(SubBytesIns_Inst_Sbox_8_L24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_L25_U1 ( .A(SubBytesIns_Inst_Sbox_8_L6), 
        .B(SubBytesIns_Inst_Sbox_8_L10), .Z(SubBytesIns_Inst_Sbox_8_L25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_L26_U1 ( .A(SubBytesIns_Inst_Sbox_8_L7), 
        .B(SubBytesIns_Inst_Sbox_8_L9), .Z(SubBytesIns_Inst_Sbox_8_L26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_L27_U1 ( .A(SubBytesIns_Inst_Sbox_8_L8), 
        .B(SubBytesIns_Inst_Sbox_8_L10), .Z(SubBytesIns_Inst_Sbox_8_L27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_L28_U1 ( .A(SubBytesIns_Inst_Sbox_8_L11), 
        .B(SubBytesIns_Inst_Sbox_8_L14), .Z(SubBytesIns_Inst_Sbox_8_L28) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_L29_U1 ( .A(SubBytesIns_Inst_Sbox_8_L11), 
        .B(SubBytesIns_Inst_Sbox_8_L17), .Z(SubBytesIns_Inst_Sbox_8_L29) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_S0_U1 ( .A(SubBytesIns_Inst_Sbox_8_L6), 
        .B(SubBytesIns_Inst_Sbox_8_L24), .Z(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_S1_U1 ( .A(SubBytesIns_Inst_Sbox_8_L16), 
        .B(SubBytesIns_Inst_Sbox_8_L26), .ZN(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[7]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_S2_U1 ( .A(SubBytesIns_Inst_Sbox_8_L19), 
        .B(SubBytesIns_Inst_Sbox_8_L28), .ZN(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[6]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_S3_U1 ( .A(SubBytesIns_Inst_Sbox_8_L6), 
        .B(SubBytesIns_Inst_Sbox_8_L21), .Z(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[5]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_S4_U1 ( .A(SubBytesIns_Inst_Sbox_8_L20), 
        .B(SubBytesIns_Inst_Sbox_8_L22), .Z(MixColumnsInput[35]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_S5_U1 ( .A(SubBytesIns_Inst_Sbox_8_L25), 
        .B(SubBytesIns_Inst_Sbox_8_L29), .Z(MixColumnsInput[34]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_S6_U1 ( .A(SubBytesIns_Inst_Sbox_8_L13), 
        .B(SubBytesIns_Inst_Sbox_8_L27), .ZN(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[2]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_8_XOR_S7_U1 ( .A(SubBytesIns_Inst_Sbox_8_L6), 
        .B(SubBytesIns_Inst_Sbox_8_L23), .ZN(MixColumnsInput[32]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_T1_U1 ( .A(SubBytesInput[79]), .B(
        SubBytesInput[76]), .Z(SubBytesIns_Inst_Sbox_9_T1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_T2_U1 ( .A(SubBytesInput[79]), .B(
        SubBytesInput[74]), .Z(SubBytesIns_Inst_Sbox_9_T2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_T3_U1 ( .A(SubBytesInput[79]), .B(
        SubBytesInput[73]), .Z(SubBytesIns_Inst_Sbox_9_T3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_T4_U1 ( .A(SubBytesInput[76]), .B(
        SubBytesInput[74]), .Z(SubBytesIns_Inst_Sbox_9_T4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_T5_U1 ( .A(SubBytesInput[75]), .B(
        SubBytesInput[73]), .Z(SubBytesIns_Inst_Sbox_9_T5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_T6_U1 ( .A(SubBytesIns_Inst_Sbox_9_T1), 
        .B(SubBytesIns_Inst_Sbox_9_T5), .Z(SubBytesIns_Inst_Sbox_9_T6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_T7_U1 ( .A(SubBytesInput[78]), .B(
        SubBytesInput[77]), .Z(SubBytesIns_Inst_Sbox_9_T7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_T8_U1 ( .A(SubBytesInput[72]), .B(
        SubBytesIns_Inst_Sbox_9_T6), .Z(SubBytesIns_Inst_Sbox_9_T8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_T9_U1 ( .A(SubBytesInput[72]), .B(
        SubBytesIns_Inst_Sbox_9_T7), .Z(SubBytesIns_Inst_Sbox_9_T9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_T10_U1 ( .A(SubBytesIns_Inst_Sbox_9_T6), 
        .B(SubBytesIns_Inst_Sbox_9_T7), .Z(SubBytesIns_Inst_Sbox_9_T10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_T11_U1 ( .A(SubBytesInput[78]), .B(
        SubBytesInput[74]), .Z(SubBytesIns_Inst_Sbox_9_T11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_T12_U1 ( .A(SubBytesInput[77]), .B(
        SubBytesInput[74]), .Z(SubBytesIns_Inst_Sbox_9_T12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_T13_U1 ( .A(SubBytesIns_Inst_Sbox_9_T3), 
        .B(SubBytesIns_Inst_Sbox_9_T4), .Z(SubBytesIns_Inst_Sbox_9_T13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_T14_U1 ( .A(SubBytesIns_Inst_Sbox_9_T6), 
        .B(SubBytesIns_Inst_Sbox_9_T11), .Z(SubBytesIns_Inst_Sbox_9_T14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_T15_U1 ( .A(SubBytesIns_Inst_Sbox_9_T5), 
        .B(SubBytesIns_Inst_Sbox_9_T11), .Z(SubBytesIns_Inst_Sbox_9_T15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_T16_U1 ( .A(SubBytesIns_Inst_Sbox_9_T5), 
        .B(SubBytesIns_Inst_Sbox_9_T12), .Z(SubBytesIns_Inst_Sbox_9_T16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_T17_U1 ( .A(SubBytesIns_Inst_Sbox_9_T9), 
        .B(SubBytesIns_Inst_Sbox_9_T16), .Z(SubBytesIns_Inst_Sbox_9_T17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_T18_U1 ( .A(SubBytesInput[76]), .B(
        SubBytesInput[72]), .Z(SubBytesIns_Inst_Sbox_9_T18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_T19_U1 ( .A(SubBytesIns_Inst_Sbox_9_T7), 
        .B(SubBytesIns_Inst_Sbox_9_T18), .Z(SubBytesIns_Inst_Sbox_9_T19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_T20_U1 ( .A(SubBytesIns_Inst_Sbox_9_T1), 
        .B(SubBytesIns_Inst_Sbox_9_T19), .Z(SubBytesIns_Inst_Sbox_9_T20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_T21_U1 ( .A(SubBytesInput[73]), .B(
        SubBytesInput[72]), .Z(SubBytesIns_Inst_Sbox_9_T21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_T22_U1 ( .A(SubBytesIns_Inst_Sbox_9_T7), 
        .B(SubBytesIns_Inst_Sbox_9_T21), .Z(SubBytesIns_Inst_Sbox_9_T22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_T23_U1 ( .A(SubBytesIns_Inst_Sbox_9_T2), 
        .B(SubBytesIns_Inst_Sbox_9_T22), .Z(SubBytesIns_Inst_Sbox_9_T23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_T24_U1 ( .A(SubBytesIns_Inst_Sbox_9_T2), 
        .B(SubBytesIns_Inst_Sbox_9_T10), .Z(SubBytesIns_Inst_Sbox_9_T24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_T25_U1 ( .A(SubBytesIns_Inst_Sbox_9_T20), 
        .B(SubBytesIns_Inst_Sbox_9_T17), .Z(SubBytesIns_Inst_Sbox_9_T25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_T26_U1 ( .A(SubBytesIns_Inst_Sbox_9_T3), 
        .B(SubBytesIns_Inst_Sbox_9_T16), .Z(SubBytesIns_Inst_Sbox_9_T26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_T27_U1 ( .A(SubBytesIns_Inst_Sbox_9_T1), 
        .B(SubBytesIns_Inst_Sbox_9_T12), .Z(SubBytesIns_Inst_Sbox_9_T27) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M1_U1 ( .A1(SubBytesIns_Inst_Sbox_9_T13), 
        .A2(SubBytesIns_Inst_Sbox_9_T6), .ZN(SubBytesIns_Inst_Sbox_9_M1) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M2_U1 ( .A1(SubBytesIns_Inst_Sbox_9_T23), 
        .A2(SubBytesIns_Inst_Sbox_9_T8), .ZN(SubBytesIns_Inst_Sbox_9_M2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_M3_U1 ( .A(SubBytesIns_Inst_Sbox_9_T14), 
        .B(SubBytesIns_Inst_Sbox_9_M1), .Z(SubBytesIns_Inst_Sbox_9_M3) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M4_U1 ( .A1(SubBytesIns_Inst_Sbox_9_T19), 
        .A2(SubBytesInput[72]), .ZN(SubBytesIns_Inst_Sbox_9_M4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_M5_U1 ( .A(SubBytesIns_Inst_Sbox_9_M4), 
        .B(SubBytesIns_Inst_Sbox_9_M1), .Z(SubBytesIns_Inst_Sbox_9_M5) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M6_U1 ( .A1(SubBytesIns_Inst_Sbox_9_T3), 
        .A2(SubBytesIns_Inst_Sbox_9_T16), .ZN(SubBytesIns_Inst_Sbox_9_M6) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M7_U1 ( .A1(SubBytesIns_Inst_Sbox_9_T22), 
        .A2(SubBytesIns_Inst_Sbox_9_T9), .ZN(SubBytesIns_Inst_Sbox_9_M7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_M8_U1 ( .A(SubBytesIns_Inst_Sbox_9_T26), 
        .B(SubBytesIns_Inst_Sbox_9_M6), .Z(SubBytesIns_Inst_Sbox_9_M8) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M9_U1 ( .A1(SubBytesIns_Inst_Sbox_9_T20), 
        .A2(SubBytesIns_Inst_Sbox_9_T17), .ZN(SubBytesIns_Inst_Sbox_9_M9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_M10_U1 ( .A(SubBytesIns_Inst_Sbox_9_M9), 
        .B(SubBytesIns_Inst_Sbox_9_M6), .Z(SubBytesIns_Inst_Sbox_9_M10) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M11_U1 ( .A1(SubBytesIns_Inst_Sbox_9_T1), 
        .A2(SubBytesIns_Inst_Sbox_9_T15), .ZN(SubBytesIns_Inst_Sbox_9_M11) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M12_U1 ( .A1(SubBytesIns_Inst_Sbox_9_T4), 
        .A2(SubBytesIns_Inst_Sbox_9_T27), .ZN(SubBytesIns_Inst_Sbox_9_M12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_M13_U1 ( .A(SubBytesIns_Inst_Sbox_9_M12), 
        .B(SubBytesIns_Inst_Sbox_9_M11), .Z(SubBytesIns_Inst_Sbox_9_M13) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M14_U1 ( .A1(SubBytesIns_Inst_Sbox_9_T2), 
        .A2(SubBytesIns_Inst_Sbox_9_T10), .ZN(SubBytesIns_Inst_Sbox_9_M14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_M15_U1 ( .A(SubBytesIns_Inst_Sbox_9_M14), 
        .B(SubBytesIns_Inst_Sbox_9_M11), .Z(SubBytesIns_Inst_Sbox_9_M15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_M16_U1 ( .A(SubBytesIns_Inst_Sbox_9_M3), 
        .B(SubBytesIns_Inst_Sbox_9_M2), .Z(SubBytesIns_Inst_Sbox_9_M16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_M17_U1 ( .A(SubBytesIns_Inst_Sbox_9_M5), 
        .B(SubBytesIns_Inst_Sbox_9_T24), .Z(SubBytesIns_Inst_Sbox_9_M17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_M18_U1 ( .A(SubBytesIns_Inst_Sbox_9_M8), 
        .B(SubBytesIns_Inst_Sbox_9_M7), .Z(SubBytesIns_Inst_Sbox_9_M18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_M19_U1 ( .A(SubBytesIns_Inst_Sbox_9_M10), 
        .B(SubBytesIns_Inst_Sbox_9_M15), .Z(SubBytesIns_Inst_Sbox_9_M19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_M20_U1 ( .A(SubBytesIns_Inst_Sbox_9_M16), 
        .B(SubBytesIns_Inst_Sbox_9_M13), .Z(SubBytesIns_Inst_Sbox_9_M20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_M21_U1 ( .A(SubBytesIns_Inst_Sbox_9_M17), 
        .B(SubBytesIns_Inst_Sbox_9_M15), .Z(SubBytesIns_Inst_Sbox_9_M21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_M22_U1 ( .A(SubBytesIns_Inst_Sbox_9_M18), 
        .B(SubBytesIns_Inst_Sbox_9_M13), .Z(SubBytesIns_Inst_Sbox_9_M22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_M23_U1 ( .A(SubBytesIns_Inst_Sbox_9_M19), 
        .B(SubBytesIns_Inst_Sbox_9_T25), .Z(SubBytesIns_Inst_Sbox_9_M23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_M24_U1 ( .A(SubBytesIns_Inst_Sbox_9_M22), 
        .B(SubBytesIns_Inst_Sbox_9_M23), .Z(SubBytesIns_Inst_Sbox_9_M24) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M25_U1 ( .A1(SubBytesIns_Inst_Sbox_9_M22), .A2(SubBytesIns_Inst_Sbox_9_M20), .ZN(SubBytesIns_Inst_Sbox_9_M25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_M26_U1 ( .A(SubBytesIns_Inst_Sbox_9_M21), 
        .B(SubBytesIns_Inst_Sbox_9_M25), .Z(SubBytesIns_Inst_Sbox_9_M26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_M27_U1 ( .A(SubBytesIns_Inst_Sbox_9_M20), 
        .B(SubBytesIns_Inst_Sbox_9_M21), .Z(SubBytesIns_Inst_Sbox_9_M27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_M28_U1 ( .A(SubBytesIns_Inst_Sbox_9_M23), 
        .B(SubBytesIns_Inst_Sbox_9_M25), .Z(SubBytesIns_Inst_Sbox_9_M28) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M29_U1 ( .A1(SubBytesIns_Inst_Sbox_9_M28), .A2(SubBytesIns_Inst_Sbox_9_M27), .ZN(SubBytesIns_Inst_Sbox_9_M29) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M30_U1 ( .A1(SubBytesIns_Inst_Sbox_9_M26), .A2(SubBytesIns_Inst_Sbox_9_M24), .ZN(SubBytesIns_Inst_Sbox_9_M30) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M31_U1 ( .A1(SubBytesIns_Inst_Sbox_9_M20), .A2(SubBytesIns_Inst_Sbox_9_M23), .ZN(SubBytesIns_Inst_Sbox_9_M31) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M32_U1 ( .A1(SubBytesIns_Inst_Sbox_9_M27), .A2(SubBytesIns_Inst_Sbox_9_M31), .ZN(SubBytesIns_Inst_Sbox_9_M32) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_M33_U1 ( .A(SubBytesIns_Inst_Sbox_9_M27), 
        .B(SubBytesIns_Inst_Sbox_9_M25), .Z(SubBytesIns_Inst_Sbox_9_M33) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M34_U1 ( .A1(SubBytesIns_Inst_Sbox_9_M21), .A2(SubBytesIns_Inst_Sbox_9_M22), .ZN(SubBytesIns_Inst_Sbox_9_M34) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M35_U1 ( .A1(SubBytesIns_Inst_Sbox_9_M24), .A2(SubBytesIns_Inst_Sbox_9_M34), .ZN(SubBytesIns_Inst_Sbox_9_M35) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_M36_U1 ( .A(SubBytesIns_Inst_Sbox_9_M24), 
        .B(SubBytesIns_Inst_Sbox_9_M25), .Z(SubBytesIns_Inst_Sbox_9_M36) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_M37_U1 ( .A(SubBytesIns_Inst_Sbox_9_M21), 
        .B(SubBytesIns_Inst_Sbox_9_M29), .Z(SubBytesIns_Inst_Sbox_9_M37) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_M38_U1 ( .A(SubBytesIns_Inst_Sbox_9_M32), 
        .B(SubBytesIns_Inst_Sbox_9_M33), .Z(SubBytesIns_Inst_Sbox_9_M38) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_M39_U1 ( .A(SubBytesIns_Inst_Sbox_9_M23), 
        .B(SubBytesIns_Inst_Sbox_9_M30), .Z(SubBytesIns_Inst_Sbox_9_M39) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_M40_U1 ( .A(SubBytesIns_Inst_Sbox_9_M35), 
        .B(SubBytesIns_Inst_Sbox_9_M36), .Z(SubBytesIns_Inst_Sbox_9_M40) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_M41_U1 ( .A(SubBytesIns_Inst_Sbox_9_M38), 
        .B(SubBytesIns_Inst_Sbox_9_M40), .Z(SubBytesIns_Inst_Sbox_9_M41) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_M42_U1 ( .A(SubBytesIns_Inst_Sbox_9_M37), 
        .B(SubBytesIns_Inst_Sbox_9_M39), .Z(SubBytesIns_Inst_Sbox_9_M42) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_M43_U1 ( .A(SubBytesIns_Inst_Sbox_9_M37), 
        .B(SubBytesIns_Inst_Sbox_9_M38), .Z(SubBytesIns_Inst_Sbox_9_M43) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_M44_U1 ( .A(SubBytesIns_Inst_Sbox_9_M39), 
        .B(SubBytesIns_Inst_Sbox_9_M40), .Z(SubBytesIns_Inst_Sbox_9_M44) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_M45_U1 ( .A(SubBytesIns_Inst_Sbox_9_M42), 
        .B(SubBytesIns_Inst_Sbox_9_M41), .Z(SubBytesIns_Inst_Sbox_9_M45) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M46_U1 ( .A1(SubBytesIns_Inst_Sbox_9_M44), .A2(SubBytesIns_Inst_Sbox_9_T6), .ZN(SubBytesIns_Inst_Sbox_9_M46) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M47_U1 ( .A1(SubBytesIns_Inst_Sbox_9_M40), .A2(SubBytesIns_Inst_Sbox_9_T8), .ZN(SubBytesIns_Inst_Sbox_9_M47) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M48_U1 ( .A1(SubBytesIns_Inst_Sbox_9_M39), .A2(SubBytesInput[72]), .ZN(SubBytesIns_Inst_Sbox_9_M48) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M49_U1 ( .A1(SubBytesIns_Inst_Sbox_9_M43), .A2(SubBytesIns_Inst_Sbox_9_T16), .ZN(SubBytesIns_Inst_Sbox_9_M49) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M50_U1 ( .A1(SubBytesIns_Inst_Sbox_9_M38), .A2(SubBytesIns_Inst_Sbox_9_T9), .ZN(SubBytesIns_Inst_Sbox_9_M50) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M51_U1 ( .A1(SubBytesIns_Inst_Sbox_9_M37), .A2(SubBytesIns_Inst_Sbox_9_T17), .ZN(SubBytesIns_Inst_Sbox_9_M51) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M52_U1 ( .A1(SubBytesIns_Inst_Sbox_9_M42), .A2(SubBytesIns_Inst_Sbox_9_T15), .ZN(SubBytesIns_Inst_Sbox_9_M52) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M53_U1 ( .A1(SubBytesIns_Inst_Sbox_9_M45), .A2(SubBytesIns_Inst_Sbox_9_T27), .ZN(SubBytesIns_Inst_Sbox_9_M53) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M54_U1 ( .A1(SubBytesIns_Inst_Sbox_9_M41), .A2(SubBytesIns_Inst_Sbox_9_T10), .ZN(SubBytesIns_Inst_Sbox_9_M54) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M55_U1 ( .A1(SubBytesIns_Inst_Sbox_9_M44), .A2(SubBytesIns_Inst_Sbox_9_T13), .ZN(SubBytesIns_Inst_Sbox_9_M55) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M56_U1 ( .A1(SubBytesIns_Inst_Sbox_9_M40), .A2(SubBytesIns_Inst_Sbox_9_T23), .ZN(SubBytesIns_Inst_Sbox_9_M56) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M57_U1 ( .A1(SubBytesIns_Inst_Sbox_9_M39), .A2(SubBytesIns_Inst_Sbox_9_T19), .ZN(SubBytesIns_Inst_Sbox_9_M57) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M58_U1 ( .A1(SubBytesIns_Inst_Sbox_9_M43), .A2(SubBytesIns_Inst_Sbox_9_T3), .ZN(SubBytesIns_Inst_Sbox_9_M58) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M59_U1 ( .A1(SubBytesIns_Inst_Sbox_9_M38), .A2(SubBytesIns_Inst_Sbox_9_T22), .ZN(SubBytesIns_Inst_Sbox_9_M59) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M60_U1 ( .A1(SubBytesIns_Inst_Sbox_9_M37), .A2(SubBytesIns_Inst_Sbox_9_T20), .ZN(SubBytesIns_Inst_Sbox_9_M60) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M61_U1 ( .A1(SubBytesIns_Inst_Sbox_9_M42), .A2(SubBytesIns_Inst_Sbox_9_T1), .ZN(SubBytesIns_Inst_Sbox_9_M61) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M62_U1 ( .A1(SubBytesIns_Inst_Sbox_9_M45), .A2(SubBytesIns_Inst_Sbox_9_T4), .ZN(SubBytesIns_Inst_Sbox_9_M62) );
  AND2_X1 SubBytesIns_Inst_Sbox_9_AND_M63_U1 ( .A1(SubBytesIns_Inst_Sbox_9_M41), .A2(SubBytesIns_Inst_Sbox_9_T2), .ZN(SubBytesIns_Inst_Sbox_9_M63) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_L0_U1 ( .A(SubBytesIns_Inst_Sbox_9_M61), 
        .B(SubBytesIns_Inst_Sbox_9_M62), .Z(SubBytesIns_Inst_Sbox_9_L0) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_L1_U1 ( .A(SubBytesIns_Inst_Sbox_9_M50), 
        .B(SubBytesIns_Inst_Sbox_9_M56), .Z(SubBytesIns_Inst_Sbox_9_L1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_L2_U1 ( .A(SubBytesIns_Inst_Sbox_9_M46), 
        .B(SubBytesIns_Inst_Sbox_9_M48), .Z(SubBytesIns_Inst_Sbox_9_L2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_L3_U1 ( .A(SubBytesIns_Inst_Sbox_9_M47), 
        .B(SubBytesIns_Inst_Sbox_9_M55), .Z(SubBytesIns_Inst_Sbox_9_L3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_L4_U1 ( .A(SubBytesIns_Inst_Sbox_9_M54), 
        .B(SubBytesIns_Inst_Sbox_9_M58), .Z(SubBytesIns_Inst_Sbox_9_L4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_L5_U1 ( .A(SubBytesIns_Inst_Sbox_9_M49), 
        .B(SubBytesIns_Inst_Sbox_9_M61), .Z(SubBytesIns_Inst_Sbox_9_L5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_L6_U1 ( .A(SubBytesIns_Inst_Sbox_9_M62), 
        .B(SubBytesIns_Inst_Sbox_9_L5), .Z(SubBytesIns_Inst_Sbox_9_L6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_L7_U1 ( .A(SubBytesIns_Inst_Sbox_9_M46), 
        .B(SubBytesIns_Inst_Sbox_9_L3), .Z(SubBytesIns_Inst_Sbox_9_L7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_L8_U1 ( .A(SubBytesIns_Inst_Sbox_9_M51), 
        .B(SubBytesIns_Inst_Sbox_9_M59), .Z(SubBytesIns_Inst_Sbox_9_L8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_L9_U1 ( .A(SubBytesIns_Inst_Sbox_9_M52), 
        .B(SubBytesIns_Inst_Sbox_9_M53), .Z(SubBytesIns_Inst_Sbox_9_L9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_L10_U1 ( .A(SubBytesIns_Inst_Sbox_9_M53), 
        .B(SubBytesIns_Inst_Sbox_9_L4), .Z(SubBytesIns_Inst_Sbox_9_L10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_L11_U1 ( .A(SubBytesIns_Inst_Sbox_9_M60), 
        .B(SubBytesIns_Inst_Sbox_9_L2), .Z(SubBytesIns_Inst_Sbox_9_L11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_L12_U1 ( .A(SubBytesIns_Inst_Sbox_9_M48), 
        .B(SubBytesIns_Inst_Sbox_9_M51), .Z(SubBytesIns_Inst_Sbox_9_L12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_L13_U1 ( .A(SubBytesIns_Inst_Sbox_9_M50), 
        .B(SubBytesIns_Inst_Sbox_9_L0), .Z(SubBytesIns_Inst_Sbox_9_L13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_L14_U1 ( .A(SubBytesIns_Inst_Sbox_9_M52), 
        .B(SubBytesIns_Inst_Sbox_9_M61), .Z(SubBytesIns_Inst_Sbox_9_L14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_L15_U1 ( .A(SubBytesIns_Inst_Sbox_9_M55), 
        .B(SubBytesIns_Inst_Sbox_9_L1), .Z(SubBytesIns_Inst_Sbox_9_L15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_L16_U1 ( .A(SubBytesIns_Inst_Sbox_9_M56), 
        .B(SubBytesIns_Inst_Sbox_9_L0), .Z(SubBytesIns_Inst_Sbox_9_L16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_L17_U1 ( .A(SubBytesIns_Inst_Sbox_9_M57), 
        .B(SubBytesIns_Inst_Sbox_9_L1), .Z(SubBytesIns_Inst_Sbox_9_L17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_L18_U1 ( .A(SubBytesIns_Inst_Sbox_9_M58), 
        .B(SubBytesIns_Inst_Sbox_9_L8), .Z(SubBytesIns_Inst_Sbox_9_L18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_L19_U1 ( .A(SubBytesIns_Inst_Sbox_9_M63), 
        .B(SubBytesIns_Inst_Sbox_9_L4), .Z(SubBytesIns_Inst_Sbox_9_L19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_L20_U1 ( .A(SubBytesIns_Inst_Sbox_9_L0), 
        .B(SubBytesIns_Inst_Sbox_9_L1), .Z(SubBytesIns_Inst_Sbox_9_L20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_L21_U1 ( .A(SubBytesIns_Inst_Sbox_9_L1), 
        .B(SubBytesIns_Inst_Sbox_9_L7), .Z(SubBytesIns_Inst_Sbox_9_L21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_L22_U1 ( .A(SubBytesIns_Inst_Sbox_9_L3), 
        .B(SubBytesIns_Inst_Sbox_9_L12), .Z(SubBytesIns_Inst_Sbox_9_L22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_L23_U1 ( .A(SubBytesIns_Inst_Sbox_9_L18), 
        .B(SubBytesIns_Inst_Sbox_9_L2), .Z(SubBytesIns_Inst_Sbox_9_L23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_L24_U1 ( .A(SubBytesIns_Inst_Sbox_9_L15), 
        .B(SubBytesIns_Inst_Sbox_9_L9), .Z(SubBytesIns_Inst_Sbox_9_L24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_L25_U1 ( .A(SubBytesIns_Inst_Sbox_9_L6), 
        .B(SubBytesIns_Inst_Sbox_9_L10), .Z(SubBytesIns_Inst_Sbox_9_L25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_L26_U1 ( .A(SubBytesIns_Inst_Sbox_9_L7), 
        .B(SubBytesIns_Inst_Sbox_9_L9), .Z(SubBytesIns_Inst_Sbox_9_L26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_L27_U1 ( .A(SubBytesIns_Inst_Sbox_9_L8), 
        .B(SubBytesIns_Inst_Sbox_9_L10), .Z(SubBytesIns_Inst_Sbox_9_L27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_L28_U1 ( .A(SubBytesIns_Inst_Sbox_9_L11), 
        .B(SubBytesIns_Inst_Sbox_9_L14), .Z(SubBytesIns_Inst_Sbox_9_L28) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_L29_U1 ( .A(SubBytesIns_Inst_Sbox_9_L11), 
        .B(SubBytesIns_Inst_Sbox_9_L17), .Z(SubBytesIns_Inst_Sbox_9_L29) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_S0_U1 ( .A(SubBytesIns_Inst_Sbox_9_L6), 
        .B(SubBytesIns_Inst_Sbox_9_L24), .Z(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_S1_U1 ( .A(SubBytesIns_Inst_Sbox_9_L16), 
        .B(SubBytesIns_Inst_Sbox_9_L26), .ZN(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[15]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_S2_U1 ( .A(SubBytesIns_Inst_Sbox_9_L19), 
        .B(SubBytesIns_Inst_Sbox_9_L28), .ZN(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[14]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_S3_U1 ( .A(SubBytesIns_Inst_Sbox_9_L6), 
        .B(SubBytesIns_Inst_Sbox_9_L21), .Z(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[13]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_S4_U1 ( .A(SubBytesIns_Inst_Sbox_9_L20), 
        .B(SubBytesIns_Inst_Sbox_9_L22), .Z(MixColumnsInput[11]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_S5_U1 ( .A(SubBytesIns_Inst_Sbox_9_L25), 
        .B(SubBytesIns_Inst_Sbox_9_L29), .Z(MixColumnsInput[10]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_S6_U1 ( .A(SubBytesIns_Inst_Sbox_9_L13), 
        .B(SubBytesIns_Inst_Sbox_9_L27), .ZN(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[10]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_9_XOR_S7_U1 ( .A(SubBytesIns_Inst_Sbox_9_L6), 
        .B(SubBytesIns_Inst_Sbox_9_L23), .ZN(MixColumnsInput[8]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_T1_U1 ( .A(SubBytesInput[87]), .B(
        SubBytesInput[84]), .Z(SubBytesIns_Inst_Sbox_10_T1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_T2_U1 ( .A(SubBytesInput[87]), .B(
        SubBytesInput[82]), .Z(SubBytesIns_Inst_Sbox_10_T2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_T3_U1 ( .A(SubBytesInput[87]), .B(
        SubBytesInput[81]), .Z(SubBytesIns_Inst_Sbox_10_T3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_T4_U1 ( .A(SubBytesInput[84]), .B(
        SubBytesInput[82]), .Z(SubBytesIns_Inst_Sbox_10_T4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_T5_U1 ( .A(SubBytesInput[83]), .B(
        SubBytesInput[81]), .Z(SubBytesIns_Inst_Sbox_10_T5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_T6_U1 ( .A(SubBytesIns_Inst_Sbox_10_T1), 
        .B(SubBytesIns_Inst_Sbox_10_T5), .Z(SubBytesIns_Inst_Sbox_10_T6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_T7_U1 ( .A(SubBytesInput[86]), .B(
        SubBytesInput[85]), .Z(SubBytesIns_Inst_Sbox_10_T7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_T8_U1 ( .A(SubBytesInput[80]), .B(
        SubBytesIns_Inst_Sbox_10_T6), .Z(SubBytesIns_Inst_Sbox_10_T8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_T9_U1 ( .A(SubBytesInput[80]), .B(
        SubBytesIns_Inst_Sbox_10_T7), .Z(SubBytesIns_Inst_Sbox_10_T9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_T10_U1 ( .A(SubBytesIns_Inst_Sbox_10_T6), .B(SubBytesIns_Inst_Sbox_10_T7), .Z(SubBytesIns_Inst_Sbox_10_T10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_T11_U1 ( .A(SubBytesInput[86]), .B(
        SubBytesInput[82]), .Z(SubBytesIns_Inst_Sbox_10_T11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_T12_U1 ( .A(SubBytesInput[85]), .B(
        SubBytesInput[82]), .Z(SubBytesIns_Inst_Sbox_10_T12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_T13_U1 ( .A(SubBytesIns_Inst_Sbox_10_T3), .B(SubBytesIns_Inst_Sbox_10_T4), .Z(SubBytesIns_Inst_Sbox_10_T13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_T14_U1 ( .A(SubBytesIns_Inst_Sbox_10_T6), .B(SubBytesIns_Inst_Sbox_10_T11), .Z(SubBytesIns_Inst_Sbox_10_T14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_T15_U1 ( .A(SubBytesIns_Inst_Sbox_10_T5), .B(SubBytesIns_Inst_Sbox_10_T11), .Z(SubBytesIns_Inst_Sbox_10_T15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_T16_U1 ( .A(SubBytesIns_Inst_Sbox_10_T5), .B(SubBytesIns_Inst_Sbox_10_T12), .Z(SubBytesIns_Inst_Sbox_10_T16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_T17_U1 ( .A(SubBytesIns_Inst_Sbox_10_T9), .B(SubBytesIns_Inst_Sbox_10_T16), .Z(SubBytesIns_Inst_Sbox_10_T17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_T18_U1 ( .A(SubBytesInput[84]), .B(
        SubBytesInput[80]), .Z(SubBytesIns_Inst_Sbox_10_T18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_T19_U1 ( .A(SubBytesIns_Inst_Sbox_10_T7), .B(SubBytesIns_Inst_Sbox_10_T18), .Z(SubBytesIns_Inst_Sbox_10_T19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_T20_U1 ( .A(SubBytesIns_Inst_Sbox_10_T1), .B(SubBytesIns_Inst_Sbox_10_T19), .Z(SubBytesIns_Inst_Sbox_10_T20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_T21_U1 ( .A(SubBytesInput[81]), .B(
        SubBytesInput[80]), .Z(SubBytesIns_Inst_Sbox_10_T21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_T22_U1 ( .A(SubBytesIns_Inst_Sbox_10_T7), .B(SubBytesIns_Inst_Sbox_10_T21), .Z(SubBytesIns_Inst_Sbox_10_T22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_T23_U1 ( .A(SubBytesIns_Inst_Sbox_10_T2), .B(SubBytesIns_Inst_Sbox_10_T22), .Z(SubBytesIns_Inst_Sbox_10_T23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_T24_U1 ( .A(SubBytesIns_Inst_Sbox_10_T2), .B(SubBytesIns_Inst_Sbox_10_T10), .Z(SubBytesIns_Inst_Sbox_10_T24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_T25_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_T20), .B(SubBytesIns_Inst_Sbox_10_T17), .Z(
        SubBytesIns_Inst_Sbox_10_T25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_T26_U1 ( .A(SubBytesIns_Inst_Sbox_10_T3), .B(SubBytesIns_Inst_Sbox_10_T16), .Z(SubBytesIns_Inst_Sbox_10_T26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_T27_U1 ( .A(SubBytesIns_Inst_Sbox_10_T1), .B(SubBytesIns_Inst_Sbox_10_T12), .Z(SubBytesIns_Inst_Sbox_10_T27) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M1_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_T13), .A2(SubBytesIns_Inst_Sbox_10_T6), .ZN(
        SubBytesIns_Inst_Sbox_10_M1) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M2_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_T23), .A2(SubBytesIns_Inst_Sbox_10_T8), .ZN(
        SubBytesIns_Inst_Sbox_10_M2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_M3_U1 ( .A(SubBytesIns_Inst_Sbox_10_T14), .B(SubBytesIns_Inst_Sbox_10_M1), .Z(SubBytesIns_Inst_Sbox_10_M3) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M4_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_T19), .A2(SubBytesInput[80]), .ZN(
        SubBytesIns_Inst_Sbox_10_M4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_M5_U1 ( .A(SubBytesIns_Inst_Sbox_10_M4), 
        .B(SubBytesIns_Inst_Sbox_10_M1), .Z(SubBytesIns_Inst_Sbox_10_M5) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M6_U1 ( .A1(SubBytesIns_Inst_Sbox_10_T3), .A2(SubBytesIns_Inst_Sbox_10_T16), .ZN(SubBytesIns_Inst_Sbox_10_M6) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M7_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_T22), .A2(SubBytesIns_Inst_Sbox_10_T9), .ZN(
        SubBytesIns_Inst_Sbox_10_M7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_M8_U1 ( .A(SubBytesIns_Inst_Sbox_10_T26), .B(SubBytesIns_Inst_Sbox_10_M6), .Z(SubBytesIns_Inst_Sbox_10_M8) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M9_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_T20), .A2(SubBytesIns_Inst_Sbox_10_T17), .ZN(
        SubBytesIns_Inst_Sbox_10_M9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_M10_U1 ( .A(SubBytesIns_Inst_Sbox_10_M9), .B(SubBytesIns_Inst_Sbox_10_M6), .Z(SubBytesIns_Inst_Sbox_10_M10) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M11_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_T1), .A2(SubBytesIns_Inst_Sbox_10_T15), .ZN(
        SubBytesIns_Inst_Sbox_10_M11) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M12_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_T4), .A2(SubBytesIns_Inst_Sbox_10_T27), .ZN(
        SubBytesIns_Inst_Sbox_10_M12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_M13_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_M12), .B(SubBytesIns_Inst_Sbox_10_M11), .Z(
        SubBytesIns_Inst_Sbox_10_M13) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M14_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_T2), .A2(SubBytesIns_Inst_Sbox_10_T10), .ZN(
        SubBytesIns_Inst_Sbox_10_M14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_M15_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_M14), .B(SubBytesIns_Inst_Sbox_10_M11), .Z(
        SubBytesIns_Inst_Sbox_10_M15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_M16_U1 ( .A(SubBytesIns_Inst_Sbox_10_M3), .B(SubBytesIns_Inst_Sbox_10_M2), .Z(SubBytesIns_Inst_Sbox_10_M16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_M17_U1 ( .A(SubBytesIns_Inst_Sbox_10_M5), .B(SubBytesIns_Inst_Sbox_10_T24), .Z(SubBytesIns_Inst_Sbox_10_M17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_M18_U1 ( .A(SubBytesIns_Inst_Sbox_10_M8), .B(SubBytesIns_Inst_Sbox_10_M7), .Z(SubBytesIns_Inst_Sbox_10_M18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_M19_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_M10), .B(SubBytesIns_Inst_Sbox_10_M15), .Z(
        SubBytesIns_Inst_Sbox_10_M19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_M20_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_M16), .B(SubBytesIns_Inst_Sbox_10_M13), .Z(
        SubBytesIns_Inst_Sbox_10_M20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_M21_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_M17), .B(SubBytesIns_Inst_Sbox_10_M15), .Z(
        SubBytesIns_Inst_Sbox_10_M21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_M22_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_M18), .B(SubBytesIns_Inst_Sbox_10_M13), .Z(
        SubBytesIns_Inst_Sbox_10_M22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_M23_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_M19), .B(SubBytesIns_Inst_Sbox_10_T25), .Z(
        SubBytesIns_Inst_Sbox_10_M23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_M24_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_M22), .B(SubBytesIns_Inst_Sbox_10_M23), .Z(
        SubBytesIns_Inst_Sbox_10_M24) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M25_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_M22), .A2(SubBytesIns_Inst_Sbox_10_M20), .ZN(
        SubBytesIns_Inst_Sbox_10_M25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_M26_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_M21), .B(SubBytesIns_Inst_Sbox_10_M25), .Z(
        SubBytesIns_Inst_Sbox_10_M26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_M27_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_M20), .B(SubBytesIns_Inst_Sbox_10_M21), .Z(
        SubBytesIns_Inst_Sbox_10_M27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_M28_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_M23), .B(SubBytesIns_Inst_Sbox_10_M25), .Z(
        SubBytesIns_Inst_Sbox_10_M28) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M29_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_M28), .A2(SubBytesIns_Inst_Sbox_10_M27), .ZN(
        SubBytesIns_Inst_Sbox_10_M29) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M30_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_M26), .A2(SubBytesIns_Inst_Sbox_10_M24), .ZN(
        SubBytesIns_Inst_Sbox_10_M30) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M31_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_M20), .A2(SubBytesIns_Inst_Sbox_10_M23), .ZN(
        SubBytesIns_Inst_Sbox_10_M31) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M32_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_M27), .A2(SubBytesIns_Inst_Sbox_10_M31), .ZN(
        SubBytesIns_Inst_Sbox_10_M32) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_M33_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_M27), .B(SubBytesIns_Inst_Sbox_10_M25), .Z(
        SubBytesIns_Inst_Sbox_10_M33) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M34_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_M21), .A2(SubBytesIns_Inst_Sbox_10_M22), .ZN(
        SubBytesIns_Inst_Sbox_10_M34) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M35_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_M24), .A2(SubBytesIns_Inst_Sbox_10_M34), .ZN(
        SubBytesIns_Inst_Sbox_10_M35) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_M36_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_M24), .B(SubBytesIns_Inst_Sbox_10_M25), .Z(
        SubBytesIns_Inst_Sbox_10_M36) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_M37_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_M21), .B(SubBytesIns_Inst_Sbox_10_M29), .Z(
        SubBytesIns_Inst_Sbox_10_M37) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_M38_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_M32), .B(SubBytesIns_Inst_Sbox_10_M33), .Z(
        SubBytesIns_Inst_Sbox_10_M38) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_M39_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_M23), .B(SubBytesIns_Inst_Sbox_10_M30), .Z(
        SubBytesIns_Inst_Sbox_10_M39) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_M40_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_M35), .B(SubBytesIns_Inst_Sbox_10_M36), .Z(
        SubBytesIns_Inst_Sbox_10_M40) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_M41_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_M38), .B(SubBytesIns_Inst_Sbox_10_M40), .Z(
        SubBytesIns_Inst_Sbox_10_M41) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_M42_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_M37), .B(SubBytesIns_Inst_Sbox_10_M39), .Z(
        SubBytesIns_Inst_Sbox_10_M42) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_M43_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_M37), .B(SubBytesIns_Inst_Sbox_10_M38), .Z(
        SubBytesIns_Inst_Sbox_10_M43) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_M44_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_M39), .B(SubBytesIns_Inst_Sbox_10_M40), .Z(
        SubBytesIns_Inst_Sbox_10_M44) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_M45_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_M42), .B(SubBytesIns_Inst_Sbox_10_M41), .Z(
        SubBytesIns_Inst_Sbox_10_M45) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M46_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_M44), .A2(SubBytesIns_Inst_Sbox_10_T6), .ZN(
        SubBytesIns_Inst_Sbox_10_M46) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M47_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_M40), .A2(SubBytesIns_Inst_Sbox_10_T8), .ZN(
        SubBytesIns_Inst_Sbox_10_M47) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M48_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_M39), .A2(SubBytesInput[80]), .ZN(
        SubBytesIns_Inst_Sbox_10_M48) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M49_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_M43), .A2(SubBytesIns_Inst_Sbox_10_T16), .ZN(
        SubBytesIns_Inst_Sbox_10_M49) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M50_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_M38), .A2(SubBytesIns_Inst_Sbox_10_T9), .ZN(
        SubBytesIns_Inst_Sbox_10_M50) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M51_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_M37), .A2(SubBytesIns_Inst_Sbox_10_T17), .ZN(
        SubBytesIns_Inst_Sbox_10_M51) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M52_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_M42), .A2(SubBytesIns_Inst_Sbox_10_T15), .ZN(
        SubBytesIns_Inst_Sbox_10_M52) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M53_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_M45), .A2(SubBytesIns_Inst_Sbox_10_T27), .ZN(
        SubBytesIns_Inst_Sbox_10_M53) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M54_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_M41), .A2(SubBytesIns_Inst_Sbox_10_T10), .ZN(
        SubBytesIns_Inst_Sbox_10_M54) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M55_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_M44), .A2(SubBytesIns_Inst_Sbox_10_T13), .ZN(
        SubBytesIns_Inst_Sbox_10_M55) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M56_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_M40), .A2(SubBytesIns_Inst_Sbox_10_T23), .ZN(
        SubBytesIns_Inst_Sbox_10_M56) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M57_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_M39), .A2(SubBytesIns_Inst_Sbox_10_T19), .ZN(
        SubBytesIns_Inst_Sbox_10_M57) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M58_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_M43), .A2(SubBytesIns_Inst_Sbox_10_T3), .ZN(
        SubBytesIns_Inst_Sbox_10_M58) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M59_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_M38), .A2(SubBytesIns_Inst_Sbox_10_T22), .ZN(
        SubBytesIns_Inst_Sbox_10_M59) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M60_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_M37), .A2(SubBytesIns_Inst_Sbox_10_T20), .ZN(
        SubBytesIns_Inst_Sbox_10_M60) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M61_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_M42), .A2(SubBytesIns_Inst_Sbox_10_T1), .ZN(
        SubBytesIns_Inst_Sbox_10_M61) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M62_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_M45), .A2(SubBytesIns_Inst_Sbox_10_T4), .ZN(
        SubBytesIns_Inst_Sbox_10_M62) );
  AND2_X1 SubBytesIns_Inst_Sbox_10_AND_M63_U1 ( .A1(
        SubBytesIns_Inst_Sbox_10_M41), .A2(SubBytesIns_Inst_Sbox_10_T2), .ZN(
        SubBytesIns_Inst_Sbox_10_M63) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_L0_U1 ( .A(SubBytesIns_Inst_Sbox_10_M61), .B(SubBytesIns_Inst_Sbox_10_M62), .Z(SubBytesIns_Inst_Sbox_10_L0) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_L1_U1 ( .A(SubBytesIns_Inst_Sbox_10_M50), .B(SubBytesIns_Inst_Sbox_10_M56), .Z(SubBytesIns_Inst_Sbox_10_L1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_L2_U1 ( .A(SubBytesIns_Inst_Sbox_10_M46), .B(SubBytesIns_Inst_Sbox_10_M48), .Z(SubBytesIns_Inst_Sbox_10_L2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_L3_U1 ( .A(SubBytesIns_Inst_Sbox_10_M47), .B(SubBytesIns_Inst_Sbox_10_M55), .Z(SubBytesIns_Inst_Sbox_10_L3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_L4_U1 ( .A(SubBytesIns_Inst_Sbox_10_M54), .B(SubBytesIns_Inst_Sbox_10_M58), .Z(SubBytesIns_Inst_Sbox_10_L4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_L5_U1 ( .A(SubBytesIns_Inst_Sbox_10_M49), .B(SubBytesIns_Inst_Sbox_10_M61), .Z(SubBytesIns_Inst_Sbox_10_L5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_L6_U1 ( .A(SubBytesIns_Inst_Sbox_10_M62), .B(SubBytesIns_Inst_Sbox_10_L5), .Z(SubBytesIns_Inst_Sbox_10_L6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_L7_U1 ( .A(SubBytesIns_Inst_Sbox_10_M46), .B(SubBytesIns_Inst_Sbox_10_L3), .Z(SubBytesIns_Inst_Sbox_10_L7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_L8_U1 ( .A(SubBytesIns_Inst_Sbox_10_M51), .B(SubBytesIns_Inst_Sbox_10_M59), .Z(SubBytesIns_Inst_Sbox_10_L8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_L9_U1 ( .A(SubBytesIns_Inst_Sbox_10_M52), .B(SubBytesIns_Inst_Sbox_10_M53), .Z(SubBytesIns_Inst_Sbox_10_L9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_L10_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_M53), .B(SubBytesIns_Inst_Sbox_10_L4), .Z(
        SubBytesIns_Inst_Sbox_10_L10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_L11_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_M60), .B(SubBytesIns_Inst_Sbox_10_L2), .Z(
        SubBytesIns_Inst_Sbox_10_L11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_L12_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_M48), .B(SubBytesIns_Inst_Sbox_10_M51), .Z(
        SubBytesIns_Inst_Sbox_10_L12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_L13_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_M50), .B(SubBytesIns_Inst_Sbox_10_L0), .Z(
        SubBytesIns_Inst_Sbox_10_L13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_L14_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_M52), .B(SubBytesIns_Inst_Sbox_10_M61), .Z(
        SubBytesIns_Inst_Sbox_10_L14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_L15_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_M55), .B(SubBytesIns_Inst_Sbox_10_L1), .Z(
        SubBytesIns_Inst_Sbox_10_L15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_L16_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_M56), .B(SubBytesIns_Inst_Sbox_10_L0), .Z(
        SubBytesIns_Inst_Sbox_10_L16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_L17_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_M57), .B(SubBytesIns_Inst_Sbox_10_L1), .Z(
        SubBytesIns_Inst_Sbox_10_L17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_L18_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_M58), .B(SubBytesIns_Inst_Sbox_10_L8), .Z(
        SubBytesIns_Inst_Sbox_10_L18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_L19_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_M63), .B(SubBytesIns_Inst_Sbox_10_L4), .Z(
        SubBytesIns_Inst_Sbox_10_L19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_L20_U1 ( .A(SubBytesIns_Inst_Sbox_10_L0), .B(SubBytesIns_Inst_Sbox_10_L1), .Z(SubBytesIns_Inst_Sbox_10_L20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_L21_U1 ( .A(SubBytesIns_Inst_Sbox_10_L1), .B(SubBytesIns_Inst_Sbox_10_L7), .Z(SubBytesIns_Inst_Sbox_10_L21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_L22_U1 ( .A(SubBytesIns_Inst_Sbox_10_L3), .B(SubBytesIns_Inst_Sbox_10_L12), .Z(SubBytesIns_Inst_Sbox_10_L22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_L23_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_L18), .B(SubBytesIns_Inst_Sbox_10_L2), .Z(
        SubBytesIns_Inst_Sbox_10_L23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_L24_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_L15), .B(SubBytesIns_Inst_Sbox_10_L9), .Z(
        SubBytesIns_Inst_Sbox_10_L24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_L25_U1 ( .A(SubBytesIns_Inst_Sbox_10_L6), .B(SubBytesIns_Inst_Sbox_10_L10), .Z(SubBytesIns_Inst_Sbox_10_L25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_L26_U1 ( .A(SubBytesIns_Inst_Sbox_10_L7), .B(SubBytesIns_Inst_Sbox_10_L9), .Z(SubBytesIns_Inst_Sbox_10_L26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_L27_U1 ( .A(SubBytesIns_Inst_Sbox_10_L8), .B(SubBytesIns_Inst_Sbox_10_L10), .Z(SubBytesIns_Inst_Sbox_10_L27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_L28_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_L11), .B(SubBytesIns_Inst_Sbox_10_L14), .Z(
        SubBytesIns_Inst_Sbox_10_L28) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_L29_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_L11), .B(SubBytesIns_Inst_Sbox_10_L17), .Z(
        SubBytesIns_Inst_Sbox_10_L29) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_S0_U1 ( .A(SubBytesIns_Inst_Sbox_10_L6), 
        .B(SubBytesIns_Inst_Sbox_10_L24), .Z(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_S1_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_L16), .B(SubBytesIns_Inst_Sbox_10_L26), .ZN(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[23]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_S2_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_L19), .B(SubBytesIns_Inst_Sbox_10_L28), .ZN(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[22]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_S3_U1 ( .A(SubBytesIns_Inst_Sbox_10_L6), 
        .B(SubBytesIns_Inst_Sbox_10_L21), .Z(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[21]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_S4_U1 ( .A(SubBytesIns_Inst_Sbox_10_L20), .B(SubBytesIns_Inst_Sbox_10_L22), .Z(MixColumnsInput[115]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_S5_U1 ( .A(SubBytesIns_Inst_Sbox_10_L25), .B(SubBytesIns_Inst_Sbox_10_L29), .Z(MixColumnsInput[114]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_S6_U1 ( .A(
        SubBytesIns_Inst_Sbox_10_L13), .B(SubBytesIns_Inst_Sbox_10_L27), .ZN(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[18]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_10_XOR_S7_U1 ( .A(SubBytesIns_Inst_Sbox_10_L6), .B(SubBytesIns_Inst_Sbox_10_L23), .ZN(MixColumnsInput[112]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_T1_U1 ( .A(SubBytesInput[95]), .B(
        SubBytesInput[92]), .Z(SubBytesIns_Inst_Sbox_11_T1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_T2_U1 ( .A(SubBytesInput[95]), .B(
        SubBytesInput[90]), .Z(SubBytesIns_Inst_Sbox_11_T2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_T3_U1 ( .A(SubBytesInput[95]), .B(
        SubBytesInput[89]), .Z(SubBytesIns_Inst_Sbox_11_T3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_T4_U1 ( .A(SubBytesInput[92]), .B(
        SubBytesInput[90]), .Z(SubBytesIns_Inst_Sbox_11_T4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_T5_U1 ( .A(SubBytesInput[91]), .B(
        SubBytesInput[89]), .Z(SubBytesIns_Inst_Sbox_11_T5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_T6_U1 ( .A(SubBytesIns_Inst_Sbox_11_T1), 
        .B(SubBytesIns_Inst_Sbox_11_T5), .Z(SubBytesIns_Inst_Sbox_11_T6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_T7_U1 ( .A(SubBytesInput[94]), .B(
        SubBytesInput[93]), .Z(SubBytesIns_Inst_Sbox_11_T7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_T8_U1 ( .A(SubBytesInput[88]), .B(
        SubBytesIns_Inst_Sbox_11_T6), .Z(SubBytesIns_Inst_Sbox_11_T8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_T9_U1 ( .A(SubBytesInput[88]), .B(
        SubBytesIns_Inst_Sbox_11_T7), .Z(SubBytesIns_Inst_Sbox_11_T9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_T10_U1 ( .A(SubBytesIns_Inst_Sbox_11_T6), .B(SubBytesIns_Inst_Sbox_11_T7), .Z(SubBytesIns_Inst_Sbox_11_T10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_T11_U1 ( .A(SubBytesInput[94]), .B(
        SubBytesInput[90]), .Z(SubBytesIns_Inst_Sbox_11_T11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_T12_U1 ( .A(SubBytesInput[93]), .B(
        SubBytesInput[90]), .Z(SubBytesIns_Inst_Sbox_11_T12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_T13_U1 ( .A(SubBytesIns_Inst_Sbox_11_T3), .B(SubBytesIns_Inst_Sbox_11_T4), .Z(SubBytesIns_Inst_Sbox_11_T13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_T14_U1 ( .A(SubBytesIns_Inst_Sbox_11_T6), .B(SubBytesIns_Inst_Sbox_11_T11), .Z(SubBytesIns_Inst_Sbox_11_T14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_T15_U1 ( .A(SubBytesIns_Inst_Sbox_11_T5), .B(SubBytesIns_Inst_Sbox_11_T11), .Z(SubBytesIns_Inst_Sbox_11_T15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_T16_U1 ( .A(SubBytesIns_Inst_Sbox_11_T5), .B(SubBytesIns_Inst_Sbox_11_T12), .Z(SubBytesIns_Inst_Sbox_11_T16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_T17_U1 ( .A(SubBytesIns_Inst_Sbox_11_T9), .B(SubBytesIns_Inst_Sbox_11_T16), .Z(SubBytesIns_Inst_Sbox_11_T17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_T18_U1 ( .A(SubBytesInput[92]), .B(
        SubBytesInput[88]), .Z(SubBytesIns_Inst_Sbox_11_T18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_T19_U1 ( .A(SubBytesIns_Inst_Sbox_11_T7), .B(SubBytesIns_Inst_Sbox_11_T18), .Z(SubBytesIns_Inst_Sbox_11_T19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_T20_U1 ( .A(SubBytesIns_Inst_Sbox_11_T1), .B(SubBytesIns_Inst_Sbox_11_T19), .Z(SubBytesIns_Inst_Sbox_11_T20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_T21_U1 ( .A(SubBytesInput[89]), .B(
        SubBytesInput[88]), .Z(SubBytesIns_Inst_Sbox_11_T21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_T22_U1 ( .A(SubBytesIns_Inst_Sbox_11_T7), .B(SubBytesIns_Inst_Sbox_11_T21), .Z(SubBytesIns_Inst_Sbox_11_T22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_T23_U1 ( .A(SubBytesIns_Inst_Sbox_11_T2), .B(SubBytesIns_Inst_Sbox_11_T22), .Z(SubBytesIns_Inst_Sbox_11_T23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_T24_U1 ( .A(SubBytesIns_Inst_Sbox_11_T2), .B(SubBytesIns_Inst_Sbox_11_T10), .Z(SubBytesIns_Inst_Sbox_11_T24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_T25_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_T20), .B(SubBytesIns_Inst_Sbox_11_T17), .Z(
        SubBytesIns_Inst_Sbox_11_T25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_T26_U1 ( .A(SubBytesIns_Inst_Sbox_11_T3), .B(SubBytesIns_Inst_Sbox_11_T16), .Z(SubBytesIns_Inst_Sbox_11_T26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_T27_U1 ( .A(SubBytesIns_Inst_Sbox_11_T1), .B(SubBytesIns_Inst_Sbox_11_T12), .Z(SubBytesIns_Inst_Sbox_11_T27) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M1_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_T13), .A2(SubBytesIns_Inst_Sbox_11_T6), .ZN(
        SubBytesIns_Inst_Sbox_11_M1) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M2_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_T23), .A2(SubBytesIns_Inst_Sbox_11_T8), .ZN(
        SubBytesIns_Inst_Sbox_11_M2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_M3_U1 ( .A(SubBytesIns_Inst_Sbox_11_T14), .B(SubBytesIns_Inst_Sbox_11_M1), .Z(SubBytesIns_Inst_Sbox_11_M3) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M4_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_T19), .A2(SubBytesInput[88]), .ZN(
        SubBytesIns_Inst_Sbox_11_M4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_M5_U1 ( .A(SubBytesIns_Inst_Sbox_11_M4), 
        .B(SubBytesIns_Inst_Sbox_11_M1), .Z(SubBytesIns_Inst_Sbox_11_M5) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M6_U1 ( .A1(SubBytesIns_Inst_Sbox_11_T3), .A2(SubBytesIns_Inst_Sbox_11_T16), .ZN(SubBytesIns_Inst_Sbox_11_M6) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M7_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_T22), .A2(SubBytesIns_Inst_Sbox_11_T9), .ZN(
        SubBytesIns_Inst_Sbox_11_M7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_M8_U1 ( .A(SubBytesIns_Inst_Sbox_11_T26), .B(SubBytesIns_Inst_Sbox_11_M6), .Z(SubBytesIns_Inst_Sbox_11_M8) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M9_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_T20), .A2(SubBytesIns_Inst_Sbox_11_T17), .ZN(
        SubBytesIns_Inst_Sbox_11_M9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_M10_U1 ( .A(SubBytesIns_Inst_Sbox_11_M9), .B(SubBytesIns_Inst_Sbox_11_M6), .Z(SubBytesIns_Inst_Sbox_11_M10) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M11_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_T1), .A2(SubBytesIns_Inst_Sbox_11_T15), .ZN(
        SubBytesIns_Inst_Sbox_11_M11) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M12_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_T4), .A2(SubBytesIns_Inst_Sbox_11_T27), .ZN(
        SubBytesIns_Inst_Sbox_11_M12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_M13_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_M12), .B(SubBytesIns_Inst_Sbox_11_M11), .Z(
        SubBytesIns_Inst_Sbox_11_M13) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M14_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_T2), .A2(SubBytesIns_Inst_Sbox_11_T10), .ZN(
        SubBytesIns_Inst_Sbox_11_M14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_M15_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_M14), .B(SubBytesIns_Inst_Sbox_11_M11), .Z(
        SubBytesIns_Inst_Sbox_11_M15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_M16_U1 ( .A(SubBytesIns_Inst_Sbox_11_M3), .B(SubBytesIns_Inst_Sbox_11_M2), .Z(SubBytesIns_Inst_Sbox_11_M16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_M17_U1 ( .A(SubBytesIns_Inst_Sbox_11_M5), .B(SubBytesIns_Inst_Sbox_11_T24), .Z(SubBytesIns_Inst_Sbox_11_M17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_M18_U1 ( .A(SubBytesIns_Inst_Sbox_11_M8), .B(SubBytesIns_Inst_Sbox_11_M7), .Z(SubBytesIns_Inst_Sbox_11_M18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_M19_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_M10), .B(SubBytesIns_Inst_Sbox_11_M15), .Z(
        SubBytesIns_Inst_Sbox_11_M19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_M20_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_M16), .B(SubBytesIns_Inst_Sbox_11_M13), .Z(
        SubBytesIns_Inst_Sbox_11_M20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_M21_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_M17), .B(SubBytesIns_Inst_Sbox_11_M15), .Z(
        SubBytesIns_Inst_Sbox_11_M21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_M22_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_M18), .B(SubBytesIns_Inst_Sbox_11_M13), .Z(
        SubBytesIns_Inst_Sbox_11_M22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_M23_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_M19), .B(SubBytesIns_Inst_Sbox_11_T25), .Z(
        SubBytesIns_Inst_Sbox_11_M23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_M24_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_M22), .B(SubBytesIns_Inst_Sbox_11_M23), .Z(
        SubBytesIns_Inst_Sbox_11_M24) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M25_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_M22), .A2(SubBytesIns_Inst_Sbox_11_M20), .ZN(
        SubBytesIns_Inst_Sbox_11_M25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_M26_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_M21), .B(SubBytesIns_Inst_Sbox_11_M25), .Z(
        SubBytesIns_Inst_Sbox_11_M26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_M27_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_M20), .B(SubBytesIns_Inst_Sbox_11_M21), .Z(
        SubBytesIns_Inst_Sbox_11_M27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_M28_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_M23), .B(SubBytesIns_Inst_Sbox_11_M25), .Z(
        SubBytesIns_Inst_Sbox_11_M28) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M29_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_M28), .A2(SubBytesIns_Inst_Sbox_11_M27), .ZN(
        SubBytesIns_Inst_Sbox_11_M29) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M30_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_M26), .A2(SubBytesIns_Inst_Sbox_11_M24), .ZN(
        SubBytesIns_Inst_Sbox_11_M30) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M31_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_M20), .A2(SubBytesIns_Inst_Sbox_11_M23), .ZN(
        SubBytesIns_Inst_Sbox_11_M31) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M32_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_M27), .A2(SubBytesIns_Inst_Sbox_11_M31), .ZN(
        SubBytesIns_Inst_Sbox_11_M32) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_M33_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_M27), .B(SubBytesIns_Inst_Sbox_11_M25), .Z(
        SubBytesIns_Inst_Sbox_11_M33) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M34_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_M21), .A2(SubBytesIns_Inst_Sbox_11_M22), .ZN(
        SubBytesIns_Inst_Sbox_11_M34) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M35_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_M24), .A2(SubBytesIns_Inst_Sbox_11_M34), .ZN(
        SubBytesIns_Inst_Sbox_11_M35) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_M36_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_M24), .B(SubBytesIns_Inst_Sbox_11_M25), .Z(
        SubBytesIns_Inst_Sbox_11_M36) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_M37_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_M21), .B(SubBytesIns_Inst_Sbox_11_M29), .Z(
        SubBytesIns_Inst_Sbox_11_M37) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_M38_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_M32), .B(SubBytesIns_Inst_Sbox_11_M33), .Z(
        SubBytesIns_Inst_Sbox_11_M38) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_M39_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_M23), .B(SubBytesIns_Inst_Sbox_11_M30), .Z(
        SubBytesIns_Inst_Sbox_11_M39) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_M40_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_M35), .B(SubBytesIns_Inst_Sbox_11_M36), .Z(
        SubBytesIns_Inst_Sbox_11_M40) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_M41_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_M38), .B(SubBytesIns_Inst_Sbox_11_M40), .Z(
        SubBytesIns_Inst_Sbox_11_M41) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_M42_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_M37), .B(SubBytesIns_Inst_Sbox_11_M39), .Z(
        SubBytesIns_Inst_Sbox_11_M42) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_M43_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_M37), .B(SubBytesIns_Inst_Sbox_11_M38), .Z(
        SubBytesIns_Inst_Sbox_11_M43) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_M44_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_M39), .B(SubBytesIns_Inst_Sbox_11_M40), .Z(
        SubBytesIns_Inst_Sbox_11_M44) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_M45_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_M42), .B(SubBytesIns_Inst_Sbox_11_M41), .Z(
        SubBytesIns_Inst_Sbox_11_M45) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M46_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_M44), .A2(SubBytesIns_Inst_Sbox_11_T6), .ZN(
        SubBytesIns_Inst_Sbox_11_M46) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M47_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_M40), .A2(SubBytesIns_Inst_Sbox_11_T8), .ZN(
        SubBytesIns_Inst_Sbox_11_M47) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M48_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_M39), .A2(SubBytesInput[88]), .ZN(
        SubBytesIns_Inst_Sbox_11_M48) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M49_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_M43), .A2(SubBytesIns_Inst_Sbox_11_T16), .ZN(
        SubBytesIns_Inst_Sbox_11_M49) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M50_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_M38), .A2(SubBytesIns_Inst_Sbox_11_T9), .ZN(
        SubBytesIns_Inst_Sbox_11_M50) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M51_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_M37), .A2(SubBytesIns_Inst_Sbox_11_T17), .ZN(
        SubBytesIns_Inst_Sbox_11_M51) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M52_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_M42), .A2(SubBytesIns_Inst_Sbox_11_T15), .ZN(
        SubBytesIns_Inst_Sbox_11_M52) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M53_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_M45), .A2(SubBytesIns_Inst_Sbox_11_T27), .ZN(
        SubBytesIns_Inst_Sbox_11_M53) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M54_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_M41), .A2(SubBytesIns_Inst_Sbox_11_T10), .ZN(
        SubBytesIns_Inst_Sbox_11_M54) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M55_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_M44), .A2(SubBytesIns_Inst_Sbox_11_T13), .ZN(
        SubBytesIns_Inst_Sbox_11_M55) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M56_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_M40), .A2(SubBytesIns_Inst_Sbox_11_T23), .ZN(
        SubBytesIns_Inst_Sbox_11_M56) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M57_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_M39), .A2(SubBytesIns_Inst_Sbox_11_T19), .ZN(
        SubBytesIns_Inst_Sbox_11_M57) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M58_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_M43), .A2(SubBytesIns_Inst_Sbox_11_T3), .ZN(
        SubBytesIns_Inst_Sbox_11_M58) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M59_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_M38), .A2(SubBytesIns_Inst_Sbox_11_T22), .ZN(
        SubBytesIns_Inst_Sbox_11_M59) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M60_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_M37), .A2(SubBytesIns_Inst_Sbox_11_T20), .ZN(
        SubBytesIns_Inst_Sbox_11_M60) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M61_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_M42), .A2(SubBytesIns_Inst_Sbox_11_T1), .ZN(
        SubBytesIns_Inst_Sbox_11_M61) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M62_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_M45), .A2(SubBytesIns_Inst_Sbox_11_T4), .ZN(
        SubBytesIns_Inst_Sbox_11_M62) );
  AND2_X1 SubBytesIns_Inst_Sbox_11_AND_M63_U1 ( .A1(
        SubBytesIns_Inst_Sbox_11_M41), .A2(SubBytesIns_Inst_Sbox_11_T2), .ZN(
        SubBytesIns_Inst_Sbox_11_M63) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_L0_U1 ( .A(SubBytesIns_Inst_Sbox_11_M61), .B(SubBytesIns_Inst_Sbox_11_M62), .Z(SubBytesIns_Inst_Sbox_11_L0) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_L1_U1 ( .A(SubBytesIns_Inst_Sbox_11_M50), .B(SubBytesIns_Inst_Sbox_11_M56), .Z(SubBytesIns_Inst_Sbox_11_L1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_L2_U1 ( .A(SubBytesIns_Inst_Sbox_11_M46), .B(SubBytesIns_Inst_Sbox_11_M48), .Z(SubBytesIns_Inst_Sbox_11_L2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_L3_U1 ( .A(SubBytesIns_Inst_Sbox_11_M47), .B(SubBytesIns_Inst_Sbox_11_M55), .Z(SubBytesIns_Inst_Sbox_11_L3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_L4_U1 ( .A(SubBytesIns_Inst_Sbox_11_M54), .B(SubBytesIns_Inst_Sbox_11_M58), .Z(SubBytesIns_Inst_Sbox_11_L4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_L5_U1 ( .A(SubBytesIns_Inst_Sbox_11_M49), .B(SubBytesIns_Inst_Sbox_11_M61), .Z(SubBytesIns_Inst_Sbox_11_L5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_L6_U1 ( .A(SubBytesIns_Inst_Sbox_11_M62), .B(SubBytesIns_Inst_Sbox_11_L5), .Z(SubBytesIns_Inst_Sbox_11_L6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_L7_U1 ( .A(SubBytesIns_Inst_Sbox_11_M46), .B(SubBytesIns_Inst_Sbox_11_L3), .Z(SubBytesIns_Inst_Sbox_11_L7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_L8_U1 ( .A(SubBytesIns_Inst_Sbox_11_M51), .B(SubBytesIns_Inst_Sbox_11_M59), .Z(SubBytesIns_Inst_Sbox_11_L8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_L9_U1 ( .A(SubBytesIns_Inst_Sbox_11_M52), .B(SubBytesIns_Inst_Sbox_11_M53), .Z(SubBytesIns_Inst_Sbox_11_L9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_L10_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_M53), .B(SubBytesIns_Inst_Sbox_11_L4), .Z(
        SubBytesIns_Inst_Sbox_11_L10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_L11_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_M60), .B(SubBytesIns_Inst_Sbox_11_L2), .Z(
        SubBytesIns_Inst_Sbox_11_L11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_L12_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_M48), .B(SubBytesIns_Inst_Sbox_11_M51), .Z(
        SubBytesIns_Inst_Sbox_11_L12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_L13_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_M50), .B(SubBytesIns_Inst_Sbox_11_L0), .Z(
        SubBytesIns_Inst_Sbox_11_L13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_L14_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_M52), .B(SubBytesIns_Inst_Sbox_11_M61), .Z(
        SubBytesIns_Inst_Sbox_11_L14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_L15_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_M55), .B(SubBytesIns_Inst_Sbox_11_L1), .Z(
        SubBytesIns_Inst_Sbox_11_L15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_L16_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_M56), .B(SubBytesIns_Inst_Sbox_11_L0), .Z(
        SubBytesIns_Inst_Sbox_11_L16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_L17_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_M57), .B(SubBytesIns_Inst_Sbox_11_L1), .Z(
        SubBytesIns_Inst_Sbox_11_L17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_L18_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_M58), .B(SubBytesIns_Inst_Sbox_11_L8), .Z(
        SubBytesIns_Inst_Sbox_11_L18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_L19_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_M63), .B(SubBytesIns_Inst_Sbox_11_L4), .Z(
        SubBytesIns_Inst_Sbox_11_L19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_L20_U1 ( .A(SubBytesIns_Inst_Sbox_11_L0), .B(SubBytesIns_Inst_Sbox_11_L1), .Z(SubBytesIns_Inst_Sbox_11_L20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_L21_U1 ( .A(SubBytesIns_Inst_Sbox_11_L1), .B(SubBytesIns_Inst_Sbox_11_L7), .Z(SubBytesIns_Inst_Sbox_11_L21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_L22_U1 ( .A(SubBytesIns_Inst_Sbox_11_L3), .B(SubBytesIns_Inst_Sbox_11_L12), .Z(SubBytesIns_Inst_Sbox_11_L22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_L23_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_L18), .B(SubBytesIns_Inst_Sbox_11_L2), .Z(
        SubBytesIns_Inst_Sbox_11_L23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_L24_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_L15), .B(SubBytesIns_Inst_Sbox_11_L9), .Z(
        SubBytesIns_Inst_Sbox_11_L24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_L25_U1 ( .A(SubBytesIns_Inst_Sbox_11_L6), .B(SubBytesIns_Inst_Sbox_11_L10), .Z(SubBytesIns_Inst_Sbox_11_L25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_L26_U1 ( .A(SubBytesIns_Inst_Sbox_11_L7), .B(SubBytesIns_Inst_Sbox_11_L9), .Z(SubBytesIns_Inst_Sbox_11_L26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_L27_U1 ( .A(SubBytesIns_Inst_Sbox_11_L8), .B(SubBytesIns_Inst_Sbox_11_L10), .Z(SubBytesIns_Inst_Sbox_11_L27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_L28_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_L11), .B(SubBytesIns_Inst_Sbox_11_L14), .Z(
        SubBytesIns_Inst_Sbox_11_L28) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_L29_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_L11), .B(SubBytesIns_Inst_Sbox_11_L17), .Z(
        SubBytesIns_Inst_Sbox_11_L29) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_S0_U1 ( .A(SubBytesIns_Inst_Sbox_11_L6), 
        .B(SubBytesIns_Inst_Sbox_11_L24), .Z(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_S1_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_L16), .B(SubBytesIns_Inst_Sbox_11_L26), .ZN(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[31]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_S2_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_L19), .B(SubBytesIns_Inst_Sbox_11_L28), .ZN(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[30]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_S3_U1 ( .A(SubBytesIns_Inst_Sbox_11_L6), 
        .B(SubBytesIns_Inst_Sbox_11_L21), .Z(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[29]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_S4_U1 ( .A(SubBytesIns_Inst_Sbox_11_L20), .B(SubBytesIns_Inst_Sbox_11_L22), .Z(MixColumnsInput[91]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_S5_U1 ( .A(SubBytesIns_Inst_Sbox_11_L25), .B(SubBytesIns_Inst_Sbox_11_L29), .Z(MixColumnsInput[90]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_S6_U1 ( .A(
        SubBytesIns_Inst_Sbox_11_L13), .B(SubBytesIns_Inst_Sbox_11_L27), .ZN(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[26]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_11_XOR_S7_U1 ( .A(SubBytesIns_Inst_Sbox_11_L6), .B(SubBytesIns_Inst_Sbox_11_L23), .ZN(MixColumnsInput[88]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_T1_U1 ( .A(SubBytesInput[103]), .B(
        SubBytesInput[100]), .Z(SubBytesIns_Inst_Sbox_12_T1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_T2_U1 ( .A(SubBytesInput[103]), .B(
        SubBytesInput[98]), .Z(SubBytesIns_Inst_Sbox_12_T2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_T3_U1 ( .A(SubBytesInput[103]), .B(
        SubBytesInput[97]), .Z(SubBytesIns_Inst_Sbox_12_T3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_T4_U1 ( .A(SubBytesInput[100]), .B(
        SubBytesInput[98]), .Z(SubBytesIns_Inst_Sbox_12_T4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_T5_U1 ( .A(SubBytesInput[99]), .B(
        SubBytesInput[97]), .Z(SubBytesIns_Inst_Sbox_12_T5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_T6_U1 ( .A(SubBytesIns_Inst_Sbox_12_T1), 
        .B(SubBytesIns_Inst_Sbox_12_T5), .Z(SubBytesIns_Inst_Sbox_12_T6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_T7_U1 ( .A(SubBytesInput[102]), .B(
        SubBytesInput[101]), .Z(SubBytesIns_Inst_Sbox_12_T7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_T8_U1 ( .A(SubBytesInput[96]), .B(
        SubBytesIns_Inst_Sbox_12_T6), .Z(SubBytesIns_Inst_Sbox_12_T8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_T9_U1 ( .A(SubBytesInput[96]), .B(
        SubBytesIns_Inst_Sbox_12_T7), .Z(SubBytesIns_Inst_Sbox_12_T9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_T10_U1 ( .A(SubBytesIns_Inst_Sbox_12_T6), .B(SubBytesIns_Inst_Sbox_12_T7), .Z(SubBytesIns_Inst_Sbox_12_T10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_T11_U1 ( .A(SubBytesInput[102]), .B(
        SubBytesInput[98]), .Z(SubBytesIns_Inst_Sbox_12_T11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_T12_U1 ( .A(SubBytesInput[101]), .B(
        SubBytesInput[98]), .Z(SubBytesIns_Inst_Sbox_12_T12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_T13_U1 ( .A(SubBytesIns_Inst_Sbox_12_T3), .B(SubBytesIns_Inst_Sbox_12_T4), .Z(SubBytesIns_Inst_Sbox_12_T13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_T14_U1 ( .A(SubBytesIns_Inst_Sbox_12_T6), .B(SubBytesIns_Inst_Sbox_12_T11), .Z(SubBytesIns_Inst_Sbox_12_T14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_T15_U1 ( .A(SubBytesIns_Inst_Sbox_12_T5), .B(SubBytesIns_Inst_Sbox_12_T11), .Z(SubBytesIns_Inst_Sbox_12_T15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_T16_U1 ( .A(SubBytesIns_Inst_Sbox_12_T5), .B(SubBytesIns_Inst_Sbox_12_T12), .Z(SubBytesIns_Inst_Sbox_12_T16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_T17_U1 ( .A(SubBytesIns_Inst_Sbox_12_T9), .B(SubBytesIns_Inst_Sbox_12_T16), .Z(SubBytesIns_Inst_Sbox_12_T17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_T18_U1 ( .A(SubBytesInput[100]), .B(
        SubBytesInput[96]), .Z(SubBytesIns_Inst_Sbox_12_T18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_T19_U1 ( .A(SubBytesIns_Inst_Sbox_12_T7), .B(SubBytesIns_Inst_Sbox_12_T18), .Z(SubBytesIns_Inst_Sbox_12_T19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_T20_U1 ( .A(SubBytesIns_Inst_Sbox_12_T1), .B(SubBytesIns_Inst_Sbox_12_T19), .Z(SubBytesIns_Inst_Sbox_12_T20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_T21_U1 ( .A(SubBytesInput[97]), .B(
        SubBytesInput[96]), .Z(SubBytesIns_Inst_Sbox_12_T21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_T22_U1 ( .A(SubBytesIns_Inst_Sbox_12_T7), .B(SubBytesIns_Inst_Sbox_12_T21), .Z(SubBytesIns_Inst_Sbox_12_T22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_T23_U1 ( .A(SubBytesIns_Inst_Sbox_12_T2), .B(SubBytesIns_Inst_Sbox_12_T22), .Z(SubBytesIns_Inst_Sbox_12_T23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_T24_U1 ( .A(SubBytesIns_Inst_Sbox_12_T2), .B(SubBytesIns_Inst_Sbox_12_T10), .Z(SubBytesIns_Inst_Sbox_12_T24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_T25_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_T20), .B(SubBytesIns_Inst_Sbox_12_T17), .Z(
        SubBytesIns_Inst_Sbox_12_T25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_T26_U1 ( .A(SubBytesIns_Inst_Sbox_12_T3), .B(SubBytesIns_Inst_Sbox_12_T16), .Z(SubBytesIns_Inst_Sbox_12_T26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_T27_U1 ( .A(SubBytesIns_Inst_Sbox_12_T1), .B(SubBytesIns_Inst_Sbox_12_T12), .Z(SubBytesIns_Inst_Sbox_12_T27) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M1_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_T13), .A2(SubBytesIns_Inst_Sbox_12_T6), .ZN(
        SubBytesIns_Inst_Sbox_12_M1) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M2_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_T23), .A2(SubBytesIns_Inst_Sbox_12_T8), .ZN(
        SubBytesIns_Inst_Sbox_12_M2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_M3_U1 ( .A(SubBytesIns_Inst_Sbox_12_T14), .B(SubBytesIns_Inst_Sbox_12_M1), .Z(SubBytesIns_Inst_Sbox_12_M3) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M4_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_T19), .A2(SubBytesInput[96]), .ZN(
        SubBytesIns_Inst_Sbox_12_M4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_M5_U1 ( .A(SubBytesIns_Inst_Sbox_12_M4), 
        .B(SubBytesIns_Inst_Sbox_12_M1), .Z(SubBytesIns_Inst_Sbox_12_M5) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M6_U1 ( .A1(SubBytesIns_Inst_Sbox_12_T3), .A2(SubBytesIns_Inst_Sbox_12_T16), .ZN(SubBytesIns_Inst_Sbox_12_M6) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M7_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_T22), .A2(SubBytesIns_Inst_Sbox_12_T9), .ZN(
        SubBytesIns_Inst_Sbox_12_M7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_M8_U1 ( .A(SubBytesIns_Inst_Sbox_12_T26), .B(SubBytesIns_Inst_Sbox_12_M6), .Z(SubBytesIns_Inst_Sbox_12_M8) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M9_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_T20), .A2(SubBytesIns_Inst_Sbox_12_T17), .ZN(
        SubBytesIns_Inst_Sbox_12_M9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_M10_U1 ( .A(SubBytesIns_Inst_Sbox_12_M9), .B(SubBytesIns_Inst_Sbox_12_M6), .Z(SubBytesIns_Inst_Sbox_12_M10) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M11_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_T1), .A2(SubBytesIns_Inst_Sbox_12_T15), .ZN(
        SubBytesIns_Inst_Sbox_12_M11) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M12_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_T4), .A2(SubBytesIns_Inst_Sbox_12_T27), .ZN(
        SubBytesIns_Inst_Sbox_12_M12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_M13_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_M12), .B(SubBytesIns_Inst_Sbox_12_M11), .Z(
        SubBytesIns_Inst_Sbox_12_M13) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M14_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_T2), .A2(SubBytesIns_Inst_Sbox_12_T10), .ZN(
        SubBytesIns_Inst_Sbox_12_M14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_M15_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_M14), .B(SubBytesIns_Inst_Sbox_12_M11), .Z(
        SubBytesIns_Inst_Sbox_12_M15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_M16_U1 ( .A(SubBytesIns_Inst_Sbox_12_M3), .B(SubBytesIns_Inst_Sbox_12_M2), .Z(SubBytesIns_Inst_Sbox_12_M16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_M17_U1 ( .A(SubBytesIns_Inst_Sbox_12_M5), .B(SubBytesIns_Inst_Sbox_12_T24), .Z(SubBytesIns_Inst_Sbox_12_M17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_M18_U1 ( .A(SubBytesIns_Inst_Sbox_12_M8), .B(SubBytesIns_Inst_Sbox_12_M7), .Z(SubBytesIns_Inst_Sbox_12_M18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_M19_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_M10), .B(SubBytesIns_Inst_Sbox_12_M15), .Z(
        SubBytesIns_Inst_Sbox_12_M19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_M20_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_M16), .B(SubBytesIns_Inst_Sbox_12_M13), .Z(
        SubBytesIns_Inst_Sbox_12_M20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_M21_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_M17), .B(SubBytesIns_Inst_Sbox_12_M15), .Z(
        SubBytesIns_Inst_Sbox_12_M21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_M22_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_M18), .B(SubBytesIns_Inst_Sbox_12_M13), .Z(
        SubBytesIns_Inst_Sbox_12_M22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_M23_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_M19), .B(SubBytesIns_Inst_Sbox_12_T25), .Z(
        SubBytesIns_Inst_Sbox_12_M23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_M24_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_M22), .B(SubBytesIns_Inst_Sbox_12_M23), .Z(
        SubBytesIns_Inst_Sbox_12_M24) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M25_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_M22), .A2(SubBytesIns_Inst_Sbox_12_M20), .ZN(
        SubBytesIns_Inst_Sbox_12_M25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_M26_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_M21), .B(SubBytesIns_Inst_Sbox_12_M25), .Z(
        SubBytesIns_Inst_Sbox_12_M26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_M27_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_M20), .B(SubBytesIns_Inst_Sbox_12_M21), .Z(
        SubBytesIns_Inst_Sbox_12_M27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_M28_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_M23), .B(SubBytesIns_Inst_Sbox_12_M25), .Z(
        SubBytesIns_Inst_Sbox_12_M28) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M29_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_M28), .A2(SubBytesIns_Inst_Sbox_12_M27), .ZN(
        SubBytesIns_Inst_Sbox_12_M29) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M30_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_M26), .A2(SubBytesIns_Inst_Sbox_12_M24), .ZN(
        SubBytesIns_Inst_Sbox_12_M30) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M31_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_M20), .A2(SubBytesIns_Inst_Sbox_12_M23), .ZN(
        SubBytesIns_Inst_Sbox_12_M31) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M32_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_M27), .A2(SubBytesIns_Inst_Sbox_12_M31), .ZN(
        SubBytesIns_Inst_Sbox_12_M32) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_M33_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_M27), .B(SubBytesIns_Inst_Sbox_12_M25), .Z(
        SubBytesIns_Inst_Sbox_12_M33) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M34_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_M21), .A2(SubBytesIns_Inst_Sbox_12_M22), .ZN(
        SubBytesIns_Inst_Sbox_12_M34) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M35_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_M24), .A2(SubBytesIns_Inst_Sbox_12_M34), .ZN(
        SubBytesIns_Inst_Sbox_12_M35) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_M36_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_M24), .B(SubBytesIns_Inst_Sbox_12_M25), .Z(
        SubBytesIns_Inst_Sbox_12_M36) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_M37_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_M21), .B(SubBytesIns_Inst_Sbox_12_M29), .Z(
        SubBytesIns_Inst_Sbox_12_M37) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_M38_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_M32), .B(SubBytesIns_Inst_Sbox_12_M33), .Z(
        SubBytesIns_Inst_Sbox_12_M38) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_M39_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_M23), .B(SubBytesIns_Inst_Sbox_12_M30), .Z(
        SubBytesIns_Inst_Sbox_12_M39) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_M40_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_M35), .B(SubBytesIns_Inst_Sbox_12_M36), .Z(
        SubBytesIns_Inst_Sbox_12_M40) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_M41_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_M38), .B(SubBytesIns_Inst_Sbox_12_M40), .Z(
        SubBytesIns_Inst_Sbox_12_M41) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_M42_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_M37), .B(SubBytesIns_Inst_Sbox_12_M39), .Z(
        SubBytesIns_Inst_Sbox_12_M42) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_M43_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_M37), .B(SubBytesIns_Inst_Sbox_12_M38), .Z(
        SubBytesIns_Inst_Sbox_12_M43) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_M44_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_M39), .B(SubBytesIns_Inst_Sbox_12_M40), .Z(
        SubBytesIns_Inst_Sbox_12_M44) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_M45_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_M42), .B(SubBytesIns_Inst_Sbox_12_M41), .Z(
        SubBytesIns_Inst_Sbox_12_M45) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M46_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_M44), .A2(SubBytesIns_Inst_Sbox_12_T6), .ZN(
        SubBytesIns_Inst_Sbox_12_M46) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M47_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_M40), .A2(SubBytesIns_Inst_Sbox_12_T8), .ZN(
        SubBytesIns_Inst_Sbox_12_M47) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M48_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_M39), .A2(SubBytesInput[96]), .ZN(
        SubBytesIns_Inst_Sbox_12_M48) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M49_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_M43), .A2(SubBytesIns_Inst_Sbox_12_T16), .ZN(
        SubBytesIns_Inst_Sbox_12_M49) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M50_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_M38), .A2(SubBytesIns_Inst_Sbox_12_T9), .ZN(
        SubBytesIns_Inst_Sbox_12_M50) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M51_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_M37), .A2(SubBytesIns_Inst_Sbox_12_T17), .ZN(
        SubBytesIns_Inst_Sbox_12_M51) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M52_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_M42), .A2(SubBytesIns_Inst_Sbox_12_T15), .ZN(
        SubBytesIns_Inst_Sbox_12_M52) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M53_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_M45), .A2(SubBytesIns_Inst_Sbox_12_T27), .ZN(
        SubBytesIns_Inst_Sbox_12_M53) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M54_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_M41), .A2(SubBytesIns_Inst_Sbox_12_T10), .ZN(
        SubBytesIns_Inst_Sbox_12_M54) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M55_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_M44), .A2(SubBytesIns_Inst_Sbox_12_T13), .ZN(
        SubBytesIns_Inst_Sbox_12_M55) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M56_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_M40), .A2(SubBytesIns_Inst_Sbox_12_T23), .ZN(
        SubBytesIns_Inst_Sbox_12_M56) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M57_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_M39), .A2(SubBytesIns_Inst_Sbox_12_T19), .ZN(
        SubBytesIns_Inst_Sbox_12_M57) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M58_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_M43), .A2(SubBytesIns_Inst_Sbox_12_T3), .ZN(
        SubBytesIns_Inst_Sbox_12_M58) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M59_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_M38), .A2(SubBytesIns_Inst_Sbox_12_T22), .ZN(
        SubBytesIns_Inst_Sbox_12_M59) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M60_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_M37), .A2(SubBytesIns_Inst_Sbox_12_T20), .ZN(
        SubBytesIns_Inst_Sbox_12_M60) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M61_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_M42), .A2(SubBytesIns_Inst_Sbox_12_T1), .ZN(
        SubBytesIns_Inst_Sbox_12_M61) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M62_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_M45), .A2(SubBytesIns_Inst_Sbox_12_T4), .ZN(
        SubBytesIns_Inst_Sbox_12_M62) );
  AND2_X1 SubBytesIns_Inst_Sbox_12_AND_M63_U1 ( .A1(
        SubBytesIns_Inst_Sbox_12_M41), .A2(SubBytesIns_Inst_Sbox_12_T2), .ZN(
        SubBytesIns_Inst_Sbox_12_M63) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_L0_U1 ( .A(SubBytesIns_Inst_Sbox_12_M61), .B(SubBytesIns_Inst_Sbox_12_M62), .Z(SubBytesIns_Inst_Sbox_12_L0) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_L1_U1 ( .A(SubBytesIns_Inst_Sbox_12_M50), .B(SubBytesIns_Inst_Sbox_12_M56), .Z(SubBytesIns_Inst_Sbox_12_L1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_L2_U1 ( .A(SubBytesIns_Inst_Sbox_12_M46), .B(SubBytesIns_Inst_Sbox_12_M48), .Z(SubBytesIns_Inst_Sbox_12_L2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_L3_U1 ( .A(SubBytesIns_Inst_Sbox_12_M47), .B(SubBytesIns_Inst_Sbox_12_M55), .Z(SubBytesIns_Inst_Sbox_12_L3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_L4_U1 ( .A(SubBytesIns_Inst_Sbox_12_M54), .B(SubBytesIns_Inst_Sbox_12_M58), .Z(SubBytesIns_Inst_Sbox_12_L4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_L5_U1 ( .A(SubBytesIns_Inst_Sbox_12_M49), .B(SubBytesIns_Inst_Sbox_12_M61), .Z(SubBytesIns_Inst_Sbox_12_L5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_L6_U1 ( .A(SubBytesIns_Inst_Sbox_12_M62), .B(SubBytesIns_Inst_Sbox_12_L5), .Z(SubBytesIns_Inst_Sbox_12_L6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_L7_U1 ( .A(SubBytesIns_Inst_Sbox_12_M46), .B(SubBytesIns_Inst_Sbox_12_L3), .Z(SubBytesIns_Inst_Sbox_12_L7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_L8_U1 ( .A(SubBytesIns_Inst_Sbox_12_M51), .B(SubBytesIns_Inst_Sbox_12_M59), .Z(SubBytesIns_Inst_Sbox_12_L8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_L9_U1 ( .A(SubBytesIns_Inst_Sbox_12_M52), .B(SubBytesIns_Inst_Sbox_12_M53), .Z(SubBytesIns_Inst_Sbox_12_L9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_L10_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_M53), .B(SubBytesIns_Inst_Sbox_12_L4), .Z(
        SubBytesIns_Inst_Sbox_12_L10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_L11_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_M60), .B(SubBytesIns_Inst_Sbox_12_L2), .Z(
        SubBytesIns_Inst_Sbox_12_L11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_L12_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_M48), .B(SubBytesIns_Inst_Sbox_12_M51), .Z(
        SubBytesIns_Inst_Sbox_12_L12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_L13_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_M50), .B(SubBytesIns_Inst_Sbox_12_L0), .Z(
        SubBytesIns_Inst_Sbox_12_L13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_L14_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_M52), .B(SubBytesIns_Inst_Sbox_12_M61), .Z(
        SubBytesIns_Inst_Sbox_12_L14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_L15_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_M55), .B(SubBytesIns_Inst_Sbox_12_L1), .Z(
        SubBytesIns_Inst_Sbox_12_L15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_L16_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_M56), .B(SubBytesIns_Inst_Sbox_12_L0), .Z(
        SubBytesIns_Inst_Sbox_12_L16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_L17_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_M57), .B(SubBytesIns_Inst_Sbox_12_L1), .Z(
        SubBytesIns_Inst_Sbox_12_L17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_L18_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_M58), .B(SubBytesIns_Inst_Sbox_12_L8), .Z(
        SubBytesIns_Inst_Sbox_12_L18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_L19_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_M63), .B(SubBytesIns_Inst_Sbox_12_L4), .Z(
        SubBytesIns_Inst_Sbox_12_L19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_L20_U1 ( .A(SubBytesIns_Inst_Sbox_12_L0), .B(SubBytesIns_Inst_Sbox_12_L1), .Z(SubBytesIns_Inst_Sbox_12_L20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_L21_U1 ( .A(SubBytesIns_Inst_Sbox_12_L1), .B(SubBytesIns_Inst_Sbox_12_L7), .Z(SubBytesIns_Inst_Sbox_12_L21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_L22_U1 ( .A(SubBytesIns_Inst_Sbox_12_L3), .B(SubBytesIns_Inst_Sbox_12_L12), .Z(SubBytesIns_Inst_Sbox_12_L22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_L23_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_L18), .B(SubBytesIns_Inst_Sbox_12_L2), .Z(
        SubBytesIns_Inst_Sbox_12_L23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_L24_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_L15), .B(SubBytesIns_Inst_Sbox_12_L9), .Z(
        SubBytesIns_Inst_Sbox_12_L24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_L25_U1 ( .A(SubBytesIns_Inst_Sbox_12_L6), .B(SubBytesIns_Inst_Sbox_12_L10), .Z(SubBytesIns_Inst_Sbox_12_L25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_L26_U1 ( .A(SubBytesIns_Inst_Sbox_12_L7), .B(SubBytesIns_Inst_Sbox_12_L9), .Z(SubBytesIns_Inst_Sbox_12_L26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_L27_U1 ( .A(SubBytesIns_Inst_Sbox_12_L8), .B(SubBytesIns_Inst_Sbox_12_L10), .Z(SubBytesIns_Inst_Sbox_12_L27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_L28_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_L11), .B(SubBytesIns_Inst_Sbox_12_L14), .Z(
        SubBytesIns_Inst_Sbox_12_L28) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_L29_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_L11), .B(SubBytesIns_Inst_Sbox_12_L17), .Z(
        SubBytesIns_Inst_Sbox_12_L29) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_S0_U1 ( .A(SubBytesIns_Inst_Sbox_12_L6), 
        .B(SubBytesIns_Inst_Sbox_12_L24), .Z(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_S1_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_L16), .B(SubBytesIns_Inst_Sbox_12_L26), .ZN(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[7]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_S2_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_L19), .B(SubBytesIns_Inst_Sbox_12_L28), .ZN(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[6]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_S3_U1 ( .A(SubBytesIns_Inst_Sbox_12_L6), 
        .B(SubBytesIns_Inst_Sbox_12_L21), .Z(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[5]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_S4_U1 ( .A(SubBytesIns_Inst_Sbox_12_L20), .B(SubBytesIns_Inst_Sbox_12_L22), .Z(MixColumnsInput[67]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_S5_U1 ( .A(SubBytesIns_Inst_Sbox_12_L25), .B(SubBytesIns_Inst_Sbox_12_L29), .Z(MixColumnsInput[66]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_S6_U1 ( .A(
        SubBytesIns_Inst_Sbox_12_L13), .B(SubBytesIns_Inst_Sbox_12_L27), .ZN(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[2]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_12_XOR_S7_U1 ( .A(SubBytesIns_Inst_Sbox_12_L6), .B(SubBytesIns_Inst_Sbox_12_L23), .ZN(MixColumnsInput[64]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_T1_U1 ( .A(SubBytesInput[111]), .B(
        SubBytesInput[108]), .Z(SubBytesIns_Inst_Sbox_13_T1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_T2_U1 ( .A(SubBytesInput[111]), .B(
        SubBytesInput[106]), .Z(SubBytesIns_Inst_Sbox_13_T2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_T3_U1 ( .A(SubBytesInput[111]), .B(
        SubBytesInput[105]), .Z(SubBytesIns_Inst_Sbox_13_T3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_T4_U1 ( .A(SubBytesInput[108]), .B(
        SubBytesInput[106]), .Z(SubBytesIns_Inst_Sbox_13_T4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_T5_U1 ( .A(SubBytesInput[107]), .B(
        SubBytesInput[105]), .Z(SubBytesIns_Inst_Sbox_13_T5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_T6_U1 ( .A(SubBytesIns_Inst_Sbox_13_T1), 
        .B(SubBytesIns_Inst_Sbox_13_T5), .Z(SubBytesIns_Inst_Sbox_13_T6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_T7_U1 ( .A(SubBytesInput[110]), .B(
        SubBytesInput[109]), .Z(SubBytesIns_Inst_Sbox_13_T7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_T8_U1 ( .A(SubBytesInput[104]), .B(
        SubBytesIns_Inst_Sbox_13_T6), .Z(SubBytesIns_Inst_Sbox_13_T8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_T9_U1 ( .A(SubBytesInput[104]), .B(
        SubBytesIns_Inst_Sbox_13_T7), .Z(SubBytesIns_Inst_Sbox_13_T9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_T10_U1 ( .A(SubBytesIns_Inst_Sbox_13_T6), .B(SubBytesIns_Inst_Sbox_13_T7), .Z(SubBytesIns_Inst_Sbox_13_T10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_T11_U1 ( .A(SubBytesInput[110]), .B(
        SubBytesInput[106]), .Z(SubBytesIns_Inst_Sbox_13_T11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_T12_U1 ( .A(SubBytesInput[109]), .B(
        SubBytesInput[106]), .Z(SubBytesIns_Inst_Sbox_13_T12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_T13_U1 ( .A(SubBytesIns_Inst_Sbox_13_T3), .B(SubBytesIns_Inst_Sbox_13_T4), .Z(SubBytesIns_Inst_Sbox_13_T13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_T14_U1 ( .A(SubBytesIns_Inst_Sbox_13_T6), .B(SubBytesIns_Inst_Sbox_13_T11), .Z(SubBytesIns_Inst_Sbox_13_T14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_T15_U1 ( .A(SubBytesIns_Inst_Sbox_13_T5), .B(SubBytesIns_Inst_Sbox_13_T11), .Z(SubBytesIns_Inst_Sbox_13_T15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_T16_U1 ( .A(SubBytesIns_Inst_Sbox_13_T5), .B(SubBytesIns_Inst_Sbox_13_T12), .Z(SubBytesIns_Inst_Sbox_13_T16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_T17_U1 ( .A(SubBytesIns_Inst_Sbox_13_T9), .B(SubBytesIns_Inst_Sbox_13_T16), .Z(SubBytesIns_Inst_Sbox_13_T17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_T18_U1 ( .A(SubBytesInput[108]), .B(
        SubBytesInput[104]), .Z(SubBytesIns_Inst_Sbox_13_T18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_T19_U1 ( .A(SubBytesIns_Inst_Sbox_13_T7), .B(SubBytesIns_Inst_Sbox_13_T18), .Z(SubBytesIns_Inst_Sbox_13_T19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_T20_U1 ( .A(SubBytesIns_Inst_Sbox_13_T1), .B(SubBytesIns_Inst_Sbox_13_T19), .Z(SubBytesIns_Inst_Sbox_13_T20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_T21_U1 ( .A(SubBytesInput[105]), .B(
        SubBytesInput[104]), .Z(SubBytesIns_Inst_Sbox_13_T21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_T22_U1 ( .A(SubBytesIns_Inst_Sbox_13_T7), .B(SubBytesIns_Inst_Sbox_13_T21), .Z(SubBytesIns_Inst_Sbox_13_T22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_T23_U1 ( .A(SubBytesIns_Inst_Sbox_13_T2), .B(SubBytesIns_Inst_Sbox_13_T22), .Z(SubBytesIns_Inst_Sbox_13_T23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_T24_U1 ( .A(SubBytesIns_Inst_Sbox_13_T2), .B(SubBytesIns_Inst_Sbox_13_T10), .Z(SubBytesIns_Inst_Sbox_13_T24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_T25_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_T20), .B(SubBytesIns_Inst_Sbox_13_T17), .Z(
        SubBytesIns_Inst_Sbox_13_T25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_T26_U1 ( .A(SubBytesIns_Inst_Sbox_13_T3), .B(SubBytesIns_Inst_Sbox_13_T16), .Z(SubBytesIns_Inst_Sbox_13_T26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_T27_U1 ( .A(SubBytesIns_Inst_Sbox_13_T1), .B(SubBytesIns_Inst_Sbox_13_T12), .Z(SubBytesIns_Inst_Sbox_13_T27) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M1_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_T13), .A2(SubBytesIns_Inst_Sbox_13_T6), .ZN(
        SubBytesIns_Inst_Sbox_13_M1) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M2_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_T23), .A2(SubBytesIns_Inst_Sbox_13_T8), .ZN(
        SubBytesIns_Inst_Sbox_13_M2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_M3_U1 ( .A(SubBytesIns_Inst_Sbox_13_T14), .B(SubBytesIns_Inst_Sbox_13_M1), .Z(SubBytesIns_Inst_Sbox_13_M3) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M4_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_T19), .A2(SubBytesInput[104]), .ZN(
        SubBytesIns_Inst_Sbox_13_M4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_M5_U1 ( .A(SubBytesIns_Inst_Sbox_13_M4), 
        .B(SubBytesIns_Inst_Sbox_13_M1), .Z(SubBytesIns_Inst_Sbox_13_M5) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M6_U1 ( .A1(SubBytesIns_Inst_Sbox_13_T3), .A2(SubBytesIns_Inst_Sbox_13_T16), .ZN(SubBytesIns_Inst_Sbox_13_M6) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M7_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_T22), .A2(SubBytesIns_Inst_Sbox_13_T9), .ZN(
        SubBytesIns_Inst_Sbox_13_M7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_M8_U1 ( .A(SubBytesIns_Inst_Sbox_13_T26), .B(SubBytesIns_Inst_Sbox_13_M6), .Z(SubBytesIns_Inst_Sbox_13_M8) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M9_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_T20), .A2(SubBytesIns_Inst_Sbox_13_T17), .ZN(
        SubBytesIns_Inst_Sbox_13_M9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_M10_U1 ( .A(SubBytesIns_Inst_Sbox_13_M9), .B(SubBytesIns_Inst_Sbox_13_M6), .Z(SubBytesIns_Inst_Sbox_13_M10) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M11_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_T1), .A2(SubBytesIns_Inst_Sbox_13_T15), .ZN(
        SubBytesIns_Inst_Sbox_13_M11) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M12_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_T4), .A2(SubBytesIns_Inst_Sbox_13_T27), .ZN(
        SubBytesIns_Inst_Sbox_13_M12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_M13_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_M12), .B(SubBytesIns_Inst_Sbox_13_M11), .Z(
        SubBytesIns_Inst_Sbox_13_M13) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M14_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_T2), .A2(SubBytesIns_Inst_Sbox_13_T10), .ZN(
        SubBytesIns_Inst_Sbox_13_M14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_M15_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_M14), .B(SubBytesIns_Inst_Sbox_13_M11), .Z(
        SubBytesIns_Inst_Sbox_13_M15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_M16_U1 ( .A(SubBytesIns_Inst_Sbox_13_M3), .B(SubBytesIns_Inst_Sbox_13_M2), .Z(SubBytesIns_Inst_Sbox_13_M16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_M17_U1 ( .A(SubBytesIns_Inst_Sbox_13_M5), .B(SubBytesIns_Inst_Sbox_13_T24), .Z(SubBytesIns_Inst_Sbox_13_M17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_M18_U1 ( .A(SubBytesIns_Inst_Sbox_13_M8), .B(SubBytesIns_Inst_Sbox_13_M7), .Z(SubBytesIns_Inst_Sbox_13_M18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_M19_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_M10), .B(SubBytesIns_Inst_Sbox_13_M15), .Z(
        SubBytesIns_Inst_Sbox_13_M19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_M20_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_M16), .B(SubBytesIns_Inst_Sbox_13_M13), .Z(
        SubBytesIns_Inst_Sbox_13_M20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_M21_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_M17), .B(SubBytesIns_Inst_Sbox_13_M15), .Z(
        SubBytesIns_Inst_Sbox_13_M21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_M22_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_M18), .B(SubBytesIns_Inst_Sbox_13_M13), .Z(
        SubBytesIns_Inst_Sbox_13_M22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_M23_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_M19), .B(SubBytesIns_Inst_Sbox_13_T25), .Z(
        SubBytesIns_Inst_Sbox_13_M23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_M24_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_M22), .B(SubBytesIns_Inst_Sbox_13_M23), .Z(
        SubBytesIns_Inst_Sbox_13_M24) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M25_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_M22), .A2(SubBytesIns_Inst_Sbox_13_M20), .ZN(
        SubBytesIns_Inst_Sbox_13_M25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_M26_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_M21), .B(SubBytesIns_Inst_Sbox_13_M25), .Z(
        SubBytesIns_Inst_Sbox_13_M26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_M27_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_M20), .B(SubBytesIns_Inst_Sbox_13_M21), .Z(
        SubBytesIns_Inst_Sbox_13_M27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_M28_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_M23), .B(SubBytesIns_Inst_Sbox_13_M25), .Z(
        SubBytesIns_Inst_Sbox_13_M28) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M29_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_M28), .A2(SubBytesIns_Inst_Sbox_13_M27), .ZN(
        SubBytesIns_Inst_Sbox_13_M29) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M30_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_M26), .A2(SubBytesIns_Inst_Sbox_13_M24), .ZN(
        SubBytesIns_Inst_Sbox_13_M30) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M31_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_M20), .A2(SubBytesIns_Inst_Sbox_13_M23), .ZN(
        SubBytesIns_Inst_Sbox_13_M31) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M32_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_M27), .A2(SubBytesIns_Inst_Sbox_13_M31), .ZN(
        SubBytesIns_Inst_Sbox_13_M32) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_M33_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_M27), .B(SubBytesIns_Inst_Sbox_13_M25), .Z(
        SubBytesIns_Inst_Sbox_13_M33) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M34_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_M21), .A2(SubBytesIns_Inst_Sbox_13_M22), .ZN(
        SubBytesIns_Inst_Sbox_13_M34) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M35_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_M24), .A2(SubBytesIns_Inst_Sbox_13_M34), .ZN(
        SubBytesIns_Inst_Sbox_13_M35) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_M36_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_M24), .B(SubBytesIns_Inst_Sbox_13_M25), .Z(
        SubBytesIns_Inst_Sbox_13_M36) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_M37_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_M21), .B(SubBytesIns_Inst_Sbox_13_M29), .Z(
        SubBytesIns_Inst_Sbox_13_M37) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_M38_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_M32), .B(SubBytesIns_Inst_Sbox_13_M33), .Z(
        SubBytesIns_Inst_Sbox_13_M38) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_M39_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_M23), .B(SubBytesIns_Inst_Sbox_13_M30), .Z(
        SubBytesIns_Inst_Sbox_13_M39) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_M40_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_M35), .B(SubBytesIns_Inst_Sbox_13_M36), .Z(
        SubBytesIns_Inst_Sbox_13_M40) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_M41_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_M38), .B(SubBytesIns_Inst_Sbox_13_M40), .Z(
        SubBytesIns_Inst_Sbox_13_M41) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_M42_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_M37), .B(SubBytesIns_Inst_Sbox_13_M39), .Z(
        SubBytesIns_Inst_Sbox_13_M42) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_M43_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_M37), .B(SubBytesIns_Inst_Sbox_13_M38), .Z(
        SubBytesIns_Inst_Sbox_13_M43) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_M44_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_M39), .B(SubBytesIns_Inst_Sbox_13_M40), .Z(
        SubBytesIns_Inst_Sbox_13_M44) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_M45_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_M42), .B(SubBytesIns_Inst_Sbox_13_M41), .Z(
        SubBytesIns_Inst_Sbox_13_M45) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M46_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_M44), .A2(SubBytesIns_Inst_Sbox_13_T6), .ZN(
        SubBytesIns_Inst_Sbox_13_M46) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M47_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_M40), .A2(SubBytesIns_Inst_Sbox_13_T8), .ZN(
        SubBytesIns_Inst_Sbox_13_M47) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M48_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_M39), .A2(SubBytesInput[104]), .ZN(
        SubBytesIns_Inst_Sbox_13_M48) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M49_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_M43), .A2(SubBytesIns_Inst_Sbox_13_T16), .ZN(
        SubBytesIns_Inst_Sbox_13_M49) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M50_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_M38), .A2(SubBytesIns_Inst_Sbox_13_T9), .ZN(
        SubBytesIns_Inst_Sbox_13_M50) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M51_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_M37), .A2(SubBytesIns_Inst_Sbox_13_T17), .ZN(
        SubBytesIns_Inst_Sbox_13_M51) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M52_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_M42), .A2(SubBytesIns_Inst_Sbox_13_T15), .ZN(
        SubBytesIns_Inst_Sbox_13_M52) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M53_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_M45), .A2(SubBytesIns_Inst_Sbox_13_T27), .ZN(
        SubBytesIns_Inst_Sbox_13_M53) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M54_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_M41), .A2(SubBytesIns_Inst_Sbox_13_T10), .ZN(
        SubBytesIns_Inst_Sbox_13_M54) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M55_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_M44), .A2(SubBytesIns_Inst_Sbox_13_T13), .ZN(
        SubBytesIns_Inst_Sbox_13_M55) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M56_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_M40), .A2(SubBytesIns_Inst_Sbox_13_T23), .ZN(
        SubBytesIns_Inst_Sbox_13_M56) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M57_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_M39), .A2(SubBytesIns_Inst_Sbox_13_T19), .ZN(
        SubBytesIns_Inst_Sbox_13_M57) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M58_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_M43), .A2(SubBytesIns_Inst_Sbox_13_T3), .ZN(
        SubBytesIns_Inst_Sbox_13_M58) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M59_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_M38), .A2(SubBytesIns_Inst_Sbox_13_T22), .ZN(
        SubBytesIns_Inst_Sbox_13_M59) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M60_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_M37), .A2(SubBytesIns_Inst_Sbox_13_T20), .ZN(
        SubBytesIns_Inst_Sbox_13_M60) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M61_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_M42), .A2(SubBytesIns_Inst_Sbox_13_T1), .ZN(
        SubBytesIns_Inst_Sbox_13_M61) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M62_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_M45), .A2(SubBytesIns_Inst_Sbox_13_T4), .ZN(
        SubBytesIns_Inst_Sbox_13_M62) );
  AND2_X1 SubBytesIns_Inst_Sbox_13_AND_M63_U1 ( .A1(
        SubBytesIns_Inst_Sbox_13_M41), .A2(SubBytesIns_Inst_Sbox_13_T2), .ZN(
        SubBytesIns_Inst_Sbox_13_M63) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_L0_U1 ( .A(SubBytesIns_Inst_Sbox_13_M61), .B(SubBytesIns_Inst_Sbox_13_M62), .Z(SubBytesIns_Inst_Sbox_13_L0) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_L1_U1 ( .A(SubBytesIns_Inst_Sbox_13_M50), .B(SubBytesIns_Inst_Sbox_13_M56), .Z(SubBytesIns_Inst_Sbox_13_L1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_L2_U1 ( .A(SubBytesIns_Inst_Sbox_13_M46), .B(SubBytesIns_Inst_Sbox_13_M48), .Z(SubBytesIns_Inst_Sbox_13_L2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_L3_U1 ( .A(SubBytesIns_Inst_Sbox_13_M47), .B(SubBytesIns_Inst_Sbox_13_M55), .Z(SubBytesIns_Inst_Sbox_13_L3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_L4_U1 ( .A(SubBytesIns_Inst_Sbox_13_M54), .B(SubBytesIns_Inst_Sbox_13_M58), .Z(SubBytesIns_Inst_Sbox_13_L4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_L5_U1 ( .A(SubBytesIns_Inst_Sbox_13_M49), .B(SubBytesIns_Inst_Sbox_13_M61), .Z(SubBytesIns_Inst_Sbox_13_L5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_L6_U1 ( .A(SubBytesIns_Inst_Sbox_13_M62), .B(SubBytesIns_Inst_Sbox_13_L5), .Z(SubBytesIns_Inst_Sbox_13_L6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_L7_U1 ( .A(SubBytesIns_Inst_Sbox_13_M46), .B(SubBytesIns_Inst_Sbox_13_L3), .Z(SubBytesIns_Inst_Sbox_13_L7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_L8_U1 ( .A(SubBytesIns_Inst_Sbox_13_M51), .B(SubBytesIns_Inst_Sbox_13_M59), .Z(SubBytesIns_Inst_Sbox_13_L8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_L9_U1 ( .A(SubBytesIns_Inst_Sbox_13_M52), .B(SubBytesIns_Inst_Sbox_13_M53), .Z(SubBytesIns_Inst_Sbox_13_L9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_L10_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_M53), .B(SubBytesIns_Inst_Sbox_13_L4), .Z(
        SubBytesIns_Inst_Sbox_13_L10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_L11_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_M60), .B(SubBytesIns_Inst_Sbox_13_L2), .Z(
        SubBytesIns_Inst_Sbox_13_L11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_L12_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_M48), .B(SubBytesIns_Inst_Sbox_13_M51), .Z(
        SubBytesIns_Inst_Sbox_13_L12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_L13_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_M50), .B(SubBytesIns_Inst_Sbox_13_L0), .Z(
        SubBytesIns_Inst_Sbox_13_L13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_L14_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_M52), .B(SubBytesIns_Inst_Sbox_13_M61), .Z(
        SubBytesIns_Inst_Sbox_13_L14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_L15_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_M55), .B(SubBytesIns_Inst_Sbox_13_L1), .Z(
        SubBytesIns_Inst_Sbox_13_L15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_L16_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_M56), .B(SubBytesIns_Inst_Sbox_13_L0), .Z(
        SubBytesIns_Inst_Sbox_13_L16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_L17_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_M57), .B(SubBytesIns_Inst_Sbox_13_L1), .Z(
        SubBytesIns_Inst_Sbox_13_L17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_L18_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_M58), .B(SubBytesIns_Inst_Sbox_13_L8), .Z(
        SubBytesIns_Inst_Sbox_13_L18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_L19_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_M63), .B(SubBytesIns_Inst_Sbox_13_L4), .Z(
        SubBytesIns_Inst_Sbox_13_L19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_L20_U1 ( .A(SubBytesIns_Inst_Sbox_13_L0), .B(SubBytesIns_Inst_Sbox_13_L1), .Z(SubBytesIns_Inst_Sbox_13_L20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_L21_U1 ( .A(SubBytesIns_Inst_Sbox_13_L1), .B(SubBytesIns_Inst_Sbox_13_L7), .Z(SubBytesIns_Inst_Sbox_13_L21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_L22_U1 ( .A(SubBytesIns_Inst_Sbox_13_L3), .B(SubBytesIns_Inst_Sbox_13_L12), .Z(SubBytesIns_Inst_Sbox_13_L22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_L23_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_L18), .B(SubBytesIns_Inst_Sbox_13_L2), .Z(
        SubBytesIns_Inst_Sbox_13_L23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_L24_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_L15), .B(SubBytesIns_Inst_Sbox_13_L9), .Z(
        SubBytesIns_Inst_Sbox_13_L24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_L25_U1 ( .A(SubBytesIns_Inst_Sbox_13_L6), .B(SubBytesIns_Inst_Sbox_13_L10), .Z(SubBytesIns_Inst_Sbox_13_L25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_L26_U1 ( .A(SubBytesIns_Inst_Sbox_13_L7), .B(SubBytesIns_Inst_Sbox_13_L9), .Z(SubBytesIns_Inst_Sbox_13_L26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_L27_U1 ( .A(SubBytesIns_Inst_Sbox_13_L8), .B(SubBytesIns_Inst_Sbox_13_L10), .Z(SubBytesIns_Inst_Sbox_13_L27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_L28_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_L11), .B(SubBytesIns_Inst_Sbox_13_L14), .Z(
        SubBytesIns_Inst_Sbox_13_L28) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_L29_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_L11), .B(SubBytesIns_Inst_Sbox_13_L17), .Z(
        SubBytesIns_Inst_Sbox_13_L29) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_S0_U1 ( .A(SubBytesIns_Inst_Sbox_13_L6), 
        .B(SubBytesIns_Inst_Sbox_13_L24), .Z(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_S1_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_L16), .B(SubBytesIns_Inst_Sbox_13_L26), .ZN(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[15]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_S2_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_L19), .B(SubBytesIns_Inst_Sbox_13_L28), .ZN(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[14]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_S3_U1 ( .A(SubBytesIns_Inst_Sbox_13_L6), 
        .B(SubBytesIns_Inst_Sbox_13_L21), .Z(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[13]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_S4_U1 ( .A(SubBytesIns_Inst_Sbox_13_L20), .B(SubBytesIns_Inst_Sbox_13_L22), .Z(MixColumnsInput[43]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_S5_U1 ( .A(SubBytesIns_Inst_Sbox_13_L25), .B(SubBytesIns_Inst_Sbox_13_L29), .Z(MixColumnsInput[42]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_S6_U1 ( .A(
        SubBytesIns_Inst_Sbox_13_L13), .B(SubBytesIns_Inst_Sbox_13_L27), .ZN(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[10]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_13_XOR_S7_U1 ( .A(SubBytesIns_Inst_Sbox_13_L6), .B(SubBytesIns_Inst_Sbox_13_L23), .ZN(MixColumnsInput[40]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_T1_U1 ( .A(SubBytesInput[119]), .B(
        SubBytesInput[116]), .Z(SubBytesIns_Inst_Sbox_14_T1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_T2_U1 ( .A(SubBytesInput[119]), .B(
        SubBytesInput[114]), .Z(SubBytesIns_Inst_Sbox_14_T2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_T3_U1 ( .A(SubBytesInput[119]), .B(
        SubBytesInput[113]), .Z(SubBytesIns_Inst_Sbox_14_T3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_T4_U1 ( .A(SubBytesInput[116]), .B(
        SubBytesInput[114]), .Z(SubBytesIns_Inst_Sbox_14_T4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_T5_U1 ( .A(SubBytesInput[115]), .B(
        SubBytesInput[113]), .Z(SubBytesIns_Inst_Sbox_14_T5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_T6_U1 ( .A(SubBytesIns_Inst_Sbox_14_T1), 
        .B(SubBytesIns_Inst_Sbox_14_T5), .Z(SubBytesIns_Inst_Sbox_14_T6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_T7_U1 ( .A(SubBytesInput[118]), .B(
        SubBytesInput[117]), .Z(SubBytesIns_Inst_Sbox_14_T7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_T8_U1 ( .A(SubBytesInput[112]), .B(
        SubBytesIns_Inst_Sbox_14_T6), .Z(SubBytesIns_Inst_Sbox_14_T8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_T9_U1 ( .A(SubBytesInput[112]), .B(
        SubBytesIns_Inst_Sbox_14_T7), .Z(SubBytesIns_Inst_Sbox_14_T9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_T10_U1 ( .A(SubBytesIns_Inst_Sbox_14_T6), .B(SubBytesIns_Inst_Sbox_14_T7), .Z(SubBytesIns_Inst_Sbox_14_T10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_T11_U1 ( .A(SubBytesInput[118]), .B(
        SubBytesInput[114]), .Z(SubBytesIns_Inst_Sbox_14_T11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_T12_U1 ( .A(SubBytesInput[117]), .B(
        SubBytesInput[114]), .Z(SubBytesIns_Inst_Sbox_14_T12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_T13_U1 ( .A(SubBytesIns_Inst_Sbox_14_T3), .B(SubBytesIns_Inst_Sbox_14_T4), .Z(SubBytesIns_Inst_Sbox_14_T13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_T14_U1 ( .A(SubBytesIns_Inst_Sbox_14_T6), .B(SubBytesIns_Inst_Sbox_14_T11), .Z(SubBytesIns_Inst_Sbox_14_T14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_T15_U1 ( .A(SubBytesIns_Inst_Sbox_14_T5), .B(SubBytesIns_Inst_Sbox_14_T11), .Z(SubBytesIns_Inst_Sbox_14_T15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_T16_U1 ( .A(SubBytesIns_Inst_Sbox_14_T5), .B(SubBytesIns_Inst_Sbox_14_T12), .Z(SubBytesIns_Inst_Sbox_14_T16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_T17_U1 ( .A(SubBytesIns_Inst_Sbox_14_T9), .B(SubBytesIns_Inst_Sbox_14_T16), .Z(SubBytesIns_Inst_Sbox_14_T17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_T18_U1 ( .A(SubBytesInput[116]), .B(
        SubBytesInput[112]), .Z(SubBytesIns_Inst_Sbox_14_T18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_T19_U1 ( .A(SubBytesIns_Inst_Sbox_14_T7), .B(SubBytesIns_Inst_Sbox_14_T18), .Z(SubBytesIns_Inst_Sbox_14_T19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_T20_U1 ( .A(SubBytesIns_Inst_Sbox_14_T1), .B(SubBytesIns_Inst_Sbox_14_T19), .Z(SubBytesIns_Inst_Sbox_14_T20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_T21_U1 ( .A(SubBytesInput[113]), .B(
        SubBytesInput[112]), .Z(SubBytesIns_Inst_Sbox_14_T21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_T22_U1 ( .A(SubBytesIns_Inst_Sbox_14_T7), .B(SubBytesIns_Inst_Sbox_14_T21), .Z(SubBytesIns_Inst_Sbox_14_T22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_T23_U1 ( .A(SubBytesIns_Inst_Sbox_14_T2), .B(SubBytesIns_Inst_Sbox_14_T22), .Z(SubBytesIns_Inst_Sbox_14_T23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_T24_U1 ( .A(SubBytesIns_Inst_Sbox_14_T2), .B(SubBytesIns_Inst_Sbox_14_T10), .Z(SubBytesIns_Inst_Sbox_14_T24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_T25_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_T20), .B(SubBytesIns_Inst_Sbox_14_T17), .Z(
        SubBytesIns_Inst_Sbox_14_T25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_T26_U1 ( .A(SubBytesIns_Inst_Sbox_14_T3), .B(SubBytesIns_Inst_Sbox_14_T16), .Z(SubBytesIns_Inst_Sbox_14_T26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_T27_U1 ( .A(SubBytesIns_Inst_Sbox_14_T1), .B(SubBytesIns_Inst_Sbox_14_T12), .Z(SubBytesIns_Inst_Sbox_14_T27) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M1_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_T13), .A2(SubBytesIns_Inst_Sbox_14_T6), .ZN(
        SubBytesIns_Inst_Sbox_14_M1) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M2_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_T23), .A2(SubBytesIns_Inst_Sbox_14_T8), .ZN(
        SubBytesIns_Inst_Sbox_14_M2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_M3_U1 ( .A(SubBytesIns_Inst_Sbox_14_T14), .B(SubBytesIns_Inst_Sbox_14_M1), .Z(SubBytesIns_Inst_Sbox_14_M3) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M4_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_T19), .A2(SubBytesInput[112]), .ZN(
        SubBytesIns_Inst_Sbox_14_M4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_M5_U1 ( .A(SubBytesIns_Inst_Sbox_14_M4), 
        .B(SubBytesIns_Inst_Sbox_14_M1), .Z(SubBytesIns_Inst_Sbox_14_M5) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M6_U1 ( .A1(SubBytesIns_Inst_Sbox_14_T3), .A2(SubBytesIns_Inst_Sbox_14_T16), .ZN(SubBytesIns_Inst_Sbox_14_M6) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M7_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_T22), .A2(SubBytesIns_Inst_Sbox_14_T9), .ZN(
        SubBytesIns_Inst_Sbox_14_M7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_M8_U1 ( .A(SubBytesIns_Inst_Sbox_14_T26), .B(SubBytesIns_Inst_Sbox_14_M6), .Z(SubBytesIns_Inst_Sbox_14_M8) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M9_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_T20), .A2(SubBytesIns_Inst_Sbox_14_T17), .ZN(
        SubBytesIns_Inst_Sbox_14_M9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_M10_U1 ( .A(SubBytesIns_Inst_Sbox_14_M9), .B(SubBytesIns_Inst_Sbox_14_M6), .Z(SubBytesIns_Inst_Sbox_14_M10) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M11_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_T1), .A2(SubBytesIns_Inst_Sbox_14_T15), .ZN(
        SubBytesIns_Inst_Sbox_14_M11) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M12_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_T4), .A2(SubBytesIns_Inst_Sbox_14_T27), .ZN(
        SubBytesIns_Inst_Sbox_14_M12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_M13_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_M12), .B(SubBytesIns_Inst_Sbox_14_M11), .Z(
        SubBytesIns_Inst_Sbox_14_M13) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M14_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_T2), .A2(SubBytesIns_Inst_Sbox_14_T10), .ZN(
        SubBytesIns_Inst_Sbox_14_M14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_M15_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_M14), .B(SubBytesIns_Inst_Sbox_14_M11), .Z(
        SubBytesIns_Inst_Sbox_14_M15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_M16_U1 ( .A(SubBytesIns_Inst_Sbox_14_M3), .B(SubBytesIns_Inst_Sbox_14_M2), .Z(SubBytesIns_Inst_Sbox_14_M16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_M17_U1 ( .A(SubBytesIns_Inst_Sbox_14_M5), .B(SubBytesIns_Inst_Sbox_14_T24), .Z(SubBytesIns_Inst_Sbox_14_M17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_M18_U1 ( .A(SubBytesIns_Inst_Sbox_14_M8), .B(SubBytesIns_Inst_Sbox_14_M7), .Z(SubBytesIns_Inst_Sbox_14_M18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_M19_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_M10), .B(SubBytesIns_Inst_Sbox_14_M15), .Z(
        SubBytesIns_Inst_Sbox_14_M19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_M20_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_M16), .B(SubBytesIns_Inst_Sbox_14_M13), .Z(
        SubBytesIns_Inst_Sbox_14_M20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_M21_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_M17), .B(SubBytesIns_Inst_Sbox_14_M15), .Z(
        SubBytesIns_Inst_Sbox_14_M21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_M22_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_M18), .B(SubBytesIns_Inst_Sbox_14_M13), .Z(
        SubBytesIns_Inst_Sbox_14_M22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_M23_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_M19), .B(SubBytesIns_Inst_Sbox_14_T25), .Z(
        SubBytesIns_Inst_Sbox_14_M23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_M24_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_M22), .B(SubBytesIns_Inst_Sbox_14_M23), .Z(
        SubBytesIns_Inst_Sbox_14_M24) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M25_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_M22), .A2(SubBytesIns_Inst_Sbox_14_M20), .ZN(
        SubBytesIns_Inst_Sbox_14_M25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_M26_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_M21), .B(SubBytesIns_Inst_Sbox_14_M25), .Z(
        SubBytesIns_Inst_Sbox_14_M26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_M27_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_M20), .B(SubBytesIns_Inst_Sbox_14_M21), .Z(
        SubBytesIns_Inst_Sbox_14_M27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_M28_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_M23), .B(SubBytesIns_Inst_Sbox_14_M25), .Z(
        SubBytesIns_Inst_Sbox_14_M28) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M29_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_M28), .A2(SubBytesIns_Inst_Sbox_14_M27), .ZN(
        SubBytesIns_Inst_Sbox_14_M29) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M30_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_M26), .A2(SubBytesIns_Inst_Sbox_14_M24), .ZN(
        SubBytesIns_Inst_Sbox_14_M30) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M31_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_M20), .A2(SubBytesIns_Inst_Sbox_14_M23), .ZN(
        SubBytesIns_Inst_Sbox_14_M31) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M32_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_M27), .A2(SubBytesIns_Inst_Sbox_14_M31), .ZN(
        SubBytesIns_Inst_Sbox_14_M32) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_M33_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_M27), .B(SubBytesIns_Inst_Sbox_14_M25), .Z(
        SubBytesIns_Inst_Sbox_14_M33) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M34_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_M21), .A2(SubBytesIns_Inst_Sbox_14_M22), .ZN(
        SubBytesIns_Inst_Sbox_14_M34) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M35_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_M24), .A2(SubBytesIns_Inst_Sbox_14_M34), .ZN(
        SubBytesIns_Inst_Sbox_14_M35) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_M36_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_M24), .B(SubBytesIns_Inst_Sbox_14_M25), .Z(
        SubBytesIns_Inst_Sbox_14_M36) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_M37_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_M21), .B(SubBytesIns_Inst_Sbox_14_M29), .Z(
        SubBytesIns_Inst_Sbox_14_M37) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_M38_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_M32), .B(SubBytesIns_Inst_Sbox_14_M33), .Z(
        SubBytesIns_Inst_Sbox_14_M38) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_M39_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_M23), .B(SubBytesIns_Inst_Sbox_14_M30), .Z(
        SubBytesIns_Inst_Sbox_14_M39) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_M40_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_M35), .B(SubBytesIns_Inst_Sbox_14_M36), .Z(
        SubBytesIns_Inst_Sbox_14_M40) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_M41_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_M38), .B(SubBytesIns_Inst_Sbox_14_M40), .Z(
        SubBytesIns_Inst_Sbox_14_M41) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_M42_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_M37), .B(SubBytesIns_Inst_Sbox_14_M39), .Z(
        SubBytesIns_Inst_Sbox_14_M42) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_M43_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_M37), .B(SubBytesIns_Inst_Sbox_14_M38), .Z(
        SubBytesIns_Inst_Sbox_14_M43) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_M44_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_M39), .B(SubBytesIns_Inst_Sbox_14_M40), .Z(
        SubBytesIns_Inst_Sbox_14_M44) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_M45_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_M42), .B(SubBytesIns_Inst_Sbox_14_M41), .Z(
        SubBytesIns_Inst_Sbox_14_M45) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M46_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_M44), .A2(SubBytesIns_Inst_Sbox_14_T6), .ZN(
        SubBytesIns_Inst_Sbox_14_M46) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M47_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_M40), .A2(SubBytesIns_Inst_Sbox_14_T8), .ZN(
        SubBytesIns_Inst_Sbox_14_M47) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M48_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_M39), .A2(SubBytesInput[112]), .ZN(
        SubBytesIns_Inst_Sbox_14_M48) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M49_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_M43), .A2(SubBytesIns_Inst_Sbox_14_T16), .ZN(
        SubBytesIns_Inst_Sbox_14_M49) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M50_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_M38), .A2(SubBytesIns_Inst_Sbox_14_T9), .ZN(
        SubBytesIns_Inst_Sbox_14_M50) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M51_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_M37), .A2(SubBytesIns_Inst_Sbox_14_T17), .ZN(
        SubBytesIns_Inst_Sbox_14_M51) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M52_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_M42), .A2(SubBytesIns_Inst_Sbox_14_T15), .ZN(
        SubBytesIns_Inst_Sbox_14_M52) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M53_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_M45), .A2(SubBytesIns_Inst_Sbox_14_T27), .ZN(
        SubBytesIns_Inst_Sbox_14_M53) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M54_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_M41), .A2(SubBytesIns_Inst_Sbox_14_T10), .ZN(
        SubBytesIns_Inst_Sbox_14_M54) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M55_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_M44), .A2(SubBytesIns_Inst_Sbox_14_T13), .ZN(
        SubBytesIns_Inst_Sbox_14_M55) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M56_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_M40), .A2(SubBytesIns_Inst_Sbox_14_T23), .ZN(
        SubBytesIns_Inst_Sbox_14_M56) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M57_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_M39), .A2(SubBytesIns_Inst_Sbox_14_T19), .ZN(
        SubBytesIns_Inst_Sbox_14_M57) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M58_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_M43), .A2(SubBytesIns_Inst_Sbox_14_T3), .ZN(
        SubBytesIns_Inst_Sbox_14_M58) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M59_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_M38), .A2(SubBytesIns_Inst_Sbox_14_T22), .ZN(
        SubBytesIns_Inst_Sbox_14_M59) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M60_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_M37), .A2(SubBytesIns_Inst_Sbox_14_T20), .ZN(
        SubBytesIns_Inst_Sbox_14_M60) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M61_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_M42), .A2(SubBytesIns_Inst_Sbox_14_T1), .ZN(
        SubBytesIns_Inst_Sbox_14_M61) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M62_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_M45), .A2(SubBytesIns_Inst_Sbox_14_T4), .ZN(
        SubBytesIns_Inst_Sbox_14_M62) );
  AND2_X1 SubBytesIns_Inst_Sbox_14_AND_M63_U1 ( .A1(
        SubBytesIns_Inst_Sbox_14_M41), .A2(SubBytesIns_Inst_Sbox_14_T2), .ZN(
        SubBytesIns_Inst_Sbox_14_M63) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_L0_U1 ( .A(SubBytesIns_Inst_Sbox_14_M61), .B(SubBytesIns_Inst_Sbox_14_M62), .Z(SubBytesIns_Inst_Sbox_14_L0) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_L1_U1 ( .A(SubBytesIns_Inst_Sbox_14_M50), .B(SubBytesIns_Inst_Sbox_14_M56), .Z(SubBytesIns_Inst_Sbox_14_L1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_L2_U1 ( .A(SubBytesIns_Inst_Sbox_14_M46), .B(SubBytesIns_Inst_Sbox_14_M48), .Z(SubBytesIns_Inst_Sbox_14_L2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_L3_U1 ( .A(SubBytesIns_Inst_Sbox_14_M47), .B(SubBytesIns_Inst_Sbox_14_M55), .Z(SubBytesIns_Inst_Sbox_14_L3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_L4_U1 ( .A(SubBytesIns_Inst_Sbox_14_M54), .B(SubBytesIns_Inst_Sbox_14_M58), .Z(SubBytesIns_Inst_Sbox_14_L4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_L5_U1 ( .A(SubBytesIns_Inst_Sbox_14_M49), .B(SubBytesIns_Inst_Sbox_14_M61), .Z(SubBytesIns_Inst_Sbox_14_L5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_L6_U1 ( .A(SubBytesIns_Inst_Sbox_14_M62), .B(SubBytesIns_Inst_Sbox_14_L5), .Z(SubBytesIns_Inst_Sbox_14_L6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_L7_U1 ( .A(SubBytesIns_Inst_Sbox_14_M46), .B(SubBytesIns_Inst_Sbox_14_L3), .Z(SubBytesIns_Inst_Sbox_14_L7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_L8_U1 ( .A(SubBytesIns_Inst_Sbox_14_M51), .B(SubBytesIns_Inst_Sbox_14_M59), .Z(SubBytesIns_Inst_Sbox_14_L8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_L9_U1 ( .A(SubBytesIns_Inst_Sbox_14_M52), .B(SubBytesIns_Inst_Sbox_14_M53), .Z(SubBytesIns_Inst_Sbox_14_L9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_L10_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_M53), .B(SubBytesIns_Inst_Sbox_14_L4), .Z(
        SubBytesIns_Inst_Sbox_14_L10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_L11_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_M60), .B(SubBytesIns_Inst_Sbox_14_L2), .Z(
        SubBytesIns_Inst_Sbox_14_L11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_L12_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_M48), .B(SubBytesIns_Inst_Sbox_14_M51), .Z(
        SubBytesIns_Inst_Sbox_14_L12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_L13_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_M50), .B(SubBytesIns_Inst_Sbox_14_L0), .Z(
        SubBytesIns_Inst_Sbox_14_L13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_L14_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_M52), .B(SubBytesIns_Inst_Sbox_14_M61), .Z(
        SubBytesIns_Inst_Sbox_14_L14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_L15_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_M55), .B(SubBytesIns_Inst_Sbox_14_L1), .Z(
        SubBytesIns_Inst_Sbox_14_L15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_L16_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_M56), .B(SubBytesIns_Inst_Sbox_14_L0), .Z(
        SubBytesIns_Inst_Sbox_14_L16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_L17_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_M57), .B(SubBytesIns_Inst_Sbox_14_L1), .Z(
        SubBytesIns_Inst_Sbox_14_L17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_L18_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_M58), .B(SubBytesIns_Inst_Sbox_14_L8), .Z(
        SubBytesIns_Inst_Sbox_14_L18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_L19_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_M63), .B(SubBytesIns_Inst_Sbox_14_L4), .Z(
        SubBytesIns_Inst_Sbox_14_L19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_L20_U1 ( .A(SubBytesIns_Inst_Sbox_14_L0), .B(SubBytesIns_Inst_Sbox_14_L1), .Z(SubBytesIns_Inst_Sbox_14_L20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_L21_U1 ( .A(SubBytesIns_Inst_Sbox_14_L1), .B(SubBytesIns_Inst_Sbox_14_L7), .Z(SubBytesIns_Inst_Sbox_14_L21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_L22_U1 ( .A(SubBytesIns_Inst_Sbox_14_L3), .B(SubBytesIns_Inst_Sbox_14_L12), .Z(SubBytesIns_Inst_Sbox_14_L22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_L23_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_L18), .B(SubBytesIns_Inst_Sbox_14_L2), .Z(
        SubBytesIns_Inst_Sbox_14_L23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_L24_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_L15), .B(SubBytesIns_Inst_Sbox_14_L9), .Z(
        SubBytesIns_Inst_Sbox_14_L24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_L25_U1 ( .A(SubBytesIns_Inst_Sbox_14_L6), .B(SubBytesIns_Inst_Sbox_14_L10), .Z(SubBytesIns_Inst_Sbox_14_L25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_L26_U1 ( .A(SubBytesIns_Inst_Sbox_14_L7), .B(SubBytesIns_Inst_Sbox_14_L9), .Z(SubBytesIns_Inst_Sbox_14_L26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_L27_U1 ( .A(SubBytesIns_Inst_Sbox_14_L8), .B(SubBytesIns_Inst_Sbox_14_L10), .Z(SubBytesIns_Inst_Sbox_14_L27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_L28_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_L11), .B(SubBytesIns_Inst_Sbox_14_L14), .Z(
        SubBytesIns_Inst_Sbox_14_L28) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_L29_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_L11), .B(SubBytesIns_Inst_Sbox_14_L17), .Z(
        SubBytesIns_Inst_Sbox_14_L29) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_S0_U1 ( .A(SubBytesIns_Inst_Sbox_14_L6), 
        .B(SubBytesIns_Inst_Sbox_14_L24), .Z(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_S1_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_L16), .B(SubBytesIns_Inst_Sbox_14_L26), .ZN(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[23]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_S2_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_L19), .B(SubBytesIns_Inst_Sbox_14_L28), .ZN(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[22]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_S3_U1 ( .A(SubBytesIns_Inst_Sbox_14_L6), 
        .B(SubBytesIns_Inst_Sbox_14_L21), .Z(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[21]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_S4_U1 ( .A(SubBytesIns_Inst_Sbox_14_L20), .B(SubBytesIns_Inst_Sbox_14_L22), .Z(MixColumnsInput[19]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_S5_U1 ( .A(SubBytesIns_Inst_Sbox_14_L25), .B(SubBytesIns_Inst_Sbox_14_L29), .Z(MixColumnsInput[18]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_S6_U1 ( .A(
        SubBytesIns_Inst_Sbox_14_L13), .B(SubBytesIns_Inst_Sbox_14_L27), .ZN(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[18]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_14_XOR_S7_U1 ( .A(SubBytesIns_Inst_Sbox_14_L6), .B(SubBytesIns_Inst_Sbox_14_L23), .ZN(MixColumnsInput[16]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_T1_U1 ( .A(port_out[7]), .B(port_out[4]), .Z(SubBytesIns_Inst_Sbox_15_T1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_T2_U1 ( .A(port_out[7]), .B(port_out[2]), .Z(SubBytesIns_Inst_Sbox_15_T2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_T3_U1 ( .A(port_out[7]), .B(port_out[1]), .Z(SubBytesIns_Inst_Sbox_15_T3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_T4_U1 ( .A(port_out[4]), .B(port_out[2]), .Z(SubBytesIns_Inst_Sbox_15_T4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_T5_U1 ( .A(port_out[3]), .B(port_out[1]), .Z(SubBytesIns_Inst_Sbox_15_T5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_T6_U1 ( .A(SubBytesIns_Inst_Sbox_15_T1), 
        .B(SubBytesIns_Inst_Sbox_15_T5), .Z(SubBytesIns_Inst_Sbox_15_T6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_T7_U1 ( .A(port_out[6]), .B(port_out[5]), .Z(SubBytesIns_Inst_Sbox_15_T7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_T8_U1 ( .A(port_out[0]), .B(
        SubBytesIns_Inst_Sbox_15_T6), .Z(SubBytesIns_Inst_Sbox_15_T8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_T9_U1 ( .A(port_out[0]), .B(
        SubBytesIns_Inst_Sbox_15_T7), .Z(SubBytesIns_Inst_Sbox_15_T9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_T10_U1 ( .A(SubBytesIns_Inst_Sbox_15_T6), .B(SubBytesIns_Inst_Sbox_15_T7), .Z(SubBytesIns_Inst_Sbox_15_T10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_T11_U1 ( .A(port_out[6]), .B(
        port_out[2]), .Z(SubBytesIns_Inst_Sbox_15_T11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_T12_U1 ( .A(port_out[5]), .B(
        port_out[2]), .Z(SubBytesIns_Inst_Sbox_15_T12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_T13_U1 ( .A(SubBytesIns_Inst_Sbox_15_T3), .B(SubBytesIns_Inst_Sbox_15_T4), .Z(SubBytesIns_Inst_Sbox_15_T13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_T14_U1 ( .A(SubBytesIns_Inst_Sbox_15_T6), .B(SubBytesIns_Inst_Sbox_15_T11), .Z(SubBytesIns_Inst_Sbox_15_T14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_T15_U1 ( .A(SubBytesIns_Inst_Sbox_15_T5), .B(SubBytesIns_Inst_Sbox_15_T11), .Z(SubBytesIns_Inst_Sbox_15_T15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_T16_U1 ( .A(SubBytesIns_Inst_Sbox_15_T5), .B(SubBytesIns_Inst_Sbox_15_T12), .Z(SubBytesIns_Inst_Sbox_15_T16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_T17_U1 ( .A(SubBytesIns_Inst_Sbox_15_T9), .B(SubBytesIns_Inst_Sbox_15_T16), .Z(SubBytesIns_Inst_Sbox_15_T17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_T18_U1 ( .A(port_out[4]), .B(
        port_out[0]), .Z(SubBytesIns_Inst_Sbox_15_T18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_T19_U1 ( .A(SubBytesIns_Inst_Sbox_15_T7), .B(SubBytesIns_Inst_Sbox_15_T18), .Z(SubBytesIns_Inst_Sbox_15_T19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_T20_U1 ( .A(SubBytesIns_Inst_Sbox_15_T1), .B(SubBytesIns_Inst_Sbox_15_T19), .Z(SubBytesIns_Inst_Sbox_15_T20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_T21_U1 ( .A(port_out[1]), .B(
        port_out[0]), .Z(SubBytesIns_Inst_Sbox_15_T21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_T22_U1 ( .A(SubBytesIns_Inst_Sbox_15_T7), .B(SubBytesIns_Inst_Sbox_15_T21), .Z(SubBytesIns_Inst_Sbox_15_T22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_T23_U1 ( .A(SubBytesIns_Inst_Sbox_15_T2), .B(SubBytesIns_Inst_Sbox_15_T22), .Z(SubBytesIns_Inst_Sbox_15_T23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_T24_U1 ( .A(SubBytesIns_Inst_Sbox_15_T2), .B(SubBytesIns_Inst_Sbox_15_T10), .Z(SubBytesIns_Inst_Sbox_15_T24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_T25_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_T20), .B(SubBytesIns_Inst_Sbox_15_T17), .Z(
        SubBytesIns_Inst_Sbox_15_T25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_T26_U1 ( .A(SubBytesIns_Inst_Sbox_15_T3), .B(SubBytesIns_Inst_Sbox_15_T16), .Z(SubBytesIns_Inst_Sbox_15_T26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_T27_U1 ( .A(SubBytesIns_Inst_Sbox_15_T1), .B(SubBytesIns_Inst_Sbox_15_T12), .Z(SubBytesIns_Inst_Sbox_15_T27) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M1_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_T13), .A2(SubBytesIns_Inst_Sbox_15_T6), .ZN(
        SubBytesIns_Inst_Sbox_15_M1) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M2_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_T23), .A2(SubBytesIns_Inst_Sbox_15_T8), .ZN(
        SubBytesIns_Inst_Sbox_15_M2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_M3_U1 ( .A(SubBytesIns_Inst_Sbox_15_T14), .B(SubBytesIns_Inst_Sbox_15_M1), .Z(SubBytesIns_Inst_Sbox_15_M3) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M4_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_T19), .A2(port_out[0]), .ZN(
        SubBytesIns_Inst_Sbox_15_M4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_M5_U1 ( .A(SubBytesIns_Inst_Sbox_15_M4), 
        .B(SubBytesIns_Inst_Sbox_15_M1), .Z(SubBytesIns_Inst_Sbox_15_M5) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M6_U1 ( .A1(SubBytesIns_Inst_Sbox_15_T3), .A2(SubBytesIns_Inst_Sbox_15_T16), .ZN(SubBytesIns_Inst_Sbox_15_M6) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M7_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_T22), .A2(SubBytesIns_Inst_Sbox_15_T9), .ZN(
        SubBytesIns_Inst_Sbox_15_M7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_M8_U1 ( .A(SubBytesIns_Inst_Sbox_15_T26), .B(SubBytesIns_Inst_Sbox_15_M6), .Z(SubBytesIns_Inst_Sbox_15_M8) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M9_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_T20), .A2(SubBytesIns_Inst_Sbox_15_T17), .ZN(
        SubBytesIns_Inst_Sbox_15_M9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_M10_U1 ( .A(SubBytesIns_Inst_Sbox_15_M9), .B(SubBytesIns_Inst_Sbox_15_M6), .Z(SubBytesIns_Inst_Sbox_15_M10) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M11_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_T1), .A2(SubBytesIns_Inst_Sbox_15_T15), .ZN(
        SubBytesIns_Inst_Sbox_15_M11) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M12_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_T4), .A2(SubBytesIns_Inst_Sbox_15_T27), .ZN(
        SubBytesIns_Inst_Sbox_15_M12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_M13_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_M12), .B(SubBytesIns_Inst_Sbox_15_M11), .Z(
        SubBytesIns_Inst_Sbox_15_M13) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M14_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_T2), .A2(SubBytesIns_Inst_Sbox_15_T10), .ZN(
        SubBytesIns_Inst_Sbox_15_M14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_M15_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_M14), .B(SubBytesIns_Inst_Sbox_15_M11), .Z(
        SubBytesIns_Inst_Sbox_15_M15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_M16_U1 ( .A(SubBytesIns_Inst_Sbox_15_M3), .B(SubBytesIns_Inst_Sbox_15_M2), .Z(SubBytesIns_Inst_Sbox_15_M16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_M17_U1 ( .A(SubBytesIns_Inst_Sbox_15_M5), .B(SubBytesIns_Inst_Sbox_15_T24), .Z(SubBytesIns_Inst_Sbox_15_M17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_M18_U1 ( .A(SubBytesIns_Inst_Sbox_15_M8), .B(SubBytesIns_Inst_Sbox_15_M7), .Z(SubBytesIns_Inst_Sbox_15_M18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_M19_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_M10), .B(SubBytesIns_Inst_Sbox_15_M15), .Z(
        SubBytesIns_Inst_Sbox_15_M19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_M20_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_M16), .B(SubBytesIns_Inst_Sbox_15_M13), .Z(
        SubBytesIns_Inst_Sbox_15_M20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_M21_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_M17), .B(SubBytesIns_Inst_Sbox_15_M15), .Z(
        SubBytesIns_Inst_Sbox_15_M21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_M22_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_M18), .B(SubBytesIns_Inst_Sbox_15_M13), .Z(
        SubBytesIns_Inst_Sbox_15_M22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_M23_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_M19), .B(SubBytesIns_Inst_Sbox_15_T25), .Z(
        SubBytesIns_Inst_Sbox_15_M23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_M24_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_M22), .B(SubBytesIns_Inst_Sbox_15_M23), .Z(
        SubBytesIns_Inst_Sbox_15_M24) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M25_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_M22), .A2(SubBytesIns_Inst_Sbox_15_M20), .ZN(
        SubBytesIns_Inst_Sbox_15_M25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_M26_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_M21), .B(SubBytesIns_Inst_Sbox_15_M25), .Z(
        SubBytesIns_Inst_Sbox_15_M26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_M27_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_M20), .B(SubBytesIns_Inst_Sbox_15_M21), .Z(
        SubBytesIns_Inst_Sbox_15_M27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_M28_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_M23), .B(SubBytesIns_Inst_Sbox_15_M25), .Z(
        SubBytesIns_Inst_Sbox_15_M28) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M29_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_M28), .A2(SubBytesIns_Inst_Sbox_15_M27), .ZN(
        SubBytesIns_Inst_Sbox_15_M29) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M30_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_M26), .A2(SubBytesIns_Inst_Sbox_15_M24), .ZN(
        SubBytesIns_Inst_Sbox_15_M30) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M31_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_M20), .A2(SubBytesIns_Inst_Sbox_15_M23), .ZN(
        SubBytesIns_Inst_Sbox_15_M31) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M32_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_M27), .A2(SubBytesIns_Inst_Sbox_15_M31), .ZN(
        SubBytesIns_Inst_Sbox_15_M32) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_M33_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_M27), .B(SubBytesIns_Inst_Sbox_15_M25), .Z(
        SubBytesIns_Inst_Sbox_15_M33) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M34_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_M21), .A2(SubBytesIns_Inst_Sbox_15_M22), .ZN(
        SubBytesIns_Inst_Sbox_15_M34) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M35_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_M24), .A2(SubBytesIns_Inst_Sbox_15_M34), .ZN(
        SubBytesIns_Inst_Sbox_15_M35) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_M36_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_M24), .B(SubBytesIns_Inst_Sbox_15_M25), .Z(
        SubBytesIns_Inst_Sbox_15_M36) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_M37_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_M21), .B(SubBytesIns_Inst_Sbox_15_M29), .Z(
        SubBytesIns_Inst_Sbox_15_M37) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_M38_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_M32), .B(SubBytesIns_Inst_Sbox_15_M33), .Z(
        SubBytesIns_Inst_Sbox_15_M38) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_M39_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_M23), .B(SubBytesIns_Inst_Sbox_15_M30), .Z(
        SubBytesIns_Inst_Sbox_15_M39) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_M40_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_M35), .B(SubBytesIns_Inst_Sbox_15_M36), .Z(
        SubBytesIns_Inst_Sbox_15_M40) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_M41_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_M38), .B(SubBytesIns_Inst_Sbox_15_M40), .Z(
        SubBytesIns_Inst_Sbox_15_M41) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_M42_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_M37), .B(SubBytesIns_Inst_Sbox_15_M39), .Z(
        SubBytesIns_Inst_Sbox_15_M42) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_M43_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_M37), .B(SubBytesIns_Inst_Sbox_15_M38), .Z(
        SubBytesIns_Inst_Sbox_15_M43) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_M44_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_M39), .B(SubBytesIns_Inst_Sbox_15_M40), .Z(
        SubBytesIns_Inst_Sbox_15_M44) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_M45_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_M42), .B(SubBytesIns_Inst_Sbox_15_M41), .Z(
        SubBytesIns_Inst_Sbox_15_M45) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M46_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_M44), .A2(SubBytesIns_Inst_Sbox_15_T6), .ZN(
        SubBytesIns_Inst_Sbox_15_M46) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M47_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_M40), .A2(SubBytesIns_Inst_Sbox_15_T8), .ZN(
        SubBytesIns_Inst_Sbox_15_M47) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M48_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_M39), .A2(port_out[0]), .ZN(
        SubBytesIns_Inst_Sbox_15_M48) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M49_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_M43), .A2(SubBytesIns_Inst_Sbox_15_T16), .ZN(
        SubBytesIns_Inst_Sbox_15_M49) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M50_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_M38), .A2(SubBytesIns_Inst_Sbox_15_T9), .ZN(
        SubBytesIns_Inst_Sbox_15_M50) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M51_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_M37), .A2(SubBytesIns_Inst_Sbox_15_T17), .ZN(
        SubBytesIns_Inst_Sbox_15_M51) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M52_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_M42), .A2(SubBytesIns_Inst_Sbox_15_T15), .ZN(
        SubBytesIns_Inst_Sbox_15_M52) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M53_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_M45), .A2(SubBytesIns_Inst_Sbox_15_T27), .ZN(
        SubBytesIns_Inst_Sbox_15_M53) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M54_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_M41), .A2(SubBytesIns_Inst_Sbox_15_T10), .ZN(
        SubBytesIns_Inst_Sbox_15_M54) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M55_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_M44), .A2(SubBytesIns_Inst_Sbox_15_T13), .ZN(
        SubBytesIns_Inst_Sbox_15_M55) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M56_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_M40), .A2(SubBytesIns_Inst_Sbox_15_T23), .ZN(
        SubBytesIns_Inst_Sbox_15_M56) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M57_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_M39), .A2(SubBytesIns_Inst_Sbox_15_T19), .ZN(
        SubBytesIns_Inst_Sbox_15_M57) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M58_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_M43), .A2(SubBytesIns_Inst_Sbox_15_T3), .ZN(
        SubBytesIns_Inst_Sbox_15_M58) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M59_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_M38), .A2(SubBytesIns_Inst_Sbox_15_T22), .ZN(
        SubBytesIns_Inst_Sbox_15_M59) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M60_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_M37), .A2(SubBytesIns_Inst_Sbox_15_T20), .ZN(
        SubBytesIns_Inst_Sbox_15_M60) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M61_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_M42), .A2(SubBytesIns_Inst_Sbox_15_T1), .ZN(
        SubBytesIns_Inst_Sbox_15_M61) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M62_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_M45), .A2(SubBytesIns_Inst_Sbox_15_T4), .ZN(
        SubBytesIns_Inst_Sbox_15_M62) );
  AND2_X1 SubBytesIns_Inst_Sbox_15_AND_M63_U1 ( .A1(
        SubBytesIns_Inst_Sbox_15_M41), .A2(SubBytesIns_Inst_Sbox_15_T2), .ZN(
        SubBytesIns_Inst_Sbox_15_M63) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_L0_U1 ( .A(SubBytesIns_Inst_Sbox_15_M61), .B(SubBytesIns_Inst_Sbox_15_M62), .Z(SubBytesIns_Inst_Sbox_15_L0) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_L1_U1 ( .A(SubBytesIns_Inst_Sbox_15_M50), .B(SubBytesIns_Inst_Sbox_15_M56), .Z(SubBytesIns_Inst_Sbox_15_L1) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_L2_U1 ( .A(SubBytesIns_Inst_Sbox_15_M46), .B(SubBytesIns_Inst_Sbox_15_M48), .Z(SubBytesIns_Inst_Sbox_15_L2) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_L3_U1 ( .A(SubBytesIns_Inst_Sbox_15_M47), .B(SubBytesIns_Inst_Sbox_15_M55), .Z(SubBytesIns_Inst_Sbox_15_L3) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_L4_U1 ( .A(SubBytesIns_Inst_Sbox_15_M54), .B(SubBytesIns_Inst_Sbox_15_M58), .Z(SubBytesIns_Inst_Sbox_15_L4) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_L5_U1 ( .A(SubBytesIns_Inst_Sbox_15_M49), .B(SubBytesIns_Inst_Sbox_15_M61), .Z(SubBytesIns_Inst_Sbox_15_L5) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_L6_U1 ( .A(SubBytesIns_Inst_Sbox_15_M62), .B(SubBytesIns_Inst_Sbox_15_L5), .Z(SubBytesIns_Inst_Sbox_15_L6) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_L7_U1 ( .A(SubBytesIns_Inst_Sbox_15_M46), .B(SubBytesIns_Inst_Sbox_15_L3), .Z(SubBytesIns_Inst_Sbox_15_L7) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_L8_U1 ( .A(SubBytesIns_Inst_Sbox_15_M51), .B(SubBytesIns_Inst_Sbox_15_M59), .Z(SubBytesIns_Inst_Sbox_15_L8) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_L9_U1 ( .A(SubBytesIns_Inst_Sbox_15_M52), .B(SubBytesIns_Inst_Sbox_15_M53), .Z(SubBytesIns_Inst_Sbox_15_L9) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_L10_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_M53), .B(SubBytesIns_Inst_Sbox_15_L4), .Z(
        SubBytesIns_Inst_Sbox_15_L10) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_L11_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_M60), .B(SubBytesIns_Inst_Sbox_15_L2), .Z(
        SubBytesIns_Inst_Sbox_15_L11) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_L12_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_M48), .B(SubBytesIns_Inst_Sbox_15_M51), .Z(
        SubBytesIns_Inst_Sbox_15_L12) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_L13_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_M50), .B(SubBytesIns_Inst_Sbox_15_L0), .Z(
        SubBytesIns_Inst_Sbox_15_L13) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_L14_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_M52), .B(SubBytesIns_Inst_Sbox_15_M61), .Z(
        SubBytesIns_Inst_Sbox_15_L14) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_L15_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_M55), .B(SubBytesIns_Inst_Sbox_15_L1), .Z(
        SubBytesIns_Inst_Sbox_15_L15) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_L16_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_M56), .B(SubBytesIns_Inst_Sbox_15_L0), .Z(
        SubBytesIns_Inst_Sbox_15_L16) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_L17_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_M57), .B(SubBytesIns_Inst_Sbox_15_L1), .Z(
        SubBytesIns_Inst_Sbox_15_L17) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_L18_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_M58), .B(SubBytesIns_Inst_Sbox_15_L8), .Z(
        SubBytesIns_Inst_Sbox_15_L18) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_L19_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_M63), .B(SubBytesIns_Inst_Sbox_15_L4), .Z(
        SubBytesIns_Inst_Sbox_15_L19) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_L20_U1 ( .A(SubBytesIns_Inst_Sbox_15_L0), .B(SubBytesIns_Inst_Sbox_15_L1), .Z(SubBytesIns_Inst_Sbox_15_L20) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_L21_U1 ( .A(SubBytesIns_Inst_Sbox_15_L1), .B(SubBytesIns_Inst_Sbox_15_L7), .Z(SubBytesIns_Inst_Sbox_15_L21) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_L22_U1 ( .A(SubBytesIns_Inst_Sbox_15_L3), .B(SubBytesIns_Inst_Sbox_15_L12), .Z(SubBytesIns_Inst_Sbox_15_L22) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_L23_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_L18), .B(SubBytesIns_Inst_Sbox_15_L2), .Z(
        SubBytesIns_Inst_Sbox_15_L23) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_L24_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_L15), .B(SubBytesIns_Inst_Sbox_15_L9), .Z(
        SubBytesIns_Inst_Sbox_15_L24) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_L25_U1 ( .A(SubBytesIns_Inst_Sbox_15_L6), .B(SubBytesIns_Inst_Sbox_15_L10), .Z(SubBytesIns_Inst_Sbox_15_L25) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_L26_U1 ( .A(SubBytesIns_Inst_Sbox_15_L7), .B(SubBytesIns_Inst_Sbox_15_L9), .Z(SubBytesIns_Inst_Sbox_15_L26) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_L27_U1 ( .A(SubBytesIns_Inst_Sbox_15_L8), .B(SubBytesIns_Inst_Sbox_15_L10), .Z(SubBytesIns_Inst_Sbox_15_L27) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_L28_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_L11), .B(SubBytesIns_Inst_Sbox_15_L14), .Z(
        SubBytesIns_Inst_Sbox_15_L28) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_L29_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_L11), .B(SubBytesIns_Inst_Sbox_15_L17), .Z(
        SubBytesIns_Inst_Sbox_15_L29) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_S0_U1 ( .A(SubBytesIns_Inst_Sbox_15_L6), 
        .B(SubBytesIns_Inst_Sbox_15_L24), .Z(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_S1_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_L16), .B(SubBytesIns_Inst_Sbox_15_L26), .ZN(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[31]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_S2_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_L19), .B(SubBytesIns_Inst_Sbox_15_L28), .ZN(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[30]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_S3_U1 ( .A(SubBytesIns_Inst_Sbox_15_L6), 
        .B(SubBytesIns_Inst_Sbox_15_L21), .Z(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[29]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_S4_U1 ( .A(SubBytesIns_Inst_Sbox_15_L20), .B(SubBytesIns_Inst_Sbox_15_L22), .Z(MixColumnsInput[123]) );
  XOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_S5_U1 ( .A(SubBytesIns_Inst_Sbox_15_L25), .B(SubBytesIns_Inst_Sbox_15_L29), .Z(MixColumnsInput[122]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_S6_U1 ( .A(
        SubBytesIns_Inst_Sbox_15_L13), .B(SubBytesIns_Inst_Sbox_15_L27), .ZN(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[26]) );
  XNOR2_X1 SubBytesIns_Inst_Sbox_15_XOR_S7_U1 ( .A(SubBytesIns_Inst_Sbox_15_L6), .B(SubBytesIns_Inst_Sbox_15_L23), .ZN(MixColumnsInput[120]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U96 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n64), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[18]), .ZN(
        MixColumnsOutput[105]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U95 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n63), .B(
        MixColumnsIns_MixOneColumnInst_0_n62), .ZN(
        MixColumnsIns_MixOneColumnInst_0_n64) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U94 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n61), .B(
        MixColumnsIns_MixOneColumnInst_0_n60), .ZN(MixColumnsOutput[104]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U93 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n59), .B(MixColumnsInput[112]), .ZN(
        MixColumnsIns_MixOneColumnInst_0_n61) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U92 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n58), .B(
        MixColumnsIns_MixOneColumnInst_0_n57), .ZN(MixColumnsOutput[103]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U91 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n56), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]), .ZN(
        MixColumnsIns_MixOneColumnInst_0_n58) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U90 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n55), .B(
        MixColumnsIns_MixOneColumnInst_0_n54), .ZN(MixColumnsOutput[102]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U89 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n53), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[15]), .ZN(
        MixColumnsIns_MixOneColumnInst_0_n55) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U88 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n52), .B(
        MixColumnsIns_MixOneColumnInst_0_n51), .ZN(MixColumnsOutput[101]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U87 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n50), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[14]), .ZN(
        MixColumnsIns_MixOneColumnInst_0_n52) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U86 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n49), .B(
        MixColumnsIns_MixOneColumnInst_0_n48), .ZN(MixColumnsOutput[100]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U85 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n47), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[13]), .ZN(
        MixColumnsIns_MixOneColumnInst_0_n49) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U84 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n46), .B(
        MixColumnsIns_MixOneColumnInst_0_n45), .ZN(MixColumnsOutput[99]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U83 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n44), .B(MixColumnsInput[107]), .ZN(
        MixColumnsIns_MixOneColumnInst_0_n46) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U82 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n43), .B(
        MixColumnsIns_MixOneColumnInst_0_n57), .ZN(MixColumnsOutput[127]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_U81 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[31]), .Z(
        MixColumnsIns_MixOneColumnInst_0_n57) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U80 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]), .B(
        MixColumnsIns_MixOneColumnInst_0_n42), .ZN(
        MixColumnsIns_MixOneColumnInst_0_n43) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U79 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n41), .B(
        MixColumnsIns_MixOneColumnInst_0_n54), .ZN(MixColumnsOutput[126]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_U78 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[23]), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[30]), .Z(
        MixColumnsIns_MixOneColumnInst_0_n54) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U77 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[7]), .B(
        MixColumnsIns_MixOneColumnInst_0_n40), .ZN(
        MixColumnsIns_MixOneColumnInst_0_n41) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U76 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n39), .B(
        MixColumnsIns_MixOneColumnInst_0_n38), .ZN(MixColumnsOutput[98]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U75 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n37), .B(MixColumnsInput[106]), .ZN(
        MixColumnsIns_MixOneColumnInst_0_n39) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U74 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n36), .B(
        MixColumnsIns_MixOneColumnInst_0_n51), .ZN(MixColumnsOutput[125]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_U73 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[22]), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[29]), .Z(
        MixColumnsIns_MixOneColumnInst_0_n51) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U72 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[6]), .B(
        MixColumnsIns_MixOneColumnInst_0_n35), .ZN(
        MixColumnsIns_MixOneColumnInst_0_n36) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U71 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n34), .B(
        MixColumnsIns_MixOneColumnInst_0_n48), .ZN(MixColumnsOutput[124]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_U70 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[21]), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[28]), .Z(
        MixColumnsIns_MixOneColumnInst_0_n48) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U69 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[5]), .B(
        MixColumnsIns_MixOneColumnInst_0_n33), .ZN(
        MixColumnsIns_MixOneColumnInst_0_n34) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U68 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n32), .B(
        MixColumnsIns_MixOneColumnInst_0_n45), .ZN(MixColumnsOutput[123]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_U67 ( .A(MixColumnsInput[115]), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[27]), .Z(
        MixColumnsIns_MixOneColumnInst_0_n45) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U66 ( .A(MixColumnsInput[99]), .B(
        MixColumnsIns_MixOneColumnInst_0_n31), .ZN(
        MixColumnsIns_MixOneColumnInst_0_n32) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U65 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n30), .B(
        MixColumnsIns_MixOneColumnInst_0_n38), .ZN(MixColumnsOutput[122]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_U64 ( .A(MixColumnsInput[114]), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[26]), .Z(
        MixColumnsIns_MixOneColumnInst_0_n38) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U63 ( .A(MixColumnsInput[98]), .B(
        MixColumnsIns_MixOneColumnInst_0_n29), .ZN(
        MixColumnsIns_MixOneColumnInst_0_n30) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U62 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n28), .B(
        MixColumnsIns_MixOneColumnInst_0_n27), .ZN(MixColumnsOutput[121]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U61 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[2]), .B(
        MixColumnsIns_MixOneColumnInst_0_n26), .ZN(
        MixColumnsIns_MixOneColumnInst_0_n28) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U60 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n25), .B(
        MixColumnsIns_MixOneColumnInst_0_n24), .ZN(MixColumnsOutput[120]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U59 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n23), .B(MixColumnsInput[96]), .ZN(
        MixColumnsIns_MixOneColumnInst_0_n25) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U58 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n22), .B(
        MixColumnsIns_MixOneColumnInst_0_n42), .ZN(MixColumnsOutput[119]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_U57 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[23]), .Z(
        MixColumnsIns_MixOneColumnInst_0_n42) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U56 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]), .B(
        MixColumnsIns_MixOneColumnInst_0_n21), .ZN(
        MixColumnsIns_MixOneColumnInst_0_n22) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U55 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n20), .B(
        MixColumnsIns_MixOneColumnInst_0_n40), .ZN(MixColumnsOutput[118]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_U54 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[15]), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[22]), .Z(
        MixColumnsIns_MixOneColumnInst_0_n40) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U53 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[31]), .B(
        MixColumnsIns_MixOneColumnInst_0_n19), .ZN(
        MixColumnsIns_MixOneColumnInst_0_n20) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U52 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n18), .B(
        MixColumnsIns_MixOneColumnInst_0_n35), .ZN(MixColumnsOutput[117]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_U51 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[14]), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[21]), .Z(
        MixColumnsIns_MixOneColumnInst_0_n35) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U50 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[30]), .B(
        MixColumnsIns_MixOneColumnInst_0_n17), .ZN(
        MixColumnsIns_MixOneColumnInst_0_n18) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U49 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n16), .B(
        MixColumnsIns_MixOneColumnInst_0_n33), .ZN(MixColumnsOutput[116]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_U48 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[13]), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[20]), .Z(
        MixColumnsIns_MixOneColumnInst_0_n33) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U47 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[29]), .B(
        MixColumnsIns_MixOneColumnInst_0_n15), .ZN(
        MixColumnsIns_MixOneColumnInst_0_n16) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U46 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n14), .B(
        MixColumnsIns_MixOneColumnInst_0_n27), .ZN(MixColumnsOutput[97]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_U45 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[18]), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[25]), .Z(
        MixColumnsIns_MixOneColumnInst_0_n27) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U44 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[10]), .B(
        MixColumnsIns_MixOneColumnInst_0_n62), .ZN(
        MixColumnsIns_MixOneColumnInst_0_n14) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_U43 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[26]), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[1]), .Z(
        MixColumnsIns_MixOneColumnInst_0_n62) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U42 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n13), .B(
        MixColumnsIns_MixOneColumnInst_0_n31), .ZN(MixColumnsOutput[115]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_U41 ( .A(MixColumnsInput[107]), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[19]), .Z(
        MixColumnsIns_MixOneColumnInst_0_n31) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U40 ( .A(MixColumnsInput[123]), 
        .B(MixColumnsIns_MixOneColumnInst_0_n12), .ZN(
        MixColumnsIns_MixOneColumnInst_0_n13) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U39 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n11), .B(
        MixColumnsIns_MixOneColumnInst_0_n29), .ZN(MixColumnsOutput[114]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_U38 ( .A(MixColumnsInput[106]), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[18]), .Z(
        MixColumnsIns_MixOneColumnInst_0_n29) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U37 ( .A(MixColumnsInput[122]), 
        .B(MixColumnsIns_MixOneColumnInst_0_n10), .ZN(
        MixColumnsIns_MixOneColumnInst_0_n11) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U36 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n9), .B(
        MixColumnsIns_MixOneColumnInst_0_n26), .ZN(MixColumnsOutput[113]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_U35 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[17]), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[10]), .Z(
        MixColumnsIns_MixOneColumnInst_0_n26) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U34 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n63), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[26]), .ZN(
        MixColumnsIns_MixOneColumnInst_0_n9) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_U33 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[9]), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[2]), .Z(
        MixColumnsIns_MixOneColumnInst_0_n63) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U32 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n8), .B(
        MixColumnsIns_MixOneColumnInst_0_n24), .ZN(MixColumnsOutput[112]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_U31 ( .A(MixColumnsInput[104]), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]), .Z(
        MixColumnsIns_MixOneColumnInst_0_n24) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U30 ( .A(MixColumnsInput[120]), 
        .B(MixColumnsIns_MixOneColumnInst_0_n60), .ZN(
        MixColumnsIns_MixOneColumnInst_0_n8) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_U29 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]), .B(
        MixColumnsInput[96]), .Z(MixColumnsIns_MixOneColumnInst_0_n60) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U28 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n7), .B(
        MixColumnsIns_MixOneColumnInst_0_n21), .ZN(MixColumnsOutput[111]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_U27 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[15]), .Z(
        MixColumnsIns_MixOneColumnInst_0_n21) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U26 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n56), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]), .ZN(
        MixColumnsIns_MixOneColumnInst_0_n7) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_U25 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[7]), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]), .Z(
        MixColumnsIns_MixOneColumnInst_0_n56) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U24 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n6), .B(
        MixColumnsIns_MixOneColumnInst_0_n19), .ZN(MixColumnsOutput[110]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_U23 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[7]), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[14]), .Z(
        MixColumnsIns_MixOneColumnInst_0_n19) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U22 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n53), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[23]), .ZN(
        MixColumnsIns_MixOneColumnInst_0_n6) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_U21 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[6]), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[31]), .Z(
        MixColumnsIns_MixOneColumnInst_0_n53) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U20 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n5), .B(
        MixColumnsIns_MixOneColumnInst_0_n17), .ZN(MixColumnsOutput[109]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_U19 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[6]), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[13]), .Z(
        MixColumnsIns_MixOneColumnInst_0_n17) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U18 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n50), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[22]), .ZN(
        MixColumnsIns_MixOneColumnInst_0_n5) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_U17 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[5]), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[30]), .Z(
        MixColumnsIns_MixOneColumnInst_0_n50) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U16 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n4), .B(
        MixColumnsIns_MixOneColumnInst_0_n15), .ZN(MixColumnsOutput[108]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_U15 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[5]), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[12]), .Z(
        MixColumnsIns_MixOneColumnInst_0_n15) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U14 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n47), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[21]), .ZN(
        MixColumnsIns_MixOneColumnInst_0_n4) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_U13 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[4]), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[29]), .Z(
        MixColumnsIns_MixOneColumnInst_0_n47) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U12 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n3), .B(
        MixColumnsIns_MixOneColumnInst_0_n12), .ZN(MixColumnsOutput[107]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_U11 ( .A(MixColumnsInput[99]), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[11]), .Z(
        MixColumnsIns_MixOneColumnInst_0_n12) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U10 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n44), .B(MixColumnsInput[115]), .ZN(
        MixColumnsIns_MixOneColumnInst_0_n3) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_U9 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[3]), .B(
        MixColumnsInput[123]), .Z(MixColumnsIns_MixOneColumnInst_0_n44) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U8 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n2), .B(
        MixColumnsIns_MixOneColumnInst_0_n10), .ZN(MixColumnsOutput[106]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_U7 ( .A(MixColumnsInput[98]), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[10]), .Z(
        MixColumnsIns_MixOneColumnInst_0_n10) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U6 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n37), .B(MixColumnsInput[114]), .ZN(
        MixColumnsIns_MixOneColumnInst_0_n2) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_U5 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[2]), .B(
        MixColumnsInput[122]), .Z(MixColumnsIns_MixOneColumnInst_0_n37) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U4 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n1), .B(MixColumnsInput[104]), .ZN(
        MixColumnsOutput[96]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_0_U3 ( .A(
        MixColumnsIns_MixOneColumnInst_0_n59), .B(
        MixColumnsIns_MixOneColumnInst_0_n23), .ZN(
        MixColumnsIns_MixOneColumnInst_0_n1) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_U2 ( .A(MixColumnsInput[112]), .B(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]), .Z(
        MixColumnsIns_MixOneColumnInst_0_n23) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_U1 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]), .B(
        MixColumnsInput[120]), .Z(MixColumnsIns_MixOneColumnInst_0_n59) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_Mul2Inst_0_U3 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]), .B(
        MixColumnsInput[123]), .Z(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[28]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_Mul2Inst_0_U2 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]), .B(
        MixColumnsInput[122]), .Z(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[27]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_Mul2Inst_0_U1 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]), .B(
        MixColumnsInput[120]), .Z(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[25]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_Mul2Inst_1_U3 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]), .B(
        MixColumnsInput[115]), .Z(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[20]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_Mul2Inst_1_U2 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]), .B(
        MixColumnsInput[114]), .Z(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[19]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_Mul2Inst_1_U1 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]), .B(
        MixColumnsInput[112]), .Z(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[17]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_Mul2Inst_2_U3 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]), .B(
        MixColumnsInput[107]), .Z(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[12]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_Mul2Inst_2_U2 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]), .B(
        MixColumnsInput[106]), .Z(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[11]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_Mul2Inst_2_U1 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]), .B(
        MixColumnsInput[104]), .Z(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[9]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_Mul2Inst_3_U3 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]), .B(
        MixColumnsInput[99]), .Z(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[4]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_Mul2Inst_3_U2 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]), .B(
        MixColumnsInput[98]), .Z(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[3]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_0_Mul2Inst_3_U1 ( .A(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]), .B(
        MixColumnsInput[96]), .Z(
        MixColumnsIns_MixOneColumnInst_0_DoubleBytes[1]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U96 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n64), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[18]), .ZN(
        MixColumnsOutput[73]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U95 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n63), .B(
        MixColumnsIns_MixOneColumnInst_1_n62), .ZN(
        MixColumnsIns_MixOneColumnInst_1_n64) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U94 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n61), .B(
        MixColumnsIns_MixOneColumnInst_1_n60), .ZN(MixColumnsOutput[72]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U93 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n59), .B(MixColumnsInput[80]), .ZN(
        MixColumnsIns_MixOneColumnInst_1_n61) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U92 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n58), .B(
        MixColumnsIns_MixOneColumnInst_1_n57), .ZN(MixColumnsOutput[71]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U91 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n56), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]), .ZN(
        MixColumnsIns_MixOneColumnInst_1_n58) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U90 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n55), .B(
        MixColumnsIns_MixOneColumnInst_1_n54), .ZN(MixColumnsOutput[70]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U89 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n53), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[15]), .ZN(
        MixColumnsIns_MixOneColumnInst_1_n55) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U88 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n52), .B(
        MixColumnsIns_MixOneColumnInst_1_n51), .ZN(MixColumnsOutput[69]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U87 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n50), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[14]), .ZN(
        MixColumnsIns_MixOneColumnInst_1_n52) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U86 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n49), .B(
        MixColumnsIns_MixOneColumnInst_1_n48), .ZN(MixColumnsOutput[68]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U85 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n47), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[13]), .ZN(
        MixColumnsIns_MixOneColumnInst_1_n49) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U84 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n46), .B(
        MixColumnsIns_MixOneColumnInst_1_n45), .ZN(MixColumnsOutput[67]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U83 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n44), .B(MixColumnsInput[75]), .ZN(
        MixColumnsIns_MixOneColumnInst_1_n46) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U82 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n43), .B(
        MixColumnsIns_MixOneColumnInst_1_n57), .ZN(MixColumnsOutput[95]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_U81 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[31]), .Z(
        MixColumnsIns_MixOneColumnInst_1_n57) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U80 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]), .B(
        MixColumnsIns_MixOneColumnInst_1_n42), .ZN(
        MixColumnsIns_MixOneColumnInst_1_n43) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U79 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n41), .B(
        MixColumnsIns_MixOneColumnInst_1_n54), .ZN(MixColumnsOutput[94]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_U78 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[23]), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[30]), .Z(
        MixColumnsIns_MixOneColumnInst_1_n54) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U77 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[7]), .B(
        MixColumnsIns_MixOneColumnInst_1_n40), .ZN(
        MixColumnsIns_MixOneColumnInst_1_n41) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U76 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n39), .B(
        MixColumnsIns_MixOneColumnInst_1_n38), .ZN(MixColumnsOutput[66]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U75 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n37), .B(MixColumnsInput[74]), .ZN(
        MixColumnsIns_MixOneColumnInst_1_n39) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U74 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n36), .B(
        MixColumnsIns_MixOneColumnInst_1_n51), .ZN(MixColumnsOutput[93]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_U73 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[22]), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[29]), .Z(
        MixColumnsIns_MixOneColumnInst_1_n51) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U72 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[6]), .B(
        MixColumnsIns_MixOneColumnInst_1_n35), .ZN(
        MixColumnsIns_MixOneColumnInst_1_n36) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U71 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n34), .B(
        MixColumnsIns_MixOneColumnInst_1_n48), .ZN(MixColumnsOutput[92]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_U70 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[21]), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[28]), .Z(
        MixColumnsIns_MixOneColumnInst_1_n48) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U69 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[5]), .B(
        MixColumnsIns_MixOneColumnInst_1_n33), .ZN(
        MixColumnsIns_MixOneColumnInst_1_n34) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U68 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n32), .B(
        MixColumnsIns_MixOneColumnInst_1_n45), .ZN(MixColumnsOutput[91]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_U67 ( .A(MixColumnsInput[83]), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[27]), .Z(
        MixColumnsIns_MixOneColumnInst_1_n45) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U66 ( .A(MixColumnsInput[67]), .B(
        MixColumnsIns_MixOneColumnInst_1_n31), .ZN(
        MixColumnsIns_MixOneColumnInst_1_n32) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U65 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n30), .B(
        MixColumnsIns_MixOneColumnInst_1_n38), .ZN(MixColumnsOutput[90]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_U64 ( .A(MixColumnsInput[82]), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[26]), .Z(
        MixColumnsIns_MixOneColumnInst_1_n38) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U63 ( .A(MixColumnsInput[66]), .B(
        MixColumnsIns_MixOneColumnInst_1_n29), .ZN(
        MixColumnsIns_MixOneColumnInst_1_n30) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U62 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n28), .B(
        MixColumnsIns_MixOneColumnInst_1_n27), .ZN(MixColumnsOutput[89]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U61 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[2]), .B(
        MixColumnsIns_MixOneColumnInst_1_n26), .ZN(
        MixColumnsIns_MixOneColumnInst_1_n28) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U60 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n25), .B(
        MixColumnsIns_MixOneColumnInst_1_n24), .ZN(MixColumnsOutput[88]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U59 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n23), .B(MixColumnsInput[64]), .ZN(
        MixColumnsIns_MixOneColumnInst_1_n25) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U58 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n22), .B(
        MixColumnsIns_MixOneColumnInst_1_n42), .ZN(MixColumnsOutput[87]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_U57 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[23]), .Z(
        MixColumnsIns_MixOneColumnInst_1_n42) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U56 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]), .B(
        MixColumnsIns_MixOneColumnInst_1_n21), .ZN(
        MixColumnsIns_MixOneColumnInst_1_n22) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U55 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n20), .B(
        MixColumnsIns_MixOneColumnInst_1_n40), .ZN(MixColumnsOutput[86]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_U54 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[15]), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[22]), .Z(
        MixColumnsIns_MixOneColumnInst_1_n40) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U53 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[31]), .B(
        MixColumnsIns_MixOneColumnInst_1_n19), .ZN(
        MixColumnsIns_MixOneColumnInst_1_n20) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U52 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n18), .B(
        MixColumnsIns_MixOneColumnInst_1_n35), .ZN(MixColumnsOutput[85]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_U51 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[14]), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[21]), .Z(
        MixColumnsIns_MixOneColumnInst_1_n35) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U50 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[30]), .B(
        MixColumnsIns_MixOneColumnInst_1_n17), .ZN(
        MixColumnsIns_MixOneColumnInst_1_n18) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U49 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n16), .B(
        MixColumnsIns_MixOneColumnInst_1_n33), .ZN(MixColumnsOutput[84]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_U48 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[13]), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[20]), .Z(
        MixColumnsIns_MixOneColumnInst_1_n33) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U47 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[29]), .B(
        MixColumnsIns_MixOneColumnInst_1_n15), .ZN(
        MixColumnsIns_MixOneColumnInst_1_n16) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U46 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n14), .B(
        MixColumnsIns_MixOneColumnInst_1_n27), .ZN(MixColumnsOutput[65]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_U45 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[18]), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[25]), .Z(
        MixColumnsIns_MixOneColumnInst_1_n27) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U44 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[10]), .B(
        MixColumnsIns_MixOneColumnInst_1_n62), .ZN(
        MixColumnsIns_MixOneColumnInst_1_n14) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_U43 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[26]), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[1]), .Z(
        MixColumnsIns_MixOneColumnInst_1_n62) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U42 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n13), .B(
        MixColumnsIns_MixOneColumnInst_1_n31), .ZN(MixColumnsOutput[83]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_U41 ( .A(MixColumnsInput[75]), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[19]), .Z(
        MixColumnsIns_MixOneColumnInst_1_n31) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U40 ( .A(MixColumnsInput[91]), .B(
        MixColumnsIns_MixOneColumnInst_1_n12), .ZN(
        MixColumnsIns_MixOneColumnInst_1_n13) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U39 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n11), .B(
        MixColumnsIns_MixOneColumnInst_1_n29), .ZN(MixColumnsOutput[82]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_U38 ( .A(MixColumnsInput[74]), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[18]), .Z(
        MixColumnsIns_MixOneColumnInst_1_n29) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U37 ( .A(MixColumnsInput[90]), .B(
        MixColumnsIns_MixOneColumnInst_1_n10), .ZN(
        MixColumnsIns_MixOneColumnInst_1_n11) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U36 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n9), .B(
        MixColumnsIns_MixOneColumnInst_1_n26), .ZN(MixColumnsOutput[81]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_U35 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[17]), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[10]), .Z(
        MixColumnsIns_MixOneColumnInst_1_n26) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U34 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n63), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[26]), .ZN(
        MixColumnsIns_MixOneColumnInst_1_n9) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_U33 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[9]), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[2]), .Z(
        MixColumnsIns_MixOneColumnInst_1_n63) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U32 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n8), .B(
        MixColumnsIns_MixOneColumnInst_1_n24), .ZN(MixColumnsOutput[80]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_U31 ( .A(MixColumnsInput[72]), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]), .Z(
        MixColumnsIns_MixOneColumnInst_1_n24) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U30 ( .A(MixColumnsInput[88]), .B(
        MixColumnsIns_MixOneColumnInst_1_n60), .ZN(
        MixColumnsIns_MixOneColumnInst_1_n8) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_U29 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]), .B(
        MixColumnsInput[64]), .Z(MixColumnsIns_MixOneColumnInst_1_n60) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U28 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n7), .B(
        MixColumnsIns_MixOneColumnInst_1_n21), .ZN(MixColumnsOutput[79]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_U27 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[15]), .Z(
        MixColumnsIns_MixOneColumnInst_1_n21) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U26 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n56), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]), .ZN(
        MixColumnsIns_MixOneColumnInst_1_n7) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_U25 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[7]), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]), .Z(
        MixColumnsIns_MixOneColumnInst_1_n56) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U24 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n6), .B(
        MixColumnsIns_MixOneColumnInst_1_n19), .ZN(MixColumnsOutput[78]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_U23 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[7]), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[14]), .Z(
        MixColumnsIns_MixOneColumnInst_1_n19) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U22 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n53), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[23]), .ZN(
        MixColumnsIns_MixOneColumnInst_1_n6) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_U21 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[6]), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[31]), .Z(
        MixColumnsIns_MixOneColumnInst_1_n53) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U20 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n5), .B(
        MixColumnsIns_MixOneColumnInst_1_n17), .ZN(MixColumnsOutput[77]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_U19 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[6]), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[13]), .Z(
        MixColumnsIns_MixOneColumnInst_1_n17) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U18 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n50), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[22]), .ZN(
        MixColumnsIns_MixOneColumnInst_1_n5) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_U17 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[5]), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[30]), .Z(
        MixColumnsIns_MixOneColumnInst_1_n50) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U16 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n4), .B(
        MixColumnsIns_MixOneColumnInst_1_n15), .ZN(MixColumnsOutput[76]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_U15 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[5]), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[12]), .Z(
        MixColumnsIns_MixOneColumnInst_1_n15) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U14 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n47), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[21]), .ZN(
        MixColumnsIns_MixOneColumnInst_1_n4) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_U13 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[4]), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[29]), .Z(
        MixColumnsIns_MixOneColumnInst_1_n47) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U12 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n3), .B(
        MixColumnsIns_MixOneColumnInst_1_n12), .ZN(MixColumnsOutput[75]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_U11 ( .A(MixColumnsInput[67]), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[11]), .Z(
        MixColumnsIns_MixOneColumnInst_1_n12) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U10 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n44), .B(MixColumnsInput[83]), .ZN(
        MixColumnsIns_MixOneColumnInst_1_n3) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_U9 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[3]), .B(
        MixColumnsInput[91]), .Z(MixColumnsIns_MixOneColumnInst_1_n44) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U8 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n2), .B(
        MixColumnsIns_MixOneColumnInst_1_n10), .ZN(MixColumnsOutput[74]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_U7 ( .A(MixColumnsInput[66]), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[10]), .Z(
        MixColumnsIns_MixOneColumnInst_1_n10) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U6 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n37), .B(MixColumnsInput[82]), .ZN(
        MixColumnsIns_MixOneColumnInst_1_n2) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_U5 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[2]), .B(
        MixColumnsInput[90]), .Z(MixColumnsIns_MixOneColumnInst_1_n37) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U4 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n1), .B(MixColumnsInput[72]), .ZN(
        MixColumnsOutput[64]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_1_U3 ( .A(
        MixColumnsIns_MixOneColumnInst_1_n59), .B(
        MixColumnsIns_MixOneColumnInst_1_n23), .ZN(
        MixColumnsIns_MixOneColumnInst_1_n1) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_U2 ( .A(MixColumnsInput[80]), .B(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]), .Z(
        MixColumnsIns_MixOneColumnInst_1_n23) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_U1 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]), .B(
        MixColumnsInput[88]), .Z(MixColumnsIns_MixOneColumnInst_1_n59) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_Mul2Inst_0_U3 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]), .B(
        MixColumnsInput[91]), .Z(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[28]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_Mul2Inst_0_U2 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]), .B(
        MixColumnsInput[90]), .Z(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[27]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_Mul2Inst_0_U1 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]), .B(
        MixColumnsInput[88]), .Z(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[25]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_Mul2Inst_1_U3 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]), .B(
        MixColumnsInput[83]), .Z(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[20]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_Mul2Inst_1_U2 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]), .B(
        MixColumnsInput[82]), .Z(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[19]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_Mul2Inst_1_U1 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]), .B(
        MixColumnsInput[80]), .Z(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[17]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_Mul2Inst_2_U3 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]), .B(
        MixColumnsInput[75]), .Z(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[12]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_Mul2Inst_2_U2 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]), .B(
        MixColumnsInput[74]), .Z(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[11]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_Mul2Inst_2_U1 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]), .B(
        MixColumnsInput[72]), .Z(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[9]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_Mul2Inst_3_U3 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]), .B(
        MixColumnsInput[67]), .Z(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[4]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_Mul2Inst_3_U2 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]), .B(
        MixColumnsInput[66]), .Z(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[3]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_1_Mul2Inst_3_U1 ( .A(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]), .B(
        MixColumnsInput[64]), .Z(
        MixColumnsIns_MixOneColumnInst_1_DoubleBytes[1]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U96 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n64), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[18]), .ZN(
        MixColumnsOutput[41]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U95 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n63), .B(
        MixColumnsIns_MixOneColumnInst_2_n62), .ZN(
        MixColumnsIns_MixOneColumnInst_2_n64) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U94 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n61), .B(
        MixColumnsIns_MixOneColumnInst_2_n60), .ZN(MixColumnsOutput[40]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U93 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n59), .B(MixColumnsInput[48]), .ZN(
        MixColumnsIns_MixOneColumnInst_2_n61) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U92 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n58), .B(
        MixColumnsIns_MixOneColumnInst_2_n57), .ZN(MixColumnsOutput[39]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U91 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n56), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]), .ZN(
        MixColumnsIns_MixOneColumnInst_2_n58) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U90 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n55), .B(
        MixColumnsIns_MixOneColumnInst_2_n54), .ZN(MixColumnsOutput[38]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U89 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n53), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[15]), .ZN(
        MixColumnsIns_MixOneColumnInst_2_n55) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U88 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n52), .B(
        MixColumnsIns_MixOneColumnInst_2_n51), .ZN(MixColumnsOutput[37]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U87 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n50), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[14]), .ZN(
        MixColumnsIns_MixOneColumnInst_2_n52) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U86 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n49), .B(
        MixColumnsIns_MixOneColumnInst_2_n48), .ZN(MixColumnsOutput[36]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U85 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n47), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[13]), .ZN(
        MixColumnsIns_MixOneColumnInst_2_n49) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U84 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n46), .B(
        MixColumnsIns_MixOneColumnInst_2_n45), .ZN(MixColumnsOutput[35]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U83 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n44), .B(MixColumnsInput[43]), .ZN(
        MixColumnsIns_MixOneColumnInst_2_n46) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U82 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n43), .B(
        MixColumnsIns_MixOneColumnInst_2_n57), .ZN(MixColumnsOutput[63]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_U81 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[31]), .Z(
        MixColumnsIns_MixOneColumnInst_2_n57) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U80 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]), .B(
        MixColumnsIns_MixOneColumnInst_2_n42), .ZN(
        MixColumnsIns_MixOneColumnInst_2_n43) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U79 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n41), .B(
        MixColumnsIns_MixOneColumnInst_2_n54), .ZN(MixColumnsOutput[62]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_U78 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[23]), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[30]), .Z(
        MixColumnsIns_MixOneColumnInst_2_n54) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U77 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[7]), .B(
        MixColumnsIns_MixOneColumnInst_2_n40), .ZN(
        MixColumnsIns_MixOneColumnInst_2_n41) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U76 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n39), .B(
        MixColumnsIns_MixOneColumnInst_2_n38), .ZN(MixColumnsOutput[34]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U75 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n37), .B(MixColumnsInput[42]), .ZN(
        MixColumnsIns_MixOneColumnInst_2_n39) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U74 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n36), .B(
        MixColumnsIns_MixOneColumnInst_2_n51), .ZN(MixColumnsOutput[61]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_U73 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[22]), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[29]), .Z(
        MixColumnsIns_MixOneColumnInst_2_n51) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U72 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[6]), .B(
        MixColumnsIns_MixOneColumnInst_2_n35), .ZN(
        MixColumnsIns_MixOneColumnInst_2_n36) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U71 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n34), .B(
        MixColumnsIns_MixOneColumnInst_2_n48), .ZN(MixColumnsOutput[60]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_U70 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[21]), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[28]), .Z(
        MixColumnsIns_MixOneColumnInst_2_n48) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U69 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[5]), .B(
        MixColumnsIns_MixOneColumnInst_2_n33), .ZN(
        MixColumnsIns_MixOneColumnInst_2_n34) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U68 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n32), .B(
        MixColumnsIns_MixOneColumnInst_2_n45), .ZN(MixColumnsOutput[59]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_U67 ( .A(MixColumnsInput[51]), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[27]), .Z(
        MixColumnsIns_MixOneColumnInst_2_n45) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U66 ( .A(MixColumnsInput[35]), .B(
        MixColumnsIns_MixOneColumnInst_2_n31), .ZN(
        MixColumnsIns_MixOneColumnInst_2_n32) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U65 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n30), .B(
        MixColumnsIns_MixOneColumnInst_2_n38), .ZN(MixColumnsOutput[58]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_U64 ( .A(MixColumnsInput[50]), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[26]), .Z(
        MixColumnsIns_MixOneColumnInst_2_n38) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U63 ( .A(MixColumnsInput[34]), .B(
        MixColumnsIns_MixOneColumnInst_2_n29), .ZN(
        MixColumnsIns_MixOneColumnInst_2_n30) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U62 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n28), .B(
        MixColumnsIns_MixOneColumnInst_2_n27), .ZN(MixColumnsOutput[57]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U61 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[2]), .B(
        MixColumnsIns_MixOneColumnInst_2_n26), .ZN(
        MixColumnsIns_MixOneColumnInst_2_n28) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U60 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n25), .B(
        MixColumnsIns_MixOneColumnInst_2_n24), .ZN(MixColumnsOutput[56]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U59 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n23), .B(MixColumnsInput[32]), .ZN(
        MixColumnsIns_MixOneColumnInst_2_n25) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U58 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n22), .B(
        MixColumnsIns_MixOneColumnInst_2_n42), .ZN(MixColumnsOutput[55]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_U57 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[23]), .Z(
        MixColumnsIns_MixOneColumnInst_2_n42) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U56 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]), .B(
        MixColumnsIns_MixOneColumnInst_2_n21), .ZN(
        MixColumnsIns_MixOneColumnInst_2_n22) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U55 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n20), .B(
        MixColumnsIns_MixOneColumnInst_2_n40), .ZN(MixColumnsOutput[54]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_U54 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[15]), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[22]), .Z(
        MixColumnsIns_MixOneColumnInst_2_n40) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U53 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[31]), .B(
        MixColumnsIns_MixOneColumnInst_2_n19), .ZN(
        MixColumnsIns_MixOneColumnInst_2_n20) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U52 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n18), .B(
        MixColumnsIns_MixOneColumnInst_2_n35), .ZN(MixColumnsOutput[53]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_U51 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[14]), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[21]), .Z(
        MixColumnsIns_MixOneColumnInst_2_n35) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U50 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[30]), .B(
        MixColumnsIns_MixOneColumnInst_2_n17), .ZN(
        MixColumnsIns_MixOneColumnInst_2_n18) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U49 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n16), .B(
        MixColumnsIns_MixOneColumnInst_2_n33), .ZN(MixColumnsOutput[52]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_U48 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[13]), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[20]), .Z(
        MixColumnsIns_MixOneColumnInst_2_n33) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U47 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[29]), .B(
        MixColumnsIns_MixOneColumnInst_2_n15), .ZN(
        MixColumnsIns_MixOneColumnInst_2_n16) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U46 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n14), .B(
        MixColumnsIns_MixOneColumnInst_2_n27), .ZN(MixColumnsOutput[33]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_U45 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[18]), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[25]), .Z(
        MixColumnsIns_MixOneColumnInst_2_n27) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U44 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[10]), .B(
        MixColumnsIns_MixOneColumnInst_2_n62), .ZN(
        MixColumnsIns_MixOneColumnInst_2_n14) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_U43 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[26]), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[1]), .Z(
        MixColumnsIns_MixOneColumnInst_2_n62) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U42 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n13), .B(
        MixColumnsIns_MixOneColumnInst_2_n31), .ZN(MixColumnsOutput[51]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_U41 ( .A(MixColumnsInput[43]), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[19]), .Z(
        MixColumnsIns_MixOneColumnInst_2_n31) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U40 ( .A(MixColumnsInput[59]), .B(
        MixColumnsIns_MixOneColumnInst_2_n12), .ZN(
        MixColumnsIns_MixOneColumnInst_2_n13) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U39 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n11), .B(
        MixColumnsIns_MixOneColumnInst_2_n29), .ZN(MixColumnsOutput[50]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_U38 ( .A(MixColumnsInput[42]), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[18]), .Z(
        MixColumnsIns_MixOneColumnInst_2_n29) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U37 ( .A(MixColumnsInput[58]), .B(
        MixColumnsIns_MixOneColumnInst_2_n10), .ZN(
        MixColumnsIns_MixOneColumnInst_2_n11) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U36 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n9), .B(
        MixColumnsIns_MixOneColumnInst_2_n26), .ZN(MixColumnsOutput[49]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_U35 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[17]), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[10]), .Z(
        MixColumnsIns_MixOneColumnInst_2_n26) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U34 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n63), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[26]), .ZN(
        MixColumnsIns_MixOneColumnInst_2_n9) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_U33 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[9]), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[2]), .Z(
        MixColumnsIns_MixOneColumnInst_2_n63) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U32 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n8), .B(
        MixColumnsIns_MixOneColumnInst_2_n24), .ZN(MixColumnsOutput[48]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_U31 ( .A(MixColumnsInput[40]), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]), .Z(
        MixColumnsIns_MixOneColumnInst_2_n24) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U30 ( .A(MixColumnsInput[56]), .B(
        MixColumnsIns_MixOneColumnInst_2_n60), .ZN(
        MixColumnsIns_MixOneColumnInst_2_n8) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_U29 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]), .B(
        MixColumnsInput[32]), .Z(MixColumnsIns_MixOneColumnInst_2_n60) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U28 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n7), .B(
        MixColumnsIns_MixOneColumnInst_2_n21), .ZN(MixColumnsOutput[47]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_U27 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[15]), .Z(
        MixColumnsIns_MixOneColumnInst_2_n21) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U26 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n56), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]), .ZN(
        MixColumnsIns_MixOneColumnInst_2_n7) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_U25 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[7]), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]), .Z(
        MixColumnsIns_MixOneColumnInst_2_n56) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U24 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n6), .B(
        MixColumnsIns_MixOneColumnInst_2_n19), .ZN(MixColumnsOutput[46]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_U23 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[7]), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[14]), .Z(
        MixColumnsIns_MixOneColumnInst_2_n19) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U22 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n53), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[23]), .ZN(
        MixColumnsIns_MixOneColumnInst_2_n6) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_U21 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[6]), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[31]), .Z(
        MixColumnsIns_MixOneColumnInst_2_n53) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U20 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n5), .B(
        MixColumnsIns_MixOneColumnInst_2_n17), .ZN(MixColumnsOutput[45]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_U19 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[6]), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[13]), .Z(
        MixColumnsIns_MixOneColumnInst_2_n17) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U18 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n50), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[22]), .ZN(
        MixColumnsIns_MixOneColumnInst_2_n5) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_U17 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[5]), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[30]), .Z(
        MixColumnsIns_MixOneColumnInst_2_n50) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U16 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n4), .B(
        MixColumnsIns_MixOneColumnInst_2_n15), .ZN(MixColumnsOutput[44]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_U15 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[5]), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[12]), .Z(
        MixColumnsIns_MixOneColumnInst_2_n15) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U14 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n47), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[21]), .ZN(
        MixColumnsIns_MixOneColumnInst_2_n4) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_U13 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[4]), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[29]), .Z(
        MixColumnsIns_MixOneColumnInst_2_n47) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U12 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n3), .B(
        MixColumnsIns_MixOneColumnInst_2_n12), .ZN(MixColumnsOutput[43]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_U11 ( .A(MixColumnsInput[35]), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[11]), .Z(
        MixColumnsIns_MixOneColumnInst_2_n12) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U10 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n44), .B(MixColumnsInput[51]), .ZN(
        MixColumnsIns_MixOneColumnInst_2_n3) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_U9 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[3]), .B(
        MixColumnsInput[59]), .Z(MixColumnsIns_MixOneColumnInst_2_n44) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U8 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n2), .B(
        MixColumnsIns_MixOneColumnInst_2_n10), .ZN(MixColumnsOutput[42]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_U7 ( .A(MixColumnsInput[34]), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[10]), .Z(
        MixColumnsIns_MixOneColumnInst_2_n10) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U6 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n37), .B(MixColumnsInput[50]), .ZN(
        MixColumnsIns_MixOneColumnInst_2_n2) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_U5 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[2]), .B(
        MixColumnsInput[58]), .Z(MixColumnsIns_MixOneColumnInst_2_n37) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U4 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n1), .B(MixColumnsInput[40]), .ZN(
        MixColumnsOutput[32]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_2_U3 ( .A(
        MixColumnsIns_MixOneColumnInst_2_n59), .B(
        MixColumnsIns_MixOneColumnInst_2_n23), .ZN(
        MixColumnsIns_MixOneColumnInst_2_n1) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_U2 ( .A(MixColumnsInput[48]), .B(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]), .Z(
        MixColumnsIns_MixOneColumnInst_2_n23) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_U1 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]), .B(
        MixColumnsInput[56]), .Z(MixColumnsIns_MixOneColumnInst_2_n59) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_Mul2Inst_0_U3 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]), .B(
        MixColumnsInput[59]), .Z(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[28]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_Mul2Inst_0_U2 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]), .B(
        MixColumnsInput[58]), .Z(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[27]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_Mul2Inst_0_U1 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]), .B(
        MixColumnsInput[56]), .Z(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[25]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_Mul2Inst_1_U3 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]), .B(
        MixColumnsInput[51]), .Z(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[20]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_Mul2Inst_1_U2 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]), .B(
        MixColumnsInput[50]), .Z(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[19]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_Mul2Inst_1_U1 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]), .B(
        MixColumnsInput[48]), .Z(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[17]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_Mul2Inst_2_U3 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]), .B(
        MixColumnsInput[43]), .Z(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[12]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_Mul2Inst_2_U2 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]), .B(
        MixColumnsInput[42]), .Z(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[11]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_Mul2Inst_2_U1 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]), .B(
        MixColumnsInput[40]), .Z(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[9]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_Mul2Inst_3_U3 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]), .B(
        MixColumnsInput[35]), .Z(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[4]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_Mul2Inst_3_U2 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]), .B(
        MixColumnsInput[34]), .Z(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[3]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_2_Mul2Inst_3_U1 ( .A(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]), .B(
        MixColumnsInput[32]), .Z(
        MixColumnsIns_MixOneColumnInst_2_DoubleBytes[1]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U96 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n64), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[18]), .ZN(
        MixColumnsOutput[9]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U95 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n63), .B(
        MixColumnsIns_MixOneColumnInst_3_n62), .ZN(
        MixColumnsIns_MixOneColumnInst_3_n64) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U94 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n61), .B(
        MixColumnsIns_MixOneColumnInst_3_n60), .ZN(MixColumnsOutput[8]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U93 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n59), .B(MixColumnsInput[16]), .ZN(
        MixColumnsIns_MixOneColumnInst_3_n61) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U92 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n58), .B(
        MixColumnsIns_MixOneColumnInst_3_n57), .ZN(MixColumnsOutput[7]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U91 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n56), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]), .ZN(
        MixColumnsIns_MixOneColumnInst_3_n58) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U90 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n55), .B(
        MixColumnsIns_MixOneColumnInst_3_n54), .ZN(MixColumnsOutput[6]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U89 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n53), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[15]), .ZN(
        MixColumnsIns_MixOneColumnInst_3_n55) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U88 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n52), .B(
        MixColumnsIns_MixOneColumnInst_3_n51), .ZN(MixColumnsOutput[5]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U87 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n50), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[14]), .ZN(
        MixColumnsIns_MixOneColumnInst_3_n52) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U86 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n49), .B(
        MixColumnsIns_MixOneColumnInst_3_n48), .ZN(MixColumnsOutput[4]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U85 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n47), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[13]), .ZN(
        MixColumnsIns_MixOneColumnInst_3_n49) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U84 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n46), .B(
        MixColumnsIns_MixOneColumnInst_3_n45), .ZN(MixColumnsOutput[3]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U83 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n44), .B(MixColumnsInput[11]), .ZN(
        MixColumnsIns_MixOneColumnInst_3_n46) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U82 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n43), .B(
        MixColumnsIns_MixOneColumnInst_3_n57), .ZN(MixColumnsOutput[31]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_U81 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[31]), .Z(
        MixColumnsIns_MixOneColumnInst_3_n57) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U80 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]), .B(
        MixColumnsIns_MixOneColumnInst_3_n42), .ZN(
        MixColumnsIns_MixOneColumnInst_3_n43) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U79 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n41), .B(
        MixColumnsIns_MixOneColumnInst_3_n54), .ZN(MixColumnsOutput[30]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_U78 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[23]), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[30]), .Z(
        MixColumnsIns_MixOneColumnInst_3_n54) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U77 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[7]), .B(
        MixColumnsIns_MixOneColumnInst_3_n40), .ZN(
        MixColumnsIns_MixOneColumnInst_3_n41) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U76 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n39), .B(
        MixColumnsIns_MixOneColumnInst_3_n38), .ZN(MixColumnsOutput[2]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U75 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n37), .B(MixColumnsInput[10]), .ZN(
        MixColumnsIns_MixOneColumnInst_3_n39) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U74 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n36), .B(
        MixColumnsIns_MixOneColumnInst_3_n51), .ZN(MixColumnsOutput[29]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_U73 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[22]), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[29]), .Z(
        MixColumnsIns_MixOneColumnInst_3_n51) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U72 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[6]), .B(
        MixColumnsIns_MixOneColumnInst_3_n35), .ZN(
        MixColumnsIns_MixOneColumnInst_3_n36) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U71 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n34), .B(
        MixColumnsIns_MixOneColumnInst_3_n48), .ZN(MixColumnsOutput[28]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_U70 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[21]), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[28]), .Z(
        MixColumnsIns_MixOneColumnInst_3_n48) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U69 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[5]), .B(
        MixColumnsIns_MixOneColumnInst_3_n33), .ZN(
        MixColumnsIns_MixOneColumnInst_3_n34) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U68 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n32), .B(
        MixColumnsIns_MixOneColumnInst_3_n45), .ZN(MixColumnsOutput[27]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_U67 ( .A(MixColumnsInput[19]), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[27]), .Z(
        MixColumnsIns_MixOneColumnInst_3_n45) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U66 ( .A(MixColumnsInput[3]), .B(
        MixColumnsIns_MixOneColumnInst_3_n31), .ZN(
        MixColumnsIns_MixOneColumnInst_3_n32) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U65 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n30), .B(
        MixColumnsIns_MixOneColumnInst_3_n38), .ZN(MixColumnsOutput[26]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_U64 ( .A(MixColumnsInput[18]), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[26]), .Z(
        MixColumnsIns_MixOneColumnInst_3_n38) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U63 ( .A(MixColumnsInput[2]), .B(
        MixColumnsIns_MixOneColumnInst_3_n29), .ZN(
        MixColumnsIns_MixOneColumnInst_3_n30) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U62 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n28), .B(
        MixColumnsIns_MixOneColumnInst_3_n27), .ZN(MixColumnsOutput[25]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U61 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[2]), .B(
        MixColumnsIns_MixOneColumnInst_3_n26), .ZN(
        MixColumnsIns_MixOneColumnInst_3_n28) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U60 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n25), .B(
        MixColumnsIns_MixOneColumnInst_3_n24), .ZN(MixColumnsOutput[24]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U59 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n23), .B(MixColumnsInput[0]), .ZN(
        MixColumnsIns_MixOneColumnInst_3_n25) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U58 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n22), .B(
        MixColumnsIns_MixOneColumnInst_3_n42), .ZN(MixColumnsOutput[23]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_U57 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[23]), .Z(
        MixColumnsIns_MixOneColumnInst_3_n42) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U56 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]), .B(
        MixColumnsIns_MixOneColumnInst_3_n21), .ZN(
        MixColumnsIns_MixOneColumnInst_3_n22) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U55 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n20), .B(
        MixColumnsIns_MixOneColumnInst_3_n40), .ZN(MixColumnsOutput[22]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_U54 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[15]), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[22]), .Z(
        MixColumnsIns_MixOneColumnInst_3_n40) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U53 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[31]), .B(
        MixColumnsIns_MixOneColumnInst_3_n19), .ZN(
        MixColumnsIns_MixOneColumnInst_3_n20) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U52 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n18), .B(
        MixColumnsIns_MixOneColumnInst_3_n35), .ZN(MixColumnsOutput[21]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_U51 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[14]), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[21]), .Z(
        MixColumnsIns_MixOneColumnInst_3_n35) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U50 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[30]), .B(
        MixColumnsIns_MixOneColumnInst_3_n17), .ZN(
        MixColumnsIns_MixOneColumnInst_3_n18) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U49 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n16), .B(
        MixColumnsIns_MixOneColumnInst_3_n33), .ZN(MixColumnsOutput[20]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_U48 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[13]), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[20]), .Z(
        MixColumnsIns_MixOneColumnInst_3_n33) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U47 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[29]), .B(
        MixColumnsIns_MixOneColumnInst_3_n15), .ZN(
        MixColumnsIns_MixOneColumnInst_3_n16) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U46 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n14), .B(
        MixColumnsIns_MixOneColumnInst_3_n27), .ZN(MixColumnsOutput[1]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_U45 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[18]), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[25]), .Z(
        MixColumnsIns_MixOneColumnInst_3_n27) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U44 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[10]), .B(
        MixColumnsIns_MixOneColumnInst_3_n62), .ZN(
        MixColumnsIns_MixOneColumnInst_3_n14) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_U43 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[26]), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[1]), .Z(
        MixColumnsIns_MixOneColumnInst_3_n62) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U42 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n13), .B(
        MixColumnsIns_MixOneColumnInst_3_n31), .ZN(MixColumnsOutput[19]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_U41 ( .A(MixColumnsInput[11]), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[19]), .Z(
        MixColumnsIns_MixOneColumnInst_3_n31) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U40 ( .A(MixColumnsInput[27]), .B(
        MixColumnsIns_MixOneColumnInst_3_n12), .ZN(
        MixColumnsIns_MixOneColumnInst_3_n13) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U39 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n11), .B(
        MixColumnsIns_MixOneColumnInst_3_n29), .ZN(MixColumnsOutput[18]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_U38 ( .A(MixColumnsInput[10]), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[18]), .Z(
        MixColumnsIns_MixOneColumnInst_3_n29) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U37 ( .A(MixColumnsInput[26]), .B(
        MixColumnsIns_MixOneColumnInst_3_n10), .ZN(
        MixColumnsIns_MixOneColumnInst_3_n11) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U36 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n9), .B(
        MixColumnsIns_MixOneColumnInst_3_n26), .ZN(MixColumnsOutput[17]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_U35 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[17]), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[10]), .Z(
        MixColumnsIns_MixOneColumnInst_3_n26) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U34 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n63), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[26]), .ZN(
        MixColumnsIns_MixOneColumnInst_3_n9) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_U33 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[9]), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[2]), .Z(
        MixColumnsIns_MixOneColumnInst_3_n63) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U32 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n8), .B(
        MixColumnsIns_MixOneColumnInst_3_n24), .ZN(MixColumnsOutput[16]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_U31 ( .A(MixColumnsInput[8]), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]), .Z(
        MixColumnsIns_MixOneColumnInst_3_n24) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U30 ( .A(MixColumnsInput[24]), .B(
        MixColumnsIns_MixOneColumnInst_3_n60), .ZN(
        MixColumnsIns_MixOneColumnInst_3_n8) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_U29 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]), .B(
        MixColumnsInput[0]), .Z(MixColumnsIns_MixOneColumnInst_3_n60) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U28 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n7), .B(
        MixColumnsIns_MixOneColumnInst_3_n21), .ZN(MixColumnsOutput[15]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_U27 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[15]), .Z(
        MixColumnsIns_MixOneColumnInst_3_n21) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U26 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n56), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]), .ZN(
        MixColumnsIns_MixOneColumnInst_3_n7) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_U25 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[7]), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]), .Z(
        MixColumnsIns_MixOneColumnInst_3_n56) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U24 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n6), .B(
        MixColumnsIns_MixOneColumnInst_3_n19), .ZN(MixColumnsOutput[14]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_U23 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[7]), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[14]), .Z(
        MixColumnsIns_MixOneColumnInst_3_n19) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U22 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n53), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[23]), .ZN(
        MixColumnsIns_MixOneColumnInst_3_n6) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_U21 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[6]), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[31]), .Z(
        MixColumnsIns_MixOneColumnInst_3_n53) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U20 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n5), .B(
        MixColumnsIns_MixOneColumnInst_3_n17), .ZN(MixColumnsOutput[13]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_U19 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[6]), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[13]), .Z(
        MixColumnsIns_MixOneColumnInst_3_n17) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U18 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n50), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[22]), .ZN(
        MixColumnsIns_MixOneColumnInst_3_n5) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_U17 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[5]), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[30]), .Z(
        MixColumnsIns_MixOneColumnInst_3_n50) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U16 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n4), .B(
        MixColumnsIns_MixOneColumnInst_3_n15), .ZN(MixColumnsOutput[12]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_U15 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[5]), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[12]), .Z(
        MixColumnsIns_MixOneColumnInst_3_n15) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U14 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n47), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[21]), .ZN(
        MixColumnsIns_MixOneColumnInst_3_n4) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_U13 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[4]), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[29]), .Z(
        MixColumnsIns_MixOneColumnInst_3_n47) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U12 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n3), .B(
        MixColumnsIns_MixOneColumnInst_3_n12), .ZN(MixColumnsOutput[11]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_U11 ( .A(MixColumnsInput[3]), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[11]), .Z(
        MixColumnsIns_MixOneColumnInst_3_n12) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U10 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n44), .B(MixColumnsInput[19]), .ZN(
        MixColumnsIns_MixOneColumnInst_3_n3) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_U9 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[3]), .B(
        MixColumnsInput[27]), .Z(MixColumnsIns_MixOneColumnInst_3_n44) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U8 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n2), .B(
        MixColumnsIns_MixOneColumnInst_3_n10), .ZN(MixColumnsOutput[10]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_U7 ( .A(MixColumnsInput[2]), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[10]), .Z(
        MixColumnsIns_MixOneColumnInst_3_n10) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U6 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n37), .B(MixColumnsInput[18]), .ZN(
        MixColumnsIns_MixOneColumnInst_3_n2) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_U5 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[2]), .B(
        MixColumnsInput[26]), .Z(MixColumnsIns_MixOneColumnInst_3_n37) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U4 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n1), .B(MixColumnsInput[8]), .ZN(
        MixColumnsOutput[0]) );
  XNOR2_X1 MixColumnsIns_MixOneColumnInst_3_U3 ( .A(
        MixColumnsIns_MixOneColumnInst_3_n59), .B(
        MixColumnsIns_MixOneColumnInst_3_n23), .ZN(
        MixColumnsIns_MixOneColumnInst_3_n1) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_U2 ( .A(MixColumnsInput[16]), .B(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]), .Z(
        MixColumnsIns_MixOneColumnInst_3_n23) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_U1 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]), .B(
        MixColumnsInput[24]), .Z(MixColumnsIns_MixOneColumnInst_3_n59) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_Mul2Inst_0_U3 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]), .B(
        MixColumnsInput[27]), .Z(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[28]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_Mul2Inst_0_U2 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]), .B(
        MixColumnsInput[26]), .Z(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[27]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_Mul2Inst_0_U1 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]), .B(
        MixColumnsInput[24]), .Z(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[25]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_Mul2Inst_1_U3 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]), .B(
        MixColumnsInput[19]), .Z(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[20]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_Mul2Inst_1_U2 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]), .B(
        MixColumnsInput[18]), .Z(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[19]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_Mul2Inst_1_U1 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]), .B(
        MixColumnsInput[16]), .Z(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[17]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_Mul2Inst_2_U3 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]), .B(
        MixColumnsInput[11]), .Z(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[12]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_Mul2Inst_2_U2 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]), .B(
        MixColumnsInput[10]), .Z(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[11]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_Mul2Inst_2_U1 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]), .B(
        MixColumnsInput[8]), .Z(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[9]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_Mul2Inst_3_U3 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]), .B(
        MixColumnsInput[3]), .Z(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[4]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_Mul2Inst_3_U2 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]), .B(
        MixColumnsInput[2]), .Z(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[3]) );
  XOR2_X1 MixColumnsIns_MixOneColumnInst_3_Mul2Inst_3_U1 ( .A(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]), .B(
        MixColumnsInput[0]), .Z(
        MixColumnsIns_MixOneColumnInst_3_DoubleBytes[1]) );
  INV_X1 KeyReg_U5 ( .A(start_done), .ZN(KeyReg_n10) );
  INV_X1 KeyReg_U4 ( .A(KeyReg_n10), .ZN(KeyReg_n9) );
  INV_X1 KeyReg_U3 ( .A(KeyReg_n10), .ZN(KeyReg_n8) );
  INV_X1 KeyReg_U2 ( .A(KeyReg_n10), .ZN(KeyReg_n7) );
  INV_X1 KeyReg_U1 ( .A(KeyReg_n10), .ZN(KeyReg_n6) );
  XOR2_X1 KeyReg_Inst_ff_SDE_0_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[0]), 
        .B(RoundInput[120]), .Z(KeyReg_Inst_ff_SDE_0_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_0_MUX_inst_AND1_U1 ( .A1(KeyReg_n8), .A2(
        KeyReg_Inst_ff_SDE_0_MUX_inst_X), .ZN(KeyReg_Inst_ff_SDE_0_MUX_inst_Y)
         );
  XOR2_X1 KeyReg_Inst_ff_SDE_0_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_0_MUX_inst_Y), .B(KeyExpansionOutput[0]), .Z(
        KeyReg_Inst_ff_SDE_0_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_0_current_state_reg_U1 ( .A(key_shifted[8]), .ZN(
        KeyReg_Inst_ff_SDE_0_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_0_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_0_next_state), .CK(clk), .Q(key_shifted[8]), .QN()
         );
  XOR2_X1 KeyReg_Inst_ff_SDE_1_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[1]), 
        .B(RoundInput[121]), .Z(KeyReg_Inst_ff_SDE_1_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_1_MUX_inst_AND1_U1 ( .A1(KeyReg_n9), .A2(
        KeyReg_Inst_ff_SDE_1_MUX_inst_X), .ZN(KeyReg_Inst_ff_SDE_1_MUX_inst_Y)
         );
  XOR2_X1 KeyReg_Inst_ff_SDE_1_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_1_MUX_inst_Y), .B(KeyExpansionOutput[1]), .Z(
        KeyReg_Inst_ff_SDE_1_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_1_current_state_reg_U1 ( .A(key_shifted[9]), .ZN(
        KeyReg_Inst_ff_SDE_1_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_1_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_1_next_state), .CK(clk), .Q(key_shifted[9]), .QN()
         );
  XOR2_X1 KeyReg_Inst_ff_SDE_2_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[2]), 
        .B(RoundInput[122]), .Z(KeyReg_Inst_ff_SDE_2_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_2_MUX_inst_AND1_U1 ( .A1(KeyReg_n6), .A2(
        KeyReg_Inst_ff_SDE_2_MUX_inst_X), .ZN(KeyReg_Inst_ff_SDE_2_MUX_inst_Y)
         );
  XOR2_X1 KeyReg_Inst_ff_SDE_2_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_2_MUX_inst_Y), .B(KeyExpansionOutput[2]), .Z(
        KeyReg_Inst_ff_SDE_2_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_2_current_state_reg_U1 ( .A(key_shifted[10]), .ZN(
        KeyReg_Inst_ff_SDE_2_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_2_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_2_next_state), .CK(clk), .Q(key_shifted[10]), .QN()
         );
  XOR2_X1 KeyReg_Inst_ff_SDE_3_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[3]), 
        .B(RoundInput[123]), .Z(KeyReg_Inst_ff_SDE_3_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_3_MUX_inst_AND1_U1 ( .A1(KeyReg_n7), .A2(
        KeyReg_Inst_ff_SDE_3_MUX_inst_X), .ZN(KeyReg_Inst_ff_SDE_3_MUX_inst_Y)
         );
  XOR2_X1 KeyReg_Inst_ff_SDE_3_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_3_MUX_inst_Y), .B(KeyExpansionOutput[3]), .Z(
        KeyReg_Inst_ff_SDE_3_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_3_current_state_reg_U1 ( .A(key_shifted[11]), .ZN(
        KeyReg_Inst_ff_SDE_3_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_3_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_3_next_state), .CK(clk), .Q(key_shifted[11]), .QN()
         );
  XOR2_X1 KeyReg_Inst_ff_SDE_4_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[4]), 
        .B(RoundInput[124]), .Z(KeyReg_Inst_ff_SDE_4_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_4_MUX_inst_AND1_U1 ( .A1(KeyReg_n6), .A2(
        KeyReg_Inst_ff_SDE_4_MUX_inst_X), .ZN(KeyReg_Inst_ff_SDE_4_MUX_inst_Y)
         );
  XOR2_X1 KeyReg_Inst_ff_SDE_4_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_4_MUX_inst_Y), .B(KeyExpansionOutput[4]), .Z(
        KeyReg_Inst_ff_SDE_4_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_4_current_state_reg_U1 ( .A(key_shifted[12]), .ZN(
        KeyReg_Inst_ff_SDE_4_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_4_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_4_next_state), .CK(clk), .Q(key_shifted[12]), .QN()
         );
  XOR2_X1 KeyReg_Inst_ff_SDE_5_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[5]), 
        .B(RoundInput[125]), .Z(KeyReg_Inst_ff_SDE_5_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_5_MUX_inst_AND1_U1 ( .A1(KeyReg_n7), .A2(
        KeyReg_Inst_ff_SDE_5_MUX_inst_X), .ZN(KeyReg_Inst_ff_SDE_5_MUX_inst_Y)
         );
  XOR2_X1 KeyReg_Inst_ff_SDE_5_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_5_MUX_inst_Y), .B(KeyExpansionOutput[5]), .Z(
        KeyReg_Inst_ff_SDE_5_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_5_current_state_reg_U1 ( .A(key_shifted[13]), .ZN(
        KeyReg_Inst_ff_SDE_5_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_5_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_5_next_state), .CK(clk), .Q(key_shifted[13]), .QN()
         );
  XOR2_X1 KeyReg_Inst_ff_SDE_6_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[6]), 
        .B(RoundInput[126]), .Z(KeyReg_Inst_ff_SDE_6_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_6_MUX_inst_AND1_U1 ( .A1(KeyReg_n8), .A2(
        KeyReg_Inst_ff_SDE_6_MUX_inst_X), .ZN(KeyReg_Inst_ff_SDE_6_MUX_inst_Y)
         );
  XOR2_X1 KeyReg_Inst_ff_SDE_6_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_6_MUX_inst_Y), .B(KeyExpansionOutput[6]), .Z(
        KeyReg_Inst_ff_SDE_6_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_6_current_state_reg_U1 ( .A(key_shifted[14]), .ZN(
        KeyReg_Inst_ff_SDE_6_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_6_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_6_next_state), .CK(clk), .Q(key_shifted[14]), .QN()
         );
  XOR2_X1 KeyReg_Inst_ff_SDE_7_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[7]), 
        .B(RoundInput[127]), .Z(KeyReg_Inst_ff_SDE_7_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_7_MUX_inst_AND1_U1 ( .A1(KeyReg_n6), .A2(
        KeyReg_Inst_ff_SDE_7_MUX_inst_X), .ZN(KeyReg_Inst_ff_SDE_7_MUX_inst_Y)
         );
  XOR2_X1 KeyReg_Inst_ff_SDE_7_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_7_MUX_inst_Y), .B(KeyExpansionOutput[7]), .Z(
        KeyReg_Inst_ff_SDE_7_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_7_current_state_reg_U1 ( .A(key_shifted[15]), .ZN(
        KeyReg_Inst_ff_SDE_7_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_7_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_7_next_state), .CK(clk), .Q(key_shifted[15]), .QN()
         );
  XOR2_X1 KeyReg_Inst_ff_SDE_8_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[8]), 
        .B(key_shifted[8]), .Z(KeyReg_Inst_ff_SDE_8_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_8_MUX_inst_AND1_U1 ( .A1(KeyReg_n7), .A2(
        KeyReg_Inst_ff_SDE_8_MUX_inst_X), .ZN(KeyReg_Inst_ff_SDE_8_MUX_inst_Y)
         );
  XOR2_X1 KeyReg_Inst_ff_SDE_8_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_8_MUX_inst_Y), .B(KeyExpansionOutput[8]), .Z(
        KeyReg_Inst_ff_SDE_8_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_8_current_state_reg_U1 ( .A(key_shifted[16]), .ZN(
        KeyReg_Inst_ff_SDE_8_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_8_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_8_next_state), .CK(clk), .Q(key_shifted[16]), .QN()
         );
  XOR2_X1 KeyReg_Inst_ff_SDE_9_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[9]), 
        .B(key_shifted[9]), .Z(KeyReg_Inst_ff_SDE_9_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_9_MUX_inst_AND1_U1 ( .A1(KeyReg_n8), .A2(
        KeyReg_Inst_ff_SDE_9_MUX_inst_X), .ZN(KeyReg_Inst_ff_SDE_9_MUX_inst_Y)
         );
  XOR2_X1 KeyReg_Inst_ff_SDE_9_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_9_MUX_inst_Y), .B(KeyExpansionOutput[9]), .Z(
        KeyReg_Inst_ff_SDE_9_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_9_current_state_reg_U1 ( .A(key_shifted[17]), .ZN(
        KeyReg_Inst_ff_SDE_9_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_9_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_9_next_state), .CK(clk), .Q(key_shifted[17]), .QN()
         );
  XOR2_X1 KeyReg_Inst_ff_SDE_10_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[10]), 
        .B(key_shifted[10]), .Z(KeyReg_Inst_ff_SDE_10_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_10_MUX_inst_AND1_U1 ( .A1(KeyReg_n9), .A2(
        KeyReg_Inst_ff_SDE_10_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_10_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_10_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_10_MUX_inst_Y), .B(KeyExpansionOutput[10]), .Z(
        KeyReg_Inst_ff_SDE_10_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_10_current_state_reg_U1 ( .A(key_shifted[18]), 
        .ZN(KeyReg_Inst_ff_SDE_10_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_10_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_10_next_state), .CK(clk), .Q(key_shifted[18]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_11_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[11]), 
        .B(key_shifted[11]), .Z(KeyReg_Inst_ff_SDE_11_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_11_MUX_inst_AND1_U1 ( .A1(KeyReg_n7), .A2(
        KeyReg_Inst_ff_SDE_11_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_11_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_11_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_11_MUX_inst_Y), .B(KeyExpansionOutput[11]), .Z(
        KeyReg_Inst_ff_SDE_11_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_11_current_state_reg_U1 ( .A(key_shifted[19]), 
        .ZN(KeyReg_Inst_ff_SDE_11_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_11_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_11_next_state), .CK(clk), .Q(key_shifted[19]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_12_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[12]), 
        .B(key_shifted[12]), .Z(KeyReg_Inst_ff_SDE_12_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_12_MUX_inst_AND1_U1 ( .A1(KeyReg_n6), .A2(
        KeyReg_Inst_ff_SDE_12_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_12_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_12_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_12_MUX_inst_Y), .B(KeyExpansionOutput[12]), .Z(
        KeyReg_Inst_ff_SDE_12_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_12_current_state_reg_U1 ( .A(key_shifted[20]), 
        .ZN(KeyReg_Inst_ff_SDE_12_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_12_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_12_next_state), .CK(clk), .Q(key_shifted[20]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_13_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[13]), 
        .B(key_shifted[13]), .Z(KeyReg_Inst_ff_SDE_13_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_13_MUX_inst_AND1_U1 ( .A1(KeyReg_n6), .A2(
        KeyReg_Inst_ff_SDE_13_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_13_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_13_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_13_MUX_inst_Y), .B(KeyExpansionOutput[13]), .Z(
        KeyReg_Inst_ff_SDE_13_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_13_current_state_reg_U1 ( .A(key_shifted[21]), 
        .ZN(KeyReg_Inst_ff_SDE_13_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_13_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_13_next_state), .CK(clk), .Q(key_shifted[21]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_14_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[14]), 
        .B(key_shifted[14]), .Z(KeyReg_Inst_ff_SDE_14_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_14_MUX_inst_AND1_U1 ( .A1(KeyReg_n9), .A2(
        KeyReg_Inst_ff_SDE_14_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_14_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_14_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_14_MUX_inst_Y), .B(KeyExpansionOutput[14]), .Z(
        KeyReg_Inst_ff_SDE_14_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_14_current_state_reg_U1 ( .A(key_shifted[22]), 
        .ZN(KeyReg_Inst_ff_SDE_14_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_14_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_14_next_state), .CK(clk), .Q(key_shifted[22]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_15_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[15]), 
        .B(key_shifted[15]), .Z(KeyReg_Inst_ff_SDE_15_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_15_MUX_inst_AND1_U1 ( .A1(KeyReg_n8), .A2(
        KeyReg_Inst_ff_SDE_15_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_15_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_15_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_15_MUX_inst_Y), .B(KeyExpansionOutput[15]), .Z(
        KeyReg_Inst_ff_SDE_15_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_15_current_state_reg_U1 ( .A(key_shifted[23]), 
        .ZN(KeyReg_Inst_ff_SDE_15_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_15_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_15_next_state), .CK(clk), .Q(key_shifted[23]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_16_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[16]), 
        .B(key_shifted[16]), .Z(KeyReg_Inst_ff_SDE_16_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_16_MUX_inst_AND1_U1 ( .A1(KeyReg_n7), .A2(
        KeyReg_Inst_ff_SDE_16_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_16_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_16_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_16_MUX_inst_Y), .B(KeyExpansionOutput[16]), .Z(
        KeyReg_Inst_ff_SDE_16_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_16_current_state_reg_U1 ( .A(key_shifted[24]), 
        .ZN(KeyReg_Inst_ff_SDE_16_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_16_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_16_next_state), .CK(clk), .Q(key_shifted[24]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_17_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[17]), 
        .B(key_shifted[17]), .Z(KeyReg_Inst_ff_SDE_17_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_17_MUX_inst_AND1_U1 ( .A1(KeyReg_n8), .A2(
        KeyReg_Inst_ff_SDE_17_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_17_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_17_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_17_MUX_inst_Y), .B(KeyExpansionOutput[17]), .Z(
        KeyReg_Inst_ff_SDE_17_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_17_current_state_reg_U1 ( .A(key_shifted[25]), 
        .ZN(KeyReg_Inst_ff_SDE_17_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_17_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_17_next_state), .CK(clk), .Q(key_shifted[25]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_18_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[18]), 
        .B(key_shifted[18]), .Z(KeyReg_Inst_ff_SDE_18_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_18_MUX_inst_AND1_U1 ( .A1(KeyReg_n9), .A2(
        KeyReg_Inst_ff_SDE_18_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_18_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_18_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_18_MUX_inst_Y), .B(KeyExpansionOutput[18]), .Z(
        KeyReg_Inst_ff_SDE_18_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_18_current_state_reg_U1 ( .A(key_shifted[26]), 
        .ZN(KeyReg_Inst_ff_SDE_18_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_18_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_18_next_state), .CK(clk), .Q(key_shifted[26]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_19_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[19]), 
        .B(key_shifted[19]), .Z(KeyReg_Inst_ff_SDE_19_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_19_MUX_inst_AND1_U1 ( .A1(KeyReg_n8), .A2(
        KeyReg_Inst_ff_SDE_19_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_19_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_19_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_19_MUX_inst_Y), .B(KeyExpansionOutput[19]), .Z(
        KeyReg_Inst_ff_SDE_19_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_19_current_state_reg_U1 ( .A(key_shifted[27]), 
        .ZN(KeyReg_Inst_ff_SDE_19_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_19_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_19_next_state), .CK(clk), .Q(key_shifted[27]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_20_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[20]), 
        .B(key_shifted[20]), .Z(KeyReg_Inst_ff_SDE_20_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_20_MUX_inst_AND1_U1 ( .A1(KeyReg_n9), .A2(
        KeyReg_Inst_ff_SDE_20_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_20_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_20_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_20_MUX_inst_Y), .B(KeyExpansionOutput[20]), .Z(
        KeyReg_Inst_ff_SDE_20_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_20_current_state_reg_U1 ( .A(key_shifted[28]), 
        .ZN(KeyReg_Inst_ff_SDE_20_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_20_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_20_next_state), .CK(clk), .Q(key_shifted[28]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_21_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[21]), 
        .B(key_shifted[21]), .Z(KeyReg_Inst_ff_SDE_21_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_21_MUX_inst_AND1_U1 ( .A1(KeyReg_n6), .A2(
        KeyReg_Inst_ff_SDE_21_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_21_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_21_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_21_MUX_inst_Y), .B(KeyExpansionOutput[21]), .Z(
        KeyReg_Inst_ff_SDE_21_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_21_current_state_reg_U1 ( .A(key_shifted[29]), 
        .ZN(KeyReg_Inst_ff_SDE_21_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_21_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_21_next_state), .CK(clk), .Q(key_shifted[29]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_22_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[22]), 
        .B(key_shifted[22]), .Z(KeyReg_Inst_ff_SDE_22_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_22_MUX_inst_AND1_U1 ( .A1(KeyReg_n7), .A2(
        KeyReg_Inst_ff_SDE_22_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_22_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_22_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_22_MUX_inst_Y), .B(KeyExpansionOutput[22]), .Z(
        KeyReg_Inst_ff_SDE_22_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_22_current_state_reg_U1 ( .A(key_shifted[30]), 
        .ZN(KeyReg_Inst_ff_SDE_22_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_22_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_22_next_state), .CK(clk), .Q(key_shifted[30]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_23_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[23]), 
        .B(key_shifted[23]), .Z(KeyReg_Inst_ff_SDE_23_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_23_MUX_inst_AND1_U1 ( .A1(KeyReg_n6), .A2(
        KeyReg_Inst_ff_SDE_23_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_23_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_23_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_23_MUX_inst_Y), .B(KeyExpansionOutput[23]), .Z(
        KeyReg_Inst_ff_SDE_23_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_23_current_state_reg_U1 ( .A(key_shifted[31]), 
        .ZN(KeyReg_Inst_ff_SDE_23_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_23_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_23_next_state), .CK(clk), .Q(key_shifted[31]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_24_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[24]), 
        .B(key_shifted[24]), .Z(KeyReg_Inst_ff_SDE_24_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_24_MUX_inst_AND1_U1 ( .A1(KeyReg_n7), .A2(
        KeyReg_Inst_ff_SDE_24_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_24_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_24_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_24_MUX_inst_Y), .B(KeyExpansionOutput[24]), .Z(
        KeyReg_Inst_ff_SDE_24_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_24_current_state_reg_U1 ( .A(key_shifted[32]), 
        .ZN(KeyReg_Inst_ff_SDE_24_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_24_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_24_next_state), .CK(clk), .Q(key_shifted[32]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_25_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[25]), 
        .B(key_shifted[25]), .Z(KeyReg_Inst_ff_SDE_25_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_25_MUX_inst_AND1_U1 ( .A1(KeyReg_n8), .A2(
        KeyReg_Inst_ff_SDE_25_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_25_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_25_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_25_MUX_inst_Y), .B(KeyExpansionOutput[25]), .Z(
        KeyReg_Inst_ff_SDE_25_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_25_current_state_reg_U1 ( .A(key_shifted[33]), 
        .ZN(KeyReg_Inst_ff_SDE_25_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_25_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_25_next_state), .CK(clk), .Q(key_shifted[33]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_26_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[26]), 
        .B(key_shifted[26]), .Z(KeyReg_Inst_ff_SDE_26_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_26_MUX_inst_AND1_U1 ( .A1(KeyReg_n9), .A2(
        KeyReg_Inst_ff_SDE_26_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_26_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_26_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_26_MUX_inst_Y), .B(KeyExpansionOutput[26]), .Z(
        KeyReg_Inst_ff_SDE_26_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_26_current_state_reg_U1 ( .A(key_shifted[34]), 
        .ZN(KeyReg_Inst_ff_SDE_26_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_26_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_26_next_state), .CK(clk), .Q(key_shifted[34]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_27_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[27]), 
        .B(key_shifted[27]), .Z(KeyReg_Inst_ff_SDE_27_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_27_MUX_inst_AND1_U1 ( .A1(KeyReg_n7), .A2(
        KeyReg_Inst_ff_SDE_27_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_27_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_27_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_27_MUX_inst_Y), .B(KeyExpansionOutput[27]), .Z(
        KeyReg_Inst_ff_SDE_27_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_27_current_state_reg_U1 ( .A(key_shifted[35]), 
        .ZN(KeyReg_Inst_ff_SDE_27_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_27_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_27_next_state), .CK(clk), .Q(key_shifted[35]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_28_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[28]), 
        .B(key_shifted[28]), .Z(KeyReg_Inst_ff_SDE_28_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_28_MUX_inst_AND1_U1 ( .A1(KeyReg_n6), .A2(
        KeyReg_Inst_ff_SDE_28_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_28_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_28_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_28_MUX_inst_Y), .B(KeyExpansionOutput[28]), .Z(
        KeyReg_Inst_ff_SDE_28_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_28_current_state_reg_U1 ( .A(key_shifted[36]), 
        .ZN(KeyReg_Inst_ff_SDE_28_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_28_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_28_next_state), .CK(clk), .Q(key_shifted[36]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_29_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[29]), 
        .B(key_shifted[29]), .Z(KeyReg_Inst_ff_SDE_29_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_29_MUX_inst_AND1_U1 ( .A1(KeyReg_n8), .A2(
        KeyReg_Inst_ff_SDE_29_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_29_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_29_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_29_MUX_inst_Y), .B(KeyExpansionOutput[29]), .Z(
        KeyReg_Inst_ff_SDE_29_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_29_current_state_reg_U1 ( .A(key_shifted[37]), 
        .ZN(KeyReg_Inst_ff_SDE_29_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_29_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_29_next_state), .CK(clk), .Q(key_shifted[37]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_30_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[30]), 
        .B(key_shifted[30]), .Z(KeyReg_Inst_ff_SDE_30_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_30_MUX_inst_AND1_U1 ( .A1(KeyReg_n9), .A2(
        KeyReg_Inst_ff_SDE_30_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_30_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_30_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_30_MUX_inst_Y), .B(KeyExpansionOutput[30]), .Z(
        KeyReg_Inst_ff_SDE_30_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_30_current_state_reg_U1 ( .A(key_shifted[38]), 
        .ZN(KeyReg_Inst_ff_SDE_30_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_30_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_30_next_state), .CK(clk), .Q(key_shifted[38]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_31_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[31]), 
        .B(key_shifted[31]), .Z(KeyReg_Inst_ff_SDE_31_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_31_MUX_inst_AND1_U1 ( .A1(KeyReg_n7), .A2(
        KeyReg_Inst_ff_SDE_31_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_31_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_31_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_31_MUX_inst_Y), .B(KeyExpansionOutput[31]), .Z(
        KeyReg_Inst_ff_SDE_31_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_31_current_state_reg_U1 ( .A(key_shifted[39]), 
        .ZN(KeyReg_Inst_ff_SDE_31_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_31_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_31_next_state), .CK(clk), .Q(key_shifted[39]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_32_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[32]), 
        .B(key_shifted[32]), .Z(KeyReg_Inst_ff_SDE_32_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_32_MUX_inst_AND1_U1 ( .A1(KeyReg_n9), .A2(
        KeyReg_Inst_ff_SDE_32_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_32_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_32_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_32_MUX_inst_Y), .B(KeyExpansionOutput[32]), .Z(
        KeyReg_Inst_ff_SDE_32_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_32_current_state_reg_U1 ( .A(key_shifted[40]), 
        .ZN(KeyReg_Inst_ff_SDE_32_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_32_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_32_next_state), .CK(clk), .Q(key_shifted[40]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_33_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[33]), 
        .B(key_shifted[33]), .Z(KeyReg_Inst_ff_SDE_33_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_33_MUX_inst_AND1_U1 ( .A1(KeyReg_n7), .A2(
        KeyReg_Inst_ff_SDE_33_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_33_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_33_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_33_MUX_inst_Y), .B(KeyExpansionOutput[33]), .Z(
        KeyReg_Inst_ff_SDE_33_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_33_current_state_reg_U1 ( .A(key_shifted[41]), 
        .ZN(KeyReg_Inst_ff_SDE_33_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_33_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_33_next_state), .CK(clk), .Q(key_shifted[41]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_34_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[34]), 
        .B(key_shifted[34]), .Z(KeyReg_Inst_ff_SDE_34_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_34_MUX_inst_AND1_U1 ( .A1(KeyReg_n8), .A2(
        KeyReg_Inst_ff_SDE_34_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_34_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_34_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_34_MUX_inst_Y), .B(KeyExpansionOutput[34]), .Z(
        KeyReg_Inst_ff_SDE_34_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_34_current_state_reg_U1 ( .A(key_shifted[42]), 
        .ZN(KeyReg_Inst_ff_SDE_34_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_34_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_34_next_state), .CK(clk), .Q(key_shifted[42]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_35_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[35]), 
        .B(key_shifted[35]), .Z(KeyReg_Inst_ff_SDE_35_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_35_MUX_inst_AND1_U1 ( .A1(KeyReg_n7), .A2(
        KeyReg_Inst_ff_SDE_35_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_35_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_35_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_35_MUX_inst_Y), .B(KeyExpansionOutput[35]), .Z(
        KeyReg_Inst_ff_SDE_35_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_35_current_state_reg_U1 ( .A(key_shifted[43]), 
        .ZN(KeyReg_Inst_ff_SDE_35_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_35_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_35_next_state), .CK(clk), .Q(key_shifted[43]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_36_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[36]), 
        .B(key_shifted[36]), .Z(KeyReg_Inst_ff_SDE_36_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_36_MUX_inst_AND1_U1 ( .A1(KeyReg_n8), .A2(
        KeyReg_Inst_ff_SDE_36_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_36_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_36_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_36_MUX_inst_Y), .B(KeyExpansionOutput[36]), .Z(
        KeyReg_Inst_ff_SDE_36_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_36_current_state_reg_U1 ( .A(key_shifted[44]), 
        .ZN(KeyReg_Inst_ff_SDE_36_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_36_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_36_next_state), .CK(clk), .Q(key_shifted[44]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_37_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[37]), 
        .B(key_shifted[37]), .Z(KeyReg_Inst_ff_SDE_37_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_37_MUX_inst_AND1_U1 ( .A1(KeyReg_n9), .A2(
        KeyReg_Inst_ff_SDE_37_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_37_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_37_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_37_MUX_inst_Y), .B(KeyExpansionOutput[37]), .Z(
        KeyReg_Inst_ff_SDE_37_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_37_current_state_reg_U1 ( .A(key_shifted[45]), 
        .ZN(KeyReg_Inst_ff_SDE_37_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_37_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_37_next_state), .CK(clk), .Q(key_shifted[45]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_38_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[38]), 
        .B(key_shifted[38]), .Z(KeyReg_Inst_ff_SDE_38_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_38_MUX_inst_AND1_U1 ( .A1(KeyReg_n8), .A2(
        KeyReg_Inst_ff_SDE_38_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_38_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_38_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_38_MUX_inst_Y), .B(KeyExpansionOutput[38]), .Z(
        KeyReg_Inst_ff_SDE_38_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_38_current_state_reg_U1 ( .A(key_shifted[46]), 
        .ZN(KeyReg_Inst_ff_SDE_38_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_38_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_38_next_state), .CK(clk), .Q(key_shifted[46]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_39_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[39]), 
        .B(key_shifted[39]), .Z(KeyReg_Inst_ff_SDE_39_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_39_MUX_inst_AND1_U1 ( .A1(KeyReg_n9), .A2(
        KeyReg_Inst_ff_SDE_39_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_39_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_39_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_39_MUX_inst_Y), .B(KeyExpansionOutput[39]), .Z(
        KeyReg_Inst_ff_SDE_39_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_39_current_state_reg_U1 ( .A(key_shifted[47]), 
        .ZN(KeyReg_Inst_ff_SDE_39_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_39_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_39_next_state), .CK(clk), .Q(key_shifted[47]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_40_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[40]), 
        .B(key_shifted[40]), .Z(KeyReg_Inst_ff_SDE_40_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_40_MUX_inst_AND1_U1 ( .A1(KeyReg_n7), .A2(
        KeyReg_Inst_ff_SDE_40_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_40_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_40_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_40_MUX_inst_Y), .B(KeyExpansionOutput[40]), .Z(
        KeyReg_Inst_ff_SDE_40_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_40_current_state_reg_U1 ( .A(key_shifted[48]), 
        .ZN(KeyReg_Inst_ff_SDE_40_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_40_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_40_next_state), .CK(clk), .Q(key_shifted[48]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_41_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[41]), 
        .B(key_shifted[41]), .Z(KeyReg_Inst_ff_SDE_41_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_41_MUX_inst_AND1_U1 ( .A1(KeyReg_n8), .A2(
        KeyReg_Inst_ff_SDE_41_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_41_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_41_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_41_MUX_inst_Y), .B(KeyExpansionOutput[41]), .Z(
        KeyReg_Inst_ff_SDE_41_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_41_current_state_reg_U1 ( .A(key_shifted[49]), 
        .ZN(KeyReg_Inst_ff_SDE_41_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_41_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_41_next_state), .CK(clk), .Q(key_shifted[49]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_42_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[42]), 
        .B(key_shifted[42]), .Z(KeyReg_Inst_ff_SDE_42_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_42_MUX_inst_AND1_U1 ( .A1(KeyReg_n9), .A2(
        KeyReg_Inst_ff_SDE_42_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_42_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_42_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_42_MUX_inst_Y), .B(KeyExpansionOutput[42]), .Z(
        KeyReg_Inst_ff_SDE_42_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_42_current_state_reg_U1 ( .A(key_shifted[50]), 
        .ZN(KeyReg_Inst_ff_SDE_42_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_42_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_42_next_state), .CK(clk), .Q(key_shifted[50]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_43_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[43]), 
        .B(key_shifted[43]), .Z(KeyReg_Inst_ff_SDE_43_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_43_MUX_inst_AND1_U1 ( .A1(KeyReg_n9), .A2(
        KeyReg_Inst_ff_SDE_43_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_43_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_43_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_43_MUX_inst_Y), .B(KeyExpansionOutput[43]), .Z(
        KeyReg_Inst_ff_SDE_43_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_43_current_state_reg_U1 ( .A(key_shifted[51]), 
        .ZN(KeyReg_Inst_ff_SDE_43_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_43_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_43_next_state), .CK(clk), .Q(key_shifted[51]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_44_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[44]), 
        .B(key_shifted[44]), .Z(KeyReg_Inst_ff_SDE_44_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_44_MUX_inst_AND1_U1 ( .A1(KeyReg_n7), .A2(
        KeyReg_Inst_ff_SDE_44_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_44_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_44_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_44_MUX_inst_Y), .B(KeyExpansionOutput[44]), .Z(
        KeyReg_Inst_ff_SDE_44_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_44_current_state_reg_U1 ( .A(key_shifted[52]), 
        .ZN(KeyReg_Inst_ff_SDE_44_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_44_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_44_next_state), .CK(clk), .Q(key_shifted[52]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_45_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[45]), 
        .B(key_shifted[45]), .Z(KeyReg_Inst_ff_SDE_45_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_45_MUX_inst_AND1_U1 ( .A1(KeyReg_n7), .A2(
        KeyReg_Inst_ff_SDE_45_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_45_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_45_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_45_MUX_inst_Y), .B(KeyExpansionOutput[45]), .Z(
        KeyReg_Inst_ff_SDE_45_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_45_current_state_reg_U1 ( .A(key_shifted[53]), 
        .ZN(KeyReg_Inst_ff_SDE_45_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_45_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_45_next_state), .CK(clk), .Q(key_shifted[53]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_46_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[46]), 
        .B(key_shifted[46]), .Z(KeyReg_Inst_ff_SDE_46_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_46_MUX_inst_AND1_U1 ( .A1(KeyReg_n8), .A2(
        KeyReg_Inst_ff_SDE_46_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_46_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_46_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_46_MUX_inst_Y), .B(KeyExpansionOutput[46]), .Z(
        KeyReg_Inst_ff_SDE_46_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_46_current_state_reg_U1 ( .A(key_shifted[54]), 
        .ZN(KeyReg_Inst_ff_SDE_46_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_46_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_46_next_state), .CK(clk), .Q(key_shifted[54]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_47_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[47]), 
        .B(key_shifted[47]), .Z(KeyReg_Inst_ff_SDE_47_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_47_MUX_inst_AND1_U1 ( .A1(KeyReg_n9), .A2(
        KeyReg_Inst_ff_SDE_47_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_47_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_47_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_47_MUX_inst_Y), .B(KeyExpansionOutput[47]), .Z(
        KeyReg_Inst_ff_SDE_47_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_47_current_state_reg_U1 ( .A(key_shifted[55]), 
        .ZN(KeyReg_Inst_ff_SDE_47_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_47_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_47_next_state), .CK(clk), .Q(key_shifted[55]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_48_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[48]), 
        .B(key_shifted[48]), .Z(KeyReg_Inst_ff_SDE_48_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_48_MUX_inst_AND1_U1 ( .A1(KeyReg_n8), .A2(
        KeyReg_Inst_ff_SDE_48_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_48_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_48_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_48_MUX_inst_Y), .B(KeyExpansionOutput[48]), .Z(
        KeyReg_Inst_ff_SDE_48_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_48_current_state_reg_U1 ( .A(key_shifted[56]), 
        .ZN(KeyReg_Inst_ff_SDE_48_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_48_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_48_next_state), .CK(clk), .Q(key_shifted[56]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_49_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[49]), 
        .B(key_shifted[49]), .Z(KeyReg_Inst_ff_SDE_49_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_49_MUX_inst_AND1_U1 ( .A1(KeyReg_n7), .A2(
        KeyReg_Inst_ff_SDE_49_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_49_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_49_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_49_MUX_inst_Y), .B(KeyExpansionOutput[49]), .Z(
        KeyReg_Inst_ff_SDE_49_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_49_current_state_reg_U1 ( .A(key_shifted[57]), 
        .ZN(KeyReg_Inst_ff_SDE_49_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_49_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_49_next_state), .CK(clk), .Q(key_shifted[57]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_50_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[50]), 
        .B(key_shifted[50]), .Z(KeyReg_Inst_ff_SDE_50_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_50_MUX_inst_AND1_U1 ( .A1(KeyReg_n8), .A2(
        KeyReg_Inst_ff_SDE_50_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_50_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_50_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_50_MUX_inst_Y), .B(KeyExpansionOutput[50]), .Z(
        KeyReg_Inst_ff_SDE_50_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_50_current_state_reg_U1 ( .A(key_shifted[58]), 
        .ZN(KeyReg_Inst_ff_SDE_50_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_50_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_50_next_state), .CK(clk), .Q(key_shifted[58]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_51_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[51]), 
        .B(key_shifted[51]), .Z(KeyReg_Inst_ff_SDE_51_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_51_MUX_inst_AND1_U1 ( .A1(KeyReg_n9), .A2(
        KeyReg_Inst_ff_SDE_51_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_51_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_51_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_51_MUX_inst_Y), .B(KeyExpansionOutput[51]), .Z(
        KeyReg_Inst_ff_SDE_51_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_51_current_state_reg_U1 ( .A(key_shifted[59]), 
        .ZN(KeyReg_Inst_ff_SDE_51_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_51_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_51_next_state), .CK(clk), .Q(key_shifted[59]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_52_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[52]), 
        .B(key_shifted[52]), .Z(KeyReg_Inst_ff_SDE_52_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_52_MUX_inst_AND1_U1 ( .A1(KeyReg_n9), .A2(
        KeyReg_Inst_ff_SDE_52_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_52_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_52_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_52_MUX_inst_Y), .B(KeyExpansionOutput[52]), .Z(
        KeyReg_Inst_ff_SDE_52_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_52_current_state_reg_U1 ( .A(key_shifted[60]), 
        .ZN(KeyReg_Inst_ff_SDE_52_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_52_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_52_next_state), .CK(clk), .Q(key_shifted[60]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_53_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[53]), 
        .B(key_shifted[53]), .Z(KeyReg_Inst_ff_SDE_53_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_53_MUX_inst_AND1_U1 ( .A1(KeyReg_n7), .A2(
        KeyReg_Inst_ff_SDE_53_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_53_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_53_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_53_MUX_inst_Y), .B(KeyExpansionOutput[53]), .Z(
        KeyReg_Inst_ff_SDE_53_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_53_current_state_reg_U1 ( .A(key_shifted[61]), 
        .ZN(KeyReg_Inst_ff_SDE_53_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_53_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_53_next_state), .CK(clk), .Q(key_shifted[61]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_54_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[54]), 
        .B(key_shifted[54]), .Z(KeyReg_Inst_ff_SDE_54_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_54_MUX_inst_AND1_U1 ( .A1(KeyReg_n8), .A2(
        KeyReg_Inst_ff_SDE_54_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_54_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_54_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_54_MUX_inst_Y), .B(KeyExpansionOutput[54]), .Z(
        KeyReg_Inst_ff_SDE_54_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_54_current_state_reg_U1 ( .A(key_shifted[62]), 
        .ZN(KeyReg_Inst_ff_SDE_54_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_54_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_54_next_state), .CK(clk), .Q(key_shifted[62]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_55_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[55]), 
        .B(key_shifted[55]), .Z(KeyReg_Inst_ff_SDE_55_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_55_MUX_inst_AND1_U1 ( .A1(KeyReg_n9), .A2(
        KeyReg_Inst_ff_SDE_55_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_55_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_55_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_55_MUX_inst_Y), .B(KeyExpansionOutput[55]), .Z(
        KeyReg_Inst_ff_SDE_55_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_55_current_state_reg_U1 ( .A(key_shifted[63]), 
        .ZN(KeyReg_Inst_ff_SDE_55_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_55_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_55_next_state), .CK(clk), .Q(key_shifted[63]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_56_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[56]), 
        .B(key_shifted[56]), .Z(KeyReg_Inst_ff_SDE_56_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_56_MUX_inst_AND1_U1 ( .A1(KeyReg_n7), .A2(
        KeyReg_Inst_ff_SDE_56_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_56_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_56_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_56_MUX_inst_Y), .B(KeyExpansionOutput[56]), .Z(
        KeyReg_Inst_ff_SDE_56_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_56_current_state_reg_U1 ( .A(key_shifted[64]), 
        .ZN(KeyReg_Inst_ff_SDE_56_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_56_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_56_next_state), .CK(clk), .Q(key_shifted[64]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_57_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[57]), 
        .B(key_shifted[57]), .Z(KeyReg_Inst_ff_SDE_57_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_57_MUX_inst_AND1_U1 ( .A1(KeyReg_n8), .A2(
        KeyReg_Inst_ff_SDE_57_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_57_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_57_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_57_MUX_inst_Y), .B(KeyExpansionOutput[57]), .Z(
        KeyReg_Inst_ff_SDE_57_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_57_current_state_reg_U1 ( .A(key_shifted[65]), 
        .ZN(KeyReg_Inst_ff_SDE_57_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_57_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_57_next_state), .CK(clk), .Q(key_shifted[65]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_58_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[58]), 
        .B(key_shifted[58]), .Z(KeyReg_Inst_ff_SDE_58_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_58_MUX_inst_AND1_U1 ( .A1(KeyReg_n9), .A2(
        KeyReg_Inst_ff_SDE_58_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_58_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_58_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_58_MUX_inst_Y), .B(KeyExpansionOutput[58]), .Z(
        KeyReg_Inst_ff_SDE_58_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_58_current_state_reg_U1 ( .A(key_shifted[66]), 
        .ZN(KeyReg_Inst_ff_SDE_58_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_58_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_58_next_state), .CK(clk), .Q(key_shifted[66]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_59_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[59]), 
        .B(key_shifted[59]), .Z(KeyReg_Inst_ff_SDE_59_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_59_MUX_inst_AND1_U1 ( .A1(KeyReg_n6), .A2(
        KeyReg_Inst_ff_SDE_59_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_59_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_59_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_59_MUX_inst_Y), .B(KeyExpansionOutput[59]), .Z(
        KeyReg_Inst_ff_SDE_59_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_59_current_state_reg_U1 ( .A(key_shifted[67]), 
        .ZN(KeyReg_Inst_ff_SDE_59_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_59_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_59_next_state), .CK(clk), .Q(key_shifted[67]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_60_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[60]), 
        .B(key_shifted[60]), .Z(KeyReg_Inst_ff_SDE_60_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_60_MUX_inst_AND1_U1 ( .A1(start_done), .A2(
        KeyReg_Inst_ff_SDE_60_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_60_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_60_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_60_MUX_inst_Y), .B(KeyExpansionOutput[60]), .Z(
        KeyReg_Inst_ff_SDE_60_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_60_current_state_reg_U1 ( .A(key_shifted[68]), 
        .ZN(KeyReg_Inst_ff_SDE_60_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_60_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_60_next_state), .CK(clk), .Q(key_shifted[68]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_61_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[61]), 
        .B(key_shifted[61]), .Z(KeyReg_Inst_ff_SDE_61_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_61_MUX_inst_AND1_U1 ( .A1(start_done), .A2(
        KeyReg_Inst_ff_SDE_61_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_61_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_61_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_61_MUX_inst_Y), .B(KeyExpansionOutput[61]), .Z(
        KeyReg_Inst_ff_SDE_61_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_61_current_state_reg_U1 ( .A(key_shifted[69]), 
        .ZN(KeyReg_Inst_ff_SDE_61_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_61_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_61_next_state), .CK(clk), .Q(key_shifted[69]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_62_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[62]), 
        .B(key_shifted[62]), .Z(KeyReg_Inst_ff_SDE_62_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_62_MUX_inst_AND1_U1 ( .A1(KeyReg_n6), .A2(
        KeyReg_Inst_ff_SDE_62_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_62_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_62_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_62_MUX_inst_Y), .B(KeyExpansionOutput[62]), .Z(
        KeyReg_Inst_ff_SDE_62_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_62_current_state_reg_U1 ( .A(key_shifted[70]), 
        .ZN(KeyReg_Inst_ff_SDE_62_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_62_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_62_next_state), .CK(clk), .Q(key_shifted[70]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_63_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[63]), 
        .B(key_shifted[63]), .Z(KeyReg_Inst_ff_SDE_63_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_63_MUX_inst_AND1_U1 ( .A1(KeyReg_n6), .A2(
        KeyReg_Inst_ff_SDE_63_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_63_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_63_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_63_MUX_inst_Y), .B(KeyExpansionOutput[63]), .Z(
        KeyReg_Inst_ff_SDE_63_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_63_current_state_reg_U1 ( .A(key_shifted[71]), 
        .ZN(KeyReg_Inst_ff_SDE_63_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_63_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_63_next_state), .CK(clk), .Q(key_shifted[71]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_64_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[64]), 
        .B(key_shifted[64]), .Z(KeyReg_Inst_ff_SDE_64_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_64_MUX_inst_AND1_U1 ( .A1(KeyReg_n6), .A2(
        KeyReg_Inst_ff_SDE_64_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_64_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_64_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_64_MUX_inst_Y), .B(KeyExpansionOutput[64]), .Z(
        KeyReg_Inst_ff_SDE_64_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_64_current_state_reg_U1 ( .A(key_shifted[72]), 
        .ZN(KeyReg_Inst_ff_SDE_64_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_64_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_64_next_state), .CK(clk), .Q(key_shifted[72]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_65_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[65]), 
        .B(key_shifted[65]), .Z(KeyReg_Inst_ff_SDE_65_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_65_MUX_inst_AND1_U1 ( .A1(KeyReg_n6), .A2(
        KeyReg_Inst_ff_SDE_65_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_65_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_65_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_65_MUX_inst_Y), .B(KeyExpansionOutput[65]), .Z(
        KeyReg_Inst_ff_SDE_65_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_65_current_state_reg_U1 ( .A(key_shifted[73]), 
        .ZN(KeyReg_Inst_ff_SDE_65_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_65_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_65_next_state), .CK(clk), .Q(key_shifted[73]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_66_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[66]), 
        .B(key_shifted[66]), .Z(KeyReg_Inst_ff_SDE_66_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_66_MUX_inst_AND1_U1 ( .A1(KeyReg_n6), .A2(
        KeyReg_Inst_ff_SDE_66_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_66_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_66_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_66_MUX_inst_Y), .B(KeyExpansionOutput[66]), .Z(
        KeyReg_Inst_ff_SDE_66_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_66_current_state_reg_U1 ( .A(key_shifted[74]), 
        .ZN(KeyReg_Inst_ff_SDE_66_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_66_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_66_next_state), .CK(clk), .Q(key_shifted[74]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_67_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[67]), 
        .B(key_shifted[67]), .Z(KeyReg_Inst_ff_SDE_67_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_67_MUX_inst_AND1_U1 ( .A1(KeyReg_n6), .A2(
        KeyReg_Inst_ff_SDE_67_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_67_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_67_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_67_MUX_inst_Y), .B(KeyExpansionOutput[67]), .Z(
        KeyReg_Inst_ff_SDE_67_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_67_current_state_reg_U1 ( .A(key_shifted[75]), 
        .ZN(KeyReg_Inst_ff_SDE_67_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_67_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_67_next_state), .CK(clk), .Q(key_shifted[75]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_68_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[68]), 
        .B(key_shifted[68]), .Z(KeyReg_Inst_ff_SDE_68_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_68_MUX_inst_AND1_U1 ( .A1(KeyReg_n9), .A2(
        KeyReg_Inst_ff_SDE_68_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_68_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_68_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_68_MUX_inst_Y), .B(KeyExpansionOutput[68]), .Z(
        KeyReg_Inst_ff_SDE_68_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_68_current_state_reg_U1 ( .A(key_shifted[76]), 
        .ZN(KeyReg_Inst_ff_SDE_68_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_68_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_68_next_state), .CK(clk), .Q(key_shifted[76]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_69_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[69]), 
        .B(key_shifted[69]), .Z(KeyReg_Inst_ff_SDE_69_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_69_MUX_inst_AND1_U1 ( .A1(KeyReg_n9), .A2(
        KeyReg_Inst_ff_SDE_69_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_69_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_69_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_69_MUX_inst_Y), .B(KeyExpansionOutput[69]), .Z(
        KeyReg_Inst_ff_SDE_69_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_69_current_state_reg_U1 ( .A(key_shifted[77]), 
        .ZN(KeyReg_Inst_ff_SDE_69_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_69_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_69_next_state), .CK(clk), .Q(key_shifted[77]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_70_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[70]), 
        .B(key_shifted[70]), .Z(KeyReg_Inst_ff_SDE_70_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_70_MUX_inst_AND1_U1 ( .A1(KeyReg_n9), .A2(
        KeyReg_Inst_ff_SDE_70_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_70_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_70_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_70_MUX_inst_Y), .B(KeyExpansionOutput[70]), .Z(
        KeyReg_Inst_ff_SDE_70_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_70_current_state_reg_U1 ( .A(key_shifted[78]), 
        .ZN(KeyReg_Inst_ff_SDE_70_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_70_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_70_next_state), .CK(clk), .Q(key_shifted[78]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_71_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[71]), 
        .B(key_shifted[71]), .Z(KeyReg_Inst_ff_SDE_71_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_71_MUX_inst_AND1_U1 ( .A1(KeyReg_n9), .A2(
        KeyReg_Inst_ff_SDE_71_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_71_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_71_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_71_MUX_inst_Y), .B(KeyExpansionOutput[71]), .Z(
        KeyReg_Inst_ff_SDE_71_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_71_current_state_reg_U1 ( .A(key_shifted[79]), 
        .ZN(KeyReg_Inst_ff_SDE_71_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_71_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_71_next_state), .CK(clk), .Q(key_shifted[79]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_72_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[72]), 
        .B(key_shifted[72]), .Z(KeyReg_Inst_ff_SDE_72_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_72_MUX_inst_AND1_U1 ( .A1(KeyReg_n9), .A2(
        KeyReg_Inst_ff_SDE_72_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_72_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_72_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_72_MUX_inst_Y), .B(KeyExpansionOutput[72]), .Z(
        KeyReg_Inst_ff_SDE_72_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_72_current_state_reg_U1 ( .A(key_shifted[80]), 
        .ZN(KeyReg_Inst_ff_SDE_72_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_72_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_72_next_state), .CK(clk), .Q(key_shifted[80]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_73_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[73]), 
        .B(key_shifted[73]), .Z(KeyReg_Inst_ff_SDE_73_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_73_MUX_inst_AND1_U1 ( .A1(KeyReg_n9), .A2(
        KeyReg_Inst_ff_SDE_73_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_73_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_73_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_73_MUX_inst_Y), .B(KeyExpansionOutput[73]), .Z(
        KeyReg_Inst_ff_SDE_73_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_73_current_state_reg_U1 ( .A(key_shifted[81]), 
        .ZN(KeyReg_Inst_ff_SDE_73_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_73_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_73_next_state), .CK(clk), .Q(key_shifted[81]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_74_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[74]), 
        .B(key_shifted[74]), .Z(KeyReg_Inst_ff_SDE_74_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_74_MUX_inst_AND1_U1 ( .A1(KeyReg_n9), .A2(
        KeyReg_Inst_ff_SDE_74_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_74_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_74_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_74_MUX_inst_Y), .B(KeyExpansionOutput[74]), .Z(
        KeyReg_Inst_ff_SDE_74_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_74_current_state_reg_U1 ( .A(key_shifted[82]), 
        .ZN(KeyReg_Inst_ff_SDE_74_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_74_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_74_next_state), .CK(clk), .Q(key_shifted[82]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_75_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[75]), 
        .B(key_shifted[75]), .Z(KeyReg_Inst_ff_SDE_75_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_75_MUX_inst_AND1_U1 ( .A1(KeyReg_n9), .A2(
        KeyReg_Inst_ff_SDE_75_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_75_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_75_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_75_MUX_inst_Y), .B(KeyExpansionOutput[75]), .Z(
        KeyReg_Inst_ff_SDE_75_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_75_current_state_reg_U1 ( .A(key_shifted[83]), 
        .ZN(KeyReg_Inst_ff_SDE_75_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_75_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_75_next_state), .CK(clk), .Q(key_shifted[83]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_76_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[76]), 
        .B(key_shifted[76]), .Z(KeyReg_Inst_ff_SDE_76_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_76_MUX_inst_AND1_U1 ( .A1(KeyReg_n9), .A2(
        KeyReg_Inst_ff_SDE_76_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_76_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_76_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_76_MUX_inst_Y), .B(KeyExpansionOutput[76]), .Z(
        KeyReg_Inst_ff_SDE_76_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_76_current_state_reg_U1 ( .A(key_shifted[84]), 
        .ZN(KeyReg_Inst_ff_SDE_76_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_76_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_76_next_state), .CK(clk), .Q(key_shifted[84]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_77_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[77]), 
        .B(key_shifted[77]), .Z(KeyReg_Inst_ff_SDE_77_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_77_MUX_inst_AND1_U1 ( .A1(KeyReg_n9), .A2(
        KeyReg_Inst_ff_SDE_77_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_77_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_77_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_77_MUX_inst_Y), .B(KeyExpansionOutput[77]), .Z(
        KeyReg_Inst_ff_SDE_77_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_77_current_state_reg_U1 ( .A(key_shifted[85]), 
        .ZN(KeyReg_Inst_ff_SDE_77_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_77_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_77_next_state), .CK(clk), .Q(key_shifted[85]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_78_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[78]), 
        .B(key_shifted[78]), .Z(KeyReg_Inst_ff_SDE_78_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_78_MUX_inst_AND1_U1 ( .A1(KeyReg_n9), .A2(
        KeyReg_Inst_ff_SDE_78_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_78_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_78_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_78_MUX_inst_Y), .B(KeyExpansionOutput[78]), .Z(
        KeyReg_Inst_ff_SDE_78_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_78_current_state_reg_U1 ( .A(key_shifted[86]), 
        .ZN(KeyReg_Inst_ff_SDE_78_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_78_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_78_next_state), .CK(clk), .Q(key_shifted[86]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_79_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[79]), 
        .B(key_shifted[79]), .Z(KeyReg_Inst_ff_SDE_79_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_79_MUX_inst_AND1_U1 ( .A1(KeyReg_n9), .A2(
        KeyReg_Inst_ff_SDE_79_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_79_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_79_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_79_MUX_inst_Y), .B(KeyExpansionOutput[79]), .Z(
        KeyReg_Inst_ff_SDE_79_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_79_current_state_reg_U1 ( .A(key_shifted[87]), 
        .ZN(KeyReg_Inst_ff_SDE_79_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_79_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_79_next_state), .CK(clk), .Q(key_shifted[87]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_80_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[80]), 
        .B(key_shifted[80]), .Z(KeyReg_Inst_ff_SDE_80_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_80_MUX_inst_AND1_U1 ( .A1(KeyReg_n8), .A2(
        KeyReg_Inst_ff_SDE_80_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_80_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_80_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_80_MUX_inst_Y), .B(KeyExpansionOutput[80]), .Z(
        KeyReg_Inst_ff_SDE_80_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_80_current_state_reg_U1 ( .A(key_shifted[88]), 
        .ZN(KeyReg_Inst_ff_SDE_80_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_80_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_80_next_state), .CK(clk), .Q(key_shifted[88]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_81_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[81]), 
        .B(key_shifted[81]), .Z(KeyReg_Inst_ff_SDE_81_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_81_MUX_inst_AND1_U1 ( .A1(KeyReg_n8), .A2(
        KeyReg_Inst_ff_SDE_81_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_81_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_81_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_81_MUX_inst_Y), .B(KeyExpansionOutput[81]), .Z(
        KeyReg_Inst_ff_SDE_81_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_81_current_state_reg_U1 ( .A(key_shifted[89]), 
        .ZN(KeyReg_Inst_ff_SDE_81_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_81_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_81_next_state), .CK(clk), .Q(key_shifted[89]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_82_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[82]), 
        .B(key_shifted[82]), .Z(KeyReg_Inst_ff_SDE_82_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_82_MUX_inst_AND1_U1 ( .A1(KeyReg_n8), .A2(
        KeyReg_Inst_ff_SDE_82_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_82_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_82_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_82_MUX_inst_Y), .B(KeyExpansionOutput[82]), .Z(
        KeyReg_Inst_ff_SDE_82_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_82_current_state_reg_U1 ( .A(key_shifted[90]), 
        .ZN(KeyReg_Inst_ff_SDE_82_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_82_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_82_next_state), .CK(clk), .Q(key_shifted[90]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_83_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[83]), 
        .B(key_shifted[83]), .Z(KeyReg_Inst_ff_SDE_83_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_83_MUX_inst_AND1_U1 ( .A1(KeyReg_n8), .A2(
        KeyReg_Inst_ff_SDE_83_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_83_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_83_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_83_MUX_inst_Y), .B(KeyExpansionOutput[83]), .Z(
        KeyReg_Inst_ff_SDE_83_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_83_current_state_reg_U1 ( .A(key_shifted[91]), 
        .ZN(KeyReg_Inst_ff_SDE_83_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_83_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_83_next_state), .CK(clk), .Q(key_shifted[91]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_84_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[84]), 
        .B(key_shifted[84]), .Z(KeyReg_Inst_ff_SDE_84_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_84_MUX_inst_AND1_U1 ( .A1(KeyReg_n8), .A2(
        KeyReg_Inst_ff_SDE_84_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_84_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_84_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_84_MUX_inst_Y), .B(KeyExpansionOutput[84]), .Z(
        KeyReg_Inst_ff_SDE_84_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_84_current_state_reg_U1 ( .A(key_shifted[92]), 
        .ZN(KeyReg_Inst_ff_SDE_84_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_84_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_84_next_state), .CK(clk), .Q(key_shifted[92]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_85_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[85]), 
        .B(key_shifted[85]), .Z(KeyReg_Inst_ff_SDE_85_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_85_MUX_inst_AND1_U1 ( .A1(KeyReg_n8), .A2(
        KeyReg_Inst_ff_SDE_85_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_85_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_85_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_85_MUX_inst_Y), .B(KeyExpansionOutput[85]), .Z(
        KeyReg_Inst_ff_SDE_85_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_85_current_state_reg_U1 ( .A(key_shifted[93]), 
        .ZN(KeyReg_Inst_ff_SDE_85_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_85_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_85_next_state), .CK(clk), .Q(key_shifted[93]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_86_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[86]), 
        .B(key_shifted[86]), .Z(KeyReg_Inst_ff_SDE_86_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_86_MUX_inst_AND1_U1 ( .A1(KeyReg_n8), .A2(
        KeyReg_Inst_ff_SDE_86_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_86_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_86_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_86_MUX_inst_Y), .B(KeyExpansionOutput[86]), .Z(
        KeyReg_Inst_ff_SDE_86_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_86_current_state_reg_U1 ( .A(key_shifted[94]), 
        .ZN(KeyReg_Inst_ff_SDE_86_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_86_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_86_next_state), .CK(clk), .Q(key_shifted[94]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_87_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[87]), 
        .B(key_shifted[87]), .Z(KeyReg_Inst_ff_SDE_87_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_87_MUX_inst_AND1_U1 ( .A1(KeyReg_n8), .A2(
        KeyReg_Inst_ff_SDE_87_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_87_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_87_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_87_MUX_inst_Y), .B(KeyExpansionOutput[87]), .Z(
        KeyReg_Inst_ff_SDE_87_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_87_current_state_reg_U1 ( .A(key_shifted[95]), 
        .ZN(KeyReg_Inst_ff_SDE_87_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_87_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_87_next_state), .CK(clk), .Q(key_shifted[95]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_88_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[88]), 
        .B(key_shifted[88]), .Z(KeyReg_Inst_ff_SDE_88_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_88_MUX_inst_AND1_U1 ( .A1(KeyReg_n8), .A2(
        KeyReg_Inst_ff_SDE_88_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_88_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_88_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_88_MUX_inst_Y), .B(KeyExpansionOutput[88]), .Z(
        KeyReg_Inst_ff_SDE_88_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_88_current_state_reg_U1 ( .A(key_shifted[96]), 
        .ZN(KeyReg_Inst_ff_SDE_88_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_88_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_88_next_state), .CK(clk), .Q(key_shifted[96]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_89_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[89]), 
        .B(key_shifted[89]), .Z(KeyReg_Inst_ff_SDE_89_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_89_MUX_inst_AND1_U1 ( .A1(KeyReg_n8), .A2(
        KeyReg_Inst_ff_SDE_89_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_89_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_89_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_89_MUX_inst_Y), .B(KeyExpansionOutput[89]), .Z(
        KeyReg_Inst_ff_SDE_89_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_89_current_state_reg_U1 ( .A(key_shifted[97]), 
        .ZN(KeyReg_Inst_ff_SDE_89_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_89_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_89_next_state), .CK(clk), .Q(key_shifted[97]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_90_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[90]), 
        .B(key_shifted[90]), .Z(KeyReg_Inst_ff_SDE_90_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_90_MUX_inst_AND1_U1 ( .A1(KeyReg_n8), .A2(
        KeyReg_Inst_ff_SDE_90_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_90_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_90_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_90_MUX_inst_Y), .B(KeyExpansionOutput[90]), .Z(
        KeyReg_Inst_ff_SDE_90_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_90_current_state_reg_U1 ( .A(key_shifted[98]), 
        .ZN(KeyReg_Inst_ff_SDE_90_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_90_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_90_next_state), .CK(clk), .Q(key_shifted[98]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_91_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[91]), 
        .B(key_shifted[91]), .Z(KeyReg_Inst_ff_SDE_91_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_91_MUX_inst_AND1_U1 ( .A1(KeyReg_n8), .A2(
        KeyReg_Inst_ff_SDE_91_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_91_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_91_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_91_MUX_inst_Y), .B(KeyExpansionOutput[91]), .Z(
        KeyReg_Inst_ff_SDE_91_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_91_current_state_reg_U1 ( .A(key_shifted[99]), 
        .ZN(KeyReg_Inst_ff_SDE_91_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_91_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_91_next_state), .CK(clk), .Q(key_shifted[99]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_92_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[92]), 
        .B(key_shifted[92]), .Z(KeyReg_Inst_ff_SDE_92_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_92_MUX_inst_AND1_U1 ( .A1(KeyReg_n7), .A2(
        KeyReg_Inst_ff_SDE_92_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_92_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_92_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_92_MUX_inst_Y), .B(KeyExpansionOutput[92]), .Z(
        KeyReg_Inst_ff_SDE_92_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_92_current_state_reg_U1 ( .A(key_shifted[100]), 
        .ZN(KeyReg_Inst_ff_SDE_92_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_92_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_92_next_state), .CK(clk), .Q(key_shifted[100]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_93_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[93]), 
        .B(key_shifted[93]), .Z(KeyReg_Inst_ff_SDE_93_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_93_MUX_inst_AND1_U1 ( .A1(KeyReg_n7), .A2(
        KeyReg_Inst_ff_SDE_93_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_93_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_93_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_93_MUX_inst_Y), .B(KeyExpansionOutput[93]), .Z(
        KeyReg_Inst_ff_SDE_93_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_93_current_state_reg_U1 ( .A(key_shifted[101]), 
        .ZN(KeyReg_Inst_ff_SDE_93_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_93_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_93_next_state), .CK(clk), .Q(key_shifted[101]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_94_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[94]), 
        .B(key_shifted[94]), .Z(KeyReg_Inst_ff_SDE_94_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_94_MUX_inst_AND1_U1 ( .A1(KeyReg_n7), .A2(
        KeyReg_Inst_ff_SDE_94_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_94_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_94_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_94_MUX_inst_Y), .B(KeyExpansionOutput[94]), .Z(
        KeyReg_Inst_ff_SDE_94_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_94_current_state_reg_U1 ( .A(key_shifted[102]), 
        .ZN(KeyReg_Inst_ff_SDE_94_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_94_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_94_next_state), .CK(clk), .Q(key_shifted[102]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_95_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[95]), 
        .B(key_shifted[95]), .Z(KeyReg_Inst_ff_SDE_95_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_95_MUX_inst_AND1_U1 ( .A1(KeyReg_n7), .A2(
        KeyReg_Inst_ff_SDE_95_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_95_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_95_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_95_MUX_inst_Y), .B(KeyExpansionOutput[95]), .Z(
        KeyReg_Inst_ff_SDE_95_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_95_current_state_reg_U1 ( .A(key_shifted[103]), 
        .ZN(KeyReg_Inst_ff_SDE_95_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_95_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_95_next_state), .CK(clk), .Q(key_shifted[103]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_96_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[96]), 
        .B(key_shifted[96]), .Z(KeyReg_Inst_ff_SDE_96_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_96_MUX_inst_AND1_U1 ( .A1(KeyReg_n7), .A2(
        KeyReg_Inst_ff_SDE_96_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_96_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_96_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_96_MUX_inst_Y), .B(KeyExpansionOutput[96]), .Z(
        KeyReg_Inst_ff_SDE_96_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_96_current_state_reg_U1 ( .A(key_shifted[104]), 
        .ZN(KeyReg_Inst_ff_SDE_96_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_96_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_96_next_state), .CK(clk), .Q(key_shifted[104]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_97_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[97]), 
        .B(key_shifted[97]), .Z(KeyReg_Inst_ff_SDE_97_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_97_MUX_inst_AND1_U1 ( .A1(KeyReg_n7), .A2(
        KeyReg_Inst_ff_SDE_97_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_97_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_97_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_97_MUX_inst_Y), .B(KeyExpansionOutput[97]), .Z(
        KeyReg_Inst_ff_SDE_97_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_97_current_state_reg_U1 ( .A(key_shifted[105]), 
        .ZN(KeyReg_Inst_ff_SDE_97_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_97_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_97_next_state), .CK(clk), .Q(key_shifted[105]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_98_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[98]), 
        .B(key_shifted[98]), .Z(KeyReg_Inst_ff_SDE_98_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_98_MUX_inst_AND1_U1 ( .A1(KeyReg_n7), .A2(
        KeyReg_Inst_ff_SDE_98_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_98_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_98_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_98_MUX_inst_Y), .B(KeyExpansionOutput[98]), .Z(
        KeyReg_Inst_ff_SDE_98_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_98_current_state_reg_U1 ( .A(key_shifted[106]), 
        .ZN(KeyReg_Inst_ff_SDE_98_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_98_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_98_next_state), .CK(clk), .Q(key_shifted[106]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_99_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[99]), 
        .B(key_shifted[99]), .Z(KeyReg_Inst_ff_SDE_99_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_99_MUX_inst_AND1_U1 ( .A1(KeyReg_n7), .A2(
        KeyReg_Inst_ff_SDE_99_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_99_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_99_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_99_MUX_inst_Y), .B(KeyExpansionOutput[99]), .Z(
        KeyReg_Inst_ff_SDE_99_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_99_current_state_reg_U1 ( .A(key_shifted[107]), 
        .ZN(KeyReg_Inst_ff_SDE_99_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_99_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_99_next_state), .CK(clk), .Q(key_shifted[107]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_100_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[100]), .B(key_shifted[100]), .Z(KeyReg_Inst_ff_SDE_100_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_100_MUX_inst_AND1_U1 ( .A1(KeyReg_n7), .A2(
        KeyReg_Inst_ff_SDE_100_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_100_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_100_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_100_MUX_inst_Y), .B(KeyExpansionOutput[100]), .Z(
        KeyReg_Inst_ff_SDE_100_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_100_current_state_reg_U1 ( .A(key_shifted[108]), 
        .ZN(KeyReg_Inst_ff_SDE_100_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_100_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_100_next_state), .CK(clk), .Q(key_shifted[108]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_101_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[101]), .B(key_shifted[101]), .Z(KeyReg_Inst_ff_SDE_101_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_101_MUX_inst_AND1_U1 ( .A1(KeyReg_n7), .A2(
        KeyReg_Inst_ff_SDE_101_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_101_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_101_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_101_MUX_inst_Y), .B(KeyExpansionOutput[101]), .Z(
        KeyReg_Inst_ff_SDE_101_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_101_current_state_reg_U1 ( .A(key_shifted[109]), 
        .ZN(KeyReg_Inst_ff_SDE_101_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_101_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_101_next_state), .CK(clk), .Q(key_shifted[109]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_102_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[102]), .B(key_shifted[102]), .Z(KeyReg_Inst_ff_SDE_102_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_102_MUX_inst_AND1_U1 ( .A1(KeyReg_n7), .A2(
        KeyReg_Inst_ff_SDE_102_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_102_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_102_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_102_MUX_inst_Y), .B(KeyExpansionOutput[102]), .Z(
        KeyReg_Inst_ff_SDE_102_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_102_current_state_reg_U1 ( .A(key_shifted[110]), 
        .ZN(KeyReg_Inst_ff_SDE_102_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_102_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_102_next_state), .CK(clk), .Q(key_shifted[110]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_103_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[103]), .B(key_shifted[103]), .Z(KeyReg_Inst_ff_SDE_103_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_103_MUX_inst_AND1_U1 ( .A1(KeyReg_n7), .A2(
        KeyReg_Inst_ff_SDE_103_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_103_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_103_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_103_MUX_inst_Y), .B(KeyExpansionOutput[103]), .Z(
        KeyReg_Inst_ff_SDE_103_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_103_current_state_reg_U1 ( .A(key_shifted[111]), 
        .ZN(KeyReg_Inst_ff_SDE_103_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_103_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_103_next_state), .CK(clk), .Q(key_shifted[111]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_104_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[104]), .B(key_shifted[104]), .Z(KeyReg_Inst_ff_SDE_104_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_104_MUX_inst_AND1_U1 ( .A1(KeyReg_n7), .A2(
        KeyReg_Inst_ff_SDE_104_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_104_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_104_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_104_MUX_inst_Y), .B(KeyExpansionOutput[104]), .Z(
        KeyReg_Inst_ff_SDE_104_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_104_current_state_reg_U1 ( .A(key_shifted[112]), 
        .ZN(KeyReg_Inst_ff_SDE_104_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_104_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_104_next_state), .CK(clk), .Q(key_shifted[112]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_105_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[105]), .B(key_shifted[105]), .Z(KeyReg_Inst_ff_SDE_105_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_105_MUX_inst_AND1_U1 ( .A1(KeyReg_n8), .A2(
        KeyReg_Inst_ff_SDE_105_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_105_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_105_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_105_MUX_inst_Y), .B(KeyExpansionOutput[105]), .Z(
        KeyReg_Inst_ff_SDE_105_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_105_current_state_reg_U1 ( .A(key_shifted[113]), 
        .ZN(KeyReg_Inst_ff_SDE_105_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_105_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_105_next_state), .CK(clk), .Q(key_shifted[113]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_106_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[106]), .B(key_shifted[106]), .Z(KeyReg_Inst_ff_SDE_106_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_106_MUX_inst_AND1_U1 ( .A1(KeyReg_n9), .A2(
        KeyReg_Inst_ff_SDE_106_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_106_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_106_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_106_MUX_inst_Y), .B(KeyExpansionOutput[106]), .Z(
        KeyReg_Inst_ff_SDE_106_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_106_current_state_reg_U1 ( .A(key_shifted[114]), 
        .ZN(KeyReg_Inst_ff_SDE_106_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_106_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_106_next_state), .CK(clk), .Q(key_shifted[114]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_107_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[107]), .B(key_shifted[107]), .Z(KeyReg_Inst_ff_SDE_107_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_107_MUX_inst_AND1_U1 ( .A1(KeyReg_n6), .A2(
        KeyReg_Inst_ff_SDE_107_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_107_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_107_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_107_MUX_inst_Y), .B(KeyExpansionOutput[107]), .Z(
        KeyReg_Inst_ff_SDE_107_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_107_current_state_reg_U1 ( .A(key_shifted[115]), 
        .ZN(KeyReg_Inst_ff_SDE_107_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_107_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_107_next_state), .CK(clk), .Q(key_shifted[115]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_108_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[108]), .B(key_shifted[108]), .Z(KeyReg_Inst_ff_SDE_108_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_108_MUX_inst_AND1_U1 ( .A1(KeyReg_n6), .A2(
        KeyReg_Inst_ff_SDE_108_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_108_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_108_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_108_MUX_inst_Y), .B(KeyExpansionOutput[108]), .Z(
        KeyReg_Inst_ff_SDE_108_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_108_current_state_reg_U1 ( .A(key_shifted[116]), 
        .ZN(KeyReg_Inst_ff_SDE_108_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_108_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_108_next_state), .CK(clk), .Q(key_shifted[116]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_109_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[109]), .B(key_shifted[109]), .Z(KeyReg_Inst_ff_SDE_109_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_109_MUX_inst_AND1_U1 ( .A1(KeyReg_n7), .A2(
        KeyReg_Inst_ff_SDE_109_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_109_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_109_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_109_MUX_inst_Y), .B(KeyExpansionOutput[109]), .Z(
        KeyReg_Inst_ff_SDE_109_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_109_current_state_reg_U1 ( .A(key_shifted[117]), 
        .ZN(KeyReg_Inst_ff_SDE_109_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_109_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_109_next_state), .CK(clk), .Q(key_shifted[117]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_110_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[110]), .B(key_shifted[110]), .Z(KeyReg_Inst_ff_SDE_110_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_110_MUX_inst_AND1_U1 ( .A1(KeyReg_n8), .A2(
        KeyReg_Inst_ff_SDE_110_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_110_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_110_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_110_MUX_inst_Y), .B(KeyExpansionOutput[110]), .Z(
        KeyReg_Inst_ff_SDE_110_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_110_current_state_reg_U1 ( .A(key_shifted[118]), 
        .ZN(KeyReg_Inst_ff_SDE_110_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_110_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_110_next_state), .CK(clk), .Q(key_shifted[118]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_111_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[111]), .B(key_shifted[111]), .Z(KeyReg_Inst_ff_SDE_111_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_111_MUX_inst_AND1_U1 ( .A1(KeyReg_n9), .A2(
        KeyReg_Inst_ff_SDE_111_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_111_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_111_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_111_MUX_inst_Y), .B(KeyExpansionOutput[111]), .Z(
        KeyReg_Inst_ff_SDE_111_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_111_current_state_reg_U1 ( .A(key_shifted[119]), 
        .ZN(KeyReg_Inst_ff_SDE_111_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_111_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_111_next_state), .CK(clk), .Q(key_shifted[119]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_112_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[112]), .B(key_shifted[112]), .Z(KeyReg_Inst_ff_SDE_112_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_112_MUX_inst_AND1_U1 ( .A1(KeyReg_n7), .A2(
        KeyReg_Inst_ff_SDE_112_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_112_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_112_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_112_MUX_inst_Y), .B(KeyExpansionOutput[112]), .Z(
        KeyReg_Inst_ff_SDE_112_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_112_current_state_reg_U1 ( .A(key_shifted[120]), 
        .ZN(KeyReg_Inst_ff_SDE_112_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_112_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_112_next_state), .CK(clk), .Q(key_shifted[120]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_113_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[113]), .B(key_shifted[113]), .Z(KeyReg_Inst_ff_SDE_113_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_113_MUX_inst_AND1_U1 ( .A1(KeyReg_n8), .A2(
        KeyReg_Inst_ff_SDE_113_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_113_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_113_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_113_MUX_inst_Y), .B(KeyExpansionOutput[113]), .Z(
        KeyReg_Inst_ff_SDE_113_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_113_current_state_reg_U1 ( .A(key_shifted[121]), 
        .ZN(KeyReg_Inst_ff_SDE_113_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_113_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_113_next_state), .CK(clk), .Q(key_shifted[121]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_114_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[114]), .B(key_shifted[114]), .Z(KeyReg_Inst_ff_SDE_114_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_114_MUX_inst_AND1_U1 ( .A1(KeyReg_n9), .A2(
        KeyReg_Inst_ff_SDE_114_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_114_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_114_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_114_MUX_inst_Y), .B(KeyExpansionOutput[114]), .Z(
        KeyReg_Inst_ff_SDE_114_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_114_current_state_reg_U1 ( .A(key_shifted[122]), 
        .ZN(KeyReg_Inst_ff_SDE_114_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_114_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_114_next_state), .CK(clk), .Q(key_shifted[122]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_115_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[115]), .B(key_shifted[115]), .Z(KeyReg_Inst_ff_SDE_115_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_115_MUX_inst_AND1_U1 ( .A1(KeyReg_n6), .A2(
        KeyReg_Inst_ff_SDE_115_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_115_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_115_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_115_MUX_inst_Y), .B(KeyExpansionOutput[115]), .Z(
        KeyReg_Inst_ff_SDE_115_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_115_current_state_reg_U1 ( .A(key_shifted[123]), 
        .ZN(KeyReg_Inst_ff_SDE_115_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_115_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_115_next_state), .CK(clk), .Q(key_shifted[123]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_116_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[116]), .B(key_shifted[116]), .Z(KeyReg_Inst_ff_SDE_116_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_116_MUX_inst_AND1_U1 ( .A1(KeyReg_n6), .A2(
        KeyReg_Inst_ff_SDE_116_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_116_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_116_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_116_MUX_inst_Y), .B(KeyExpansionOutput[116]), .Z(
        KeyReg_Inst_ff_SDE_116_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_116_current_state_reg_U1 ( .A(key_shifted[124]), 
        .ZN(KeyReg_Inst_ff_SDE_116_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_116_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_116_next_state), .CK(clk), .Q(key_shifted[124]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_117_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[117]), .B(key_shifted[117]), .Z(KeyReg_Inst_ff_SDE_117_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_117_MUX_inst_AND1_U1 ( .A1(KeyReg_n6), .A2(
        KeyReg_Inst_ff_SDE_117_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_117_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_117_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_117_MUX_inst_Y), .B(KeyExpansionOutput[117]), .Z(
        KeyReg_Inst_ff_SDE_117_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_117_current_state_reg_U1 ( .A(key_shifted[125]), 
        .ZN(KeyReg_Inst_ff_SDE_117_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_117_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_117_next_state), .CK(clk), .Q(key_shifted[125]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_118_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[118]), .B(key_shifted[118]), .Z(KeyReg_Inst_ff_SDE_118_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_118_MUX_inst_AND1_U1 ( .A1(KeyReg_n6), .A2(
        KeyReg_Inst_ff_SDE_118_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_118_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_118_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_118_MUX_inst_Y), .B(KeyExpansionOutput[118]), .Z(
        KeyReg_Inst_ff_SDE_118_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_118_current_state_reg_U1 ( .A(key_shifted[126]), 
        .ZN(KeyReg_Inst_ff_SDE_118_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_118_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_118_next_state), .CK(clk), .Q(key_shifted[126]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_119_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[119]), .B(key_shifted[119]), .Z(KeyReg_Inst_ff_SDE_119_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_119_MUX_inst_AND1_U1 ( .A1(KeyReg_n6), .A2(
        KeyReg_Inst_ff_SDE_119_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_119_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_119_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_119_MUX_inst_Y), .B(KeyExpansionOutput[119]), .Z(
        KeyReg_Inst_ff_SDE_119_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_119_current_state_reg_U1 ( .A(key_shifted[127]), 
        .ZN(KeyReg_Inst_ff_SDE_119_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_119_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_119_next_state), .CK(clk), .Q(key_shifted[127]), 
        .QN() );
  XOR2_X1 KeyReg_Inst_ff_SDE_120_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[120]), .B(key_shifted[120]), .Z(KeyReg_Inst_ff_SDE_120_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_120_MUX_inst_AND1_U1 ( .A1(KeyReg_n6), .A2(
        KeyReg_Inst_ff_SDE_120_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_120_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_120_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_120_MUX_inst_Y), .B(KeyExpansionOutput[120]), .Z(
        KeyReg_Inst_ff_SDE_120_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_120_current_state_reg_U1 ( .A(RoundKey[120]), .ZN(
        KeyReg_Inst_ff_SDE_120_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_120_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_120_next_state), .CK(clk), .Q(RoundKey[120]), .QN()
         );
  XOR2_X1 KeyReg_Inst_ff_SDE_121_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[121]), .B(key_shifted[121]), .Z(KeyReg_Inst_ff_SDE_121_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_121_MUX_inst_AND1_U1 ( .A1(KeyReg_n6), .A2(
        KeyReg_Inst_ff_SDE_121_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_121_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_121_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_121_MUX_inst_Y), .B(KeyExpansionOutput[121]), .Z(
        KeyReg_Inst_ff_SDE_121_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_121_current_state_reg_U1 ( .A(RoundKey[121]), .ZN(
        KeyReg_Inst_ff_SDE_121_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_121_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_121_next_state), .CK(clk), .Q(RoundKey[121]), .QN()
         );
  XOR2_X1 KeyReg_Inst_ff_SDE_122_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[122]), .B(key_shifted[122]), .Z(KeyReg_Inst_ff_SDE_122_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_122_MUX_inst_AND1_U1 ( .A1(KeyReg_n6), .A2(
        KeyReg_Inst_ff_SDE_122_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_122_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_122_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_122_MUX_inst_Y), .B(KeyExpansionOutput[122]), .Z(
        KeyReg_Inst_ff_SDE_122_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_122_current_state_reg_U1 ( .A(RoundKey[122]), .ZN(
        KeyReg_Inst_ff_SDE_122_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_122_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_122_next_state), .CK(clk), .Q(RoundKey[122]), .QN()
         );
  XOR2_X1 KeyReg_Inst_ff_SDE_123_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[123]), .B(key_shifted[123]), .Z(KeyReg_Inst_ff_SDE_123_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_123_MUX_inst_AND1_U1 ( .A1(KeyReg_n6), .A2(
        KeyReg_Inst_ff_SDE_123_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_123_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_123_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_123_MUX_inst_Y), .B(KeyExpansionOutput[123]), .Z(
        KeyReg_Inst_ff_SDE_123_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_123_current_state_reg_U1 ( .A(RoundKey[123]), .ZN(
        KeyReg_Inst_ff_SDE_123_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_123_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_123_next_state), .CK(clk), .Q(RoundKey[123]), .QN()
         );
  XOR2_X1 KeyReg_Inst_ff_SDE_124_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[124]), .B(key_shifted[124]), .Z(KeyReg_Inst_ff_SDE_124_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_124_MUX_inst_AND1_U1 ( .A1(KeyReg_n6), .A2(
        KeyReg_Inst_ff_SDE_124_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_124_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_124_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_124_MUX_inst_Y), .B(KeyExpansionOutput[124]), .Z(
        KeyReg_Inst_ff_SDE_124_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_124_current_state_reg_U1 ( .A(RoundKey[124]), .ZN(
        KeyReg_Inst_ff_SDE_124_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_124_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_124_next_state), .CK(clk), .Q(RoundKey[124]), .QN()
         );
  XOR2_X1 KeyReg_Inst_ff_SDE_125_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[125]), .B(key_shifted[125]), .Z(KeyReg_Inst_ff_SDE_125_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_125_MUX_inst_AND1_U1 ( .A1(KeyReg_n6), .A2(
        KeyReg_Inst_ff_SDE_125_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_125_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_125_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_125_MUX_inst_Y), .B(KeyExpansionOutput[125]), .Z(
        KeyReg_Inst_ff_SDE_125_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_125_current_state_reg_U1 ( .A(RoundKey[125]), .ZN(
        KeyReg_Inst_ff_SDE_125_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_125_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_125_next_state), .CK(clk), .Q(RoundKey[125]), .QN()
         );
  XOR2_X1 KeyReg_Inst_ff_SDE_126_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[126]), .B(key_shifted[126]), .Z(KeyReg_Inst_ff_SDE_126_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_126_MUX_inst_AND1_U1 ( .A1(KeyReg_n6), .A2(
        KeyReg_Inst_ff_SDE_126_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_126_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_126_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_126_MUX_inst_Y), .B(KeyExpansionOutput[126]), .Z(
        KeyReg_Inst_ff_SDE_126_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_126_current_state_reg_U1 ( .A(RoundKey[126]), .ZN(
        KeyReg_Inst_ff_SDE_126_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_126_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_126_next_state), .CK(clk), .Q(RoundKey[126]), .QN()
         );
  XOR2_X1 KeyReg_Inst_ff_SDE_127_MUX_inst_XOR1_U1 ( .A(KeyExpansionOutput[127]), .B(key_shifted[127]), .Z(KeyReg_Inst_ff_SDE_127_MUX_inst_X) );
  AND2_X1 KeyReg_Inst_ff_SDE_127_MUX_inst_AND1_U1 ( .A1(KeyReg_n6), .A2(
        KeyReg_Inst_ff_SDE_127_MUX_inst_X), .ZN(
        KeyReg_Inst_ff_SDE_127_MUX_inst_Y) );
  XOR2_X1 KeyReg_Inst_ff_SDE_127_MUX_inst_XOR2_U1 ( .A(
        KeyReg_Inst_ff_SDE_127_MUX_inst_Y), .B(KeyExpansionOutput[127]), .Z(
        KeyReg_Inst_ff_SDE_127_next_state) );
  INV_X1 KeyReg_Inst_ff_SDE_127_current_state_reg_U1 ( .A(RoundKey[127]), .ZN(
        KeyReg_Inst_ff_SDE_127_current_state_reg_QN) );
  DFF_X1 KeyReg_Inst_ff_SDE_127_current_state_reg_FF_FF ( .D(
        KeyReg_Inst_ff_SDE_127_next_state), .CK(clk), .Q(RoundKey[127]), .QN()
         );
  XOR2_X1 KeyExpansionIns_U128 ( .A(key_shifted[17]), .B(
        KeyExpansionOutput[41]), .Z(KeyExpansionOutput[9]) );
  XOR2_X1 KeyExpansionIns_U127 ( .A(key_shifted[16]), .B(
        KeyExpansionOutput[40]), .Z(KeyExpansionOutput[8]) );
  XOR2_X1 KeyExpansionIns_U126 ( .A(key_shifted[15]), .B(
        KeyExpansionOutput[39]), .Z(KeyExpansionOutput[7]) );
  XOR2_X1 KeyExpansionIns_U125 ( .A(key_shifted[14]), .B(
        KeyExpansionOutput[38]), .Z(KeyExpansionOutput[6]) );
  XOR2_X1 KeyExpansionIns_U124 ( .A(key_shifted[13]), .B(
        KeyExpansionOutput[37]), .Z(KeyExpansionOutput[5]) );
  XOR2_X1 KeyExpansionIns_U123 ( .A(key_shifted[12]), .B(
        KeyExpansionOutput[36]), .Z(KeyExpansionOutput[4]) );
  XOR2_X1 KeyExpansionIns_U122 ( .A(key_shifted[49]), .B(
        KeyExpansionOutput[73]), .Z(KeyExpansionOutput[41]) );
  XOR2_X1 KeyExpansionIns_U121 ( .A(key_shifted[81]), .B(
        KeyExpansionOutput[105]), .Z(KeyExpansionOutput[73]) );
  XOR2_X1 KeyExpansionIns_U120 ( .A(key_shifted[48]), .B(
        KeyExpansionOutput[72]), .Z(KeyExpansionOutput[40]) );
  XOR2_X1 KeyExpansionIns_U119 ( .A(key_shifted[80]), .B(
        KeyExpansionOutput[104]), .Z(KeyExpansionOutput[72]) );
  XOR2_X1 KeyExpansionIns_U118 ( .A(key_shifted[11]), .B(
        KeyExpansionOutput[35]), .Z(KeyExpansionOutput[3]) );
  XOR2_X1 KeyExpansionIns_U117 ( .A(key_shifted[47]), .B(
        KeyExpansionOutput[71]), .Z(KeyExpansionOutput[39]) );
  XOR2_X1 KeyExpansionIns_U116 ( .A(key_shifted[79]), .B(
        KeyExpansionOutput[103]), .Z(KeyExpansionOutput[71]) );
  XOR2_X1 KeyExpansionIns_U115 ( .A(key_shifted[46]), .B(
        KeyExpansionOutput[70]), .Z(KeyExpansionOutput[38]) );
  XOR2_X1 KeyExpansionIns_U114 ( .A(key_shifted[78]), .B(
        KeyExpansionOutput[102]), .Z(KeyExpansionOutput[70]) );
  XOR2_X1 KeyExpansionIns_U113 ( .A(key_shifted[45]), .B(
        KeyExpansionOutput[69]), .Z(KeyExpansionOutput[37]) );
  XOR2_X1 KeyExpansionIns_U112 ( .A(key_shifted[77]), .B(
        KeyExpansionOutput[101]), .Z(KeyExpansionOutput[69]) );
  XOR2_X1 KeyExpansionIns_U111 ( .A(key_shifted[44]), .B(
        KeyExpansionOutput[68]), .Z(KeyExpansionOutput[36]) );
  XOR2_X1 KeyExpansionIns_U110 ( .A(key_shifted[76]), .B(
        KeyExpansionOutput[100]), .Z(KeyExpansionOutput[68]) );
  XOR2_X1 KeyExpansionIns_U109 ( .A(key_shifted[43]), .B(
        KeyExpansionOutput[67]), .Z(KeyExpansionOutput[35]) );
  XOR2_X1 KeyExpansionIns_U108 ( .A(key_shifted[75]), .B(
        KeyExpansionOutput[99]), .Z(KeyExpansionOutput[67]) );
  XOR2_X1 KeyExpansionIns_U107 ( .A(key_shifted[107]), .B(
        KeyExpansionIns_tmp[3]), .Z(KeyExpansionOutput[99]) );
  XOR2_X1 KeyExpansionIns_U106 ( .A(key_shifted[39]), .B(
        KeyExpansionOutput[63]), .Z(KeyExpansionOutput[31]) );
  XOR2_X1 KeyExpansionIns_U105 ( .A(key_shifted[71]), .B(
        KeyExpansionOutput[95]), .Z(KeyExpansionOutput[63]) );
  XOR2_X1 KeyExpansionIns_U104 ( .A(key_shifted[103]), .B(
        KeyExpansionOutput[127]), .Z(KeyExpansionOutput[95]) );
  XOR2_X1 KeyExpansionIns_U103 ( .A(key_shifted[38]), .B(
        KeyExpansionOutput[62]), .Z(KeyExpansionOutput[30]) );
  XOR2_X1 KeyExpansionIns_U102 ( .A(key_shifted[70]), .B(
        KeyExpansionOutput[94]), .Z(KeyExpansionOutput[62]) );
  XOR2_X1 KeyExpansionIns_U101 ( .A(key_shifted[102]), .B(
        KeyExpansionOutput[126]), .Z(KeyExpansionOutput[94]) );
  XOR2_X1 KeyExpansionIns_U100 ( .A(key_shifted[10]), .B(
        KeyExpansionOutput[34]), .Z(KeyExpansionOutput[2]) );
  XOR2_X1 KeyExpansionIns_U99 ( .A(key_shifted[42]), .B(KeyExpansionOutput[66]), .Z(KeyExpansionOutput[34]) );
  XOR2_X1 KeyExpansionIns_U98 ( .A(key_shifted[74]), .B(KeyExpansionOutput[98]), .Z(KeyExpansionOutput[66]) );
  XOR2_X1 KeyExpansionIns_U97 ( .A(key_shifted[106]), .B(
        KeyExpansionIns_tmp[2]), .Z(KeyExpansionOutput[98]) );
  XOR2_X1 KeyExpansionIns_U96 ( .A(key_shifted[37]), .B(KeyExpansionOutput[61]), .Z(KeyExpansionOutput[29]) );
  XOR2_X1 KeyExpansionIns_U95 ( .A(key_shifted[69]), .B(KeyExpansionOutput[93]), .Z(KeyExpansionOutput[61]) );
  XOR2_X1 KeyExpansionIns_U94 ( .A(key_shifted[101]), .B(
        KeyExpansionOutput[125]), .Z(KeyExpansionOutput[93]) );
  XOR2_X1 KeyExpansionIns_U93 ( .A(key_shifted[36]), .B(KeyExpansionOutput[60]), .Z(KeyExpansionOutput[28]) );
  XOR2_X1 KeyExpansionIns_U92 ( .A(key_shifted[68]), .B(KeyExpansionOutput[92]), .Z(KeyExpansionOutput[60]) );
  XOR2_X1 KeyExpansionIns_U91 ( .A(key_shifted[100]), .B(
        KeyExpansionOutput[124]), .Z(KeyExpansionOutput[92]) );
  XOR2_X1 KeyExpansionIns_U90 ( .A(key_shifted[35]), .B(KeyExpansionOutput[59]), .Z(KeyExpansionOutput[27]) );
  XOR2_X1 KeyExpansionIns_U89 ( .A(key_shifted[67]), .B(KeyExpansionOutput[91]), .Z(KeyExpansionOutput[59]) );
  XOR2_X1 KeyExpansionIns_U88 ( .A(key_shifted[99]), .B(
        KeyExpansionOutput[123]), .Z(KeyExpansionOutput[91]) );
  XOR2_X1 KeyExpansionIns_U87 ( .A(key_shifted[34]), .B(KeyExpansionOutput[58]), .Z(KeyExpansionOutput[26]) );
  XOR2_X1 KeyExpansionIns_U86 ( .A(key_shifted[66]), .B(KeyExpansionOutput[90]), .Z(KeyExpansionOutput[58]) );
  XOR2_X1 KeyExpansionIns_U85 ( .A(key_shifted[98]), .B(
        KeyExpansionOutput[122]), .Z(KeyExpansionOutput[90]) );
  XOR2_X1 KeyExpansionIns_U84 ( .A(key_shifted[33]), .B(KeyExpansionOutput[57]), .Z(KeyExpansionOutput[25]) );
  XOR2_X1 KeyExpansionIns_U83 ( .A(key_shifted[65]), .B(KeyExpansionOutput[89]), .Z(KeyExpansionOutput[57]) );
  XOR2_X1 KeyExpansionIns_U82 ( .A(key_shifted[97]), .B(
        KeyExpansionOutput[121]), .Z(KeyExpansionOutput[89]) );
  XOR2_X1 KeyExpansionIns_U81 ( .A(key_shifted[32]), .B(KeyExpansionOutput[56]), .Z(KeyExpansionOutput[24]) );
  XOR2_X1 KeyExpansionIns_U80 ( .A(key_shifted[64]), .B(KeyExpansionOutput[88]), .Z(KeyExpansionOutput[56]) );
  XOR2_X1 KeyExpansionIns_U79 ( .A(key_shifted[96]), .B(
        KeyExpansionOutput[120]), .Z(KeyExpansionOutput[88]) );
  XOR2_X1 KeyExpansionIns_U78 ( .A(key_shifted[31]), .B(KeyExpansionOutput[55]), .Z(KeyExpansionOutput[23]) );
  XOR2_X1 KeyExpansionIns_U77 ( .A(key_shifted[63]), .B(KeyExpansionOutput[87]), .Z(KeyExpansionOutput[55]) );
  XOR2_X1 KeyExpansionIns_U76 ( .A(key_shifted[95]), .B(
        KeyExpansionOutput[119]), .Z(KeyExpansionOutput[87]) );
  XOR2_X1 KeyExpansionIns_U75 ( .A(key_shifted[30]), .B(KeyExpansionOutput[54]), .Z(KeyExpansionOutput[22]) );
  XOR2_X1 KeyExpansionIns_U74 ( .A(key_shifted[62]), .B(KeyExpansionOutput[86]), .Z(KeyExpansionOutput[54]) );
  XOR2_X1 KeyExpansionIns_U73 ( .A(key_shifted[94]), .B(
        KeyExpansionOutput[118]), .Z(KeyExpansionOutput[86]) );
  XOR2_X1 KeyExpansionIns_U72 ( .A(key_shifted[29]), .B(KeyExpansionOutput[53]), .Z(KeyExpansionOutput[21]) );
  XOR2_X1 KeyExpansionIns_U71 ( .A(key_shifted[61]), .B(KeyExpansionOutput[85]), .Z(KeyExpansionOutput[53]) );
  XOR2_X1 KeyExpansionIns_U70 ( .A(key_shifted[93]), .B(
        KeyExpansionOutput[117]), .Z(KeyExpansionOutput[85]) );
  XOR2_X1 KeyExpansionIns_U69 ( .A(key_shifted[28]), .B(KeyExpansionOutput[52]), .Z(KeyExpansionOutput[20]) );
  XOR2_X1 KeyExpansionIns_U68 ( .A(key_shifted[60]), .B(KeyExpansionOutput[84]), .Z(KeyExpansionOutput[52]) );
  XOR2_X1 KeyExpansionIns_U67 ( .A(key_shifted[92]), .B(
        KeyExpansionOutput[116]), .Z(KeyExpansionOutput[84]) );
  XOR2_X1 KeyExpansionIns_U66 ( .A(key_shifted[9]), .B(KeyExpansionOutput[33]), 
        .Z(KeyExpansionOutput[1]) );
  XOR2_X1 KeyExpansionIns_U65 ( .A(key_shifted[41]), .B(KeyExpansionOutput[65]), .Z(KeyExpansionOutput[33]) );
  XOR2_X1 KeyExpansionIns_U64 ( .A(key_shifted[73]), .B(KeyExpansionOutput[97]), .Z(KeyExpansionOutput[65]) );
  XOR2_X1 KeyExpansionIns_U63 ( .A(key_shifted[105]), .B(
        KeyExpansionIns_tmp[1]), .Z(KeyExpansionOutput[97]) );
  XOR2_X1 KeyExpansionIns_U62 ( .A(key_shifted[27]), .B(KeyExpansionOutput[51]), .Z(KeyExpansionOutput[19]) );
  XOR2_X1 KeyExpansionIns_U61 ( .A(key_shifted[59]), .B(KeyExpansionOutput[83]), .Z(KeyExpansionOutput[51]) );
  XOR2_X1 KeyExpansionIns_U60 ( .A(key_shifted[91]), .B(
        KeyExpansionOutput[115]), .Z(KeyExpansionOutput[83]) );
  XOR2_X1 KeyExpansionIns_U59 ( .A(key_shifted[26]), .B(KeyExpansionOutput[50]), .Z(KeyExpansionOutput[18]) );
  XOR2_X1 KeyExpansionIns_U58 ( .A(key_shifted[58]), .B(KeyExpansionOutput[82]), .Z(KeyExpansionOutput[50]) );
  XOR2_X1 KeyExpansionIns_U57 ( .A(key_shifted[90]), .B(
        KeyExpansionOutput[114]), .Z(KeyExpansionOutput[82]) );
  XOR2_X1 KeyExpansionIns_U56 ( .A(key_shifted[25]), .B(KeyExpansionOutput[49]), .Z(KeyExpansionOutput[17]) );
  XOR2_X1 KeyExpansionIns_U55 ( .A(key_shifted[57]), .B(KeyExpansionOutput[81]), .Z(KeyExpansionOutput[49]) );
  XOR2_X1 KeyExpansionIns_U54 ( .A(key_shifted[89]), .B(
        KeyExpansionOutput[113]), .Z(KeyExpansionOutput[81]) );
  XOR2_X1 KeyExpansionIns_U53 ( .A(key_shifted[24]), .B(KeyExpansionOutput[48]), .Z(KeyExpansionOutput[16]) );
  XOR2_X1 KeyExpansionIns_U52 ( .A(key_shifted[56]), .B(KeyExpansionOutput[80]), .Z(KeyExpansionOutput[48]) );
  XOR2_X1 KeyExpansionIns_U51 ( .A(key_shifted[88]), .B(
        KeyExpansionOutput[112]), .Z(KeyExpansionOutput[80]) );
  XOR2_X1 KeyExpansionIns_U50 ( .A(key_shifted[23]), .B(KeyExpansionOutput[47]), .Z(KeyExpansionOutput[15]) );
  XOR2_X1 KeyExpansionIns_U49 ( .A(key_shifted[55]), .B(KeyExpansionOutput[79]), .Z(KeyExpansionOutput[47]) );
  XOR2_X1 KeyExpansionIns_U48 ( .A(key_shifted[87]), .B(
        KeyExpansionOutput[111]), .Z(KeyExpansionOutput[79]) );
  XOR2_X1 KeyExpansionIns_U47 ( .A(key_shifted[22]), .B(KeyExpansionOutput[46]), .Z(KeyExpansionOutput[14]) );
  XOR2_X1 KeyExpansionIns_U46 ( .A(key_shifted[54]), .B(KeyExpansionOutput[78]), .Z(KeyExpansionOutput[46]) );
  XOR2_X1 KeyExpansionIns_U45 ( .A(key_shifted[86]), .B(
        KeyExpansionOutput[110]), .Z(KeyExpansionOutput[78]) );
  XOR2_X1 KeyExpansionIns_U44 ( .A(key_shifted[21]), .B(KeyExpansionOutput[45]), .Z(KeyExpansionOutput[13]) );
  XOR2_X1 KeyExpansionIns_U43 ( .A(key_shifted[53]), .B(KeyExpansionOutput[77]), .Z(KeyExpansionOutput[45]) );
  XOR2_X1 KeyExpansionIns_U42 ( .A(key_shifted[85]), .B(
        KeyExpansionOutput[109]), .Z(KeyExpansionOutput[77]) );
  XOR2_X1 KeyExpansionIns_U41 ( .A(key_shifted[20]), .B(KeyExpansionOutput[44]), .Z(KeyExpansionOutput[12]) );
  XOR2_X1 KeyExpansionIns_U40 ( .A(key_shifted[52]), .B(KeyExpansionOutput[76]), .Z(KeyExpansionOutput[44]) );
  XOR2_X1 KeyExpansionIns_U39 ( .A(key_shifted[84]), .B(
        KeyExpansionOutput[108]), .Z(KeyExpansionOutput[76]) );
  XOR2_X1 KeyExpansionIns_U38 ( .A(RoundKey[127]), .B(KeyExpansionIns_tmp[31]), 
        .Z(KeyExpansionOutput[127]) );
  XOR2_X1 KeyExpansionIns_U37 ( .A(RoundKey[126]), .B(KeyExpansionIns_tmp[30]), 
        .Z(KeyExpansionOutput[126]) );
  XOR2_X1 KeyExpansionIns_U36 ( .A(RoundKey[125]), .B(KeyExpansionIns_tmp[29]), 
        .Z(KeyExpansionOutput[125]) );
  XOR2_X1 KeyExpansionIns_U35 ( .A(RoundKey[124]), .B(KeyExpansionIns_tmp[28]), 
        .Z(KeyExpansionOutput[124]) );
  XOR2_X1 KeyExpansionIns_U34 ( .A(RoundKey[123]), .B(KeyExpansionIns_tmp[27]), 
        .Z(KeyExpansionOutput[123]) );
  XOR2_X1 KeyExpansionIns_U33 ( .A(RoundKey[122]), .B(KeyExpansionIns_tmp[26]), 
        .Z(KeyExpansionOutput[122]) );
  XOR2_X1 KeyExpansionIns_U32 ( .A(RoundKey[121]), .B(KeyExpansionIns_tmp[25]), 
        .Z(KeyExpansionOutput[121]) );
  XOR2_X1 KeyExpansionIns_U31 ( .A(RoundKey[120]), .B(KeyExpansionIns_tmp[24]), 
        .Z(KeyExpansionOutput[120]) );
  XOR2_X1 KeyExpansionIns_U30 ( .A(key_shifted[19]), .B(KeyExpansionOutput[43]), .Z(KeyExpansionOutput[11]) );
  XOR2_X1 KeyExpansionIns_U29 ( .A(key_shifted[51]), .B(KeyExpansionOutput[75]), .Z(KeyExpansionOutput[43]) );
  XOR2_X1 KeyExpansionIns_U28 ( .A(key_shifted[83]), .B(
        KeyExpansionOutput[107]), .Z(KeyExpansionOutput[75]) );
  XOR2_X1 KeyExpansionIns_U27 ( .A(key_shifted[127]), .B(
        KeyExpansionIns_tmp[23]), .Z(KeyExpansionOutput[119]) );
  XOR2_X1 KeyExpansionIns_U26 ( .A(key_shifted[126]), .B(
        KeyExpansionIns_tmp[22]), .Z(KeyExpansionOutput[118]) );
  XOR2_X1 KeyExpansionIns_U25 ( .A(key_shifted[125]), .B(
        KeyExpansionIns_tmp[21]), .Z(KeyExpansionOutput[117]) );
  XOR2_X1 KeyExpansionIns_U24 ( .A(key_shifted[124]), .B(
        KeyExpansionIns_tmp[20]), .Z(KeyExpansionOutput[116]) );
  XOR2_X1 KeyExpansionIns_U23 ( .A(key_shifted[123]), .B(
        KeyExpansionIns_tmp[19]), .Z(KeyExpansionOutput[115]) );
  XOR2_X1 KeyExpansionIns_U22 ( .A(key_shifted[122]), .B(
        KeyExpansionIns_tmp[18]), .Z(KeyExpansionOutput[114]) );
  XOR2_X1 KeyExpansionIns_U21 ( .A(key_shifted[121]), .B(
        KeyExpansionIns_tmp[17]), .Z(KeyExpansionOutput[113]) );
  XOR2_X1 KeyExpansionIns_U20 ( .A(key_shifted[120]), .B(
        KeyExpansionIns_tmp[16]), .Z(KeyExpansionOutput[112]) );
  XOR2_X1 KeyExpansionIns_U19 ( .A(key_shifted[119]), .B(
        KeyExpansionIns_tmp[15]), .Z(KeyExpansionOutput[111]) );
  XOR2_X1 KeyExpansionIns_U18 ( .A(key_shifted[118]), .B(
        KeyExpansionIns_tmp[14]), .Z(KeyExpansionOutput[110]) );
  XOR2_X1 KeyExpansionIns_U17 ( .A(key_shifted[18]), .B(KeyExpansionOutput[42]), .Z(KeyExpansionOutput[10]) );
  XOR2_X1 KeyExpansionIns_U16 ( .A(key_shifted[50]), .B(KeyExpansionOutput[74]), .Z(KeyExpansionOutput[42]) );
  XOR2_X1 KeyExpansionIns_U15 ( .A(key_shifted[82]), .B(
        KeyExpansionOutput[106]), .Z(KeyExpansionOutput[74]) );
  XOR2_X1 KeyExpansionIns_U14 ( .A(key_shifted[117]), .B(
        KeyExpansionIns_tmp[13]), .Z(KeyExpansionOutput[109]) );
  XOR2_X1 KeyExpansionIns_U13 ( .A(key_shifted[116]), .B(
        KeyExpansionIns_tmp[12]), .Z(KeyExpansionOutput[108]) );
  XOR2_X1 KeyExpansionIns_U12 ( .A(key_shifted[115]), .B(
        KeyExpansionIns_tmp[11]), .Z(KeyExpansionOutput[107]) );
  XOR2_X1 KeyExpansionIns_U11 ( .A(key_shifted[114]), .B(
        KeyExpansionIns_tmp[10]), .Z(KeyExpansionOutput[106]) );
  XOR2_X1 KeyExpansionIns_U10 ( .A(key_shifted[113]), .B(
        KeyExpansionIns_tmp[9]), .Z(KeyExpansionOutput[105]) );
  XOR2_X1 KeyExpansionIns_U9 ( .A(key_shifted[112]), .B(KeyExpansionIns_tmp[8]), .Z(KeyExpansionOutput[104]) );
  XOR2_X1 KeyExpansionIns_U8 ( .A(key_shifted[111]), .B(KeyExpansionIns_tmp[7]), .Z(KeyExpansionOutput[103]) );
  XOR2_X1 KeyExpansionIns_U7 ( .A(key_shifted[110]), .B(KeyExpansionIns_tmp[6]), .Z(KeyExpansionOutput[102]) );
  XOR2_X1 KeyExpansionIns_U6 ( .A(key_shifted[109]), .B(KeyExpansionIns_tmp[5]), .Z(KeyExpansionOutput[101]) );
  XOR2_X1 KeyExpansionIns_U5 ( .A(key_shifted[108]), .B(KeyExpansionIns_tmp[4]), .Z(KeyExpansionOutput[100]) );
  XOR2_X1 KeyExpansionIns_U4 ( .A(key_shifted[8]), .B(KeyExpansionOutput[32]), 
        .Z(KeyExpansionOutput[0]) );
  XOR2_X1 KeyExpansionIns_U3 ( .A(key_shifted[40]), .B(KeyExpansionOutput[64]), 
        .Z(KeyExpansionOutput[32]) );
  XOR2_X1 KeyExpansionIns_U2 ( .A(key_shifted[72]), .B(KeyExpansionOutput[96]), 
        .Z(KeyExpansionOutput[64]) );
  XOR2_X1 KeyExpansionIns_U1 ( .A(key_shifted[104]), .B(KeyExpansionIns_tmp[0]), .Z(KeyExpansionOutput[96]) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_U8 ( .A(
        KeyExpansionIns_KeySchedCoreInst_OutBytes_0__7_), .B(n286), .Z(
        KeyExpansionIns_tmp[31]) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_U7 ( .A(
        KeyExpansionIns_KeySchedCoreInst_OutBytes_0__6_), .B(n287), .Z(
        KeyExpansionIns_tmp[30]) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_U6 ( .A(
        KeyExpansionIns_KeySchedCoreInst_OutBytes_0__5_), .B(Rcon[5]), .Z(
        KeyExpansionIns_tmp[29]) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_U5 ( .A(
        KeyExpansionIns_KeySchedCoreInst_OutBytes_0__4_), .B(Rcon[4]), .Z(
        KeyExpansionIns_tmp[28]) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_U4 ( .A(
        KeyExpansionIns_KeySchedCoreInst_OutBytes_0__3_), .B(Rcon[3]), .Z(
        KeyExpansionIns_tmp[27]) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_U3 ( .A(
        KeyExpansionIns_KeySchedCoreInst_OutBytes_0__2_), .B(Rcon[2]), .Z(
        KeyExpansionIns_tmp[26]) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_U2 ( .A(
        KeyExpansionIns_KeySchedCoreInst_OutBytes_0__1_), .B(Rcon[1]), .Z(
        KeyExpansionIns_tmp[25]) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_OutBytes_0__0_), .B(Rcon[0]), .Z(
        KeyExpansionIns_tmp[24]) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T1_U1 ( .A(
        key_shifted[31]), .B(key_shifted[28]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T2_U1 ( .A(
        key_shifted[31]), .B(key_shifted[26]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T2) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T3_U1 ( .A(
        key_shifted[31]), .B(key_shifted[25]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T3) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T4_U1 ( .A(
        key_shifted[28]), .B(key_shifted[26]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T4) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T5_U1 ( .A(
        key_shifted[27]), .B(key_shifted[25]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T5) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T6_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T5), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T7_U1 ( .A(
        key_shifted[30]), .B(key_shifted[29]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T7) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T8_U1 ( .A(
        key_shifted[24]), .B(KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6), 
        .Z(KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T8) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T9_U1 ( .A(
        key_shifted[24]), .B(KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T7), 
        .Z(KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T9) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T10_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T7), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T10) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T11_U1 ( .A(
        key_shifted[30]), .B(key_shifted[26]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T11) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T12_U1 ( .A(
        key_shifted[29]), .B(key_shifted[26]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T12) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T13_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T3), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T4), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T13) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T14_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T11), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T14) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T15_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T5), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T11), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T15) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T16_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T5), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T12), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T16) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T17_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T9), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T16), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T17) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T18_U1 ( .A(
        key_shifted[28]), .B(key_shifted[24]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T18) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T19_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T7), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T18), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T19) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T20_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T19), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T20) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T21_U1 ( .A(
        key_shifted[25]), .B(key_shifted[24]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T21) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T22_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T7), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T21), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T22) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T23_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T2), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T22), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T23) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T24_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T2), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T10), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T24) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T25_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T20), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T17), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T25) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T26_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T3), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T16), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T26) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T27_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T12), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T27) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M1_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T13), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M1) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M2_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T23), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T8), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M2) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M3_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T14), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M1), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M3) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M4_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T19), .A2(key_shifted[24]), .ZN(KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M4) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M5_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M4), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M1), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M5) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M6_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T3), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T16), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M6) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M7_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T22), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T9), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M7) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M8_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T26), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M6), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M8) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M9_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T20), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T17), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M9) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M10_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M9), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M6), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M10) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M11_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T15), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M11) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M12_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T4), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T27), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M12) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M13_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M12), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M11), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M13) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M14_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T2), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T10), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M14) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M15_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M14), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M11), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M15) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M16_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M3), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M2), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M16) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M17_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M5), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T24), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M17) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M18_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M8), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M7), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M18) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M19_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M10), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M15), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M19) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M20_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M16), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M13), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M20) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M21_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M17), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M15), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M21) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M22_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M18), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M13), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M22) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M23_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M19), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T25), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M23) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M24_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M22), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M23), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M24) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M25_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M22), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M20), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M25) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M26_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M21), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M25), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M26) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M27_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M20), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M21), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M27) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M28_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M23), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M25), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M28) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M29_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M28), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M27), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M29) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M30_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M26), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M24), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M30) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M31_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M20), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M23), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M31) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M32_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M27), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M31), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M32) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M33_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M27), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M25), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M33) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M34_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M21), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M22), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M34) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M35_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M24), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M34), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M35) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M36_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M24), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M25), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M36) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M37_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M21), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M29), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M37) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M38_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M32), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M33), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M38) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M39_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M23), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M30), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M39) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M40_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M35), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M36), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M40) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M41_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M38), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M40), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M41) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M42_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M37), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M39), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M42) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M43_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M37), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M38), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M43) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M44_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M39), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M40), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M44) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M45_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M42), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M41), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M45) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M46_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M44), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M46) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M47_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M40), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T8), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M47) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M48_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M39), .A2(key_shifted[24]), .ZN(KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M48) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M49_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M43), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T16), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M49) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M50_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M38), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T9), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M50) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M51_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M37), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T17), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M51) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M52_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M42), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T15), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M52) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M53_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M45), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T27), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M53) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M54_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M41), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T10), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M54) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M55_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M44), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T13), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M55) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M56_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M40), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T23), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M56) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M57_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M39), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T19), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M57) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M58_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M43), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T3), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M58) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M59_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M38), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T22), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M59) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M60_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M37), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T20), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M60) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M61_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M42), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M61) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M62_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M45), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T4), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M62) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M63_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M41), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T2), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M63) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L0_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M61), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M62), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L0) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L1_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M50), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M56), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L1) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L2_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M46), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M48), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L2) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L3_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M47), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M55), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L3) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L4_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M54), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M58), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L4) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L5_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M49), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M61), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L5) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L6_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M62), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L5), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L6) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L7_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M46), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L3), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L7) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L8_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M51), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M59), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L8) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L9_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M52), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M53), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L9) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L10_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M53), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L4), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L10) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L11_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M60), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L2), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L11) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L12_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M48), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M51), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L12) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L13_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M50), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L0), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L13) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L14_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M52), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M61), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L14) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L15_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M55), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L1), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L15) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L16_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M56), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L0), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L16) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L17_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M57), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L1), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L17) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L18_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M58), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L8), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L18) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L19_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M63), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L4), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L19) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L20_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L0), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L1), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L20) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L21_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L1), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L7), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L21) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L22_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L3), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L12), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L22) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L23_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L18), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L2), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L23) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L24_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L15), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L9), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L24) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L25_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L6), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L10), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L25) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L26_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L7), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L9), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L26) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L27_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L8), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L10), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L27) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L28_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L11), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L14), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L28) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L29_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L11), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L17), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L29) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S0_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L6), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L24), .Z(
        KeyExpansionIns_KeySchedCoreInst_OutBytes_0__7_) );
  XNOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S1_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L16), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L26), .ZN(
        KeyExpansionIns_KeySchedCoreInst_OutBytes_0__6_) );
  XNOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S2_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L19), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L28), .ZN(
        KeyExpansionIns_KeySchedCoreInst_OutBytes_0__5_) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S3_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L6), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L21), .Z(
        KeyExpansionIns_KeySchedCoreInst_OutBytes_0__4_) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S4_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L20), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L22), .Z(
        KeyExpansionIns_KeySchedCoreInst_OutBytes_0__3_) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S5_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L25), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L29), .Z(
        KeyExpansionIns_KeySchedCoreInst_OutBytes_0__2_) );
  XNOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S6_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L13), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L27), .ZN(
        KeyExpansionIns_KeySchedCoreInst_OutBytes_0__1_) );
  XNOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S7_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L6), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L23), .ZN(
        KeyExpansionIns_KeySchedCoreInst_OutBytes_0__0_) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T1_U1 ( .A(
        key_shifted[23]), .B(key_shifted[20]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T2_U1 ( .A(
        key_shifted[23]), .B(key_shifted[18]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T2) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T3_U1 ( .A(
        key_shifted[23]), .B(key_shifted[17]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T3) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T4_U1 ( .A(
        key_shifted[20]), .B(key_shifted[18]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T4) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T5_U1 ( .A(
        key_shifted[19]), .B(key_shifted[17]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T5) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T6_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T5), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T7_U1 ( .A(
        key_shifted[22]), .B(key_shifted[21]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T7) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T8_U1 ( .A(
        key_shifted[16]), .B(KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6), 
        .Z(KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T8) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T9_U1 ( .A(
        key_shifted[16]), .B(KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T7), 
        .Z(KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T9) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T10_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T7), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T10) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T11_U1 ( .A(
        key_shifted[22]), .B(key_shifted[18]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T11) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T12_U1 ( .A(
        key_shifted[21]), .B(key_shifted[18]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T12) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T13_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T3), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T4), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T13) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T14_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T11), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T14) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T15_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T5), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T11), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T15) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T16_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T5), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T12), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T16) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T17_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T9), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T16), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T17) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T18_U1 ( .A(
        key_shifted[20]), .B(key_shifted[16]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T18) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T19_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T7), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T18), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T19) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T20_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T19), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T20) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T21_U1 ( .A(
        key_shifted[17]), .B(key_shifted[16]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T21) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T22_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T7), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T21), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T22) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T23_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T2), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T22), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T23) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T24_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T2), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T10), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T24) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T25_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T20), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T17), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T25) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T26_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T3), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T16), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T26) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T27_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T12), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T27) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M1_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T13), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M1) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M2_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T23), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T8), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M2) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M3_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T14), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M1), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M3) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M4_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T19), .A2(key_shifted[16]), .ZN(KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M4) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M5_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M4), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M1), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M5) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M6_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T3), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T16), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M6) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M7_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T22), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T9), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M7) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M8_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T26), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M6), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M8) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M9_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T20), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T17), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M9) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M10_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M9), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M6), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M10) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M11_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T15), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M11) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M12_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T4), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T27), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M12) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M13_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M12), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M11), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M13) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M14_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T2), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T10), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M14) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M15_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M14), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M11), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M15) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M16_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M3), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M2), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M16) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M17_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M5), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T24), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M17) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M18_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M8), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M7), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M18) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M19_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M10), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M15), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M19) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M20_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M16), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M13), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M20) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M21_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M17), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M15), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M21) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M22_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M18), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M13), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M22) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M23_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M19), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T25), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M23) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M24_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M22), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M23), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M24) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M25_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M22), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M20), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M25) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M26_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M21), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M25), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M26) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M27_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M20), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M21), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M27) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M28_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M23), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M25), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M28) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M29_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M28), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M27), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M29) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M30_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M26), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M24), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M30) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M31_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M20), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M23), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M31) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M32_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M27), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M31), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M32) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M33_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M27), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M25), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M33) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M34_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M21), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M22), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M34) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M35_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M24), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M34), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M35) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M36_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M24), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M25), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M36) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M37_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M21), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M29), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M37) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M38_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M32), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M33), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M38) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M39_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M23), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M30), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M39) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M40_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M35), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M36), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M40) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M41_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M38), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M40), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M41) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M42_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M37), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M39), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M42) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M43_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M37), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M38), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M43) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M44_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M39), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M40), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M44) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M45_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M42), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M41), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M45) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M46_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M44), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M46) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M47_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M40), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T8), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M47) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M48_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M39), .A2(key_shifted[16]), .ZN(KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M48) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M49_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M43), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T16), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M49) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M50_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M38), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T9), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M50) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M51_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M37), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T17), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M51) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M52_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M42), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T15), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M52) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M53_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M45), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T27), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M53) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M54_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M41), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T10), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M54) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M55_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M44), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T13), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M55) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M56_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M40), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T23), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M56) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M57_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M39), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T19), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M57) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M58_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M43), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T3), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M58) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M59_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M38), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T22), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M59) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M60_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M37), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T20), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M60) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M61_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M42), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M61) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M62_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M45), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T4), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M62) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M63_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M41), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T2), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M63) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L0_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M61), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M62), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L0) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L1_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M50), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M56), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L1) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L2_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M46), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M48), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L2) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L3_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M47), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M55), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L3) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L4_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M54), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M58), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L4) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L5_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M49), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M61), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L5) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L6_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M62), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L5), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L6) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L7_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M46), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L3), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L7) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L8_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M51), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M59), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L8) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L9_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M52), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M53), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L9) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L10_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M53), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L4), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L10) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L11_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M60), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L2), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L11) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L12_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M48), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M51), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L12) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L13_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M50), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L0), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L13) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L14_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M52), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M61), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L14) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L15_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M55), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L1), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L15) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L16_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M56), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L0), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L16) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L17_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M57), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L1), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L17) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L18_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M58), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L8), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L18) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L19_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M63), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L4), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L19) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L20_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L0), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L1), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L20) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L21_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L1), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L7), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L21) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L22_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L3), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L12), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L22) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L23_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L18), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L2), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L23) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L24_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L15), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L9), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L24) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L25_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L6), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L10), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L25) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L26_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L7), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L9), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L26) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L27_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L8), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L10), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L27) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L28_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L11), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L14), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L28) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L29_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L11), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L17), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L29) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S0_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L6), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L24), .Z(
        KeyExpansionIns_tmp[23]) );
  XNOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S1_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L16), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L26), .ZN(
        KeyExpansionIns_tmp[22]) );
  XNOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S2_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L19), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L28), .ZN(
        KeyExpansionIns_tmp[21]) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S3_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L6), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L21), .Z(
        KeyExpansionIns_tmp[20]) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S4_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L20), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L22), .Z(
        KeyExpansionIns_tmp[19]) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S5_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L25), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L29), .Z(
        KeyExpansionIns_tmp[18]) );
  XNOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S6_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L13), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L27), .ZN(
        KeyExpansionIns_tmp[17]) );
  XNOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S7_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L6), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L23), .ZN(
        KeyExpansionIns_tmp[16]) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T1_U1 ( .A(
        key_shifted[15]), .B(key_shifted[12]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T2_U1 ( .A(
        key_shifted[15]), .B(key_shifted[10]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T2) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T3_U1 ( .A(
        key_shifted[15]), .B(key_shifted[9]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T3) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T4_U1 ( .A(
        key_shifted[12]), .B(key_shifted[10]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T4) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T5_U1 ( .A(
        key_shifted[11]), .B(key_shifted[9]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T5) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T6_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T5), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T7_U1 ( .A(
        key_shifted[14]), .B(key_shifted[13]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T7) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T8_U1 ( .A(
        key_shifted[8]), .B(KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6), 
        .Z(KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T8) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T9_U1 ( .A(
        key_shifted[8]), .B(KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T7), 
        .Z(KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T9) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T10_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T7), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T10) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T11_U1 ( .A(
        key_shifted[14]), .B(key_shifted[10]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T11) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T12_U1 ( .A(
        key_shifted[13]), .B(key_shifted[10]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T12) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T13_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T3), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T4), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T13) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T14_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T11), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T14) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T15_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T5), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T11), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T15) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T16_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T5), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T12), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T16) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T17_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T9), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T16), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T17) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T18_U1 ( .A(
        key_shifted[12]), .B(key_shifted[8]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T18) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T19_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T7), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T18), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T19) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T20_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T19), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T20) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T21_U1 ( .A(
        key_shifted[9]), .B(key_shifted[8]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T21) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T22_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T7), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T21), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T22) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T23_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T2), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T22), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T23) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T24_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T2), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T10), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T24) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T25_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T20), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T17), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T25) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T26_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T3), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T16), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T26) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T27_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T12), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T27) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M1_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T13), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M1) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M2_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T23), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T8), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M2) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M3_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T14), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M1), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M3) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M4_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T19), .A2(key_shifted[8]), 
        .ZN(KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M4) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M5_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M4), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M1), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M5) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M6_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T3), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T16), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M6) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M7_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T22), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T9), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M7) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M8_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T26), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M6), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M8) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M9_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T20), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T17), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M9) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M10_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M9), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M6), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M10) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M11_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T15), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M11) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M12_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T4), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T27), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M12) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M13_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M12), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M11), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M13) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M14_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T2), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T10), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M14) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M15_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M14), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M11), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M15) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M16_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M3), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M2), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M16) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M17_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M5), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T24), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M17) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M18_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M8), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M7), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M18) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M19_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M10), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M15), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M19) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M20_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M16), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M13), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M20) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M21_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M17), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M15), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M21) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M22_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M18), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M13), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M22) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M23_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M19), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T25), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M23) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M24_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M22), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M23), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M24) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M25_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M22), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M20), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M25) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M26_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M21), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M25), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M26) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M27_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M20), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M21), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M27) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M28_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M23), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M25), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M28) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M29_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M28), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M27), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M29) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M30_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M26), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M24), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M30) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M31_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M20), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M23), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M31) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M32_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M27), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M31), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M32) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M33_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M27), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M25), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M33) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M34_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M21), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M22), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M34) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M35_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M24), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M34), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M35) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M36_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M24), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M25), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M36) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M37_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M21), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M29), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M37) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M38_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M32), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M33), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M38) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M39_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M23), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M30), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M39) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M40_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M35), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M36), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M40) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M41_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M38), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M40), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M41) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M42_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M37), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M39), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M42) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M43_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M37), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M38), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M43) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M44_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M39), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M40), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M44) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M45_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M42), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M41), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M45) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M46_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M44), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M46) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M47_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M40), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T8), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M47) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M48_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M39), .A2(key_shifted[8]), 
        .ZN(KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M48) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M49_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M43), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T16), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M49) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M50_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M38), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T9), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M50) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M51_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M37), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T17), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M51) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M52_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M42), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T15), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M52) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M53_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M45), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T27), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M53) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M54_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M41), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T10), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M54) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M55_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M44), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T13), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M55) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M56_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M40), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T23), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M56) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M57_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M39), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T19), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M57) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M58_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M43), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T3), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M58) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M59_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M38), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T22), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M59) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M60_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M37), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T20), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M60) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M61_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M42), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M61) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M62_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M45), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T4), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M62) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M63_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M41), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T2), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M63) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L0_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M61), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M62), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L0) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L1_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M50), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M56), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L1) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L2_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M46), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M48), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L2) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L3_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M47), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M55), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L3) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L4_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M54), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M58), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L4) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L5_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M49), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M61), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L5) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L6_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M62), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L5), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L6) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L7_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M46), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L3), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L7) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L8_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M51), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M59), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L8) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L9_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M52), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M53), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L9) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L10_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M53), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L4), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L10) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L11_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M60), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L2), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L11) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L12_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M48), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M51), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L12) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L13_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M50), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L0), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L13) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L14_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M52), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M61), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L14) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L15_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M55), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L1), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L15) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L16_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M56), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L0), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L16) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L17_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M57), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L1), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L17) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L18_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M58), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L8), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L18) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L19_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M63), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L4), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L19) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L20_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L0), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L1), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L20) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L21_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L1), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L7), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L21) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L22_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L3), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L12), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L22) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L23_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L18), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L2), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L23) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L24_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L15), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L9), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L24) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L25_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L6), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L10), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L25) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L26_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L7), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L9), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L26) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L27_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L8), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L10), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L27) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L28_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L11), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L14), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L28) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L29_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L11), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L17), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L29) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S0_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L6), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L24), .Z(
        KeyExpansionIns_tmp[15]) );
  XNOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S1_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L16), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L26), .ZN(
        KeyExpansionIns_tmp[14]) );
  XNOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S2_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L19), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L28), .ZN(
        KeyExpansionIns_tmp[13]) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S3_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L6), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L21), .Z(
        KeyExpansionIns_tmp[12]) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S4_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L20), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L22), .Z(
        KeyExpansionIns_tmp[11]) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S5_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L25), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L29), .Z(
        KeyExpansionIns_tmp[10]) );
  XNOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S6_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L13), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L27), .ZN(
        KeyExpansionIns_tmp[9]) );
  XNOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S7_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L6), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L23), .ZN(
        KeyExpansionIns_tmp[8]) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T1_U1 ( .A(
        key_shifted[39]), .B(key_shifted[36]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T2_U1 ( .A(
        key_shifted[39]), .B(key_shifted[34]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T2) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T3_U1 ( .A(
        key_shifted[39]), .B(key_shifted[33]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T3) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T4_U1 ( .A(
        key_shifted[36]), .B(key_shifted[34]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T4) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T5_U1 ( .A(
        key_shifted[35]), .B(key_shifted[33]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T5) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T6_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T5), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T7_U1 ( .A(
        key_shifted[38]), .B(key_shifted[37]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T7) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T8_U1 ( .A(
        key_shifted[32]), .B(KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6), 
        .Z(KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T8) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T9_U1 ( .A(
        key_shifted[32]), .B(KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T7), 
        .Z(KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T9) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T10_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T7), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T10) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T11_U1 ( .A(
        key_shifted[38]), .B(key_shifted[34]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T11) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T12_U1 ( .A(
        key_shifted[37]), .B(key_shifted[34]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T12) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T13_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T3), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T4), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T13) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T14_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T11), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T14) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T15_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T5), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T11), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T15) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T16_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T5), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T12), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T16) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T17_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T9), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T16), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T17) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T18_U1 ( .A(
        key_shifted[36]), .B(key_shifted[32]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T18) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T19_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T7), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T18), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T19) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T20_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T19), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T20) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T21_U1 ( .A(
        key_shifted[33]), .B(key_shifted[32]), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T21) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T22_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T7), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T21), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T22) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T23_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T2), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T22), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T23) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T24_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T2), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T10), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T24) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T25_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T20), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T17), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T25) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T26_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T3), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T16), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T26) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T27_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T12), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T27) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M1_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T13), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M1) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M2_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T23), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T8), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M2) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M3_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T14), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M1), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M3) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M4_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T19), .A2(key_shifted[32]), .ZN(KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M4) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M5_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M4), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M1), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M5) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M6_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T3), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T16), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M6) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M7_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T22), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T9), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M7) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M8_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T26), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M6), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M8) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M9_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T20), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T17), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M9) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M10_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M9), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M6), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M10) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M11_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T15), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M11) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M12_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T4), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T27), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M12) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M13_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M12), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M11), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M13) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M14_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T2), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T10), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M14) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M15_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M14), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M11), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M15) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M16_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M3), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M2), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M16) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M17_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M5), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T24), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M17) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M18_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M8), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M7), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M18) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M19_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M10), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M15), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M19) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M20_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M16), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M13), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M20) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M21_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M17), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M15), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M21) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M22_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M18), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M13), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M22) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M23_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M19), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T25), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M23) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M24_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M22), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M23), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M24) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M25_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M22), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M20), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M25) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M26_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M21), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M25), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M26) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M27_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M20), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M21), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M27) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M28_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M23), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M25), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M28) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M29_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M28), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M27), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M29) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M30_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M26), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M24), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M30) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M31_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M20), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M23), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M31) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M32_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M27), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M31), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M32) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M33_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M27), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M25), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M33) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M34_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M21), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M22), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M34) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M35_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M24), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M34), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M35) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M36_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M24), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M25), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M36) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M37_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M21), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M29), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M37) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M38_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M32), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M33), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M38) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M39_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M23), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M30), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M39) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M40_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M35), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M36), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M40) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M41_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M38), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M40), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M41) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M42_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M37), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M39), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M42) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M43_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M37), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M38), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M43) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M44_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M39), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M40), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M44) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M45_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M42), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M41), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M45) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M46_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M44), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M46) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M47_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M40), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T8), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M47) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M48_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M39), .A2(key_shifted[32]), .ZN(KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M48) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M49_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M43), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T16), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M49) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M50_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M38), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T9), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M50) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M51_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M37), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T17), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M51) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M52_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M42), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T15), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M52) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M53_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M45), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T27), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M53) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M54_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M41), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T10), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M54) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M55_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M44), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T13), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M55) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M56_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M40), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T23), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M56) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M57_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M39), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T19), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M57) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M58_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M43), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T3), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M58) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M59_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M38), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T22), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M59) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M60_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M37), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T20), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M60) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M61_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M42), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M61) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M62_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M45), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T4), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M62) );
  AND2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M63_U1 ( .A1(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M41), .A2(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T2), .ZN(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M63) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L0_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M61), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M62), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L0) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L1_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M50), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M56), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L1) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L2_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M46), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M48), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L2) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L3_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M47), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M55), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L3) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L4_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M54), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M58), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L4) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L5_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M49), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M61), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L5) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L6_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M62), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L5), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L6) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L7_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M46), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L3), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L7) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L8_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M51), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M59), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L8) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L9_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M52), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M53), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L9) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L10_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M53), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L4), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L10) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L11_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M60), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L2), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L11) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L12_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M48), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M51), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L12) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L13_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M50), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L0), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L13) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L14_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M52), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M61), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L14) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L15_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M55), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L1), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L15) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L16_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M56), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L0), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L16) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L17_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M57), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L1), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L17) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L18_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M58), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L8), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L18) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L19_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M63), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L4), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L19) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L20_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L0), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L1), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L20) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L21_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L1), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L7), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L21) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L22_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L3), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L12), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L22) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L23_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L18), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L2), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L23) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L24_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L15), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L9), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L24) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L25_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L6), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L10), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L25) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L26_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L7), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L9), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L26) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L27_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L8), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L10), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L27) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L28_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L11), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L14), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L28) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L29_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L11), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L17), .Z(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L29) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S0_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L6), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L24), .Z(
        KeyExpansionIns_tmp[7]) );
  XNOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S1_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L16), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L26), .ZN(
        KeyExpansionIns_tmp[6]) );
  XNOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S2_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L19), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L28), .ZN(
        KeyExpansionIns_tmp[5]) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S3_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L6), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L21), .Z(
        KeyExpansionIns_tmp[4]) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S4_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L20), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L22), .Z(
        KeyExpansionIns_tmp[3]) );
  XOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S5_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L25), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L29), .Z(
        KeyExpansionIns_tmp[2]) );
  XNOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S6_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L13), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L27), .ZN(
        KeyExpansionIns_tmp[1]) );
  XNOR2_X1 KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S7_U1 ( .A(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L6), .B(
        KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L23), .ZN(
        KeyExpansionIns_tmp[0]) );
  NOR2_X1 RoundCounterIns_U11 ( .A1(start), .A2(RoundCounterIns_n8), .ZN(
        RoundCounterIns_n27) );
  XNOR2_X1 RoundCounterIns_U10 ( .A(RoundCounter[0]), .B(notdone), .ZN(
        RoundCounterIns_n8) );
  NOR2_X1 RoundCounterIns_U9 ( .A1(start), .A2(RoundCounterIns_n7), .ZN(
        RoundCounterIns_n26) );
  XOR2_X1 RoundCounterIns_U8 ( .A(RoundCounter[1]), .B(RoundCounterIns_n6), 
        .Z(RoundCounterIns_n7) );
  NOR2_X1 RoundCounterIns_U7 ( .A1(start), .A2(RoundCounterIns_n5), .ZN(
        RoundCounterIns_n25) );
  XNOR2_X1 RoundCounterIns_U6 ( .A(RoundCounter[2]), .B(RoundCounterIns_n4), 
        .ZN(RoundCounterIns_n5) );
  NOR2_X1 RoundCounterIns_U5 ( .A1(start), .A2(RoundCounterIns_n3), .ZN(
        RoundCounterIns_n24) );
  XOR2_X1 RoundCounterIns_U4 ( .A(RoundCounter[3]), .B(RoundCounterIns_n2), 
        .Z(RoundCounterIns_n3) );
  NAND2_X1 RoundCounterIns_U3 ( .A1(RoundCounterIns_n4), .A2(RoundCounter[2]), 
        .ZN(RoundCounterIns_n2) );
  NOR2_X1 RoundCounterIns_U2 ( .A1(RoundCounterIns_n1), .A2(RoundCounterIns_n6), .ZN(RoundCounterIns_n4) );
  NAND2_X1 RoundCounterIns_U1 ( .A1(notdone), .A2(RoundCounter[0]), .ZN(
        RoundCounterIns_n6) );
  INV_X1 RoundCounterIns_count_reg_0__U1 ( .A(RoundCounter[0]), .ZN(
        RoundCounterIns_count_reg_0__QN) );
  DFF_X1 RoundCounterIns_count_reg_0__FF_FF ( .D(RoundCounterIns_n27), .CK(clk), .Q(RoundCounter[0]), .QN() );
  INV_X1 RoundCounterIns_count_reg_1__U1 ( .A(RoundCounter[1]), .ZN(
        RoundCounterIns_n1) );
  DFF_X1 RoundCounterIns_count_reg_1__FF_FF ( .D(RoundCounterIns_n26), .CK(clk), .Q(RoundCounter[1]), .QN() );
  INV_X1 RoundCounterIns_count_reg_2__U1 ( .A(RoundCounter[2]), .ZN(
        RoundCounterIns_count_reg_2__QN) );
  DFF_X1 RoundCounterIns_count_reg_2__FF_FF ( .D(RoundCounterIns_n25), .CK(clk), .Q(RoundCounter[2]), .QN() );
  INV_X1 RoundCounterIns_count_reg_3__U1 ( .A(RoundCounter[3]), .ZN(
        RoundCounterIns_count_reg_3__QN) );
  DFF_X1 RoundCounterIns_count_reg_3__FF_FF ( .D(RoundCounterIns_n24), .CK(clk), .Q(RoundCounter[3]), .QN() );
endmodule

