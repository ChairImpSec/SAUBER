// X0Y1, W_IO_custom
`define Tile_X0Y1_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000001000000000000000000000000000000000010100000100000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000001100000000000000000000000000000000000000000000000000000000000000000
// X1Y1, linear_LMDPL
`define Tile_X1Y1_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000001100000000000000000000000000000000000000000111110011000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000100010101000100000000000000000100010000000000000000000000000000000000111000000111101100001000
// X2Y1, linear_LMDPL
`define Tile_X2Y1_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001101011100000000000000000011000000000000000000010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110011000011000000000000000000001000000000000000000000000000000000000000000000000000111100000000000000000000001000100000001000000000000000001000100010101000
// X3Y1, nonlinear_LMDPL
`define Tile_X3Y1_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000001010011001000000000000000000000110100000000100100000000000000001110000000000001000000110011
// X4Y1, linear_LMDPL
`define Tile_X4Y1_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011110000000000110000110000000000000000000000000000000001010000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000101011000000000011000011000000000111000000000000000000000000000000000000000000000000010100010000000100000000000000000111110010100110
// X5Y1, linear_LMDPL
`define Tile_X5Y1_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000011000000000000000000110000000000000000000000000000000000000000000000000000000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000111111000000010001000100000000000000000000010101100110101100000000000000000000000000000000000000101100
// X6Y1, nonlinear_LMDPL
`define Tile_X6Y1_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X7Y1, linear_LMDPL
`define Tile_X7Y1_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000011000011000000000000000000000000010000000000000000000000000000000000000001010110000000000000000001010100001000110000
// X8Y1, ctrl_to_sec
`define Tile_X8Y1_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X9Y1, combined_WDDL
`define Tile_X9Y1_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010011000000000000000011000001010001000000000000000011101010
// X10Y1, ctrl_IO
`define Tile_X10Y1_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000100000000000
// X0Y2, W_IO_custom
`define Tile_X0Y2_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000000000100000000000000001000000000000000000000000000100000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000
// X1Y2, linear_LMDPL
`define Tile_X1Y2_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000110000000000000000000000000000000000001100000000000000000000000000000000000011000000000000100000000000000000000000000000000000100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000101110110110100000000000000000001010110010001001
// X2Y2, linear_LMDPL
`define Tile_X2Y2_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010010010010000000000000000000000000001100110000000000000001000000000000000011001100000000000000000000000000000000000000000000000000111100110000000000000000000010000000000000000000000011000000100000000010000000000000000000001000000000000000000000000000000100010001000100000000000000000001000100110011000000000000000000000000000000000010001001110011
// X3Y2, nonlinear_LMDPL
`define Tile_X3Y2_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100111100000000000000000000000000000000000000000000000011110000000010000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000011001000000000000000000000000000000000100111010000000000000000000000001011100000011100
// X4Y2, linear_LMDPL
`define Tile_X4Y2_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100110000000011000000000000000000000000000010000010000000000010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000010000000000000000000000110000000111000000000000000000000001000000010000010000000011000000000010001000100000000000000000000110111101110101100000000000000000000000000000001000001000010
// X5Y2, linear_LMDPL
`define Tile_X5Y2_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000101000100000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000010000000000000000000000000001100000000000000000000000000001100111100000000001010000000000000000000000000000000000000000000000000011101000111010000000000000000001010101111101101
// X6Y2, nonlinear_LMDPL
`define Tile_X6Y2_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000001100000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000100000000000000000000000010000000000000100000000000000000000000000001000000100100010000011000000000000000000001101000010
// X7Y2, linear_LMDPL
`define Tile_X7Y2_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000001111000000000000000000000000000000000000000000000000000100010001000100000000000000001000101111001001000000000000000000000000000000000010010000010011
// X8Y2, ctrl_to_sec
`define Tile_X8Y2_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X9Y2, combined_WDDL
`define Tile_X9Y2_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100110000100000000000000000100100010000000000110001000000000011111011000000000000000010001111
// X10Y2, ctrl_IO
`define Tile_X10Y2_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000100000000000
// X0Y3, W_IO_custom
`define Tile_X0Y3_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000001000011010000000000000000101100000000000000000000000000001100001000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000
// X1Y3, linear_LMDPL
`define Tile_X1Y3_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000111100000000000000000000000000000000000001001000000011000000000000000000000000000000000000000000000000000000000000000000000010000010000000000000000000000000000010110010000000100000000000001100000000000000000010001000000011000000000011000011000000000100010001000000000000000011000011011001010000000000000000011100000000000000000011010001010001
// X2Y3, linear_LMDPL
`define Tile_X2Y3_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001000000000000000000000000000000111100000000000100000000000000000000000000000000010000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000100000000010000000000000000000000000001000100000000000000000000100010100000000000000101000001010101000000000000000000001001100000000110100001100100000001001
// X3Y3, nonlinear_LMDPL
`define Tile_X3Y3_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000110000000000110000000000000010000000000000000000001100110000000000000000000000000000000000000100000000000000000000000000000000000000000000000001010000010010000000010011001000100010000000000000110100000000100100000000000000000000000000001011001110110000
// X4Y3, linear_LMDPL
`define Tile_X4Y3_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000011000000010010110010110000000000110000000000000000000000001100000000000000000000001011000011000000000000000000000000000000000000001000000010000010000000000000001010000010001010000000000000100010000000000010000000000000101011000000010001000100000000000000000000001101000111101000000000000000000000000000001100010010011101
// X5Y3, linear_LMDPL
`define Tile_X5Y3_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000011000000000000000000000000000000000011000000001100001000000000000000000000000001000000000000000000000100000100000000000000000000000000000000000000000000000000000000000010100000100000001000100000000010000000000000000000000000111100000000000000000010010001000100010000000000000011110000000000000000010011001011101010111100100011000000000000000000
// X6Y3, nonlinear_LMDPL
`define Tile_X6Y3_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100000000010000000000000000000000000100000000000000000100010000000000000000000000000000000000000000000000000000000010100001100000000000000000101011000110100
// X7Y3, linear_LMDPL
`define Tile_X7Y3_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000011110000001000110000001010000000000100010001000100000000000011001001100110001000000000000000000000000000000000000011000000000100
// X8Y3, ctrl_to_sec
`define Tile_X8Y3_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X9Y3, combined_WDDL
`define Tile_X9Y3_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000011000010010100000000000000000100001000100000011000010000000110000000000111010101101100000000000
// X10Y3, ctrl_IO
`define Tile_X10Y3_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000
// X0Y4, W_IO_custom
`define Tile_X0Y4_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011000010100010000000010000000000000000000000000000000000000000000000000000000011000000000000110000000000000000000011000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X1Y4, linear_LMDPL
`define Tile_X1Y4_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000010011000000000000000000000000000000001110110100000100000000000000000000000000000000000000000000000000000000000000000000000010000010000000000000000000000000000010000000110000100000000000000000000000100000000000000000000000000000000010000010000000000101010000000000000000000000001011110000000000000000000010001100001110000000001011000000011100
// X2Y4, linear_LMDPL
`define Tile_X2Y4_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000011110000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000010001000000000000000000010001000100000001010000000000000000000001000001000100000001100000000000100010001000100000000000000000010001100010001000000000000000000000000000000001011000001001000
// X3Y4, nonlinear_LMDPL
`define Tile_X3Y4_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000011110000000000000000000000000000000000000000001100001100000010000000000000000000000000000000001000000000000000000000000000001000000000000000000000000000000000000000000001000110100000100010000000000011001000000000000000000000000000000000100111010000000000000000000000000001100000100011
// X4Y4, linear_LMDPL
`define Tile_X4Y4_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010000000000000000000000000000000000010000001111001100001100000000000000000000000000000000000000000000001000110000000000000000001000000000000000000000000000000000001010000010000000100000001000110000000000000000000000000000001000001100000000000000101010010001000100010000000000000000110000000000000000100010101000100010001001100010000000000000000000
// X5Y4, linear_LMDPL
`define Tile_X5Y4_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000011100110000000000000000000000000001110000010101100001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000100010101000100000101000101111100010000000000000100000000000101000000000110000110010000000000000000000000000000000000000000000000000001100110010001100000000000000000100010000011010
// X6Y4, nonlinear_LMDPL
`define Tile_X6Y4_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000001111001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010000010000000000000000000000000100010000000001000101010000000000001000000000000000000000000000010010000000100000000000000000000000000000000010000100011
// X7Y4, linear_LMDPL
`define Tile_X7Y4_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100011110000000000000000000000000011001000100000001010001100010000000000000000000011001100000000000000000000001001000010001110010000000000000000000100000100
// X8Y4, ctrl_to_sec
`define Tile_X8Y4_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X9Y4, combined_WDDL
`define Tile_X9Y4_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000001000000000000000000000000000101000100010110000000000000000111101100100000110000010010000100000000000000000001010111000000000
// X10Y4, ctrl_IO
`define Tile_X10Y4_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000100000000000000000
// X0Y5, W_IO_custom
`define Tile_X0Y5_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100110000000000000000000000000000000011000000000011000000000000100000000000000000000000000000000000000000010000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X1Y5, linear_LMDPL
`define Tile_X1Y5_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000010000000000000000000000000000010001010000011100011000000000000000000000000000010001000000010000000000010000010000000000000000000000000000000000010000000000000000000001100000010000000000000000000001100101110111101
// X2Y5, linear_LMDPL
`define Tile_X2Y5_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000011000000000000000000010000110000000000001000001100000000000000000000000000000000010000000000000000000000000000000000000010001000000000000000000000000000001010000000000000000010001000001000001000000000000000001001000000001000100010000010000001000100010001000100000000000000001110111010011000000000000000000000000000000000001001101010111111
// X3Y5, nonlinear_LMDPL
`define Tile_X3Y5_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111011100001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000000000000000000000000000000000000000001100000000000000001000000000010000000000000000000000000000000010001010100000100001000100010001000100000000000000000001000000010011000000000000000000000000000000000100000100100000
// X4Y5, linear_LMDPL
`define Tile_X4Y5_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000010110011000011000000000000000000001000000000000000000000110000001000000000110011110000000000000000000000101010000010000000101100001000100010100011000000000000100000000000111010000011110000101001010001000100000000000000000000000000000000000000101101011110011010001000110000000000000000000011
// X5Y5, linear_LMDPL
`define Tile_X5Y5_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000010101000100000101011101010101110000000000000000000000000101000001010001011101011010101010101010100000000000010101001100010011000000000000000000010001010101110010000000000000000
// X6Y5, nonlinear_LMDPL
`define Tile_X6Y5_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010100010000000000000000010000000100010000000001000101010000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000
// X7Y5, linear_LMDPL
`define Tile_X7Y5_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100011000000000000000010101100000010101110100000001000010001000100010000000000001110000000000000000000101110001011101110101100100110110000000000000000
// X8Y5, ctrl_to_sec
`define Tile_X8Y5_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X9Y5, combined_WDDL
`define Tile_X9Y5_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000100001100001000000000000000000000100010000011010000000101111100011001001000000000000000011111000
// X10Y5, ctrl_IO
`define Tile_X10Y5_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000010000000000
// X0Y6, W_IO_custom
`define Tile_X0Y6_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000110000110011000000000000000000110000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X1Y6, linear_LMDPL
`define Tile_X1Y6_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100110000110011000100000001000000000000000000000000000000000000000000000000000000000000000010000010000000000000000000000000001010001010101000100000000000000000000000000000000000000000000000010000000010000010000000000000000000000000000000000000000000000000000000000001000001001000000000000000001101110111001110
// X2Y6, linear_LMDPL
`define Tile_X2Y6_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000011000000000000000000000010000010001000000000000000000000000010001010000000001000001000001000001000001011000000000000000000001000001000101110110010110010000100010001000100000000000000000010000100010000000000000000000000000000000000000101010100010010
// X3Y6, nonlinear_LMDPL
`define Tile_X3Y6_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000001100000000000000000000000000000000000000001100000010000000000000000000000000000000001000000000000000000000000000001010010000100010000000000000000000000000100110001010100000101010000000000011001000100010000000000000000000000000100111010000000000000000000000000010010000110100
// X4Y6, linear_LMDPL
`define Tile_X4Y6_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000010000000000000010000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000001010100010000000100000001000011110101110000000000000000000001000101110001110101000101010010100010001010100000000000000101000100011001011000000000000000000100000000001010000101111000000
// X5Y6, linear_LMDPL
`define Tile_X5Y6_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000000000000000000000000001001000001111000000100000000010000000000000000000000011110000000000000000000000000100000000000000000000000000000000000000000000100000000010100000100000001001000000100110000000100000100000000000100000011010001000001000010001000100010000000000000100000000000000000000100110011011101010101001100010100000000000000000
// X6Y6, nonlinear_LMDPL
`define Tile_X6Y6_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000001100000000110000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000001000101010100010000000000000000000000000110010000000011000101010000000000100000000000000000000000000000000000000100010101010100000000000101100000000001000000001
// X7Y6, linear_LMDPL
`define Tile_X7Y6_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000001000000000000000110000000000000000000010001010000000001010111110101010000000000000000000110000000010101010100000111010010001000100010000000000110000000000000000000000001100110110011010001110101011010000000000000000
// X8Y6, ctrl_to_sec
`define Tile_X8Y6_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X9Y6, combined_WDDL
`define Tile_X9Y6_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000010000000000000000000000000100010101000000000000000000000000101010100101010000000101111100010111011000000001000111100000000
// X10Y6, ctrl_IO
`define Tile_X10Y6_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X0Y7, W_IO_custom
`define Tile_X0Y7_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000011000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000110000000000000000000000000000000011000000000000000000000000000000000
// X1Y7, linear_LMDPL
`define Tile_X1Y7_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100110000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000010000000000000000000000000101010101010101000100011000000000000000000110000000010001100000000000011000011000011000000010101010101010100000000000000001100001000110000000000000000000010101011111011010000000000000000
// X2Y7, linear_LMDPL
`define Tile_X2Y7_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000011110000000000110000000000000000000000001000000000000000000000000000000000000010000010000010001110001000000000000000000000001000001011000000001000001000111000001000011000000000000000001010000000001000100010000010000010010001000100010000000000000000000000000000000000101010111100101010111010101110000000000000000000
// X3Y7, nonlinear_LMDPL
`define Tile_X3Y7_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111001100000000000000000000000000001100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000001010100000010010000000000000000000000000101010001010100100101010000101010001000100000000000000000100000000000011000000000000000000000011000000001010000011001010
// X4Y7, linear_LMDPL
`define Tile_X4Y7_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000011000000000000110000000000000000000000000000000000000000000000000000100010010000100000001000100010101110000000000000100000000011100010001110101000101010010001000100010000000000001100000000000000000000010000000011010110111100100010010000000000000000
// X5Y7, linear_LMDPL
`define Tile_X5Y7_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000010000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000100000000000011110000000000000000000000000000000000000000000010101100100000111010100100101010000000000000000000000000101000101010001000001000010000000100000000000000000010100000000000000000000100010101000100100000010000000000100000001100
// X6Y7, nonlinear_LMDPL
`define Tile_X6Y7_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000010000000110000000000000000000000000000000000000100000000000100000000000000100000100000000000000000000000000000000000000000001010001011111010000010000000000000000010000000101010000000101011101000000001000100000000000000001000000000000000000000100011001010100000001000100100000001000000000000
// X7Y7, linear_LMDPL
`define Tile_X7Y7_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000001000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000010001000000000000000101011001100000000000000000010100011100010100010100000100000010101010101010100000000001110001011111011011000000000000000000010001000101011110000000000000000
// X8Y7, ctrl_to_sec
`define Tile_X8Y7_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X9Y7, combined_WDDL
`define Tile_X9Y7_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000101110101000000000000000000000000001000111101010000000100000100000000000111110001011101100000000
// X10Y7, ctrl_IO
`define Tile_X10Y7_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X0Y8, W_IO_custom
`define Tile_X0Y8_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000011110000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X1Y8, linear_LMDPL
`define Tile_X1Y8_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000011000011000011000011000000000000000000000000000000000000000000000000000000000000000000001010000010000000000000000000101000001010101010101000100000000000000000000000000000000000001000000000000010000010100010000000000001010101000100000000000000000000000000000110011100000000000000001001101100000100000000000011
// X2Y8, linear_LMDPL
`define Tile_X2Y8_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000111000001000000000000000000000000000001100000110000011000100000000000000000000000011000000000000000000000000000000000000000011000010001000000000000000000000000010001000000000001100001100000000000000100000000000110000000000001000001000100000000010000010010001000100010000000000000000000000000000000000001000110100000110011011100010010000000000000000
// X3Y8, nonlinear_LMDPL
`define Tile_X3Y8_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000011110000000000000000000000000000000000000000000000000010000000000000001100000000000011000100000000100000000000100000101010100000100110000000000000000000000000101010001010101000101010000000010011001000000000000000000000010100000000100100000000000000000000000000000011100000101100
// X4Y8, linear_LMDPL
`define Tile_X4Y8_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000100000001011100000001010000000000000000000001000100000101010101111101010000100010001000100000000110011101000100011001011000000000000000000000000000000000001001100000001
// X5Y8, linear_LMDPL
`define Tile_X5Y8_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000001000000000000000000110000001000000000001000001000000000000000000000000000110011110000000000000000000000000000000000000000000100000000000000000000000000100000000100100000100000001001101000101010000000000000100000000000100000101010000000000000000100010001000100000000001000001011110010101011000000000000000000000000000000000010010000010111
// X6Y8, nonlinear_LMDPL
`define Tile_X6Y8_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000011000000000011110000001000000011000000000000000000000000000000000011000000000000000000000000100000100000000000000000000000000010110000000010111001001000101010000010000000000000000000000000101010000000101010101000010000000000000000000000000000000000000000000000011011101010000010110000000000000000010000100011
// X7Y8, linear_LMDPL
`define Tile_X7Y8_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000010000000000001000000000000000000000000000000000000010001000000000001100101010001000000000000000000000100000101110100010100000101110000000000000000000000000100000110000000000000000011001010110011000000000000000000010001001000000
// X8Y8, ctrl_to_sec
`define Tile_X8Y8_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000010
// X9Y8, combined_WDDL
`define Tile_X9Y8_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000011000000000000000000000000101010101100000000000000000000000101010110101010000000100000100010101110000000001111100100000000
// X10Y8, ctrl_IO
`define Tile_X10Y8_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X0Y9, W_IO_custom
`define Tile_X0Y9_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000010000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X1Y9, linear_LMDPL
`define Tile_X1Y9_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000110000000000000000000000000000000010111110000010001100000000000000000000000000000000000000000000000000000000000000000000001010000010000000000000000000000000101010101010101000100000000010000000000000000000000010000000000000000000000000000000000000000000010001000100000000000000000000111010111011011000000000000000000000000000001101110111101011
// X2Y9, linear_LMDPL
`define Tile_X2Y9_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000011000000000000000000000000000000000000000010001000000000000000000000001100001000000000000000000000000000000000100000000000000000001110000000001001100001000010000010000100000000000000000000000000000011000000000000000011001001100000000000000000000100000100010001
// X3Y9, nonlinear_LMDPL
`define Tile_X3Y9_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000001100000000000000000000110000000000000000000000000000000000110000000000001000011000000000000010000000000000000000000000000000000000000000100000000000100000101010100001101010000000000000000000000001101001001000101000101010010101010101010100100010000000000010000110000011000000000000000000110000010000100000000000000000
// X4Y9, linear_LMDPL
`define Tile_X4Y9_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000001000001111000000000000000000000000000000001100110000101000001100000000000000000000000000000000000000000000100000000000100000001010000000111010000000000000000000000010100000111010101010101010000100010001010100000000001000001100101110111000000000000000000000000000000011000010001101000000
// X5Y9, linear_LMDPL
`define Tile_X5Y9_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000100000000000000000000000000000000000000000100000000000100000000000000000000000000000000000000001100000000000000000000000000000000000000100000000000000000000000000000000000100000100000000001101011111000000000100000000000010000000011101010000001000011010101010100010100001100001100001001100000001000000000000001000011000100111011100000000000000000
// X6Y9, nonlinear_LMDPL
`define Tile_X6Y9_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000110000000000000000000000000000000000001100110000000100001000000000000000000000000000000000000000100000000000001000000000000000100000100000000000000000000000000010000000000011001000001000100010000010000000000000000010000000101010000001101000101000010000000100010000000000001000000000000000000000001110111110000100010000000100110000100100000000
// X7Y9, linear_LMDPL
`define Tile_X7Y9_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000010001000000000000000000000000000010000000000000001000010000000000000000000000000000000000000000000000000000000000000000000000001000101010001011000000000000000010111110111010100000100000101010010001000100000000111100001010000000000000000000000100100101011000010001000000000000000000000001
// X8Y9, ctrl_to_sec
`define Tile_X8Y9_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000
// X9Y9, combined_WDDL
`define Tile_X9Y9_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010100000000000000000000000000101010100101011000000101100000011111001000000001010111000000000
// X10Y9, ctrl_IO
`define Tile_X10Y9_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X0Y10, W_IO_custom
`define Tile_X0Y10_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X1Y10, linear_LMDPL
`define Tile_X1Y10_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000110000000000000000000000100000000000000000000000000000001100001100000000000000000000000000000000000000000000110000001010000010000000000000000000111100001010111010101010100000000000000000000000000000000000001100110000000000000000000000000000000100010001000100000000000000000011001001010010000000000000000000000000000000001000100111001010
// X2Y10, linear_LMDPL
`define Tile_X2Y10_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000110000000000000000000000000000000000001100000000000011000000000000000000000000000000000000000000000000000000000000000000000110001000010000000000000000000010001001000000000000000000000001000000100000000000000000000000001000001010100010000010000010000000000001000000000000000000000000000010010000010000010000000100000000000000001000110011101101
// X3Y10, nonlinear_LMDPL
`define Tile_X3Y10_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011000000001100000000000000000000000000110000000000000000000001000000000000000000000000000000000000000000010011000000100000101001100010101010000000000000000000000000101010001000101001101010000100010011001000000000000000000001010100000000000000000000000000000000000000000011000000010010
// X4Y10, linear_LMDPL
`define Tile_X4Y10_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000011000000000000000000000000000000000100000000001100011000000000000000000000001100000000000000000100000000001000000000000000000000000000000000000000000000000000100000000000100000000000000001101010000000001100000000001000100000101010101000001100010101010101010111000011001100101001101010101010000000000000000011101001111010110000000000000000
// X5Y10, linear_LMDPL
`define Tile_X5Y10_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000010000000010000000010000000001000000000000000000000000000110000000000110000000011001100000000000000000000000000000000000000100000000000100000100000000010100000001000000000000000100000000000000000101010000000000000000100010001000100000000001000001010000100011001000000000000000000000000000000001000101010001011
// X6Y10, nonlinear_LMDPL
`define Tile_X6Y10_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110011000000000000000000000000000011000000000011000000001010000000000000000000000000000000000000000000000000000000000000100000100000100000000000000000000000000010000000100000001010001000000010000010000000000000000000000000101010000010101000101000000000000000000000000000000000000000000000000000000000000100001000000000000000001100100000111010
// X7Y10, linear_LMDPL
`define Tile_X7Y10_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000010001000000000000000000000000000001000000000000000000010000000000000101010001010000000000000000011100000100010100000100000101110000100010001000100000000101100111001110010101110000000000000000000000000000000000010000001000000
// X8Y10, ctrl_to_sec
`define Tile_X8Y10_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000100000000
// X9Y10, combined_WDDL
`define Tile_X9Y10_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000100010000101010000011101011000010011000000000000000000010111111
// X10Y10, ctrl_IO
`define Tile_X10Y10_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X0Y11, W_IO_custom
`define Tile_X0Y11_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000001000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X1Y11, linear_LMDPL
`define Tile_X1Y11_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111010110010000000000000000000101000101010111010101010100000110000000000000000000000000010100000000000000000000000000000000000000100010000000100000000000000000010001000000011000000001100000000000000000000001001100110101000
// X2Y11, linear_LMDPL
`define Tile_X2Y11_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000010000000000010000000000000000000000000000000001000000000000000000000000001000000000010101000000000000000000000000000001010000000000000000000000010110000100000000000000000000000110000011000100000000010000011010100010001000100000000110000000000000000000100000000000000000000110000000000000000101110101000
// X3Y11, nonlinear_LMDPL
`define Tile_X3Y11_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000000000000000000000000000000000001111110000000000000000000000000010000011010000010100000000000000000000000000000000000000000000000000000000000000010000101010100101100110000000000000000000000010011010011000101010101010000100000000000100000000000000000001000000000000000011011100000000000000000000000101001101000010
// X4Y11, linear_LMDPL
`define Tile_X4Y11_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000011000000000000111000100000000000000011000000000011000010000000000000000010000011000000000000000000000000000000000000100011000000010000000011111100100010000000000000000000000000100000011000101000001000010101010101010100000000000000001100101110111000000000000000000010111110100011010000000000000000
// X5Y11, linear_LMDPL
`define Tile_X5Y11_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000101000000000000000000000000000000000000000000010100010000000000000100000000000000000000000000000011000000000100000000000000110011000000000000000000000000000000000000101011101100000001100001000001000000000000000000100000110001001010110000110000010101010101010100000000001000000100100110001100000000000000000000010001010000000000000000000000
// X6Y11, nonlinear_LMDPL
`define Tile_X6Y11_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000010000000000000111100001000001100000000001000000000000010001100000000000000000000010000101000100000000000000000000000001010000000000000000000100000000011000000000000000000000000000000011010000100101000000000010001000100010000000000000000000000000000000000000110100000000010011010101010000000000000000000
// X7Y11, linear_LMDPL
`define Tile_X7Y11_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000010000000110000000000000011001100000000000000000000000000000000000000000000000011000000000000101010111010000000000000000010101010100000100000110000101011010100010101010111001100001010000101011010110010000000000000000001000000110010100000001100000000
// X8Y11, ctrl_to_sec
`define Tile_X8Y11_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000
// X9Y11, combined_WDDL
`define Tile_X9Y11_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000010000000000000100000000101010100101010001100101000110011001011000000001000111100000000
// X10Y11, ctrl_IO
`define Tile_X10Y11_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X0Y12, W_IO_custom
`define Tile_X0Y12_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000001000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X1Y12, linear_LMDPL
`define Tile_X1Y12_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111010000010110000000000000000000000001010101010101010100011000000000000000000000000000000000000100000000000000000000000000000010101010100000100000000000000000010010000000100000000001010000001100011001000000000000000001000
// X2Y12, linear_LMDPL
`define Tile_X2Y12_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000011000000000000000011000010001100000000000000000000000000000000000000000000000001000000000100000000000010101000100000000000000000000010101010000000010000001001000010100001100001000000000000100000000000100000000000000000000010000100010001000100000000000000001010110011011100000000000000000000000000000000001001100110111011
// X3Y12, nonlinear_LMDPL
`define Tile_X3Y12_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000011000000001100001100000000000000000000000000010000000100000000010000000000000000000010001001000000000000000000100010000010100000011010101010101010000000000000000000111100101000001000101010101010010101010101010000000000000000000010000100110000000000000000101000000000110011000000000000000000
// X4Y12, linear_LMDPL
`define Tile_X4Y12_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000100001010000000000000000000100000000000000000000001000100000001000000000000000000000000000000000000000000010000000000000000001110101000001010000000000000000000001100100000001000101000111011010001000100010000000000001000100000000000000000010001000100001001000010001111000000000000000000
// X5Y12, linear_LMDPL
`define Tile_X5Y12_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001100000010000010001110000000000010100000000000000000000000110000000000111000111010000010100010000010000000110000110000000000001110001010110011000011000101010101010100001000001000000000000100110100000000000000000000000111010101110010000000000000
// X6Y12, nonlinear_LMDPL
`define Tile_X6Y12_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100001100000000000000000000000000000000000011000011000000000000000000101000100000000000000000000000001010000000000000001000100000010010000000000000000000000000000000101010001000101000000000000100010011001000000000000000000001010100000000000000000000000000000000000000000101001100100001
// X7Y12, linear_LMDPL
`define Tile_X7Y12_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000101010101010000000000000000000100000001100101100101110101110010101010101010100000000100000001101111010101110000000000000000011001111111110000000000000000000
// X8Y12, ctrl_to_sec
`define Tile_X8Y12_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X9Y12, combined_WDDL
`define Tile_X9Y12_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000010000000000000100000000001000100101010110000101000001100000000101111111010110100000000
// X10Y12, ctrl_IO
`define Tile_X10Y12_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X0Y13, W_IO_custom
`define Tile_X0Y13_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000001000001000000000000000000000000000000000000000000000000000110111101000000000000000000000000001001000000000000000000
// X1Y13, linear_LMDPL
`define Tile_X1Y13_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011000100000000000000000000000000000000000000000000000000000000000000001010000010010000000000000000101000101010101010101010100010001100000100000011000000000010100000110000000000000000110000000000010101010101010100000000000000000011001100100000000000000000000000000001010000110000000000000000
// X2Y13, linear_LMDPL
`define Tile_X2Y13_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000010000110000000000000000000000000000000000000000000000000000000010100010101000010000000000000000000000001010001000001010100000000000000010100010000000000000000000000000100011001111001100000000010101010101010100000000000000000000000101000011000000000000000011101101100110100000000000000000
// X3Y13, nonlinear_LMDPL
`define Tile_X3Y13_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000001100001100000100000000000000000000000000001100010100110000010000000000000000000000000000000000000100000010010010100010100010011000101010101010000000000000000000000010101000001000101000100110010101010101010100000000000100000001010000010010000000000000000010101001000000110000000000000000
// X4Y13, linear_LMDPL
`define Tile_X4Y13_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110011000000100000000000000000000000000000110000000000100000101100110000000000000000000000000000000000000000000000001100110000001010101000000010000000000000000000000000100000001000100000100010000000000100000010000010000000000000000000000000101111101011101000000000001000001000101000001000
// X5Y13, linear_LMDPL
`define Tile_X5Y13_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000100000000000000000000000110000000000000000000000000000000000000011000000001100000000000000010011000000000011110000000000100000000000000000000000001000001010000010100101000010000000000000000000000000001010001010100010000010000000000100000000000000000000000000000000000000100110111100100000000000010000001011110000001011
// X6Y13, nonlinear_LMDPL
`define Tile_X6Y13_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000100000000000000000000000000000111000000000000000000000000000000000000100000000000000000000000000101000100000000000000000000000001010000000000000000000100011100011000000000000000000000000000000000111001000100000010000000101010100010000000000000000000011000000000000000000001100110000001100110010110000000000000000
// X7Y13, linear_LMDPL
`define Tile_X7Y13_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000100000010000000011000010000000000000000000000000000000000000000000000000000000000000000000101010101000000000000000000000111110001000001000101010101010000101000101010100000000111000111101000011101100000001010000000000001101110110000100000000000000
// X8Y13, ctrl_to_sec
`define Tile_X8Y13_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X9Y13, combined_WDDL
`define Tile_X9Y13_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000011000000000000110000000101010100101010100000101000001011011010000000001011111000000000
// X10Y13, ctrl_IO
`define Tile_X10Y13_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X0Y14, W_IO_custom
`define Tile_X0Y14_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000001000001000000000000000000000000000000000000000000000000000000001101010100000000000000000000000000001101000000000000
// X1Y14, linear_LMDPL
`define Tile_X1Y14_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010000010000000000000000000000000001010101010101010101010001000111000000010000000000000000000100000111101110100100000000000010101010001010100000000000000000011001101001001000000000000000000010010000000100000000001010000
// X2Y14, linear_LMDPL
`define Tile_X2Y14_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000110000000000000000000000000000000000000000000000000011001111000000000000000000000000001100001000101001010000000010100011101100000000000000000000000011101110001000001010100000000000000010000010000000000000100000000000100010001010001000000010010001000100010000000000000000000000000000000000101110111010100101100001011000110000000000000000
// X3Y14, nonlinear_LMDPL
`define Tile_X3Y14_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000010000011110010100011001010101010101010000000001100000000101000101000001000101000101010010000000100010000000000000000000000000000000000101110001011101001000000001100000000000000000000
// X4Y14, linear_LMDPL
`define Tile_X4Y14_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000000000000000000000000000000000000000000000000101100000000001000000000000000000000100010000000000010110010001000000000100000100000000011001100000000000000000010001000000100100010100000000000000000000000000000000000000000001000000000001000010101010101010100000000001000100100001101000100000000000000000010011010110110100000000000000000
// X5Y14, linear_LMDPL
`define Tile_X5Y14_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000001000001000000000000000000000000000000000000000000000000000011001111001100000001000010000000000000100000000000000000000000000010100010100110001010001110100010011110000000000000000000000000001010111010100110110110010101010101010100000000001000000011000000100011000000000000000000000001010010010000000000000000
// X6Y14, nonlinear_LMDPL
`define Tile_X6Y14_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000001011000000000000000000000000000000001000110001110000110000000000101000100000000000000000000000001010100100000000000000101100100000000000000000000000000000000000001000000000100000100000010001000100010000000000000000100000000000000000100100110100000010110000001100100000000000000000
// X7Y14, linear_LMDPL
`define Tile_X7Y14_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000001000010000000001001000000001000000000000000000000000100000000000010000000000000000000101010001011000000000000000000100000001000001011111011101000010101010100010000000000100000001010100100000000000000000001000111111000111110100000000000000000
// X8Y14, ctrl_to_sec
`define Tile_X8Y14_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000
// X9Y14, combined_WDDL
`define Tile_X9Y14_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000000000000000000100000000000000000000000000000000000000000000000001000000000000000010000000000000000000000000000101010111101000000000100011000011011010000000001011111000000000
// X10Y14, ctrl_IO
`define Tile_X10Y14_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X0Y15, W_IO_custom
`define Tile_X0Y15_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000001000001000000000000000000000000000000000000000000000000000000001101010110000000000000000000100010001000000000000000
// X1Y15, linear_LMDPL
`define Tile_X1Y15_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000011000000000000000000000000000010001111000000000000000011000000011110000010000000000000000000101000101010011111101010101001001000001000000010000000000011100000100000000010001001100000000000000100010001000100000000000000001100110010011100000000000000000000000000000000001011100111001010
// X2Y15, linear_LMDPL
`define Tile_X2Y15_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000100000000000000000000000001100000000000000000000000000000000000000000000001000000000000011110010100000000000000000000000000000000010000110101111010010000001000010000010000000000000000000000000000010011010001001000110010101010101010100000000000000001011101111001011000000000000000000000011011001010000000000000000
// X3Y15, nonlinear_LMDPL
`define Tile_X3Y15_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000011000000001100110000000000001000000000000000000000000000000011000010001010010000100001101010101000000000000000000000000010101000001000101000101010000001000100010000000000001000000000000000000000101110001011101000001001001010000100000000000000
// X4Y15, linear_LMDPL
`define Tile_X4Y15_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000001100000000000000000000000000001100000100001100000100100000000000010000100000000000001100000000000000000010001000000000100000100000000000000000000010000000000000000000001001000000000000000100010001000100000000000000000011001001000010000000000000000000000000000000001100100110011001
// X5Y15, linear_LMDPL
`define Tile_X5Y15_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000100000000000000000000000000000000001100111000000011001110000000000000100000000000000000000000000010100010100010001010000000100000100001000000000000000000000000001001001000101010001010010101010101010100001000000000001000100111001000000000000000000010011010100011000000000000000000
// X6Y15, nonlinear_LMDPL
`define Tile_X6Y15_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000010000000101000100000000000000000000000001010100000001000000000001000100000110000000000000000000000000000111000000000101100101100010101010101010100000000000000000011110010010011000000000000000001000000010000000000000000000000
// X7Y15, linear_LMDPL
`define Tile_X7Y15_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001100000000000000000000000011001100100000100000000000000000001000000000000000000000000000000000001000000000000000000011101000000000000000000000000000101011001000001000001011101000010101010101010100000000100011101000111010001101000000000000000010101011101110000000000000000000
// X8Y15, ctrl_to_sec
`define Tile_X8Y15_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X9Y15, combined_WDDL
`define Tile_X9Y15_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000011000000000000000000000000000000111110000000000000110000000000000100010000101000000000100000000011111011000000000000000010001011
// X10Y15, ctrl_IO
`define Tile_X10Y15_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X0Y16, W_IO_custom
`define Tile_X0Y16_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000001000001000000000000000000000000000000000000000000000100000000001001010100000000000000000000000100000001000000000000
// X1Y16, linear_LMDPL
`define Tile_X1Y16_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000010000000000000000000000000000010000000000000000000000110010000010000000000000000000000000001010110011101010100100111000001000000010000000000000000000100000000010001010100000000000010101010000000000000000000000000111001000000000000000000101010100000100000000000000000011000110
// X2Y16, linear_LMDPL
`define Tile_X2Y16_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000100010000010100000000010000000111111000000000000000000100011000000000010001010001000000010010100010001010100110000001111001010100110101100000000000000000010000000000010000000010101010000
// X3Y16, nonlinear_LMDPL
`define Tile_X3Y16_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000111100110000110000000000000100000000000000000000000010100000010000000000000000000000000000001000000000000000000000000000000000000001000101000000010000100010001000000000000000000000000000001000001000101000101010010101010101010100000000000000000001001101000000000000000000000011001001000110010000000000000000
// X4Y16, linear_LMDPL
`define Tile_X4Y16_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000100000000000000000000111100000000010001110011000100101010000000011100000000000001000000001000110010001000110000101000000000000000000000000000000000000000000100001010010100000100000000000000000010000010001000100000000000000000001100100011010000000000000000001100100110011001
// X5Y16, linear_LMDPL
`define Tile_X5Y16_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000011000000000000000000000000011100001000010000000000010000000000001100000000000000000000000000000100000110000000100010000000110000100000000000000000000000000001100001100001001111100100100000100010000000000000000000000000001010000100101010000010000100010001000100000000001000000011010001000011000000000000000000000000000000001010100011011001
// X6Y16, nonlinear_LMDPL
`define Tile_X6Y16_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110011000000000000000000000000000000000000110000000000110000100000000000000000000000000000000000000000000000000000000000000010000000001000000000000000000000000000000000010001000000000000000000100000000000000000000000000000000000001000000000100000100000010001000100010000000000000000100000000000000000101011001100110011001000101010110000000000000000
// X7Y16, linear_LMDPL
`define Tile_X7Y16_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100110000110000000000000000001100000000000000000000000000000000001100000000000000000010101000000000000000000000000000100000001000001000111010101000000000000000000000000000100000000000000000000000000000100001010000000000000000001000111010111000
// X8Y16, ctrl_to_sec
`define Tile_X8Y16_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X9Y16, combined_WDDL
`define Tile_X9Y16_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000001000000000000000000000000000110010000000000000000000001000001101100100101000001100100000000000000000000000001001100100000000
// X10Y16, ctrl_IO
`define Tile_X10Y16_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X0Y17, W_IO_custom
`define Tile_X0Y17_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000001000001000000000000000000000000000000000000000000000000000000001111111110000000000000000100000000000000000000000000
// X1Y17, linear_LMDPL
`define Tile_X1Y17_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000100000000000000000000000000000000000100000000000000000000000000000000000000000001111001100000000000000000000000000000010000010000000000000001100101000111110010000111110100000001000000000000010000000000000100000100000000000000000100000000000000100010001000100000000000000001011101111001001000000000000000000000000000000001100100110101010
// X2Y17, linear_LMDPL
`define Tile_X2Y17_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000011100000000000000000000000000000000010000011110000000011000000101010000000000000000000000000000000000010001010001000000000000101010001010100000000000000000100000100100100000000000000000000001101000010100001000000110000
// X3Y17, nonlinear_LMDPL
`define Tile_X3Y17_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000001100000000000000000000000000001100000000001100000000001100000000000000000000000000000000000011000011000000000000110000000000010100000000000000000000000000000010000000000000000000000000100010001000000000000000000001000010001000001000001000011001010101010101010100000000001000000011010000110011000000000000000000011010101110100000000000000000
// X4Y17, linear_LMDPL
`define Tile_X4Y17_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000100000000111000000000000000000000000000000100000000000100000000000101010000000010000000000000000000000001000000011001100000000110000000000100000000000000011000000000000000000001000100000001000000101000001000100000000000000000001000001000000000010100000000000000001000000001011000010101011
// X5Y17, linear_LMDPL
`define Tile_X5Y17_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000110000000000000000000000000000000000000000000000000000010100000000000100000000000000001100000000000100100000000011001010000010001000100000000000000000000000001100100000101100100000111000001100100010000000000000000000000000001010000000001010000000010100010101010100000000000011001010110010111010000000000000000000110000100101100000001100000000
// X6Y17, nonlinear_LMDPL
`define Tile_X6Y17_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000010000000000000000100000000000000000000000000000000000000000000000000000000001010100000000010000000011111100000000000000000000000000000000000101010000100011100000010101010101010100000000000000000110101001010110000000000000000000111100100100110000000000000000
// X7Y17, linear_LMDPL
`define Tile_X7Y17_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000100000100000000000111111100010101100000000000000100000100000000000000000000000000000000000001000000000000010101000110000000000000000000000101010000011001100000010100011000101010101010100000000100010101011110010101011000000000000000000001010100110011110000000000000
// X8Y17, ctrl_to_sec
`define Tile_X8Y17_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X9Y17, combined_WDDL
`define Tile_X9Y17_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100010000000000000000000001000000101010100100000001000110000110011101100000000001001110100000000
// X10Y17, ctrl_IO
`define Tile_X10Y17_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X0Y18, W_IO_custom
`define Tile_X0Y18_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000001011101010000000000000000000000000000000000000010000
// X1Y18, linear_LMDPL
`define Tile_X1Y18_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000110010000010000000000000000000000000001110000000000010100011111000000000000010000000000000000000000000010000000000100000000000000101010100010000000000000000000001010000000000000000001100010100000001010000011011000000000000
// X2Y18, linear_LMDPL
`define Tile_X2Y18_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000010100010000000000000000000000000000000011010100000000000000000000000000110000000000000000000000000000110011010000000000000000000000101010000000000000000000110010000011000000000000000000111100000100010001000100000000001010001011101111001011000000000000000000000000000000001100101010101000
// X3Y18, nonlinear_LMDPL
`define Tile_X3Y18_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000001100110000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000100110000000000000000000000000000000001000001000000000101010010001010101010100000000000000000000000100100011101100000000000000110000100010110000000000000000
// X4Y18, linear_LMDPL
`define Tile_X4Y18_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000100111100100000000000010000101010110000000000000000000000000000001000000010000001000110001000000000001000000000000000001100000000001000000000101000001000000000000000000000000000001000100000000000000000001100100011000000000000000000001110101111101101
// X5Y18, linear_LMDPL
`define Tile_X5Y18_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000010011000011100010001000110000000000000000000010000000110000110000100000001000000000100010000000000000000000000000001010000000001010000000010101010101010100001000000000000110111000110001000000000000000000010100001000110000000000000000
// X6Y18, nonlinear_LMDPL
`define Tile_X6Y18_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000000000000000000000000000000000000000010000000110000000000000000000000000000000000000000110000000010110000110000000000000000000000000000000000000000000000000000000000000000000010101000000000000000000000000000010000000000000000100010100000010001000100010000000000010000100000000000000000100011001100100000111100110011000000000000000000
// X7Y18, linear_LMDPL
`define Tile_X7Y18_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000100000000000000000100000000000000000000000100000000000000000000000110000110000000010000000000000000000000000001100000000000010101000000000000000000011000000000000001000000000000010100000000101010001000100000000100000001011100011001010000000000000000000001100000000000010000000010001
// X8Y18, ctrl_to_sec
`define Tile_X8Y18_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X9Y18, combined_WDDL
`define Tile_X9Y18_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000010000000000000000000001100000100010000100000000000100000100010011101000000000000000010111001
// X10Y18, ctrl_IO
`define Tile_X10Y18_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X0Y19, W_IO_custom
`define Tile_X0Y19_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101011100000000000000000100100000000000000000000000
// X1Y19, linear_LMDPL
`define Tile_X1Y19_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000011001100000000000000000000000011000000000000000100000000000010000010000000000000001100111100000010100010000011100000001000000000000010000000000000110000100000100000000000100000000100010001000100010000000000000000000000000000000000100010111010101000010010000000010000000000000000
// X2Y19, linear_LMDPL
`define Tile_X2Y19_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000110000110000000000000000000000000000000000000000000011100010100010000000100000000000000000000000001010100000000000001010001000001000000000000000000000000000000000000000000000000000100000010001000100010000000000000000000000000000000000101110011100100110001111100110010000000000000000
// X3Y19, nonlinear_LMDPL
`define Tile_X3Y19_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001100000000000000000000000011000000000111001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000101010000000000000000000000010000010001000001000000000101000010101010101010000000000001001000011000100100000000000000000100000100100001110100000000000000000
// X4Y19, linear_LMDPL
`define Tile_X4Y19_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000010000000000000111111000000000000000000000000000000001100000001100000000001001000000100001000000000000000000000000000001000000001001000000000000000000000000010000010000000000000000000000000100101001000100100000000000000000011000101000001
// X5Y19, linear_LMDPL
`define Tile_X5Y19_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100110000000000000000000000000000000000100000011100001000010000100010001000000000000000001000000000000000000000000010100000000001110100000010000000000000000000000000110010000000000001000000010001000000010000000000000000000000000000000000010100010100000110011000000010110000000000100000
// X6Y19, nonlinear_LMDPL
`define Tile_X6Y19_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000000000000000000000000000000000000000010000000001000100000000000000000000000000000000000000000000000000000000000000000010000010000000000000000000000000001010000000000000000001101101000000000000000000000001000000000000000000000000010000000010001000101010100000000001111110000000010110001111011010000000001101010010101100000000000000000
// X7Y19, linear_LMDPL
`define Tile_X7Y19_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000001000101100001100000000100000100000000000111100000000001000000000000000000000000000000000000000000000000000000000000000000000000010101000000000000000001000000000101010001000000000000010100000000101010001000100000000100010101010100111101101000000000000000000001100000000000010000000010001
// X8Y19, ctrl_to_sec
`define Tile_X8Y19_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X9Y19, combined_WDDL
`define Tile_X9Y19_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000110000000101010100000000000000000000000010101100000000001000111100000000
// X10Y19, ctrl_IO
`define Tile_X10Y19_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X0Y20, W_IO_custom
`define Tile_X0Y20_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101010100000000000000000000100010010101000000000000
// X1Y20, linear_LMDPL
`define Tile_X1Y20_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000100000000010110010000000000000000000000000000010010001110000100011111000000000000010000000000000000000000000000000000000100000000000010100010101010100000000000000000100001100110000000000000000000000010000101110000000110100000000
// X2Y20, linear_LMDPL
`define Tile_X2Y20_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000010000000010000001100010000000110000000000000000000000001101100010000000001111000100000000000000000000000000000000000000000100000000000000000000010001000100010000000000000000000000000000000000110010101011101011011110111010010000000000000000
// X3Y20, nonlinear_LMDPL
`define Tile_X3Y20_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000100000100000000000000000000000000110000000000110000000011000000000000001100000000000000000000000011000000001111000000000000000000000000010000000000000000000000000010000000000000000000000000101000000000000000000000000000000000001001001000000000101000010100000001000100000000000000000010000000000001000010000000000010000000000000000000111001111101
// X4Y20, linear_LMDPL
`define Tile_X4Y20_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000010000000000000000000000000000111100000000000000000000000000000000000000000000000000000000110000000000110000000000000000011000000001000000001100110000000000010000000010001100000000000100010001000100000000001000101001110010001011000000000000000000000000000000000100000100110010
// X5Y20, linear_LMDPL
`define Tile_X5Y20_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000001100000100000000000000000010000000000000000100000000110010001000000000000000000000000010000000000011000011100011000010001000000000000000000000000000000000111111000000000001000000010101010101010100000000000000001010000111001000000000000000000000110000000001000000000000000000
// X6Y20, nonlinear_LMDPL
`define Tile_X6Y20_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000000000000000000000000000000000000000010000000001000000011110000000000000000000000000000000011110000001000000000000000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000000100000000000000000000000000000010100010001000100000000100000100010000000110011000000000000000001000000000000000000110010111001
// X7Y20, linear_LMDPL
`define Tile_X7Y20_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000001000000000011111100000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000010000000000101010001000100000000100000001110101010011001000000000000000000001100000000000010000000010001
// X8Y20, ctrl_to_sec
`define Tile_X8Y20_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X9Y20, combined_WDDL
`define Tile_X9Y20_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X10Y20, ctrl_IO
`define Tile_X10Y20_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X0Y21, W_IO_custom
`define Tile_X0Y21_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X1Y21, linear_LMDPL
`define Tile_X1Y21_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000010000000000000000000000000000010000000000000100000000000000011001100000000000000000000100000000000000000000000110011010101010101010100000000000000001001110110111000000000000000000000010100010000110000000000000000
// X2Y21, linear_LMDPL
`define Tile_X2Y21_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000100000000000000000000000100010000000000000000000000000000000001100100010001100001100110000000000010100000000000000000000000000010000010000000000000000010001000101010000000000000000000000000000010000110010100000110010011100010000110000000000000000
// X3Y21, nonlinear_LMDPL
`define Tile_X3Y21_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000011110000000000000000000000000011001011000000000000000011000011001011000000000000000000000000000011000000000000000000000000001000000100000000000000000010000010000000000100000000101001010101010101000100000000001010000011000000000010000000000000000010111100100100000000000000000110
// X4Y21, linear_LMDPL
`define Tile_X4Y21_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000110000100000001100000000000001000000000000000001000000000000000000000000000000000011101000000000000000000000000000000000100000000010000000000000000101010101010100000000000000000100010001001000000000000000000000000000000000011100000000000000
// X5Y21, linear_LMDPL
`define Tile_X5Y21_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001010000000000000000000000000010101000000000000000000000000010001000000000000000000000000000000000000000000000100000000000000000110011000000000000000000000000000000001101000001001100010101010101010100001000000000000101010000110001000000000000000010101001000110010000000000000000
// X6Y21, nonlinear_LMDPL
`define Tile_X6Y21_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000001100001100000000000001000000000000000000000000001000000001000000000100000000000000000000000000000000001000001000000000000000000000110000000011010101010101010100000000000000000001010000110001000000000000000010011110111011100000000000000000
// X7Y21, linear_LMDPL
`define Tile_X7Y21_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000110000000000000000000000001100000000110000000011000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000001000000000000000000000000000000000000000010101010101010100000000000000001110110111011110000000000000000010101001111011010000000000000000
// X8Y21, ctrl_to_sec
`define Tile_X8Y21_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X9Y21, combined_WDDL
`define Tile_X9Y21_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X10Y21, ctrl_IO
`define Tile_X10Y21_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X0Y22, W_IO_custom
`define Tile_X0Y22_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X1Y22, linear_LMDPL
`define Tile_X1Y22_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000011000000000000000000001000000011000000000000110000000000000000000000000000000000000000000000000000000000000000000000000101010101010100000000000000001000101010001010000000000000000000000111001100100110000000000000
// X2Y22, linear_LMDPL
`define Tile_X2Y22_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000010001000000000000000000000000000000000000000000000000000000000000000000110011000000000000000000000000000000000100110111000000000100000000000000000000000000000000000000000000010000010000000000010000000100010001000100000000000000001100100010001100000000000000000000000000000000001000101010011010
// X3Y22, nonlinear_LMDPL
`define Tile_X3Y22_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000011000000000011000000001100000100000000000000000000000000100000000000000000000000000000001000000000000000000010000000000000010011000000000000100000000100010101000100000000000000011011000110001010000000000000000000000000101000000111011000000111
// X4Y22, linear_LMDPL
`define Tile_X4Y22_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000011000000001100000000000000001011001011100000000000000100000000000000000000000000000000010000000000000000000000000000000000000000000000000000010001000100010000000000000000100000000000000000000100100001001011001011100110010000000000000000
// X5Y22, linear_LMDPL
`define Tile_X5Y22_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000011000000000000000000000000000011001111000000000000000011000011000000000000000000110000000000000000000000000000000000000000000000000011000000000000000000010101010101010100000000000000001010101100110010000000000000000010111000101010000000000000000000
// X6Y22, nonlinear_LMDPL
`define Tile_X6Y22_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000100000100000000000000000000000000000000000000000000000000000000000000000
// X7Y22, linear_LMDPL
`define Tile_X7Y22_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000
// X8Y22, ctrl_to_sec
`define Tile_X8Y22_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X9Y22, combined_WDDL
`define Tile_X9Y22_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X10Y22, ctrl_IO
`define Tile_X10Y22_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X0Y23, W_IO_custom
`define Tile_X0Y23_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X1Y23, linear_LMDPL
`define Tile_X1Y23_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X2Y23, linear_LMDPL
`define Tile_X2Y23_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100110000000000000000000000000000000000000000000000001100110000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000100000000110000000000000000000011001010010011000000000000000000
// X3Y23, nonlinear_LMDPL
`define Tile_X3Y23_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001100000000000000000000000011001000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000010101010101010000000000001000001100000001000000000000000000111011011010111010010000000000000000
// X4Y23, linear_LMDPL
`define Tile_X4Y23_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X5Y23, linear_LMDPL
`define Tile_X5Y23_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X6Y23, nonlinear_LMDPL
`define Tile_X6Y23_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000001000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X7Y23, linear_LMDPL
`define Tile_X7Y23_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X8Y23, ctrl_to_sec
`define Tile_X8Y23_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X9Y23, combined_WDDL
`define Tile_X9Y23_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
// X10Y23, ctrl_IO
`define Tile_X10Y23_Emulate_Bitstream 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000

