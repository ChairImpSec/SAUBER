//-----------------------------------------

module top(input wire [59:0] io_in_0t, io_in_0f, io_in_1t, io_in_1f, ctrl_io_in_0t, ctrl_io_in_0f,  output wire [59:0] io_out_0t, io_out_0f, io_out_1t, io_out_1f, io_oeb, ctrl_io_out_0t, ctrl_io_out_0f, ctrl_io_oeb);


    assign io_oeb      = 60'b11111111000000000000;
    assign ctrl_io_oeb = 60'b10000;

    AES_SAUBER_Pipeline_d1 generated_module (
        .port_in(io_in_0t[7:0]),

        .start(ctrl_io_in_0t[1]),

        .done(ctrl_io_out_0t[5]),

        .port_out(io_out_0t[19:12]),

    );

endmodule

/* modified netlist. Source: module AES in file /mnt/c/Users/amirm/Desktop/Papers_in_progress/SAUBER/Design for our FPGA/6-AES_EncSerial_PortSerial/4-AGEMA/AES.v */
/* 0 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 1 register stage(s) in total */

module AES_SAUBER_Pipeline_d1 (port_in, start, port_out, done);
    input [7:0] port_in ;
    input start ;
    output [7:0] port_out ;
    output done ;
    wire selMC ;
    wire selXOR ;
    wire enRCon ;
    wire intFinal ;
    wire enKS ;
    wire intselXOR ;
    wire notFirst ;
    wire ctrl_n24 ;
    wire ctrl_n19 ;
    wire ctrl_n18 ;
    wire ctrl_n17 ;
    wire ctrl_n14 ;
    wire ctrl_n13 ;
    wire ctrl_n12 ;
    wire ctrl_n11 ;
    wire ctrl_n10 ;
    wire ctrl_n9 ;
    wire ctrl_n4 ;
    wire ctrl_finalStep ;
    wire ctrl_n5 ;
    wire ctrl_seq4Out_1_ ;
    wire ctrl_seq4In_1_ ;
    wire ctrl_nRstSeq4 ;
    wire ctrl_n22 ;
    wire ctrl_seq6Out_4_ ;
    wire ctrl_seq6In_1_ ;
    wire ctrl_seq6In_2_ ;
    wire ctrl_seq6In_3_ ;
    wire ctrl_seq6In_4_ ;
    wire ctrl_seq6_SFF_0_n2 ;
    wire ctrl_seq6_SFF_0_n1 ;
    wire ctrl_seq6_SFF_0_QD ;
    wire ctrl_seq6_SFF_0_MUXInst_Y ;
    wire ctrl_seq6_SFF_0_MUXInst_X ;
    wire ctrl_seq6_SFF_1_n2 ;
    wire ctrl_seq6_SFF_1_n1 ;
    wire ctrl_seq6_SFF_1_QD ;
    wire ctrl_seq6_SFF_1_MUXInst_Y ;
    wire ctrl_seq6_SFF_1_MUXInst_X ;
    wire ctrl_seq6_SFF_2_n2 ;
    wire ctrl_seq6_SFF_2_n1 ;
    wire ctrl_seq6_SFF_2_QD ;
    wire ctrl_seq6_SFF_2_MUXInst_Y ;
    wire ctrl_seq6_SFF_2_MUXInst_X ;
    wire ctrl_seq6_SFF_3_n2 ;
    wire ctrl_seq6_SFF_3_n1 ;
    wire ctrl_seq6_SFF_3_QD ;
    wire ctrl_seq6_SFF_3_MUXInst_Y ;
    wire ctrl_seq6_SFF_3_MUXInst_X ;
    wire ctrl_seq6_SFF_4_n2 ;
    wire ctrl_seq6_SFF_4_n1 ;
    wire ctrl_seq6_SFF_4_QD ;
    wire ctrl_seq6_SFF_4_MUXInst_Y ;
    wire ctrl_seq6_SFF_4_MUXInst_X ;
    wire ctrl_seq4_SFF_0_n2 ;
    wire ctrl_seq4_SFF_0_n1 ;
    wire ctrl_seq4_SFF_0_QD ;
    wire ctrl_seq4_SFF_0_MUXInst_Y ;
    wire ctrl_seq4_SFF_0_MUXInst_X ;
    wire ctrl_seq4_SFF_1_n2 ;
    wire ctrl_seq4_SFF_1_n1 ;
    wire ctrl_seq4_SFF_1_QD ;
    wire ctrl_seq4_SFF_1_MUXInst_Y ;
    wire ctrl_seq4_SFF_1_MUXInst_X ;
    wire MUX_StateIn_mux_inst_0_Y ;
    wire MUX_StateIn_mux_inst_0_X ;
    wire MUX_StateIn_mux_inst_1_Y ;
    wire MUX_StateIn_mux_inst_1_X ;
    wire MUX_StateIn_mux_inst_2_Y ;
    wire MUX_StateIn_mux_inst_2_X ;
    wire MUX_StateIn_mux_inst_3_Y ;
    wire MUX_StateIn_mux_inst_3_X ;
    wire MUX_StateIn_mux_inst_4_Y ;
    wire MUX_StateIn_mux_inst_4_X ;
    wire MUX_StateIn_mux_inst_5_Y ;
    wire MUX_StateIn_mux_inst_5_X ;
    wire MUX_StateIn_mux_inst_6_Y ;
    wire MUX_StateIn_mux_inst_6_X ;
    wire MUX_StateIn_mux_inst_7_Y ;
    wire MUX_StateIn_mux_inst_7_X ;
    wire stateArray_nReset_selMC ;
    wire stateArray_S00reg_gff_1_SFF_0_MUXInst_Y ;
    wire stateArray_S00reg_gff_1_SFF_0_MUXInst_X ;
    wire stateArray_S00reg_gff_1_SFF_1_MUXInst_Y ;
    wire stateArray_S00reg_gff_1_SFF_1_MUXInst_X ;
    wire stateArray_S00reg_gff_1_SFF_2_MUXInst_Y ;
    wire stateArray_S00reg_gff_1_SFF_2_MUXInst_X ;
    wire stateArray_S00reg_gff_1_SFF_3_MUXInst_Y ;
    wire stateArray_S00reg_gff_1_SFF_3_MUXInst_X ;
    wire stateArray_S00reg_gff_1_SFF_4_MUXInst_Y ;
    wire stateArray_S00reg_gff_1_SFF_4_MUXInst_X ;
    wire stateArray_S00reg_gff_1_SFF_5_MUXInst_Y ;
    wire stateArray_S00reg_gff_1_SFF_5_MUXInst_X ;
    wire stateArray_S00reg_gff_1_SFF_6_MUXInst_Y ;
    wire stateArray_S00reg_gff_1_SFF_6_MUXInst_X ;
    wire stateArray_S00reg_gff_1_SFF_7_MUXInst_Y ;
    wire stateArray_S00reg_gff_1_SFF_7_MUXInst_X ;
    wire stateArray_S01reg_gff_1_SFF_0_MUXInst_Y ;
    wire stateArray_S01reg_gff_1_SFF_0_MUXInst_X ;
    wire stateArray_S01reg_gff_1_SFF_1_MUXInst_Y ;
    wire stateArray_S01reg_gff_1_SFF_1_MUXInst_X ;
    wire stateArray_S01reg_gff_1_SFF_2_MUXInst_Y ;
    wire stateArray_S01reg_gff_1_SFF_2_MUXInst_X ;
    wire stateArray_S01reg_gff_1_SFF_3_MUXInst_Y ;
    wire stateArray_S01reg_gff_1_SFF_3_MUXInst_X ;
    wire stateArray_S01reg_gff_1_SFF_4_MUXInst_Y ;
    wire stateArray_S01reg_gff_1_SFF_4_MUXInst_X ;
    wire stateArray_S01reg_gff_1_SFF_5_MUXInst_Y ;
    wire stateArray_S01reg_gff_1_SFF_5_MUXInst_X ;
    wire stateArray_S01reg_gff_1_SFF_6_MUXInst_Y ;
    wire stateArray_S01reg_gff_1_SFF_6_MUXInst_X ;
    wire stateArray_S01reg_gff_1_SFF_7_MUXInst_Y ;
    wire stateArray_S01reg_gff_1_SFF_7_MUXInst_X ;
    wire stateArray_S02reg_gff_1_SFF_0_MUXInst_Y ;
    wire stateArray_S02reg_gff_1_SFF_0_MUXInst_X ;
    wire stateArray_S02reg_gff_1_SFF_1_MUXInst_Y ;
    wire stateArray_S02reg_gff_1_SFF_1_MUXInst_X ;
    wire stateArray_S02reg_gff_1_SFF_2_MUXInst_Y ;
    wire stateArray_S02reg_gff_1_SFF_2_MUXInst_X ;
    wire stateArray_S02reg_gff_1_SFF_3_MUXInst_Y ;
    wire stateArray_S02reg_gff_1_SFF_3_MUXInst_X ;
    wire stateArray_S02reg_gff_1_SFF_4_MUXInst_Y ;
    wire stateArray_S02reg_gff_1_SFF_4_MUXInst_X ;
    wire stateArray_S02reg_gff_1_SFF_5_MUXInst_Y ;
    wire stateArray_S02reg_gff_1_SFF_5_MUXInst_X ;
    wire stateArray_S02reg_gff_1_SFF_6_MUXInst_Y ;
    wire stateArray_S02reg_gff_1_SFF_6_MUXInst_X ;
    wire stateArray_S02reg_gff_1_SFF_7_MUXInst_Y ;
    wire stateArray_S02reg_gff_1_SFF_7_MUXInst_X ;
    wire stateArray_S03reg_gff_1_SFF_0_MUXInst_Y ;
    wire stateArray_S03reg_gff_1_SFF_0_MUXInst_X ;
    wire stateArray_S03reg_gff_1_SFF_1_MUXInst_Y ;
    wire stateArray_S03reg_gff_1_SFF_1_MUXInst_X ;
    wire stateArray_S03reg_gff_1_SFF_2_MUXInst_Y ;
    wire stateArray_S03reg_gff_1_SFF_2_MUXInst_X ;
    wire stateArray_S03reg_gff_1_SFF_3_MUXInst_Y ;
    wire stateArray_S03reg_gff_1_SFF_3_MUXInst_X ;
    wire stateArray_S03reg_gff_1_SFF_4_MUXInst_Y ;
    wire stateArray_S03reg_gff_1_SFF_4_MUXInst_X ;
    wire stateArray_S03reg_gff_1_SFF_5_MUXInst_Y ;
    wire stateArray_S03reg_gff_1_SFF_5_MUXInst_X ;
    wire stateArray_S03reg_gff_1_SFF_6_MUXInst_Y ;
    wire stateArray_S03reg_gff_1_SFF_6_MUXInst_X ;
    wire stateArray_S03reg_gff_1_SFF_7_MUXInst_Y ;
    wire stateArray_S03reg_gff_1_SFF_7_MUXInst_X ;
    wire stateArray_S10reg_gff_1_SFF_0_MUXInst_Y ;
    wire stateArray_S10reg_gff_1_SFF_0_MUXInst_X ;
    wire stateArray_S10reg_gff_1_SFF_1_MUXInst_Y ;
    wire stateArray_S10reg_gff_1_SFF_1_MUXInst_X ;
    wire stateArray_S10reg_gff_1_SFF_2_MUXInst_Y ;
    wire stateArray_S10reg_gff_1_SFF_2_MUXInst_X ;
    wire stateArray_S10reg_gff_1_SFF_3_MUXInst_Y ;
    wire stateArray_S10reg_gff_1_SFF_3_MUXInst_X ;
    wire stateArray_S10reg_gff_1_SFF_4_MUXInst_Y ;
    wire stateArray_S10reg_gff_1_SFF_4_MUXInst_X ;
    wire stateArray_S10reg_gff_1_SFF_5_MUXInst_Y ;
    wire stateArray_S10reg_gff_1_SFF_5_MUXInst_X ;
    wire stateArray_S10reg_gff_1_SFF_6_MUXInst_Y ;
    wire stateArray_S10reg_gff_1_SFF_6_MUXInst_X ;
    wire stateArray_S10reg_gff_1_SFF_7_MUXInst_Y ;
    wire stateArray_S10reg_gff_1_SFF_7_MUXInst_X ;
    wire stateArray_S11reg_gff_1_SFF_0_MUXInst_Y ;
    wire stateArray_S11reg_gff_1_SFF_0_MUXInst_X ;
    wire stateArray_S11reg_gff_1_SFF_1_MUXInst_Y ;
    wire stateArray_S11reg_gff_1_SFF_1_MUXInst_X ;
    wire stateArray_S11reg_gff_1_SFF_2_MUXInst_Y ;
    wire stateArray_S11reg_gff_1_SFF_2_MUXInst_X ;
    wire stateArray_S11reg_gff_1_SFF_3_MUXInst_Y ;
    wire stateArray_S11reg_gff_1_SFF_3_MUXInst_X ;
    wire stateArray_S11reg_gff_1_SFF_4_MUXInst_Y ;
    wire stateArray_S11reg_gff_1_SFF_4_MUXInst_X ;
    wire stateArray_S11reg_gff_1_SFF_5_MUXInst_Y ;
    wire stateArray_S11reg_gff_1_SFF_5_MUXInst_X ;
    wire stateArray_S11reg_gff_1_SFF_6_MUXInst_Y ;
    wire stateArray_S11reg_gff_1_SFF_6_MUXInst_X ;
    wire stateArray_S11reg_gff_1_SFF_7_MUXInst_Y ;
    wire stateArray_S11reg_gff_1_SFF_7_MUXInst_X ;
    wire stateArray_S12reg_gff_1_SFF_0_MUXInst_Y ;
    wire stateArray_S12reg_gff_1_SFF_0_MUXInst_X ;
    wire stateArray_S12reg_gff_1_SFF_1_MUXInst_Y ;
    wire stateArray_S12reg_gff_1_SFF_1_MUXInst_X ;
    wire stateArray_S12reg_gff_1_SFF_2_MUXInst_Y ;
    wire stateArray_S12reg_gff_1_SFF_2_MUXInst_X ;
    wire stateArray_S12reg_gff_1_SFF_3_MUXInst_Y ;
    wire stateArray_S12reg_gff_1_SFF_3_MUXInst_X ;
    wire stateArray_S12reg_gff_1_SFF_4_MUXInst_Y ;
    wire stateArray_S12reg_gff_1_SFF_4_MUXInst_X ;
    wire stateArray_S12reg_gff_1_SFF_5_MUXInst_Y ;
    wire stateArray_S12reg_gff_1_SFF_5_MUXInst_X ;
    wire stateArray_S12reg_gff_1_SFF_6_MUXInst_Y ;
    wire stateArray_S12reg_gff_1_SFF_6_MUXInst_X ;
    wire stateArray_S12reg_gff_1_SFF_7_MUXInst_Y ;
    wire stateArray_S12reg_gff_1_SFF_7_MUXInst_X ;
    wire stateArray_S13reg_gff_1_SFF_0_MUXInst_Y ;
    wire stateArray_S13reg_gff_1_SFF_0_MUXInst_X ;
    wire stateArray_S13reg_gff_1_SFF_1_MUXInst_Y ;
    wire stateArray_S13reg_gff_1_SFF_1_MUXInst_X ;
    wire stateArray_S13reg_gff_1_SFF_2_MUXInst_Y ;
    wire stateArray_S13reg_gff_1_SFF_2_MUXInst_X ;
    wire stateArray_S13reg_gff_1_SFF_3_MUXInst_Y ;
    wire stateArray_S13reg_gff_1_SFF_3_MUXInst_X ;
    wire stateArray_S13reg_gff_1_SFF_4_MUXInst_Y ;
    wire stateArray_S13reg_gff_1_SFF_4_MUXInst_X ;
    wire stateArray_S13reg_gff_1_SFF_5_MUXInst_Y ;
    wire stateArray_S13reg_gff_1_SFF_5_MUXInst_X ;
    wire stateArray_S13reg_gff_1_SFF_6_MUXInst_Y ;
    wire stateArray_S13reg_gff_1_SFF_6_MUXInst_X ;
    wire stateArray_S13reg_gff_1_SFF_7_MUXInst_Y ;
    wire stateArray_S13reg_gff_1_SFF_7_MUXInst_X ;
    wire stateArray_S20reg_gff_1_SFF_0_MUXInst_Y ;
    wire stateArray_S20reg_gff_1_SFF_0_MUXInst_X ;
    wire stateArray_S20reg_gff_1_SFF_1_MUXInst_Y ;
    wire stateArray_S20reg_gff_1_SFF_1_MUXInst_X ;
    wire stateArray_S20reg_gff_1_SFF_2_MUXInst_Y ;
    wire stateArray_S20reg_gff_1_SFF_2_MUXInst_X ;
    wire stateArray_S20reg_gff_1_SFF_3_MUXInst_Y ;
    wire stateArray_S20reg_gff_1_SFF_3_MUXInst_X ;
    wire stateArray_S20reg_gff_1_SFF_4_MUXInst_Y ;
    wire stateArray_S20reg_gff_1_SFF_4_MUXInst_X ;
    wire stateArray_S20reg_gff_1_SFF_5_MUXInst_Y ;
    wire stateArray_S20reg_gff_1_SFF_5_MUXInst_X ;
    wire stateArray_S20reg_gff_1_SFF_6_MUXInst_Y ;
    wire stateArray_S20reg_gff_1_SFF_6_MUXInst_X ;
    wire stateArray_S20reg_gff_1_SFF_7_MUXInst_Y ;
    wire stateArray_S20reg_gff_1_SFF_7_MUXInst_X ;
    wire stateArray_S21reg_gff_1_SFF_0_MUXInst_Y ;
    wire stateArray_S21reg_gff_1_SFF_0_MUXInst_X ;
    wire stateArray_S21reg_gff_1_SFF_1_MUXInst_Y ;
    wire stateArray_S21reg_gff_1_SFF_1_MUXInst_X ;
    wire stateArray_S21reg_gff_1_SFF_2_MUXInst_Y ;
    wire stateArray_S21reg_gff_1_SFF_2_MUXInst_X ;
    wire stateArray_S21reg_gff_1_SFF_3_MUXInst_Y ;
    wire stateArray_S21reg_gff_1_SFF_3_MUXInst_X ;
    wire stateArray_S21reg_gff_1_SFF_4_MUXInst_Y ;
    wire stateArray_S21reg_gff_1_SFF_4_MUXInst_X ;
    wire stateArray_S21reg_gff_1_SFF_5_MUXInst_Y ;
    wire stateArray_S21reg_gff_1_SFF_5_MUXInst_X ;
    wire stateArray_S21reg_gff_1_SFF_6_MUXInst_Y ;
    wire stateArray_S21reg_gff_1_SFF_6_MUXInst_X ;
    wire stateArray_S21reg_gff_1_SFF_7_MUXInst_Y ;
    wire stateArray_S21reg_gff_1_SFF_7_MUXInst_X ;
    wire stateArray_S22reg_gff_1_SFF_0_MUXInst_Y ;
    wire stateArray_S22reg_gff_1_SFF_0_MUXInst_X ;
    wire stateArray_S22reg_gff_1_SFF_1_MUXInst_Y ;
    wire stateArray_S22reg_gff_1_SFF_1_MUXInst_X ;
    wire stateArray_S22reg_gff_1_SFF_2_MUXInst_Y ;
    wire stateArray_S22reg_gff_1_SFF_2_MUXInst_X ;
    wire stateArray_S22reg_gff_1_SFF_3_MUXInst_Y ;
    wire stateArray_S22reg_gff_1_SFF_3_MUXInst_X ;
    wire stateArray_S22reg_gff_1_SFF_4_MUXInst_Y ;
    wire stateArray_S22reg_gff_1_SFF_4_MUXInst_X ;
    wire stateArray_S22reg_gff_1_SFF_5_MUXInst_Y ;
    wire stateArray_S22reg_gff_1_SFF_5_MUXInst_X ;
    wire stateArray_S22reg_gff_1_SFF_6_MUXInst_Y ;
    wire stateArray_S22reg_gff_1_SFF_6_MUXInst_X ;
    wire stateArray_S22reg_gff_1_SFF_7_MUXInst_Y ;
    wire stateArray_S22reg_gff_1_SFF_7_MUXInst_X ;
    wire stateArray_S23reg_gff_1_SFF_0_MUXInst_Y ;
    wire stateArray_S23reg_gff_1_SFF_0_MUXInst_X ;
    wire stateArray_S23reg_gff_1_SFF_1_MUXInst_Y ;
    wire stateArray_S23reg_gff_1_SFF_1_MUXInst_X ;
    wire stateArray_S23reg_gff_1_SFF_2_MUXInst_Y ;
    wire stateArray_S23reg_gff_1_SFF_2_MUXInst_X ;
    wire stateArray_S23reg_gff_1_SFF_3_MUXInst_Y ;
    wire stateArray_S23reg_gff_1_SFF_3_MUXInst_X ;
    wire stateArray_S23reg_gff_1_SFF_4_MUXInst_Y ;
    wire stateArray_S23reg_gff_1_SFF_4_MUXInst_X ;
    wire stateArray_S23reg_gff_1_SFF_5_MUXInst_Y ;
    wire stateArray_S23reg_gff_1_SFF_5_MUXInst_X ;
    wire stateArray_S23reg_gff_1_SFF_6_MUXInst_Y ;
    wire stateArray_S23reg_gff_1_SFF_6_MUXInst_X ;
    wire stateArray_S23reg_gff_1_SFF_7_MUXInst_Y ;
    wire stateArray_S23reg_gff_1_SFF_7_MUXInst_X ;
    wire stateArray_S30reg_gff_1_SFF_0_MUXInst_Y ;
    wire stateArray_S30reg_gff_1_SFF_0_MUXInst_X ;
    wire stateArray_S30reg_gff_1_SFF_1_MUXInst_Y ;
    wire stateArray_S30reg_gff_1_SFF_1_MUXInst_X ;
    wire stateArray_S30reg_gff_1_SFF_2_MUXInst_Y ;
    wire stateArray_S30reg_gff_1_SFF_2_MUXInst_X ;
    wire stateArray_S30reg_gff_1_SFF_3_MUXInst_Y ;
    wire stateArray_S30reg_gff_1_SFF_3_MUXInst_X ;
    wire stateArray_S30reg_gff_1_SFF_4_MUXInst_Y ;
    wire stateArray_S30reg_gff_1_SFF_4_MUXInst_X ;
    wire stateArray_S30reg_gff_1_SFF_5_MUXInst_Y ;
    wire stateArray_S30reg_gff_1_SFF_5_MUXInst_X ;
    wire stateArray_S30reg_gff_1_SFF_6_MUXInst_Y ;
    wire stateArray_S30reg_gff_1_SFF_6_MUXInst_X ;
    wire stateArray_S30reg_gff_1_SFF_7_MUXInst_Y ;
    wire stateArray_S30reg_gff_1_SFF_7_MUXInst_X ;
    wire stateArray_S31reg_gff_1_SFF_0_MUXInst_Y ;
    wire stateArray_S31reg_gff_1_SFF_0_MUXInst_X ;
    wire stateArray_S31reg_gff_1_SFF_1_MUXInst_Y ;
    wire stateArray_S31reg_gff_1_SFF_1_MUXInst_X ;
    wire stateArray_S31reg_gff_1_SFF_2_MUXInst_Y ;
    wire stateArray_S31reg_gff_1_SFF_2_MUXInst_X ;
    wire stateArray_S31reg_gff_1_SFF_3_MUXInst_Y ;
    wire stateArray_S31reg_gff_1_SFF_3_MUXInst_X ;
    wire stateArray_S31reg_gff_1_SFF_4_MUXInst_Y ;
    wire stateArray_S31reg_gff_1_SFF_4_MUXInst_X ;
    wire stateArray_S31reg_gff_1_SFF_5_MUXInst_Y ;
    wire stateArray_S31reg_gff_1_SFF_5_MUXInst_X ;
    wire stateArray_S31reg_gff_1_SFF_6_MUXInst_Y ;
    wire stateArray_S31reg_gff_1_SFF_6_MUXInst_X ;
    wire stateArray_S31reg_gff_1_SFF_7_MUXInst_Y ;
    wire stateArray_S31reg_gff_1_SFF_7_MUXInst_X ;
    wire stateArray_S32reg_gff_1_SFF_0_MUXInst_Y ;
    wire stateArray_S32reg_gff_1_SFF_0_MUXInst_X ;
    wire stateArray_S32reg_gff_1_SFF_1_MUXInst_Y ;
    wire stateArray_S32reg_gff_1_SFF_1_MUXInst_X ;
    wire stateArray_S32reg_gff_1_SFF_2_MUXInst_Y ;
    wire stateArray_S32reg_gff_1_SFF_2_MUXInst_X ;
    wire stateArray_S32reg_gff_1_SFF_3_MUXInst_Y ;
    wire stateArray_S32reg_gff_1_SFF_3_MUXInst_X ;
    wire stateArray_S32reg_gff_1_SFF_4_MUXInst_Y ;
    wire stateArray_S32reg_gff_1_SFF_4_MUXInst_X ;
    wire stateArray_S32reg_gff_1_SFF_5_MUXInst_Y ;
    wire stateArray_S32reg_gff_1_SFF_5_MUXInst_X ;
    wire stateArray_S32reg_gff_1_SFF_6_MUXInst_Y ;
    wire stateArray_S32reg_gff_1_SFF_6_MUXInst_X ;
    wire stateArray_S32reg_gff_1_SFF_7_MUXInst_Y ;
    wire stateArray_S32reg_gff_1_SFF_7_MUXInst_X ;
    wire stateArray_S33reg_gff_1_SFF_0_MUXInst_Y ;
    wire stateArray_S33reg_gff_1_SFF_0_MUXInst_X ;
    wire stateArray_S33reg_gff_1_SFF_1_MUXInst_Y ;
    wire stateArray_S33reg_gff_1_SFF_1_MUXInst_X ;
    wire stateArray_S33reg_gff_1_SFF_2_MUXInst_Y ;
    wire stateArray_S33reg_gff_1_SFF_2_MUXInst_X ;
    wire stateArray_S33reg_gff_1_SFF_3_MUXInst_Y ;
    wire stateArray_S33reg_gff_1_SFF_3_MUXInst_X ;
    wire stateArray_S33reg_gff_1_SFF_4_MUXInst_Y ;
    wire stateArray_S33reg_gff_1_SFF_4_MUXInst_X ;
    wire stateArray_S33reg_gff_1_SFF_5_MUXInst_Y ;
    wire stateArray_S33reg_gff_1_SFF_5_MUXInst_X ;
    wire stateArray_S33reg_gff_1_SFF_6_MUXInst_Y ;
    wire stateArray_S33reg_gff_1_SFF_6_MUXInst_X ;
    wire stateArray_S33reg_gff_1_SFF_7_MUXInst_Y ;
    wire stateArray_S33reg_gff_1_SFF_7_MUXInst_X ;
    wire stateArray_MUX_inS03ser_mux_inst_0_Y ;
    wire stateArray_MUX_inS03ser_mux_inst_0_X ;
    wire stateArray_MUX_inS03ser_mux_inst_1_Y ;
    wire stateArray_MUX_inS03ser_mux_inst_1_X ;
    wire stateArray_MUX_inS03ser_mux_inst_2_Y ;
    wire stateArray_MUX_inS03ser_mux_inst_2_X ;
    wire stateArray_MUX_inS03ser_mux_inst_3_Y ;
    wire stateArray_MUX_inS03ser_mux_inst_3_X ;
    wire stateArray_MUX_inS03ser_mux_inst_4_Y ;
    wire stateArray_MUX_inS03ser_mux_inst_4_X ;
    wire stateArray_MUX_inS03ser_mux_inst_5_Y ;
    wire stateArray_MUX_inS03ser_mux_inst_5_X ;
    wire stateArray_MUX_inS03ser_mux_inst_6_Y ;
    wire stateArray_MUX_inS03ser_mux_inst_6_X ;
    wire stateArray_MUX_inS03ser_mux_inst_7_Y ;
    wire stateArray_MUX_inS03ser_mux_inst_7_X ;
    wire stateArray_MUX_inS13ser_mux_inst_0_Y ;
    wire stateArray_MUX_inS13ser_mux_inst_0_X ;
    wire stateArray_MUX_inS13ser_mux_inst_1_Y ;
    wire stateArray_MUX_inS13ser_mux_inst_1_X ;
    wire stateArray_MUX_inS13ser_mux_inst_2_Y ;
    wire stateArray_MUX_inS13ser_mux_inst_2_X ;
    wire stateArray_MUX_inS13ser_mux_inst_3_Y ;
    wire stateArray_MUX_inS13ser_mux_inst_3_X ;
    wire stateArray_MUX_inS13ser_mux_inst_4_Y ;
    wire stateArray_MUX_inS13ser_mux_inst_4_X ;
    wire stateArray_MUX_inS13ser_mux_inst_5_Y ;
    wire stateArray_MUX_inS13ser_mux_inst_5_X ;
    wire stateArray_MUX_inS13ser_mux_inst_6_Y ;
    wire stateArray_MUX_inS13ser_mux_inst_6_X ;
    wire stateArray_MUX_inS13ser_mux_inst_7_Y ;
    wire stateArray_MUX_inS13ser_mux_inst_7_X ;
    wire stateArray_MUX_inS23ser_mux_inst_0_Y ;
    wire stateArray_MUX_inS23ser_mux_inst_0_X ;
    wire stateArray_MUX_inS23ser_mux_inst_1_Y ;
    wire stateArray_MUX_inS23ser_mux_inst_1_X ;
    wire stateArray_MUX_inS23ser_mux_inst_2_Y ;
    wire stateArray_MUX_inS23ser_mux_inst_2_X ;
    wire stateArray_MUX_inS23ser_mux_inst_3_Y ;
    wire stateArray_MUX_inS23ser_mux_inst_3_X ;
    wire stateArray_MUX_inS23ser_mux_inst_4_Y ;
    wire stateArray_MUX_inS23ser_mux_inst_4_X ;
    wire stateArray_MUX_inS23ser_mux_inst_5_Y ;
    wire stateArray_MUX_inS23ser_mux_inst_5_X ;
    wire stateArray_MUX_inS23ser_mux_inst_6_Y ;
    wire stateArray_MUX_inS23ser_mux_inst_6_X ;
    wire stateArray_MUX_inS23ser_mux_inst_7_Y ;
    wire stateArray_MUX_inS23ser_mux_inst_7_X ;
    wire stateArray_MUX_input_MC_mux_inst_0_Y ;
    wire stateArray_MUX_input_MC_mux_inst_0_X ;
    wire stateArray_MUX_input_MC_mux_inst_1_Y ;
    wire stateArray_MUX_input_MC_mux_inst_1_X ;
    wire stateArray_MUX_input_MC_mux_inst_2_Y ;
    wire stateArray_MUX_input_MC_mux_inst_2_X ;
    wire stateArray_MUX_input_MC_mux_inst_3_Y ;
    wire stateArray_MUX_input_MC_mux_inst_3_X ;
    wire stateArray_MUX_input_MC_mux_inst_4_Y ;
    wire stateArray_MUX_input_MC_mux_inst_4_X ;
    wire stateArray_MUX_input_MC_mux_inst_5_Y ;
    wire stateArray_MUX_input_MC_mux_inst_5_X ;
    wire stateArray_MUX_input_MC_mux_inst_6_Y ;
    wire stateArray_MUX_input_MC_mux_inst_6_X ;
    wire stateArray_MUX_input_MC_mux_inst_7_Y ;
    wire stateArray_MUX_input_MC_mux_inst_7_X ;
    wire stateArray_MUX_inS33ser_mux_inst_0_Y ;
    wire stateArray_MUX_inS33ser_mux_inst_0_X ;
    wire stateArray_MUX_inS33ser_mux_inst_1_Y ;
    wire stateArray_MUX_inS33ser_mux_inst_1_X ;
    wire stateArray_MUX_inS33ser_mux_inst_2_Y ;
    wire stateArray_MUX_inS33ser_mux_inst_2_X ;
    wire stateArray_MUX_inS33ser_mux_inst_3_Y ;
    wire stateArray_MUX_inS33ser_mux_inst_3_X ;
    wire stateArray_MUX_inS33ser_mux_inst_4_Y ;
    wire stateArray_MUX_inS33ser_mux_inst_4_X ;
    wire stateArray_MUX_inS33ser_mux_inst_5_Y ;
    wire stateArray_MUX_inS33ser_mux_inst_5_X ;
    wire stateArray_MUX_inS33ser_mux_inst_6_Y ;
    wire stateArray_MUX_inS33ser_mux_inst_6_X ;
    wire stateArray_MUX_inS33ser_mux_inst_7_Y ;
    wire stateArray_MUX_inS33ser_mux_inst_7_X ;
    wire MUX_StateInMC_mux_inst_0_Y ;
    wire MUX_StateInMC_mux_inst_0_X ;
    wire MUX_StateInMC_mux_inst_1_Y ;
    wire MUX_StateInMC_mux_inst_1_X ;
    wire MUX_StateInMC_mux_inst_2_Y ;
    wire MUX_StateInMC_mux_inst_2_X ;
    wire MUX_StateInMC_mux_inst_3_Y ;
    wire MUX_StateInMC_mux_inst_3_X ;
    wire MUX_StateInMC_mux_inst_4_Y ;
    wire MUX_StateInMC_mux_inst_4_X ;
    wire MUX_StateInMC_mux_inst_5_Y ;
    wire MUX_StateInMC_mux_inst_5_X ;
    wire MUX_StateInMC_mux_inst_6_Y ;
    wire MUX_StateInMC_mux_inst_6_X ;
    wire MUX_StateInMC_mux_inst_7_Y ;
    wire MUX_StateInMC_mux_inst_7_X ;
    wire MUX_StateInMC_mux_inst_8_Y ;
    wire MUX_StateInMC_mux_inst_8_X ;
    wire MUX_StateInMC_mux_inst_9_Y ;
    wire MUX_StateInMC_mux_inst_9_X ;
    wire MUX_StateInMC_mux_inst_10_Y ;
    wire MUX_StateInMC_mux_inst_10_X ;
    wire MUX_StateInMC_mux_inst_11_Y ;
    wire MUX_StateInMC_mux_inst_11_X ;
    wire MUX_StateInMC_mux_inst_12_Y ;
    wire MUX_StateInMC_mux_inst_12_X ;
    wire MUX_StateInMC_mux_inst_13_Y ;
    wire MUX_StateInMC_mux_inst_13_X ;
    wire MUX_StateInMC_mux_inst_14_Y ;
    wire MUX_StateInMC_mux_inst_14_X ;
    wire MUX_StateInMC_mux_inst_15_Y ;
    wire MUX_StateInMC_mux_inst_15_X ;
    wire MUX_StateInMC_mux_inst_16_Y ;
    wire MUX_StateInMC_mux_inst_16_X ;
    wire MUX_StateInMC_mux_inst_17_Y ;
    wire MUX_StateInMC_mux_inst_17_X ;
    wire MUX_StateInMC_mux_inst_18_Y ;
    wire MUX_StateInMC_mux_inst_18_X ;
    wire MUX_StateInMC_mux_inst_19_Y ;
    wire MUX_StateInMC_mux_inst_19_X ;
    wire MUX_StateInMC_mux_inst_20_Y ;
    wire MUX_StateInMC_mux_inst_20_X ;
    wire MUX_StateInMC_mux_inst_21_Y ;
    wire MUX_StateInMC_mux_inst_21_X ;
    wire MUX_StateInMC_mux_inst_22_Y ;
    wire MUX_StateInMC_mux_inst_22_X ;
    wire MUX_StateInMC_mux_inst_23_Y ;
    wire MUX_StateInMC_mux_inst_23_X ;
    wire MUX_StateInMC_mux_inst_24_Y ;
    wire MUX_StateInMC_mux_inst_24_X ;
    wire MUX_StateInMC_mux_inst_25_Y ;
    wire MUX_StateInMC_mux_inst_25_X ;
    wire MUX_StateInMC_mux_inst_26_Y ;
    wire MUX_StateInMC_mux_inst_26_X ;
    wire MUX_StateInMC_mux_inst_27_Y ;
    wire MUX_StateInMC_mux_inst_27_X ;
    wire MUX_StateInMC_mux_inst_28_Y ;
    wire MUX_StateInMC_mux_inst_28_X ;
    wire MUX_StateInMC_mux_inst_29_Y ;
    wire MUX_StateInMC_mux_inst_29_X ;
    wire MUX_StateInMC_mux_inst_30_Y ;
    wire MUX_StateInMC_mux_inst_30_X ;
    wire MUX_StateInMC_mux_inst_31_Y ;
    wire MUX_StateInMC_mux_inst_31_X ;
    wire KeyArray_n32 ;
    wire KeyArray_n31 ;
    wire KeyArray_n30 ;
    wire KeyArray_n29 ;
    wire KeyArray_n28 ;
    wire KeyArray_n27 ;
    wire KeyArray_n26 ;
    wire KeyArray_n25 ;
    wire KeyArray_nReset_selXOR ;
    wire KeyArray_outS01ser_0_ ;
    wire KeyArray_outS01ser_1_ ;
    wire KeyArray_outS01ser_2_ ;
    wire KeyArray_outS01ser_3_ ;
    wire KeyArray_outS01ser_4_ ;
    wire KeyArray_outS01ser_5_ ;
    wire KeyArray_outS01ser_6_ ;
    wire KeyArray_outS01ser_7_ ;
    wire KeyArray_S00reg_gff_1_SFF_0_n2 ;
    wire KeyArray_S00reg_gff_1_SFF_0_n1 ;
    wire KeyArray_S00reg_gff_1_SFF_0_QD ;
    wire KeyArray_S00reg_gff_1_SFF_0_MUXInst_Y ;
    wire KeyArray_S00reg_gff_1_SFF_0_MUXInst_X ;
    wire KeyArray_S00reg_gff_1_SFF_1_n2 ;
    wire KeyArray_S00reg_gff_1_SFF_1_n1 ;
    wire KeyArray_S00reg_gff_1_SFF_1_QD ;
    wire KeyArray_S00reg_gff_1_SFF_1_MUXInst_Y ;
    wire KeyArray_S00reg_gff_1_SFF_1_MUXInst_X ;
    wire KeyArray_S00reg_gff_1_SFF_2_n2 ;
    wire KeyArray_S00reg_gff_1_SFF_2_n1 ;
    wire KeyArray_S00reg_gff_1_SFF_2_QD ;
    wire KeyArray_S00reg_gff_1_SFF_2_MUXInst_Y ;
    wire KeyArray_S00reg_gff_1_SFF_2_MUXInst_X ;
    wire KeyArray_S00reg_gff_1_SFF_3_n2 ;
    wire KeyArray_S00reg_gff_1_SFF_3_n1 ;
    wire KeyArray_S00reg_gff_1_SFF_3_QD ;
    wire KeyArray_S00reg_gff_1_SFF_3_MUXInst_Y ;
    wire KeyArray_S00reg_gff_1_SFF_3_MUXInst_X ;
    wire KeyArray_S00reg_gff_1_SFF_4_n2 ;
    wire KeyArray_S00reg_gff_1_SFF_4_n1 ;
    wire KeyArray_S00reg_gff_1_SFF_4_QD ;
    wire KeyArray_S00reg_gff_1_SFF_4_MUXInst_Y ;
    wire KeyArray_S00reg_gff_1_SFF_4_MUXInst_X ;
    wire KeyArray_S00reg_gff_1_SFF_5_n2 ;
    wire KeyArray_S00reg_gff_1_SFF_5_n1 ;
    wire KeyArray_S00reg_gff_1_SFF_5_QD ;
    wire KeyArray_S00reg_gff_1_SFF_5_MUXInst_Y ;
    wire KeyArray_S00reg_gff_1_SFF_5_MUXInst_X ;
    wire KeyArray_S00reg_gff_1_SFF_6_n2 ;
    wire KeyArray_S00reg_gff_1_SFF_6_n1 ;
    wire KeyArray_S00reg_gff_1_SFF_6_QD ;
    wire KeyArray_S00reg_gff_1_SFF_6_MUXInst_Y ;
    wire KeyArray_S00reg_gff_1_SFF_6_MUXInst_X ;
    wire KeyArray_S00reg_gff_1_SFF_7_n2 ;
    wire KeyArray_S00reg_gff_1_SFF_7_n1 ;
    wire KeyArray_S00reg_gff_1_SFF_7_QD ;
    wire KeyArray_S00reg_gff_1_SFF_7_MUXInst_Y ;
    wire KeyArray_S00reg_gff_1_SFF_7_MUXInst_X ;
    wire KeyArray_S01reg_gff_1_SFF_0_n2 ;
    wire KeyArray_S01reg_gff_1_SFF_0_n1 ;
    wire KeyArray_S01reg_gff_1_SFF_0_QD ;
    wire KeyArray_S01reg_gff_1_SFF_0_MUXInst_Y ;
    wire KeyArray_S01reg_gff_1_SFF_0_MUXInst_X ;
    wire KeyArray_S01reg_gff_1_SFF_1_n2 ;
    wire KeyArray_S01reg_gff_1_SFF_1_n1 ;
    wire KeyArray_S01reg_gff_1_SFF_1_QD ;
    wire KeyArray_S01reg_gff_1_SFF_1_MUXInst_Y ;
    wire KeyArray_S01reg_gff_1_SFF_1_MUXInst_X ;
    wire KeyArray_S01reg_gff_1_SFF_2_n2 ;
    wire KeyArray_S01reg_gff_1_SFF_2_n1 ;
    wire KeyArray_S01reg_gff_1_SFF_2_QD ;
    wire KeyArray_S01reg_gff_1_SFF_2_MUXInst_Y ;
    wire KeyArray_S01reg_gff_1_SFF_2_MUXInst_X ;
    wire KeyArray_S01reg_gff_1_SFF_3_n2 ;
    wire KeyArray_S01reg_gff_1_SFF_3_n1 ;
    wire KeyArray_S01reg_gff_1_SFF_3_QD ;
    wire KeyArray_S01reg_gff_1_SFF_3_MUXInst_Y ;
    wire KeyArray_S01reg_gff_1_SFF_3_MUXInst_X ;
    wire KeyArray_S01reg_gff_1_SFF_4_n2 ;
    wire KeyArray_S01reg_gff_1_SFF_4_n1 ;
    wire KeyArray_S01reg_gff_1_SFF_4_QD ;
    wire KeyArray_S01reg_gff_1_SFF_4_MUXInst_Y ;
    wire KeyArray_S01reg_gff_1_SFF_4_MUXInst_X ;
    wire KeyArray_S01reg_gff_1_SFF_5_n2 ;
    wire KeyArray_S01reg_gff_1_SFF_5_n1 ;
    wire KeyArray_S01reg_gff_1_SFF_5_QD ;
    wire KeyArray_S01reg_gff_1_SFF_5_MUXInst_Y ;
    wire KeyArray_S01reg_gff_1_SFF_5_MUXInst_X ;
    wire KeyArray_S01reg_gff_1_SFF_6_n2 ;
    wire KeyArray_S01reg_gff_1_SFF_6_n1 ;
    wire KeyArray_S01reg_gff_1_SFF_6_QD ;
    wire KeyArray_S01reg_gff_1_SFF_6_MUXInst_Y ;
    wire KeyArray_S01reg_gff_1_SFF_6_MUXInst_X ;
    wire KeyArray_S01reg_gff_1_SFF_7_n2 ;
    wire KeyArray_S01reg_gff_1_SFF_7_n1 ;
    wire KeyArray_S01reg_gff_1_SFF_7_QD ;
    wire KeyArray_S01reg_gff_1_SFF_7_MUXInst_Y ;
    wire KeyArray_S01reg_gff_1_SFF_7_MUXInst_X ;
    wire KeyArray_S02reg_gff_1_SFF_0_n2 ;
    wire KeyArray_S02reg_gff_1_SFF_0_n1 ;
    wire KeyArray_S02reg_gff_1_SFF_0_QD ;
    wire KeyArray_S02reg_gff_1_SFF_0_MUXInst_Y ;
    wire KeyArray_S02reg_gff_1_SFF_0_MUXInst_X ;
    wire KeyArray_S02reg_gff_1_SFF_1_n2 ;
    wire KeyArray_S02reg_gff_1_SFF_1_n1 ;
    wire KeyArray_S02reg_gff_1_SFF_1_QD ;
    wire KeyArray_S02reg_gff_1_SFF_1_MUXInst_Y ;
    wire KeyArray_S02reg_gff_1_SFF_1_MUXInst_X ;
    wire KeyArray_S02reg_gff_1_SFF_2_n2 ;
    wire KeyArray_S02reg_gff_1_SFF_2_n1 ;
    wire KeyArray_S02reg_gff_1_SFF_2_QD ;
    wire KeyArray_S02reg_gff_1_SFF_2_MUXInst_Y ;
    wire KeyArray_S02reg_gff_1_SFF_2_MUXInst_X ;
    wire KeyArray_S02reg_gff_1_SFF_3_n2 ;
    wire KeyArray_S02reg_gff_1_SFF_3_n1 ;
    wire KeyArray_S02reg_gff_1_SFF_3_QD ;
    wire KeyArray_S02reg_gff_1_SFF_3_MUXInst_Y ;
    wire KeyArray_S02reg_gff_1_SFF_3_MUXInst_X ;
    wire KeyArray_S02reg_gff_1_SFF_4_n2 ;
    wire KeyArray_S02reg_gff_1_SFF_4_n1 ;
    wire KeyArray_S02reg_gff_1_SFF_4_QD ;
    wire KeyArray_S02reg_gff_1_SFF_4_MUXInst_Y ;
    wire KeyArray_S02reg_gff_1_SFF_4_MUXInst_X ;
    wire KeyArray_S02reg_gff_1_SFF_5_n2 ;
    wire KeyArray_S02reg_gff_1_SFF_5_n1 ;
    wire KeyArray_S02reg_gff_1_SFF_5_QD ;
    wire KeyArray_S02reg_gff_1_SFF_5_MUXInst_Y ;
    wire KeyArray_S02reg_gff_1_SFF_5_MUXInst_X ;
    wire KeyArray_S02reg_gff_1_SFF_6_n2 ;
    wire KeyArray_S02reg_gff_1_SFF_6_n1 ;
    wire KeyArray_S02reg_gff_1_SFF_6_QD ;
    wire KeyArray_S02reg_gff_1_SFF_6_MUXInst_Y ;
    wire KeyArray_S02reg_gff_1_SFF_6_MUXInst_X ;
    wire KeyArray_S02reg_gff_1_SFF_7_n2 ;
    wire KeyArray_S02reg_gff_1_SFF_7_n1 ;
    wire KeyArray_S02reg_gff_1_SFF_7_QD ;
    wire KeyArray_S02reg_gff_1_SFF_7_MUXInst_Y ;
    wire KeyArray_S02reg_gff_1_SFF_7_MUXInst_X ;
    wire KeyArray_S03reg_gff_1_SFF_0_n2 ;
    wire KeyArray_S03reg_gff_1_SFF_0_n1 ;
    wire KeyArray_S03reg_gff_1_SFF_0_QD ;
    wire KeyArray_S03reg_gff_1_SFF_0_MUXInst_Y ;
    wire KeyArray_S03reg_gff_1_SFF_0_MUXInst_X ;
    wire KeyArray_S03reg_gff_1_SFF_1_n2 ;
    wire KeyArray_S03reg_gff_1_SFF_1_n1 ;
    wire KeyArray_S03reg_gff_1_SFF_1_QD ;
    wire KeyArray_S03reg_gff_1_SFF_1_MUXInst_Y ;
    wire KeyArray_S03reg_gff_1_SFF_1_MUXInst_X ;
    wire KeyArray_S03reg_gff_1_SFF_2_n2 ;
    wire KeyArray_S03reg_gff_1_SFF_2_n1 ;
    wire KeyArray_S03reg_gff_1_SFF_2_QD ;
    wire KeyArray_S03reg_gff_1_SFF_2_MUXInst_Y ;
    wire KeyArray_S03reg_gff_1_SFF_2_MUXInst_X ;
    wire KeyArray_S03reg_gff_1_SFF_3_n2 ;
    wire KeyArray_S03reg_gff_1_SFF_3_n1 ;
    wire KeyArray_S03reg_gff_1_SFF_3_QD ;
    wire KeyArray_S03reg_gff_1_SFF_3_MUXInst_Y ;
    wire KeyArray_S03reg_gff_1_SFF_3_MUXInst_X ;
    wire KeyArray_S03reg_gff_1_SFF_4_n2 ;
    wire KeyArray_S03reg_gff_1_SFF_4_n1 ;
    wire KeyArray_S03reg_gff_1_SFF_4_QD ;
    wire KeyArray_S03reg_gff_1_SFF_4_MUXInst_Y ;
    wire KeyArray_S03reg_gff_1_SFF_4_MUXInst_X ;
    wire KeyArray_S03reg_gff_1_SFF_5_n2 ;
    wire KeyArray_S03reg_gff_1_SFF_5_n1 ;
    wire KeyArray_S03reg_gff_1_SFF_5_QD ;
    wire KeyArray_S03reg_gff_1_SFF_5_MUXInst_Y ;
    wire KeyArray_S03reg_gff_1_SFF_5_MUXInst_X ;
    wire KeyArray_S03reg_gff_1_SFF_6_n2 ;
    wire KeyArray_S03reg_gff_1_SFF_6_n1 ;
    wire KeyArray_S03reg_gff_1_SFF_6_QD ;
    wire KeyArray_S03reg_gff_1_SFF_6_MUXInst_Y ;
    wire KeyArray_S03reg_gff_1_SFF_6_MUXInst_X ;
    wire KeyArray_S03reg_gff_1_SFF_7_n2 ;
    wire KeyArray_S03reg_gff_1_SFF_7_n1 ;
    wire KeyArray_S03reg_gff_1_SFF_7_QD ;
    wire KeyArray_S03reg_gff_1_SFF_7_MUXInst_Y ;
    wire KeyArray_S03reg_gff_1_SFF_7_MUXInst_X ;
    wire KeyArray_S10reg_gff_1_SFF_0_n2 ;
    wire KeyArray_S10reg_gff_1_SFF_0_n1 ;
    wire KeyArray_S10reg_gff_1_SFF_0_QD ;
    wire KeyArray_S10reg_gff_1_SFF_0_MUXInst_Y ;
    wire KeyArray_S10reg_gff_1_SFF_0_MUXInst_X ;
    wire KeyArray_S10reg_gff_1_SFF_1_n2 ;
    wire KeyArray_S10reg_gff_1_SFF_1_n1 ;
    wire KeyArray_S10reg_gff_1_SFF_1_QD ;
    wire KeyArray_S10reg_gff_1_SFF_1_MUXInst_Y ;
    wire KeyArray_S10reg_gff_1_SFF_1_MUXInst_X ;
    wire KeyArray_S10reg_gff_1_SFF_2_n2 ;
    wire KeyArray_S10reg_gff_1_SFF_2_n1 ;
    wire KeyArray_S10reg_gff_1_SFF_2_QD ;
    wire KeyArray_S10reg_gff_1_SFF_2_MUXInst_Y ;
    wire KeyArray_S10reg_gff_1_SFF_2_MUXInst_X ;
    wire KeyArray_S10reg_gff_1_SFF_3_n2 ;
    wire KeyArray_S10reg_gff_1_SFF_3_n1 ;
    wire KeyArray_S10reg_gff_1_SFF_3_QD ;
    wire KeyArray_S10reg_gff_1_SFF_3_MUXInst_Y ;
    wire KeyArray_S10reg_gff_1_SFF_3_MUXInst_X ;
    wire KeyArray_S10reg_gff_1_SFF_4_n2 ;
    wire KeyArray_S10reg_gff_1_SFF_4_n1 ;
    wire KeyArray_S10reg_gff_1_SFF_4_QD ;
    wire KeyArray_S10reg_gff_1_SFF_4_MUXInst_Y ;
    wire KeyArray_S10reg_gff_1_SFF_4_MUXInst_X ;
    wire KeyArray_S10reg_gff_1_SFF_5_n2 ;
    wire KeyArray_S10reg_gff_1_SFF_5_n1 ;
    wire KeyArray_S10reg_gff_1_SFF_5_QD ;
    wire KeyArray_S10reg_gff_1_SFF_5_MUXInst_Y ;
    wire KeyArray_S10reg_gff_1_SFF_5_MUXInst_X ;
    wire KeyArray_S10reg_gff_1_SFF_6_n2 ;
    wire KeyArray_S10reg_gff_1_SFF_6_n1 ;
    wire KeyArray_S10reg_gff_1_SFF_6_QD ;
    wire KeyArray_S10reg_gff_1_SFF_6_MUXInst_Y ;
    wire KeyArray_S10reg_gff_1_SFF_6_MUXInst_X ;
    wire KeyArray_S10reg_gff_1_SFF_7_n2 ;
    wire KeyArray_S10reg_gff_1_SFF_7_n1 ;
    wire KeyArray_S10reg_gff_1_SFF_7_QD ;
    wire KeyArray_S10reg_gff_1_SFF_7_MUXInst_Y ;
    wire KeyArray_S10reg_gff_1_SFF_7_MUXInst_X ;
    wire KeyArray_S11reg_gff_1_SFF_0_n2 ;
    wire KeyArray_S11reg_gff_1_SFF_0_n1 ;
    wire KeyArray_S11reg_gff_1_SFF_0_QD ;
    wire KeyArray_S11reg_gff_1_SFF_0_MUXInst_Y ;
    wire KeyArray_S11reg_gff_1_SFF_0_MUXInst_X ;
    wire KeyArray_S11reg_gff_1_SFF_1_n2 ;
    wire KeyArray_S11reg_gff_1_SFF_1_n1 ;
    wire KeyArray_S11reg_gff_1_SFF_1_QD ;
    wire KeyArray_S11reg_gff_1_SFF_1_MUXInst_Y ;
    wire KeyArray_S11reg_gff_1_SFF_1_MUXInst_X ;
    wire KeyArray_S11reg_gff_1_SFF_2_n2 ;
    wire KeyArray_S11reg_gff_1_SFF_2_n1 ;
    wire KeyArray_S11reg_gff_1_SFF_2_QD ;
    wire KeyArray_S11reg_gff_1_SFF_2_MUXInst_Y ;
    wire KeyArray_S11reg_gff_1_SFF_2_MUXInst_X ;
    wire KeyArray_S11reg_gff_1_SFF_3_n2 ;
    wire KeyArray_S11reg_gff_1_SFF_3_n1 ;
    wire KeyArray_S11reg_gff_1_SFF_3_QD ;
    wire KeyArray_S11reg_gff_1_SFF_3_MUXInst_Y ;
    wire KeyArray_S11reg_gff_1_SFF_3_MUXInst_X ;
    wire KeyArray_S11reg_gff_1_SFF_4_n2 ;
    wire KeyArray_S11reg_gff_1_SFF_4_n1 ;
    wire KeyArray_S11reg_gff_1_SFF_4_QD ;
    wire KeyArray_S11reg_gff_1_SFF_4_MUXInst_Y ;
    wire KeyArray_S11reg_gff_1_SFF_4_MUXInst_X ;
    wire KeyArray_S11reg_gff_1_SFF_5_n2 ;
    wire KeyArray_S11reg_gff_1_SFF_5_n1 ;
    wire KeyArray_S11reg_gff_1_SFF_5_QD ;
    wire KeyArray_S11reg_gff_1_SFF_5_MUXInst_Y ;
    wire KeyArray_S11reg_gff_1_SFF_5_MUXInst_X ;
    wire KeyArray_S11reg_gff_1_SFF_6_n2 ;
    wire KeyArray_S11reg_gff_1_SFF_6_n1 ;
    wire KeyArray_S11reg_gff_1_SFF_6_QD ;
    wire KeyArray_S11reg_gff_1_SFF_6_MUXInst_Y ;
    wire KeyArray_S11reg_gff_1_SFF_6_MUXInst_X ;
    wire KeyArray_S11reg_gff_1_SFF_7_n2 ;
    wire KeyArray_S11reg_gff_1_SFF_7_n1 ;
    wire KeyArray_S11reg_gff_1_SFF_7_QD ;
    wire KeyArray_S11reg_gff_1_SFF_7_MUXInst_Y ;
    wire KeyArray_S11reg_gff_1_SFF_7_MUXInst_X ;
    wire KeyArray_S12reg_gff_1_SFF_0_n2 ;
    wire KeyArray_S12reg_gff_1_SFF_0_n1 ;
    wire KeyArray_S12reg_gff_1_SFF_0_QD ;
    wire KeyArray_S12reg_gff_1_SFF_0_MUXInst_Y ;
    wire KeyArray_S12reg_gff_1_SFF_0_MUXInst_X ;
    wire KeyArray_S12reg_gff_1_SFF_1_n2 ;
    wire KeyArray_S12reg_gff_1_SFF_1_n1 ;
    wire KeyArray_S12reg_gff_1_SFF_1_QD ;
    wire KeyArray_S12reg_gff_1_SFF_1_MUXInst_Y ;
    wire KeyArray_S12reg_gff_1_SFF_1_MUXInst_X ;
    wire KeyArray_S12reg_gff_1_SFF_2_n2 ;
    wire KeyArray_S12reg_gff_1_SFF_2_n1 ;
    wire KeyArray_S12reg_gff_1_SFF_2_QD ;
    wire KeyArray_S12reg_gff_1_SFF_2_MUXInst_Y ;
    wire KeyArray_S12reg_gff_1_SFF_2_MUXInst_X ;
    wire KeyArray_S12reg_gff_1_SFF_3_n2 ;
    wire KeyArray_S12reg_gff_1_SFF_3_n1 ;
    wire KeyArray_S12reg_gff_1_SFF_3_QD ;
    wire KeyArray_S12reg_gff_1_SFF_3_MUXInst_Y ;
    wire KeyArray_S12reg_gff_1_SFF_3_MUXInst_X ;
    wire KeyArray_S12reg_gff_1_SFF_4_n2 ;
    wire KeyArray_S12reg_gff_1_SFF_4_n1 ;
    wire KeyArray_S12reg_gff_1_SFF_4_QD ;
    wire KeyArray_S12reg_gff_1_SFF_4_MUXInst_Y ;
    wire KeyArray_S12reg_gff_1_SFF_4_MUXInst_X ;
    wire KeyArray_S12reg_gff_1_SFF_5_n2 ;
    wire KeyArray_S12reg_gff_1_SFF_5_n1 ;
    wire KeyArray_S12reg_gff_1_SFF_5_QD ;
    wire KeyArray_S12reg_gff_1_SFF_5_MUXInst_Y ;
    wire KeyArray_S12reg_gff_1_SFF_5_MUXInst_X ;
    wire KeyArray_S12reg_gff_1_SFF_6_n2 ;
    wire KeyArray_S12reg_gff_1_SFF_6_n1 ;
    wire KeyArray_S12reg_gff_1_SFF_6_QD ;
    wire KeyArray_S12reg_gff_1_SFF_6_MUXInst_Y ;
    wire KeyArray_S12reg_gff_1_SFF_6_MUXInst_X ;
    wire KeyArray_S12reg_gff_1_SFF_7_n2 ;
    wire KeyArray_S12reg_gff_1_SFF_7_n1 ;
    wire KeyArray_S12reg_gff_1_SFF_7_QD ;
    wire KeyArray_S12reg_gff_1_SFF_7_MUXInst_Y ;
    wire KeyArray_S12reg_gff_1_SFF_7_MUXInst_X ;
    wire KeyArray_S13reg_gff_1_SFF_0_n2 ;
    wire KeyArray_S13reg_gff_1_SFF_0_n1 ;
    wire KeyArray_S13reg_gff_1_SFF_0_QD ;
    wire KeyArray_S13reg_gff_1_SFF_0_MUXInst_Y ;
    wire KeyArray_S13reg_gff_1_SFF_0_MUXInst_X ;
    wire KeyArray_S13reg_gff_1_SFF_1_n2 ;
    wire KeyArray_S13reg_gff_1_SFF_1_n1 ;
    wire KeyArray_S13reg_gff_1_SFF_1_QD ;
    wire KeyArray_S13reg_gff_1_SFF_1_MUXInst_Y ;
    wire KeyArray_S13reg_gff_1_SFF_1_MUXInst_X ;
    wire KeyArray_S13reg_gff_1_SFF_2_n2 ;
    wire KeyArray_S13reg_gff_1_SFF_2_n1 ;
    wire KeyArray_S13reg_gff_1_SFF_2_QD ;
    wire KeyArray_S13reg_gff_1_SFF_2_MUXInst_Y ;
    wire KeyArray_S13reg_gff_1_SFF_2_MUXInst_X ;
    wire KeyArray_S13reg_gff_1_SFF_3_n2 ;
    wire KeyArray_S13reg_gff_1_SFF_3_n1 ;
    wire KeyArray_S13reg_gff_1_SFF_3_QD ;
    wire KeyArray_S13reg_gff_1_SFF_3_MUXInst_Y ;
    wire KeyArray_S13reg_gff_1_SFF_3_MUXInst_X ;
    wire KeyArray_S13reg_gff_1_SFF_4_n2 ;
    wire KeyArray_S13reg_gff_1_SFF_4_n1 ;
    wire KeyArray_S13reg_gff_1_SFF_4_QD ;
    wire KeyArray_S13reg_gff_1_SFF_4_MUXInst_Y ;
    wire KeyArray_S13reg_gff_1_SFF_4_MUXInst_X ;
    wire KeyArray_S13reg_gff_1_SFF_5_n2 ;
    wire KeyArray_S13reg_gff_1_SFF_5_n1 ;
    wire KeyArray_S13reg_gff_1_SFF_5_QD ;
    wire KeyArray_S13reg_gff_1_SFF_5_MUXInst_Y ;
    wire KeyArray_S13reg_gff_1_SFF_5_MUXInst_X ;
    wire KeyArray_S13reg_gff_1_SFF_6_n2 ;
    wire KeyArray_S13reg_gff_1_SFF_6_n1 ;
    wire KeyArray_S13reg_gff_1_SFF_6_QD ;
    wire KeyArray_S13reg_gff_1_SFF_6_MUXInst_Y ;
    wire KeyArray_S13reg_gff_1_SFF_6_MUXInst_X ;
    wire KeyArray_S13reg_gff_1_SFF_7_n2 ;
    wire KeyArray_S13reg_gff_1_SFF_7_n1 ;
    wire KeyArray_S13reg_gff_1_SFF_7_QD ;
    wire KeyArray_S13reg_gff_1_SFF_7_MUXInst_Y ;
    wire KeyArray_S13reg_gff_1_SFF_7_MUXInst_X ;
    wire KeyArray_S20reg_gff_1_SFF_0_n2 ;
    wire KeyArray_S20reg_gff_1_SFF_0_n1 ;
    wire KeyArray_S20reg_gff_1_SFF_0_QD ;
    wire KeyArray_S20reg_gff_1_SFF_0_MUXInst_Y ;
    wire KeyArray_S20reg_gff_1_SFF_0_MUXInst_X ;
    wire KeyArray_S20reg_gff_1_SFF_1_n2 ;
    wire KeyArray_S20reg_gff_1_SFF_1_n1 ;
    wire KeyArray_S20reg_gff_1_SFF_1_QD ;
    wire KeyArray_S20reg_gff_1_SFF_1_MUXInst_Y ;
    wire KeyArray_S20reg_gff_1_SFF_1_MUXInst_X ;
    wire KeyArray_S20reg_gff_1_SFF_2_n2 ;
    wire KeyArray_S20reg_gff_1_SFF_2_n1 ;
    wire KeyArray_S20reg_gff_1_SFF_2_QD ;
    wire KeyArray_S20reg_gff_1_SFF_2_MUXInst_Y ;
    wire KeyArray_S20reg_gff_1_SFF_2_MUXInst_X ;
    wire KeyArray_S20reg_gff_1_SFF_3_n2 ;
    wire KeyArray_S20reg_gff_1_SFF_3_n1 ;
    wire KeyArray_S20reg_gff_1_SFF_3_QD ;
    wire KeyArray_S20reg_gff_1_SFF_3_MUXInst_Y ;
    wire KeyArray_S20reg_gff_1_SFF_3_MUXInst_X ;
    wire KeyArray_S20reg_gff_1_SFF_4_n2 ;
    wire KeyArray_S20reg_gff_1_SFF_4_n1 ;
    wire KeyArray_S20reg_gff_1_SFF_4_QD ;
    wire KeyArray_S20reg_gff_1_SFF_4_MUXInst_Y ;
    wire KeyArray_S20reg_gff_1_SFF_4_MUXInst_X ;
    wire KeyArray_S20reg_gff_1_SFF_5_n2 ;
    wire KeyArray_S20reg_gff_1_SFF_5_n1 ;
    wire KeyArray_S20reg_gff_1_SFF_5_QD ;
    wire KeyArray_S20reg_gff_1_SFF_5_MUXInst_Y ;
    wire KeyArray_S20reg_gff_1_SFF_5_MUXInst_X ;
    wire KeyArray_S20reg_gff_1_SFF_6_n2 ;
    wire KeyArray_S20reg_gff_1_SFF_6_n1 ;
    wire KeyArray_S20reg_gff_1_SFF_6_QD ;
    wire KeyArray_S20reg_gff_1_SFF_6_MUXInst_Y ;
    wire KeyArray_S20reg_gff_1_SFF_6_MUXInst_X ;
    wire KeyArray_S20reg_gff_1_SFF_7_n2 ;
    wire KeyArray_S20reg_gff_1_SFF_7_n1 ;
    wire KeyArray_S20reg_gff_1_SFF_7_QD ;
    wire KeyArray_S20reg_gff_1_SFF_7_MUXInst_Y ;
    wire KeyArray_S20reg_gff_1_SFF_7_MUXInst_X ;
    wire KeyArray_S21reg_gff_1_SFF_0_n2 ;
    wire KeyArray_S21reg_gff_1_SFF_0_n1 ;
    wire KeyArray_S21reg_gff_1_SFF_0_QD ;
    wire KeyArray_S21reg_gff_1_SFF_0_MUXInst_Y ;
    wire KeyArray_S21reg_gff_1_SFF_0_MUXInst_X ;
    wire KeyArray_S21reg_gff_1_SFF_1_n2 ;
    wire KeyArray_S21reg_gff_1_SFF_1_n1 ;
    wire KeyArray_S21reg_gff_1_SFF_1_QD ;
    wire KeyArray_S21reg_gff_1_SFF_1_MUXInst_Y ;
    wire KeyArray_S21reg_gff_1_SFF_1_MUXInst_X ;
    wire KeyArray_S21reg_gff_1_SFF_2_n2 ;
    wire KeyArray_S21reg_gff_1_SFF_2_n1 ;
    wire KeyArray_S21reg_gff_1_SFF_2_QD ;
    wire KeyArray_S21reg_gff_1_SFF_2_MUXInst_Y ;
    wire KeyArray_S21reg_gff_1_SFF_2_MUXInst_X ;
    wire KeyArray_S21reg_gff_1_SFF_3_n2 ;
    wire KeyArray_S21reg_gff_1_SFF_3_n1 ;
    wire KeyArray_S21reg_gff_1_SFF_3_QD ;
    wire KeyArray_S21reg_gff_1_SFF_3_MUXInst_Y ;
    wire KeyArray_S21reg_gff_1_SFF_3_MUXInst_X ;
    wire KeyArray_S21reg_gff_1_SFF_4_n2 ;
    wire KeyArray_S21reg_gff_1_SFF_4_n1 ;
    wire KeyArray_S21reg_gff_1_SFF_4_QD ;
    wire KeyArray_S21reg_gff_1_SFF_4_MUXInst_Y ;
    wire KeyArray_S21reg_gff_1_SFF_4_MUXInst_X ;
    wire KeyArray_S21reg_gff_1_SFF_5_n2 ;
    wire KeyArray_S21reg_gff_1_SFF_5_n1 ;
    wire KeyArray_S21reg_gff_1_SFF_5_QD ;
    wire KeyArray_S21reg_gff_1_SFF_5_MUXInst_Y ;
    wire KeyArray_S21reg_gff_1_SFF_5_MUXInst_X ;
    wire KeyArray_S21reg_gff_1_SFF_6_n2 ;
    wire KeyArray_S21reg_gff_1_SFF_6_n1 ;
    wire KeyArray_S21reg_gff_1_SFF_6_QD ;
    wire KeyArray_S21reg_gff_1_SFF_6_MUXInst_Y ;
    wire KeyArray_S21reg_gff_1_SFF_6_MUXInst_X ;
    wire KeyArray_S21reg_gff_1_SFF_7_n2 ;
    wire KeyArray_S21reg_gff_1_SFF_7_n1 ;
    wire KeyArray_S21reg_gff_1_SFF_7_QD ;
    wire KeyArray_S21reg_gff_1_SFF_7_MUXInst_Y ;
    wire KeyArray_S21reg_gff_1_SFF_7_MUXInst_X ;
    wire KeyArray_S22reg_gff_1_SFF_0_n2 ;
    wire KeyArray_S22reg_gff_1_SFF_0_n1 ;
    wire KeyArray_S22reg_gff_1_SFF_0_QD ;
    wire KeyArray_S22reg_gff_1_SFF_0_MUXInst_Y ;
    wire KeyArray_S22reg_gff_1_SFF_0_MUXInst_X ;
    wire KeyArray_S22reg_gff_1_SFF_1_n2 ;
    wire KeyArray_S22reg_gff_1_SFF_1_n1 ;
    wire KeyArray_S22reg_gff_1_SFF_1_QD ;
    wire KeyArray_S22reg_gff_1_SFF_1_MUXInst_Y ;
    wire KeyArray_S22reg_gff_1_SFF_1_MUXInst_X ;
    wire KeyArray_S22reg_gff_1_SFF_2_n2 ;
    wire KeyArray_S22reg_gff_1_SFF_2_n1 ;
    wire KeyArray_S22reg_gff_1_SFF_2_QD ;
    wire KeyArray_S22reg_gff_1_SFF_2_MUXInst_Y ;
    wire KeyArray_S22reg_gff_1_SFF_2_MUXInst_X ;
    wire KeyArray_S22reg_gff_1_SFF_3_n2 ;
    wire KeyArray_S22reg_gff_1_SFF_3_n1 ;
    wire KeyArray_S22reg_gff_1_SFF_3_QD ;
    wire KeyArray_S22reg_gff_1_SFF_3_MUXInst_Y ;
    wire KeyArray_S22reg_gff_1_SFF_3_MUXInst_X ;
    wire KeyArray_S22reg_gff_1_SFF_4_n2 ;
    wire KeyArray_S22reg_gff_1_SFF_4_n1 ;
    wire KeyArray_S22reg_gff_1_SFF_4_QD ;
    wire KeyArray_S22reg_gff_1_SFF_4_MUXInst_Y ;
    wire KeyArray_S22reg_gff_1_SFF_4_MUXInst_X ;
    wire KeyArray_S22reg_gff_1_SFF_5_n2 ;
    wire KeyArray_S22reg_gff_1_SFF_5_n1 ;
    wire KeyArray_S22reg_gff_1_SFF_5_QD ;
    wire KeyArray_S22reg_gff_1_SFF_5_MUXInst_Y ;
    wire KeyArray_S22reg_gff_1_SFF_5_MUXInst_X ;
    wire KeyArray_S22reg_gff_1_SFF_6_n2 ;
    wire KeyArray_S22reg_gff_1_SFF_6_n1 ;
    wire KeyArray_S22reg_gff_1_SFF_6_QD ;
    wire KeyArray_S22reg_gff_1_SFF_6_MUXInst_Y ;
    wire KeyArray_S22reg_gff_1_SFF_6_MUXInst_X ;
    wire KeyArray_S22reg_gff_1_SFF_7_n2 ;
    wire KeyArray_S22reg_gff_1_SFF_7_n1 ;
    wire KeyArray_S22reg_gff_1_SFF_7_QD ;
    wire KeyArray_S22reg_gff_1_SFF_7_MUXInst_Y ;
    wire KeyArray_S22reg_gff_1_SFF_7_MUXInst_X ;
    wire KeyArray_S23reg_gff_1_SFF_0_n2 ;
    wire KeyArray_S23reg_gff_1_SFF_0_n1 ;
    wire KeyArray_S23reg_gff_1_SFF_0_QD ;
    wire KeyArray_S23reg_gff_1_SFF_0_MUXInst_Y ;
    wire KeyArray_S23reg_gff_1_SFF_0_MUXInst_X ;
    wire KeyArray_S23reg_gff_1_SFF_1_n2 ;
    wire KeyArray_S23reg_gff_1_SFF_1_n1 ;
    wire KeyArray_S23reg_gff_1_SFF_1_QD ;
    wire KeyArray_S23reg_gff_1_SFF_1_MUXInst_Y ;
    wire KeyArray_S23reg_gff_1_SFF_1_MUXInst_X ;
    wire KeyArray_S23reg_gff_1_SFF_2_n2 ;
    wire KeyArray_S23reg_gff_1_SFF_2_n1 ;
    wire KeyArray_S23reg_gff_1_SFF_2_QD ;
    wire KeyArray_S23reg_gff_1_SFF_2_MUXInst_Y ;
    wire KeyArray_S23reg_gff_1_SFF_2_MUXInst_X ;
    wire KeyArray_S23reg_gff_1_SFF_3_n2 ;
    wire KeyArray_S23reg_gff_1_SFF_3_n1 ;
    wire KeyArray_S23reg_gff_1_SFF_3_QD ;
    wire KeyArray_S23reg_gff_1_SFF_3_MUXInst_Y ;
    wire KeyArray_S23reg_gff_1_SFF_3_MUXInst_X ;
    wire KeyArray_S23reg_gff_1_SFF_4_n2 ;
    wire KeyArray_S23reg_gff_1_SFF_4_n1 ;
    wire KeyArray_S23reg_gff_1_SFF_4_QD ;
    wire KeyArray_S23reg_gff_1_SFF_4_MUXInst_Y ;
    wire KeyArray_S23reg_gff_1_SFF_4_MUXInst_X ;
    wire KeyArray_S23reg_gff_1_SFF_5_n2 ;
    wire KeyArray_S23reg_gff_1_SFF_5_n1 ;
    wire KeyArray_S23reg_gff_1_SFF_5_QD ;
    wire KeyArray_S23reg_gff_1_SFF_5_MUXInst_Y ;
    wire KeyArray_S23reg_gff_1_SFF_5_MUXInst_X ;
    wire KeyArray_S23reg_gff_1_SFF_6_n2 ;
    wire KeyArray_S23reg_gff_1_SFF_6_n1 ;
    wire KeyArray_S23reg_gff_1_SFF_6_QD ;
    wire KeyArray_S23reg_gff_1_SFF_6_MUXInst_Y ;
    wire KeyArray_S23reg_gff_1_SFF_6_MUXInst_X ;
    wire KeyArray_S23reg_gff_1_SFF_7_n2 ;
    wire KeyArray_S23reg_gff_1_SFF_7_n1 ;
    wire KeyArray_S23reg_gff_1_SFF_7_QD ;
    wire KeyArray_S23reg_gff_1_SFF_7_MUXInst_Y ;
    wire KeyArray_S23reg_gff_1_SFF_7_MUXInst_X ;
    wire KeyArray_S30reg_gff_1_SFF_0_n2 ;
    wire KeyArray_S30reg_gff_1_SFF_0_n1 ;
    wire KeyArray_S30reg_gff_1_SFF_0_QD ;
    wire KeyArray_S30reg_gff_1_SFF_0_MUXInst_Y ;
    wire KeyArray_S30reg_gff_1_SFF_0_MUXInst_X ;
    wire KeyArray_S30reg_gff_1_SFF_1_n2 ;
    wire KeyArray_S30reg_gff_1_SFF_1_n1 ;
    wire KeyArray_S30reg_gff_1_SFF_1_QD ;
    wire KeyArray_S30reg_gff_1_SFF_1_MUXInst_Y ;
    wire KeyArray_S30reg_gff_1_SFF_1_MUXInst_X ;
    wire KeyArray_S30reg_gff_1_SFF_2_n2 ;
    wire KeyArray_S30reg_gff_1_SFF_2_n1 ;
    wire KeyArray_S30reg_gff_1_SFF_2_QD ;
    wire KeyArray_S30reg_gff_1_SFF_2_MUXInst_Y ;
    wire KeyArray_S30reg_gff_1_SFF_2_MUXInst_X ;
    wire KeyArray_S30reg_gff_1_SFF_3_n2 ;
    wire KeyArray_S30reg_gff_1_SFF_3_n1 ;
    wire KeyArray_S30reg_gff_1_SFF_3_QD ;
    wire KeyArray_S30reg_gff_1_SFF_3_MUXInst_Y ;
    wire KeyArray_S30reg_gff_1_SFF_3_MUXInst_X ;
    wire KeyArray_S30reg_gff_1_SFF_4_n2 ;
    wire KeyArray_S30reg_gff_1_SFF_4_n1 ;
    wire KeyArray_S30reg_gff_1_SFF_4_QD ;
    wire KeyArray_S30reg_gff_1_SFF_4_MUXInst_Y ;
    wire KeyArray_S30reg_gff_1_SFF_4_MUXInst_X ;
    wire KeyArray_S30reg_gff_1_SFF_5_n2 ;
    wire KeyArray_S30reg_gff_1_SFF_5_n1 ;
    wire KeyArray_S30reg_gff_1_SFF_5_QD ;
    wire KeyArray_S30reg_gff_1_SFF_5_MUXInst_Y ;
    wire KeyArray_S30reg_gff_1_SFF_5_MUXInst_X ;
    wire KeyArray_S30reg_gff_1_SFF_6_n2 ;
    wire KeyArray_S30reg_gff_1_SFF_6_n1 ;
    wire KeyArray_S30reg_gff_1_SFF_6_QD ;
    wire KeyArray_S30reg_gff_1_SFF_6_MUXInst_Y ;
    wire KeyArray_S30reg_gff_1_SFF_6_MUXInst_X ;
    wire KeyArray_S30reg_gff_1_SFF_7_n2 ;
    wire KeyArray_S30reg_gff_1_SFF_7_n1 ;
    wire KeyArray_S30reg_gff_1_SFF_7_QD ;
    wire KeyArray_S30reg_gff_1_SFF_7_MUXInst_Y ;
    wire KeyArray_S30reg_gff_1_SFF_7_MUXInst_X ;
    wire KeyArray_S31reg_gff_1_SFF_0_n2 ;
    wire KeyArray_S31reg_gff_1_SFF_0_n1 ;
    wire KeyArray_S31reg_gff_1_SFF_0_QD ;
    wire KeyArray_S31reg_gff_1_SFF_0_MUXInst_Y ;
    wire KeyArray_S31reg_gff_1_SFF_0_MUXInst_X ;
    wire KeyArray_S31reg_gff_1_SFF_1_n2 ;
    wire KeyArray_S31reg_gff_1_SFF_1_n1 ;
    wire KeyArray_S31reg_gff_1_SFF_1_QD ;
    wire KeyArray_S31reg_gff_1_SFF_1_MUXInst_Y ;
    wire KeyArray_S31reg_gff_1_SFF_1_MUXInst_X ;
    wire KeyArray_S31reg_gff_1_SFF_2_n2 ;
    wire KeyArray_S31reg_gff_1_SFF_2_n1 ;
    wire KeyArray_S31reg_gff_1_SFF_2_QD ;
    wire KeyArray_S31reg_gff_1_SFF_2_MUXInst_Y ;
    wire KeyArray_S31reg_gff_1_SFF_2_MUXInst_X ;
    wire KeyArray_S31reg_gff_1_SFF_3_n2 ;
    wire KeyArray_S31reg_gff_1_SFF_3_n1 ;
    wire KeyArray_S31reg_gff_1_SFF_3_QD ;
    wire KeyArray_S31reg_gff_1_SFF_3_MUXInst_Y ;
    wire KeyArray_S31reg_gff_1_SFF_3_MUXInst_X ;
    wire KeyArray_S31reg_gff_1_SFF_4_n2 ;
    wire KeyArray_S31reg_gff_1_SFF_4_n1 ;
    wire KeyArray_S31reg_gff_1_SFF_4_QD ;
    wire KeyArray_S31reg_gff_1_SFF_4_MUXInst_Y ;
    wire KeyArray_S31reg_gff_1_SFF_4_MUXInst_X ;
    wire KeyArray_S31reg_gff_1_SFF_5_n2 ;
    wire KeyArray_S31reg_gff_1_SFF_5_n1 ;
    wire KeyArray_S31reg_gff_1_SFF_5_QD ;
    wire KeyArray_S31reg_gff_1_SFF_5_MUXInst_Y ;
    wire KeyArray_S31reg_gff_1_SFF_5_MUXInst_X ;
    wire KeyArray_S31reg_gff_1_SFF_6_n2 ;
    wire KeyArray_S31reg_gff_1_SFF_6_n1 ;
    wire KeyArray_S31reg_gff_1_SFF_6_QD ;
    wire KeyArray_S31reg_gff_1_SFF_6_MUXInst_Y ;
    wire KeyArray_S31reg_gff_1_SFF_6_MUXInst_X ;
    wire KeyArray_S31reg_gff_1_SFF_7_n2 ;
    wire KeyArray_S31reg_gff_1_SFF_7_n1 ;
    wire KeyArray_S31reg_gff_1_SFF_7_QD ;
    wire KeyArray_S31reg_gff_1_SFF_7_MUXInst_Y ;
    wire KeyArray_S31reg_gff_1_SFF_7_MUXInst_X ;
    wire KeyArray_S32reg_gff_1_SFF_0_n2 ;
    wire KeyArray_S32reg_gff_1_SFF_0_n1 ;
    wire KeyArray_S32reg_gff_1_SFF_0_QD ;
    wire KeyArray_S32reg_gff_1_SFF_0_MUXInst_Y ;
    wire KeyArray_S32reg_gff_1_SFF_0_MUXInst_X ;
    wire KeyArray_S32reg_gff_1_SFF_1_n2 ;
    wire KeyArray_S32reg_gff_1_SFF_1_n1 ;
    wire KeyArray_S32reg_gff_1_SFF_1_QD ;
    wire KeyArray_S32reg_gff_1_SFF_1_MUXInst_Y ;
    wire KeyArray_S32reg_gff_1_SFF_1_MUXInst_X ;
    wire KeyArray_S32reg_gff_1_SFF_2_n2 ;
    wire KeyArray_S32reg_gff_1_SFF_2_n1 ;
    wire KeyArray_S32reg_gff_1_SFF_2_QD ;
    wire KeyArray_S32reg_gff_1_SFF_2_MUXInst_Y ;
    wire KeyArray_S32reg_gff_1_SFF_2_MUXInst_X ;
    wire KeyArray_S32reg_gff_1_SFF_3_n2 ;
    wire KeyArray_S32reg_gff_1_SFF_3_n1 ;
    wire KeyArray_S32reg_gff_1_SFF_3_QD ;
    wire KeyArray_S32reg_gff_1_SFF_3_MUXInst_Y ;
    wire KeyArray_S32reg_gff_1_SFF_3_MUXInst_X ;
    wire KeyArray_S32reg_gff_1_SFF_4_n2 ;
    wire KeyArray_S32reg_gff_1_SFF_4_n1 ;
    wire KeyArray_S32reg_gff_1_SFF_4_QD ;
    wire KeyArray_S32reg_gff_1_SFF_4_MUXInst_Y ;
    wire KeyArray_S32reg_gff_1_SFF_4_MUXInst_X ;
    wire KeyArray_S32reg_gff_1_SFF_5_n2 ;
    wire KeyArray_S32reg_gff_1_SFF_5_n1 ;
    wire KeyArray_S32reg_gff_1_SFF_5_QD ;
    wire KeyArray_S32reg_gff_1_SFF_5_MUXInst_Y ;
    wire KeyArray_S32reg_gff_1_SFF_5_MUXInst_X ;
    wire KeyArray_S32reg_gff_1_SFF_6_n2 ;
    wire KeyArray_S32reg_gff_1_SFF_6_n1 ;
    wire KeyArray_S32reg_gff_1_SFF_6_QD ;
    wire KeyArray_S32reg_gff_1_SFF_6_MUXInst_Y ;
    wire KeyArray_S32reg_gff_1_SFF_6_MUXInst_X ;
    wire KeyArray_S32reg_gff_1_SFF_7_n2 ;
    wire KeyArray_S32reg_gff_1_SFF_7_n1 ;
    wire KeyArray_S32reg_gff_1_SFF_7_QD ;
    wire KeyArray_S32reg_gff_1_SFF_7_MUXInst_Y ;
    wire KeyArray_S32reg_gff_1_SFF_7_MUXInst_X ;
    wire KeyArray_S33reg_gff_1_SFF_0_n2 ;
    wire KeyArray_S33reg_gff_1_SFF_0_n1 ;
    wire KeyArray_S33reg_gff_1_SFF_0_QD ;
    wire KeyArray_S33reg_gff_1_SFF_0_MUXInst_Y ;
    wire KeyArray_S33reg_gff_1_SFF_0_MUXInst_X ;
    wire KeyArray_S33reg_gff_1_SFF_1_n2 ;
    wire KeyArray_S33reg_gff_1_SFF_1_n1 ;
    wire KeyArray_S33reg_gff_1_SFF_1_QD ;
    wire KeyArray_S33reg_gff_1_SFF_1_MUXInst_Y ;
    wire KeyArray_S33reg_gff_1_SFF_1_MUXInst_X ;
    wire KeyArray_S33reg_gff_1_SFF_2_n2 ;
    wire KeyArray_S33reg_gff_1_SFF_2_n1 ;
    wire KeyArray_S33reg_gff_1_SFF_2_QD ;
    wire KeyArray_S33reg_gff_1_SFF_2_MUXInst_Y ;
    wire KeyArray_S33reg_gff_1_SFF_2_MUXInst_X ;
    wire KeyArray_S33reg_gff_1_SFF_3_n2 ;
    wire KeyArray_S33reg_gff_1_SFF_3_n1 ;
    wire KeyArray_S33reg_gff_1_SFF_3_QD ;
    wire KeyArray_S33reg_gff_1_SFF_3_MUXInst_Y ;
    wire KeyArray_S33reg_gff_1_SFF_3_MUXInst_X ;
    wire KeyArray_S33reg_gff_1_SFF_4_n2 ;
    wire KeyArray_S33reg_gff_1_SFF_4_n1 ;
    wire KeyArray_S33reg_gff_1_SFF_4_QD ;
    wire KeyArray_S33reg_gff_1_SFF_4_MUXInst_Y ;
    wire KeyArray_S33reg_gff_1_SFF_4_MUXInst_X ;
    wire KeyArray_S33reg_gff_1_SFF_5_n2 ;
    wire KeyArray_S33reg_gff_1_SFF_5_n1 ;
    wire KeyArray_S33reg_gff_1_SFF_5_QD ;
    wire KeyArray_S33reg_gff_1_SFF_5_MUXInst_Y ;
    wire KeyArray_S33reg_gff_1_SFF_5_MUXInst_X ;
    wire KeyArray_S33reg_gff_1_SFF_6_n2 ;
    wire KeyArray_S33reg_gff_1_SFF_6_n1 ;
    wire KeyArray_S33reg_gff_1_SFF_6_QD ;
    wire KeyArray_S33reg_gff_1_SFF_6_MUXInst_Y ;
    wire KeyArray_S33reg_gff_1_SFF_6_MUXInst_X ;
    wire KeyArray_S33reg_gff_1_SFF_7_n2 ;
    wire KeyArray_S33reg_gff_1_SFF_7_n1 ;
    wire KeyArray_S33reg_gff_1_SFF_7_QD ;
    wire KeyArray_S33reg_gff_1_SFF_7_MUXInst_Y ;
    wire KeyArray_S33reg_gff_1_SFF_7_MUXInst_X ;
    wire KeyArray_MUX_inS00ser_mux_inst_0_Y ;
    wire KeyArray_MUX_inS00ser_mux_inst_0_X ;
    wire KeyArray_MUX_inS00ser_mux_inst_1_Y ;
    wire KeyArray_MUX_inS00ser_mux_inst_1_X ;
    wire KeyArray_MUX_inS00ser_mux_inst_2_Y ;
    wire KeyArray_MUX_inS00ser_mux_inst_2_X ;
    wire KeyArray_MUX_inS00ser_mux_inst_3_Y ;
    wire KeyArray_MUX_inS00ser_mux_inst_3_X ;
    wire KeyArray_MUX_inS00ser_mux_inst_4_Y ;
    wire KeyArray_MUX_inS00ser_mux_inst_4_X ;
    wire KeyArray_MUX_inS00ser_mux_inst_5_Y ;
    wire KeyArray_MUX_inS00ser_mux_inst_5_X ;
    wire KeyArray_MUX_inS00ser_mux_inst_6_Y ;
    wire KeyArray_MUX_inS00ser_mux_inst_6_X ;
    wire KeyArray_MUX_inS00ser_mux_inst_7_Y ;
    wire KeyArray_MUX_inS00ser_mux_inst_7_X ;
    wire KeyArray_MUX_inS33ser_mux_inst_0_Y ;
    wire KeyArray_MUX_inS33ser_mux_inst_0_X ;
    wire KeyArray_MUX_inS33ser_mux_inst_1_Y ;
    wire KeyArray_MUX_inS33ser_mux_inst_1_X ;
    wire KeyArray_MUX_inS33ser_mux_inst_2_Y ;
    wire KeyArray_MUX_inS33ser_mux_inst_2_X ;
    wire KeyArray_MUX_inS33ser_mux_inst_3_Y ;
    wire KeyArray_MUX_inS33ser_mux_inst_3_X ;
    wire KeyArray_MUX_inS33ser_mux_inst_4_Y ;
    wire KeyArray_MUX_inS33ser_mux_inst_4_X ;
    wire KeyArray_MUX_inS33ser_mux_inst_5_Y ;
    wire KeyArray_MUX_inS33ser_mux_inst_5_X ;
    wire KeyArray_MUX_inS33ser_mux_inst_6_Y ;
    wire KeyArray_MUX_inS33ser_mux_inst_6_X ;
    wire KeyArray_MUX_inS33ser_mux_inst_7_Y ;
    wire KeyArray_MUX_inS33ser_mux_inst_7_X ;
    wire MixColumns_line0_n16 ;
    wire MixColumns_line0_n15 ;
    wire MixColumns_line0_n14 ;
    wire MixColumns_line0_n13 ;
    wire MixColumns_line0_n12 ;
    wire MixColumns_line0_n11 ;
    wire MixColumns_line0_n10 ;
    wire MixColumns_line0_n9 ;
    wire MixColumns_line0_n8 ;
    wire MixColumns_line0_n7 ;
    wire MixColumns_line0_n6 ;
    wire MixColumns_line0_n5 ;
    wire MixColumns_line0_n4 ;
    wire MixColumns_line0_n3 ;
    wire MixColumns_line0_n2 ;
    wire MixColumns_line0_n1 ;
    wire MixColumns_line1_n16 ;
    wire MixColumns_line1_n15 ;
    wire MixColumns_line1_n14 ;
    wire MixColumns_line1_n13 ;
    wire MixColumns_line1_n12 ;
    wire MixColumns_line1_n11 ;
    wire MixColumns_line1_n10 ;
    wire MixColumns_line1_n9 ;
    wire MixColumns_line1_n8 ;
    wire MixColumns_line1_n7 ;
    wire MixColumns_line1_n6 ;
    wire MixColumns_line1_n5 ;
    wire MixColumns_line1_n4 ;
    wire MixColumns_line1_n3 ;
    wire MixColumns_line1_n2 ;
    wire MixColumns_line1_n1 ;
    wire MixColumns_line2_n16 ;
    wire MixColumns_line2_n15 ;
    wire MixColumns_line2_n14 ;
    wire MixColumns_line2_n13 ;
    wire MixColumns_line2_n12 ;
    wire MixColumns_line2_n11 ;
    wire MixColumns_line2_n10 ;
    wire MixColumns_line2_n9 ;
    wire MixColumns_line2_n8 ;
    wire MixColumns_line2_n7 ;
    wire MixColumns_line2_n6 ;
    wire MixColumns_line2_n5 ;
    wire MixColumns_line2_n4 ;
    wire MixColumns_line2_n3 ;
    wire MixColumns_line2_n2 ;
    wire MixColumns_line2_n1 ;
    wire MixColumns_line3_n16 ;
    wire MixColumns_line3_n15 ;
    wire MixColumns_line3_n14 ;
    wire MixColumns_line3_n13 ;
    wire MixColumns_line3_n12 ;
    wire MixColumns_line3_n11 ;
    wire MixColumns_line3_n10 ;
    wire MixColumns_line3_n9 ;
    wire MixColumns_line3_n8 ;
    wire MixColumns_line3_n7 ;
    wire MixColumns_line3_n6 ;
    wire MixColumns_line3_n5 ;
    wire MixColumns_line3_n4 ;
    wire MixColumns_line3_n3 ;
    wire MixColumns_line3_n2 ;
    wire MixColumns_line3_n1 ;
    wire MixColumns_line3_timesTHREE_input2_1_ ;
    wire MixColumns_line3_timesTHREE_input2_3_ ;
    wire MixColumns_line3_timesTHREE_input2_4_ ;
    wire calcRCon_n42 ;
    wire calcRCon_n41 ;
    wire calcRCon_n40 ;
    wire calcRCon_n39 ;
    wire calcRCon_n38 ;
    wire calcRCon_n37 ;
    wire calcRCon_n36 ;
    wire calcRCon_n35 ;
    wire calcRCon_n34 ;
    wire calcRCon_n33 ;
    wire calcRCon_n32 ;
    wire calcRCon_n31 ;
    wire calcRCon_n30 ;
    wire calcRCon_n29 ;
    wire calcRCon_n28 ;
    wire calcRCon_n27 ;
    wire calcRCon_n26 ;
    wire calcRCon_n25 ;
    wire calcRCon_n24 ;
    wire calcRCon_n23 ;
    wire calcRCon_n22 ;
    wire calcRCon_n21 ;
    wire calcRCon_n20 ;
    wire calcRCon_n19 ;
    wire calcRCon_n18 ;
    wire calcRCon_n17 ;
    wire calcRCon_n16 ;
    wire calcRCon_n15 ;
    wire calcRCon_n14 ;
    wire calcRCon_n13 ;
    wire calcRCon_n9 ;
    wire calcRCon_n8 ;
    wire calcRCon_n7 ;
    wire calcRCon_s_current_state_0_ ;
    wire calcRCon_s_current_state_1_ ;
    wire calcRCon_s_current_state_2_ ;
    wire calcRCon_s_current_state_3_ ;
    wire calcRCon_s_current_state_4_ ;
    wire calcRCon_s_current_state_5_ ;
    wire calcRCon_s_current_state_6_ ;
    wire calcRCon_s_current_state_7_ ;
    wire MUX_SboxIn_mux_inst_0_Y ;
    wire MUX_SboxIn_mux_inst_0_X ;
    wire MUX_SboxIn_mux_inst_1_Y ;
    wire MUX_SboxIn_mux_inst_1_X ;
    wire MUX_SboxIn_mux_inst_2_Y ;
    wire MUX_SboxIn_mux_inst_2_X ;
    wire MUX_SboxIn_mux_inst_3_Y ;
    wire MUX_SboxIn_mux_inst_3_X ;
    wire MUX_SboxIn_mux_inst_4_Y ;
    wire MUX_SboxIn_mux_inst_4_X ;
    wire MUX_SboxIn_mux_inst_5_Y ;
    wire MUX_SboxIn_mux_inst_5_X ;
    wire MUX_SboxIn_mux_inst_6_Y ;
    wire MUX_SboxIn_mux_inst_6_X ;
    wire MUX_SboxIn_mux_inst_7_Y ;
    wire MUX_SboxIn_mux_inst_7_X ;
    wire Inst_bSbox_L29 ;
    wire Inst_bSbox_L28 ;
    wire Inst_bSbox_L27 ;
    wire Inst_bSbox_L26 ;
    wire Inst_bSbox_L25 ;
    wire Inst_bSbox_L24 ;
    wire Inst_bSbox_L23 ;
    wire Inst_bSbox_L22 ;
    wire Inst_bSbox_L21 ;
    wire Inst_bSbox_L20 ;
    wire Inst_bSbox_L19 ;
    wire Inst_bSbox_L18 ;
    wire Inst_bSbox_L17 ;
    wire Inst_bSbox_L16 ;
    wire Inst_bSbox_L15 ;
    wire Inst_bSbox_L14 ;
    wire Inst_bSbox_L13 ;
    wire Inst_bSbox_L12 ;
    wire Inst_bSbox_L11 ;
    wire Inst_bSbox_L10 ;
    wire Inst_bSbox_L9 ;
    wire Inst_bSbox_L8 ;
    wire Inst_bSbox_L7 ;
    wire Inst_bSbox_L6 ;
    wire Inst_bSbox_L5 ;
    wire Inst_bSbox_L4 ;
    wire Inst_bSbox_L3 ;
    wire Inst_bSbox_L2 ;
    wire Inst_bSbox_L1 ;
    wire Inst_bSbox_L0 ;
    wire Inst_bSbox_M63 ;
    wire Inst_bSbox_M62 ;
    wire Inst_bSbox_M61 ;
    wire Inst_bSbox_M60 ;
    wire Inst_bSbox_M59 ;
    wire Inst_bSbox_M58 ;
    wire Inst_bSbox_M57 ;
    wire Inst_bSbox_M56 ;
    wire Inst_bSbox_M55 ;
    wire Inst_bSbox_M54 ;
    wire Inst_bSbox_M53 ;
    wire Inst_bSbox_M52 ;
    wire Inst_bSbox_M51 ;
    wire Inst_bSbox_M50 ;
    wire Inst_bSbox_M49 ;
    wire Inst_bSbox_M48 ;
    wire Inst_bSbox_M47 ;
    wire Inst_bSbox_M46 ;
    wire Inst_bSbox_M45 ;
    wire Inst_bSbox_M44 ;
    wire Inst_bSbox_M43 ;
    wire Inst_bSbox_M42 ;
    wire Inst_bSbox_M41 ;
    wire Inst_bSbox_M40 ;
    wire Inst_bSbox_M39 ;
    wire Inst_bSbox_M38 ;
    wire Inst_bSbox_M37 ;
    wire Inst_bSbox_M36 ;
    wire Inst_bSbox_M35 ;
    wire Inst_bSbox_M34 ;
    wire Inst_bSbox_M33 ;
    wire Inst_bSbox_M32 ;
    wire Inst_bSbox_M31 ;
    wire Inst_bSbox_M30 ;
    wire Inst_bSbox_M29 ;
    wire Inst_bSbox_M28 ;
    wire Inst_bSbox_M27 ;
    wire Inst_bSbox_M26 ;
    wire Inst_bSbox_M25 ;
    wire Inst_bSbox_M24 ;
    wire Inst_bSbox_M23 ;
    wire Inst_bSbox_M22 ;
    wire Inst_bSbox_M21 ;
    wire Inst_bSbox_M20 ;
    wire Inst_bSbox_M19 ;
    wire Inst_bSbox_M18 ;
    wire Inst_bSbox_M17 ;
    wire Inst_bSbox_M16 ;
    wire Inst_bSbox_M15 ;
    wire Inst_bSbox_M14 ;
    wire Inst_bSbox_M13 ;
    wire Inst_bSbox_M12 ;
    wire Inst_bSbox_M11 ;
    wire Inst_bSbox_M10 ;
    wire Inst_bSbox_M9 ;
    wire Inst_bSbox_M8 ;
    wire Inst_bSbox_M7 ;
    wire Inst_bSbox_M6 ;
    wire Inst_bSbox_M5 ;
    wire Inst_bSbox_M4 ;
    wire Inst_bSbox_M3 ;
    wire Inst_bSbox_M2 ;
    wire Inst_bSbox_M1 ;
    wire Inst_bSbox_T27 ;
    wire Inst_bSbox_T26 ;
    wire Inst_bSbox_T25 ;
    wire Inst_bSbox_T24 ;
    wire Inst_bSbox_T23 ;
    wire Inst_bSbox_T22 ;
    wire Inst_bSbox_T21 ;
    wire Inst_bSbox_T20 ;
    wire Inst_bSbox_T19 ;
    wire Inst_bSbox_T18 ;
    wire Inst_bSbox_T17 ;
    wire Inst_bSbox_T16 ;
    wire Inst_bSbox_T15 ;
    wire Inst_bSbox_T14 ;
    wire Inst_bSbox_T13 ;
    wire Inst_bSbox_T12 ;
    wire Inst_bSbox_T11 ;
    wire Inst_bSbox_T10 ;
    wire Inst_bSbox_T9 ;
    wire Inst_bSbox_T8 ;
    wire Inst_bSbox_T7 ;
    wire Inst_bSbox_T6 ;
    wire Inst_bSbox_T5 ;
    wire Inst_bSbox_T4 ;
    wire Inst_bSbox_T3 ;
    wire Inst_bSbox_T2 ;
    wire Inst_bSbox_T1 ;
    wire [7:0] SboxOut ;
    wire [7:0] StateOutXORroundKey ;
    wire [7:0] StateIn ;
    wire [31:0] StateInMC ;
    wire [19:0] MCin ;
    wire [31:0] MCout ;
    wire [7:0] keyStateIn ;
    wire [7:0] roundConstant ;
    wire [7:0] keySBIn ;
    wire [7:0] SboxIn ;
    wire [7:0] stateArray_input_MC ;
    wire [7:0] stateArray_inS33ser ;
    wire [7:0] stateArray_outS33ser ;
    wire [7:0] stateArray_outS32ser ;
    wire [7:0] stateArray_outS31ser ;
    wire [7:0] stateArray_inS23ser ;
    wire [7:0] stateArray_outS23ser ;
    wire [7:0] stateArray_outS22ser ;
    wire [7:0] stateArray_outS21ser ;
    wire [7:0] stateArray_inS13ser ;
    wire [7:0] stateArray_outS13ser ;
    wire [7:0] stateArray_outS12ser ;
    wire [7:0] stateArray_outS11ser ;
    wire [7:0] stateArray_inS03ser ;
    wire [7:0] stateArray_outS03ser ;
    wire [7:0] stateArray_outS02ser ;
    wire [7:0] stateArray_outS01ser ;
    wire [7:0] KeyArray_outS01ser_XOR_00 ;
    wire [7:0] KeyArray_inS33ser ;
    wire [7:0] KeyArray_outS33ser ;
    wire [7:0] KeyArray_outS32ser ;
    wire [7:0] KeyArray_inS30par ;
    wire [7:0] KeyArray_outS31ser ;
    wire [7:0] KeyArray_outS30ser ;
    wire [7:0] KeyArray_outS23ser ;
    wire [7:0] KeyArray_outS22ser ;
    wire [7:0] KeyArray_outS21ser ;
    wire [7:0] KeyArray_outS20ser ;
    wire [7:0] KeyArray_outS12ser ;
    wire [7:0] KeyArray_outS11ser ;
    wire [7:0] KeyArray_outS10ser ;
    wire [7:0] KeyArray_outS03ser ;
    wire [7:0] KeyArray_outS02ser ;
    wire [7:0] KeyArray_inS00ser ;
    wire [7:0] MixColumns_line0_S13 ;
    wire [4:1] MixColumns_line0_S02 ;
    wire [4:1] MixColumns_line0_timesTHREE_input2 ;
    wire [7:0] MixColumns_line1_S13 ;
    wire [7:0] MixColumns_line1_S02 ;
    wire [4:1] MixColumns_line1_timesTHREE_input2 ;
    wire [7:0] MixColumns_line2_S13 ;
    wire [7:0] MixColumns_line2_S02 ;
    wire [4:1] MixColumns_line2_timesTHREE_input2 ;
    wire [7:0] MixColumns_line3_S13 ;
    wire [7:0] MixColumns_line3_S02 ;

    /* cells in depth 0 */
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) U23 ( .A0_t (ctrl_n4), .B0_t (start), .Z0_t (enKS) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U25 ( .A0_t (keyStateIn[0]), .B0_t (port_out[0]), .Z0_t (StateOutXORroundKey[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U26 ( .A0_t (keyStateIn[1]), .B0_t (port_out[1]), .Z0_t (StateOutXORroundKey[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U27 ( .A0_t (keyStateIn[2]), .B0_t (port_out[2]), .Z0_t (StateOutXORroundKey[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U28 ( .A0_t (keyStateIn[3]), .B0_t (port_out[3]), .Z0_t (StateOutXORroundKey[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U29 ( .A0_t (keyStateIn[4]), .B0_t (port_out[4]), .Z0_t (StateOutXORroundKey[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U30 ( .A0_t (keyStateIn[5]), .B0_t (port_out[5]), .Z0_t (StateOutXORroundKey[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U31 ( .A0_t (keyStateIn[6]), .B0_t (port_out[6]), .Z0_t (StateOutXORroundKey[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U32 ( .A0_t (keyStateIn[7]), .B0_t (port_out[7]), .Z0_t (StateOutXORroundKey[7]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) U33 ( .A0_t (notFirst), .B0_t (selXOR), .Z0_t (intselXOR) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) ctrl_U25 ( .A0_t (ctrl_n24), .B0_t (start), .Z0_t (ctrl_nRstSeq4) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b0)) ctrl_U24 ( .A0_t (ctrl_seq6Out_4_), .B0_t (ctrl_seq6In_1_), .Z0_t (ctrl_n22) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1), .NL(1'b1)) ctrl_U23 ( .A0_t (ctrl_n4), .B0_t (ctrl_n19), .Z0_t (ctrl_n5) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) ctrl_U22 ( .A0_t (selXOR), .B0_t (ctrl_n5), .Z0_t (ctrl_n19) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) ctrl_U21 ( .A0_t (start), .B0_t (ctrl_n18), .Z0_t (selXOR) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) ctrl_U20 ( .A0_t (ctrl_seq4Out_1_), .B0_t (ctrl_seq4In_1_), .Z0_t (ctrl_n18) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b1), .NL(1'b1)) ctrl_U19 ( .A0_t (ctrl_n4), .B0_t (ctrl_n17), .Z0_t (enRCon) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) ctrl_U18 ( .A0_t (enRCon), .B0_t (done), .Z0_t (ctrl_n17) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) ctrl_U17 ( .A0_t (start), .B0_t (ctrl_n24), .Z0_t (ctrl_n14) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) ctrl_U16 ( .A0_t (ctrl_seq4Out_1_), .B0_t (ctrl_n12), .Z0_t (ctrl_finalStep) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) ctrl_U15 ( .A0_t (ctrl_n24), .B0_t (ctrl_seq4In_1_), .Z0_t (ctrl_n12) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) ctrl_U14 ( .A0_t (ctrl_n10), .B0_t (ctrl_n9), .Z0_t (ctrl_n11) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) ctrl_U13 ( .A0_t (ctrl_seq6In_3_), .B0_t (ctrl_seq6Out_4_), .Z0_t (ctrl_n9) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) ctrl_U12 ( .A0_t (ctrl_seq6In_1_), .B0_t (ctrl_seq6In_4_), .Z0_t (ctrl_n10) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) ctrl_U9 ( .A0_t (ctrl_seq6In_2_), .B0_t (ctrl_n11), .Z0_t (ctrl_n24) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) ctrl_U8 ( .A0_t (start), .B0_t (ctrl_n13), .Z0_t (done) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) ctrl_U6 ( .A0_t (ctrl_finalStep), .B0_t (intFinal), .Z0_t (ctrl_n13) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) ctrl_U5 ( .A0_t (done), .B0_t (ctrl_n14), .Z0_t (ctrl_n4) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) ctrl_U3 ( .A0_t (ctrl_n5), .B0_t (start), .Z0_t (selMC) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1), .NL(1'b1)) ctrl_seq6_SFF_0_U3 ( .A0_t (ctrl_seq6_SFF_0_n2), .B0_t (ctrl_seq6_SFF_0_n1), .Z0_t (ctrl_seq6In_1_) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) ctrl_seq6_SFF_0_U2 ( .A0_t (done), .B0_t (ctrl_seq6In_1_), .Z0_t (ctrl_seq6_SFF_0_n1) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) ctrl_seq6_SFF_0_U1 ( .A0_t (ctrl_seq6_SFF_0_QD), .B0_t (done), .Z0_t (ctrl_seq6_SFF_0_n2) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) ctrl_seq6_SFF_0_MUXInst_XOR1_U1 ( .A0_t (1'b1), .B0_t (ctrl_n22), .Z0_t (ctrl_seq6_SFF_0_MUXInst_X) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) ctrl_seq6_SFF_0_MUXInst_AND1_U1 ( .A0_t (start), .B0_t (ctrl_seq6_SFF_0_MUXInst_X), .Z0_t (ctrl_seq6_SFF_0_MUXInst_Y) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) ctrl_seq6_SFF_0_MUXInst_XOR2_U1 ( .A0_t (ctrl_seq6_SFF_0_MUXInst_Y), .B0_t (1'b1), .Z0_t (ctrl_seq6_SFF_0_QD) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1), .NL(1'b1)) ctrl_seq6_SFF_1_U3 ( .A0_t (ctrl_seq6_SFF_1_n2), .B0_t (ctrl_seq6_SFF_1_n1), .Z0_t (ctrl_seq6In_2_) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) ctrl_seq6_SFF_1_U2 ( .A0_t (done), .B0_t (ctrl_seq6In_2_), .Z0_t (ctrl_seq6_SFF_1_n1) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) ctrl_seq6_SFF_1_U1 ( .A0_t (ctrl_seq6_SFF_1_QD), .B0_t (done), .Z0_t (ctrl_seq6_SFF_1_n2) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) ctrl_seq6_SFF_1_MUXInst_XOR1_U1 ( .A0_t (1'b0), .B0_t (ctrl_seq6In_1_), .Z0_t (ctrl_seq6_SFF_1_MUXInst_X) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) ctrl_seq6_SFF_1_MUXInst_AND1_U1 ( .A0_t (start), .B0_t (ctrl_seq6_SFF_1_MUXInst_X), .Z0_t (ctrl_seq6_SFF_1_MUXInst_Y) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) ctrl_seq6_SFF_1_MUXInst_XOR2_U1 ( .A0_t (ctrl_seq6_SFF_1_MUXInst_Y), .B0_t (1'b0), .Z0_t (ctrl_seq6_SFF_1_QD) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1), .NL(1'b1)) ctrl_seq6_SFF_2_U3 ( .A0_t (ctrl_seq6_SFF_2_n2), .B0_t (ctrl_seq6_SFF_2_n1), .Z0_t (ctrl_seq6In_3_) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) ctrl_seq6_SFF_2_U2 ( .A0_t (done), .B0_t (ctrl_seq6In_3_), .Z0_t (ctrl_seq6_SFF_2_n1) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) ctrl_seq6_SFF_2_U1 ( .A0_t (ctrl_seq6_SFF_2_QD), .B0_t (done), .Z0_t (ctrl_seq6_SFF_2_n2) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) ctrl_seq6_SFF_2_MUXInst_XOR1_U1 ( .A0_t (1'b1), .B0_t (ctrl_seq6In_2_), .Z0_t (ctrl_seq6_SFF_2_MUXInst_X) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) ctrl_seq6_SFF_2_MUXInst_AND1_U1 ( .A0_t (start), .B0_t (ctrl_seq6_SFF_2_MUXInst_X), .Z0_t (ctrl_seq6_SFF_2_MUXInst_Y) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) ctrl_seq6_SFF_2_MUXInst_XOR2_U1 ( .A0_t (ctrl_seq6_SFF_2_MUXInst_Y), .B0_t (1'b1), .Z0_t (ctrl_seq6_SFF_2_QD) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1), .NL(1'b1)) ctrl_seq6_SFF_3_U3 ( .A0_t (ctrl_seq6_SFF_3_n2), .B0_t (ctrl_seq6_SFF_3_n1), .Z0_t (ctrl_seq6In_4_) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) ctrl_seq6_SFF_3_U2 ( .A0_t (done), .B0_t (ctrl_seq6In_4_), .Z0_t (ctrl_seq6_SFF_3_n1) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) ctrl_seq6_SFF_3_U1 ( .A0_t (ctrl_seq6_SFF_3_QD), .B0_t (done), .Z0_t (ctrl_seq6_SFF_3_n2) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) ctrl_seq6_SFF_3_MUXInst_XOR1_U1 ( .A0_t (1'b0), .B0_t (ctrl_seq6In_3_), .Z0_t (ctrl_seq6_SFF_3_MUXInst_X) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) ctrl_seq6_SFF_3_MUXInst_AND1_U1 ( .A0_t (start), .B0_t (ctrl_seq6_SFF_3_MUXInst_X), .Z0_t (ctrl_seq6_SFF_3_MUXInst_Y) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) ctrl_seq6_SFF_3_MUXInst_XOR2_U1 ( .A0_t (ctrl_seq6_SFF_3_MUXInst_Y), .B0_t (1'b0), .Z0_t (ctrl_seq6_SFF_3_QD) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1), .NL(1'b1)) ctrl_seq6_SFF_4_U3 ( .A0_t (ctrl_seq6_SFF_4_n2), .B0_t (ctrl_seq6_SFF_4_n1), .Z0_t (ctrl_seq6Out_4_) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) ctrl_seq6_SFF_4_U2 ( .A0_t (done), .B0_t (ctrl_seq6Out_4_), .Z0_t (ctrl_seq6_SFF_4_n1) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) ctrl_seq6_SFF_4_U1 ( .A0_t (ctrl_seq6_SFF_4_QD), .B0_t (done), .Z0_t (ctrl_seq6_SFF_4_n2) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) ctrl_seq6_SFF_4_MUXInst_XOR1_U1 ( .A0_t (1'b1), .B0_t (ctrl_seq6In_4_), .Z0_t (ctrl_seq6_SFF_4_MUXInst_X) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) ctrl_seq6_SFF_4_MUXInst_AND1_U1 ( .A0_t (start), .B0_t (ctrl_seq6_SFF_4_MUXInst_X), .Z0_t (ctrl_seq6_SFF_4_MUXInst_Y) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) ctrl_seq6_SFF_4_MUXInst_XOR2_U1 ( .A0_t (ctrl_seq6_SFF_4_MUXInst_Y), .B0_t (1'b1), .Z0_t (ctrl_seq6_SFF_4_QD) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1), .NL(1'b1)) ctrl_seq4_SFF_0_U3 ( .A0_t (ctrl_seq4_SFF_0_n2), .B0_t (ctrl_seq4_SFF_0_n1), .Z0_t (ctrl_seq4In_1_) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) ctrl_seq4_SFF_0_U2 ( .A0_t (done), .B0_t (ctrl_seq4In_1_), .Z0_t (ctrl_seq4_SFF_0_n1) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) ctrl_seq4_SFF_0_U1 ( .A0_t (ctrl_seq4_SFF_0_QD), .B0_t (done), .Z0_t (ctrl_seq4_SFF_0_n2) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) ctrl_seq4_SFF_0_MUXInst_XOR1_U1 ( .A0_t (1'b1), .B0_t (ctrl_seq4Out_1_), .Z0_t (ctrl_seq4_SFF_0_MUXInst_X) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) ctrl_seq4_SFF_0_MUXInst_AND1_U1 ( .A0_t (ctrl_nRstSeq4), .B0_t (ctrl_seq4_SFF_0_MUXInst_X), .Z0_t (ctrl_seq4_SFF_0_MUXInst_Y) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) ctrl_seq4_SFF_0_MUXInst_XOR2_U1 ( .A0_t (ctrl_seq4_SFF_0_MUXInst_Y), .B0_t (1'b1), .Z0_t (ctrl_seq4_SFF_0_QD) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1), .NL(1'b1)) ctrl_seq4_SFF_1_U3 ( .A0_t (ctrl_seq4_SFF_1_n2), .B0_t (ctrl_seq4_SFF_1_n1), .Z0_t (ctrl_seq4Out_1_) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) ctrl_seq4_SFF_1_U2 ( .A0_t (done), .B0_t (ctrl_seq4Out_1_), .Z0_t (ctrl_seq4_SFF_1_n1) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) ctrl_seq4_SFF_1_U1 ( .A0_t (ctrl_seq4_SFF_1_QD), .B0_t (done), .Z0_t (ctrl_seq4_SFF_1_n2) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) ctrl_seq4_SFF_1_MUXInst_XOR1_U1 ( .A0_t (1'b0), .B0_t (ctrl_seq4In_1_), .Z0_t (ctrl_seq4_SFF_1_MUXInst_X) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) ctrl_seq4_SFF_1_MUXInst_AND1_U1 ( .A0_t (ctrl_nRstSeq4), .B0_t (ctrl_seq4_SFF_1_MUXInst_X), .Z0_t (ctrl_seq4_SFF_1_MUXInst_Y) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) ctrl_seq4_SFF_1_MUXInst_XOR2_U1 ( .A0_t (ctrl_seq4_SFF_1_MUXInst_Y), .B0_t (1'b0), .Z0_t (ctrl_seq4_SFF_1_QD) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_0_XOR1_U1 ( .A0_t (SboxOut[0]), .B0_t (StateOutXORroundKey[0]), .Z0_t (MUX_StateIn_mux_inst_0_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_0_AND1_U1 ( .A0_t (intFinal), .B0_t (MUX_StateIn_mux_inst_0_X), .Z0_t (MUX_StateIn_mux_inst_0_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_0_XOR2_U1 ( .A0_t (MUX_StateIn_mux_inst_0_Y), .B0_t (SboxOut[0]), .Z0_t (StateIn[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_1_XOR1_U1 ( .A0_t (SboxOut[1]), .B0_t (StateOutXORroundKey[1]), .Z0_t (MUX_StateIn_mux_inst_1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_1_AND1_U1 ( .A0_t (intFinal), .B0_t (MUX_StateIn_mux_inst_1_X), .Z0_t (MUX_StateIn_mux_inst_1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_1_XOR2_U1 ( .A0_t (MUX_StateIn_mux_inst_1_Y), .B0_t (SboxOut[1]), .Z0_t (StateIn[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_2_XOR1_U1 ( .A0_t (SboxOut[2]), .B0_t (StateOutXORroundKey[2]), .Z0_t (MUX_StateIn_mux_inst_2_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_2_AND1_U1 ( .A0_t (intFinal), .B0_t (MUX_StateIn_mux_inst_2_X), .Z0_t (MUX_StateIn_mux_inst_2_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_2_XOR2_U1 ( .A0_t (MUX_StateIn_mux_inst_2_Y), .B0_t (SboxOut[2]), .Z0_t (StateIn[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_3_XOR1_U1 ( .A0_t (SboxOut[3]), .B0_t (StateOutXORroundKey[3]), .Z0_t (MUX_StateIn_mux_inst_3_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_3_AND1_U1 ( .A0_t (intFinal), .B0_t (MUX_StateIn_mux_inst_3_X), .Z0_t (MUX_StateIn_mux_inst_3_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_3_XOR2_U1 ( .A0_t (MUX_StateIn_mux_inst_3_Y), .B0_t (SboxOut[3]), .Z0_t (StateIn[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_4_XOR1_U1 ( .A0_t (SboxOut[4]), .B0_t (StateOutXORroundKey[4]), .Z0_t (MUX_StateIn_mux_inst_4_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_4_AND1_U1 ( .A0_t (intFinal), .B0_t (MUX_StateIn_mux_inst_4_X), .Z0_t (MUX_StateIn_mux_inst_4_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_4_XOR2_U1 ( .A0_t (MUX_StateIn_mux_inst_4_Y), .B0_t (SboxOut[4]), .Z0_t (StateIn[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_5_XOR1_U1 ( .A0_t (SboxOut[5]), .B0_t (StateOutXORroundKey[5]), .Z0_t (MUX_StateIn_mux_inst_5_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_5_AND1_U1 ( .A0_t (intFinal), .B0_t (MUX_StateIn_mux_inst_5_X), .Z0_t (MUX_StateIn_mux_inst_5_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_5_XOR2_U1 ( .A0_t (MUX_StateIn_mux_inst_5_Y), .B0_t (SboxOut[5]), .Z0_t (StateIn[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_6_XOR1_U1 ( .A0_t (SboxOut[6]), .B0_t (StateOutXORroundKey[6]), .Z0_t (MUX_StateIn_mux_inst_6_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_6_AND1_U1 ( .A0_t (intFinal), .B0_t (MUX_StateIn_mux_inst_6_X), .Z0_t (MUX_StateIn_mux_inst_6_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_6_XOR2_U1 ( .A0_t (MUX_StateIn_mux_inst_6_Y), .B0_t (SboxOut[6]), .Z0_t (StateIn[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_7_XOR1_U1 ( .A0_t (SboxOut[7]), .B0_t (StateOutXORroundKey[7]), .Z0_t (MUX_StateIn_mux_inst_7_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_7_AND1_U1 ( .A0_t (intFinal), .B0_t (MUX_StateIn_mux_inst_7_X), .Z0_t (MUX_StateIn_mux_inst_7_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_7_XOR2_U1 ( .A0_t (MUX_StateIn_mux_inst_7_Y), .B0_t (SboxOut[7]), .Z0_t (StateIn[7]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) stateArray_U3 ( .A0_t (start), .B0_t (selMC), .Z0_t (stateArray_nReset_selMC) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S00reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS01ser[0]), .B0_t (port_out[0]), .Z0_t (stateArray_S00reg_gff_1_SFF_0_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S00reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S00reg_gff_1_SFF_0_MUXInst_X), .Z0_t (stateArray_S00reg_gff_1_SFF_0_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S00reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (stateArray_S00reg_gff_1_SFF_0_MUXInst_Y), .B0_t (stateArray_outS01ser[0]), .Z0_t (port_out[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S00reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS01ser[1]), .B0_t (port_out[1]), .Z0_t (stateArray_S00reg_gff_1_SFF_1_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S00reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S00reg_gff_1_SFF_1_MUXInst_X), .Z0_t (stateArray_S00reg_gff_1_SFF_1_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S00reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (stateArray_S00reg_gff_1_SFF_1_MUXInst_Y), .B0_t (stateArray_outS01ser[1]), .Z0_t (port_out[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S00reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS01ser[2]), .B0_t (port_out[2]), .Z0_t (stateArray_S00reg_gff_1_SFF_2_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S00reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S00reg_gff_1_SFF_2_MUXInst_X), .Z0_t (stateArray_S00reg_gff_1_SFF_2_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S00reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (stateArray_S00reg_gff_1_SFF_2_MUXInst_Y), .B0_t (stateArray_outS01ser[2]), .Z0_t (port_out[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S00reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS01ser[3]), .B0_t (port_out[3]), .Z0_t (stateArray_S00reg_gff_1_SFF_3_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S00reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S00reg_gff_1_SFF_3_MUXInst_X), .Z0_t (stateArray_S00reg_gff_1_SFF_3_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S00reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (stateArray_S00reg_gff_1_SFF_3_MUXInst_Y), .B0_t (stateArray_outS01ser[3]), .Z0_t (port_out[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S00reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS01ser[4]), .B0_t (port_out[4]), .Z0_t (stateArray_S00reg_gff_1_SFF_4_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S00reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S00reg_gff_1_SFF_4_MUXInst_X), .Z0_t (stateArray_S00reg_gff_1_SFF_4_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S00reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (stateArray_S00reg_gff_1_SFF_4_MUXInst_Y), .B0_t (stateArray_outS01ser[4]), .Z0_t (port_out[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S00reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS01ser[5]), .B0_t (port_out[5]), .Z0_t (stateArray_S00reg_gff_1_SFF_5_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S00reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S00reg_gff_1_SFF_5_MUXInst_X), .Z0_t (stateArray_S00reg_gff_1_SFF_5_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S00reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (stateArray_S00reg_gff_1_SFF_5_MUXInst_Y), .B0_t (stateArray_outS01ser[5]), .Z0_t (port_out[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S00reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS01ser[6]), .B0_t (port_out[6]), .Z0_t (stateArray_S00reg_gff_1_SFF_6_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S00reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S00reg_gff_1_SFF_6_MUXInst_X), .Z0_t (stateArray_S00reg_gff_1_SFF_6_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S00reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (stateArray_S00reg_gff_1_SFF_6_MUXInst_Y), .B0_t (stateArray_outS01ser[6]), .Z0_t (port_out[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S00reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS01ser[7]), .B0_t (port_out[7]), .Z0_t (stateArray_S00reg_gff_1_SFF_7_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S00reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S00reg_gff_1_SFF_7_MUXInst_X), .Z0_t (stateArray_S00reg_gff_1_SFF_7_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S00reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (stateArray_S00reg_gff_1_SFF_7_MUXInst_Y), .B0_t (stateArray_outS01ser[7]), .Z0_t (port_out[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S01reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS02ser[0]), .B0_t (stateArray_outS01ser[0]), .Z0_t (stateArray_S01reg_gff_1_SFF_0_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S01reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S01reg_gff_1_SFF_0_MUXInst_X), .Z0_t (stateArray_S01reg_gff_1_SFF_0_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S01reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (stateArray_S01reg_gff_1_SFF_0_MUXInst_Y), .B0_t (stateArray_outS02ser[0]), .Z0_t (stateArray_outS01ser[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S01reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS02ser[1]), .B0_t (stateArray_outS01ser[1]), .Z0_t (stateArray_S01reg_gff_1_SFF_1_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S01reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S01reg_gff_1_SFF_1_MUXInst_X), .Z0_t (stateArray_S01reg_gff_1_SFF_1_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S01reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (stateArray_S01reg_gff_1_SFF_1_MUXInst_Y), .B0_t (stateArray_outS02ser[1]), .Z0_t (stateArray_outS01ser[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S01reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS02ser[2]), .B0_t (stateArray_outS01ser[2]), .Z0_t (stateArray_S01reg_gff_1_SFF_2_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S01reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S01reg_gff_1_SFF_2_MUXInst_X), .Z0_t (stateArray_S01reg_gff_1_SFF_2_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S01reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (stateArray_S01reg_gff_1_SFF_2_MUXInst_Y), .B0_t (stateArray_outS02ser[2]), .Z0_t (stateArray_outS01ser[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S01reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS02ser[3]), .B0_t (stateArray_outS01ser[3]), .Z0_t (stateArray_S01reg_gff_1_SFF_3_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S01reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S01reg_gff_1_SFF_3_MUXInst_X), .Z0_t (stateArray_S01reg_gff_1_SFF_3_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S01reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (stateArray_S01reg_gff_1_SFF_3_MUXInst_Y), .B0_t (stateArray_outS02ser[3]), .Z0_t (stateArray_outS01ser[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S01reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS02ser[4]), .B0_t (stateArray_outS01ser[4]), .Z0_t (stateArray_S01reg_gff_1_SFF_4_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S01reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S01reg_gff_1_SFF_4_MUXInst_X), .Z0_t (stateArray_S01reg_gff_1_SFF_4_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S01reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (stateArray_S01reg_gff_1_SFF_4_MUXInst_Y), .B0_t (stateArray_outS02ser[4]), .Z0_t (stateArray_outS01ser[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S01reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS02ser[5]), .B0_t (stateArray_outS01ser[5]), .Z0_t (stateArray_S01reg_gff_1_SFF_5_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S01reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S01reg_gff_1_SFF_5_MUXInst_X), .Z0_t (stateArray_S01reg_gff_1_SFF_5_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S01reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (stateArray_S01reg_gff_1_SFF_5_MUXInst_Y), .B0_t (stateArray_outS02ser[5]), .Z0_t (stateArray_outS01ser[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S01reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS02ser[6]), .B0_t (stateArray_outS01ser[6]), .Z0_t (stateArray_S01reg_gff_1_SFF_6_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S01reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S01reg_gff_1_SFF_6_MUXInst_X), .Z0_t (stateArray_S01reg_gff_1_SFF_6_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S01reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (stateArray_S01reg_gff_1_SFF_6_MUXInst_Y), .B0_t (stateArray_outS02ser[6]), .Z0_t (stateArray_outS01ser[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S01reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS02ser[7]), .B0_t (stateArray_outS01ser[7]), .Z0_t (stateArray_S01reg_gff_1_SFF_7_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S01reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S01reg_gff_1_SFF_7_MUXInst_X), .Z0_t (stateArray_S01reg_gff_1_SFF_7_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S01reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (stateArray_S01reg_gff_1_SFF_7_MUXInst_Y), .B0_t (stateArray_outS02ser[7]), .Z0_t (stateArray_outS01ser[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S02reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS03ser[0]), .B0_t (stateArray_outS02ser[0]), .Z0_t (stateArray_S02reg_gff_1_SFF_0_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S02reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S02reg_gff_1_SFF_0_MUXInst_X), .Z0_t (stateArray_S02reg_gff_1_SFF_0_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S02reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (stateArray_S02reg_gff_1_SFF_0_MUXInst_Y), .B0_t (stateArray_outS03ser[0]), .Z0_t (stateArray_outS02ser[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S02reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS03ser[1]), .B0_t (stateArray_outS02ser[1]), .Z0_t (stateArray_S02reg_gff_1_SFF_1_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S02reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S02reg_gff_1_SFF_1_MUXInst_X), .Z0_t (stateArray_S02reg_gff_1_SFF_1_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S02reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (stateArray_S02reg_gff_1_SFF_1_MUXInst_Y), .B0_t (stateArray_outS03ser[1]), .Z0_t (stateArray_outS02ser[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S02reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS03ser[2]), .B0_t (stateArray_outS02ser[2]), .Z0_t (stateArray_S02reg_gff_1_SFF_2_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S02reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S02reg_gff_1_SFF_2_MUXInst_X), .Z0_t (stateArray_S02reg_gff_1_SFF_2_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S02reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (stateArray_S02reg_gff_1_SFF_2_MUXInst_Y), .B0_t (stateArray_outS03ser[2]), .Z0_t (stateArray_outS02ser[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S02reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS03ser[3]), .B0_t (stateArray_outS02ser[3]), .Z0_t (stateArray_S02reg_gff_1_SFF_3_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S02reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S02reg_gff_1_SFF_3_MUXInst_X), .Z0_t (stateArray_S02reg_gff_1_SFF_3_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S02reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (stateArray_S02reg_gff_1_SFF_3_MUXInst_Y), .B0_t (stateArray_outS03ser[3]), .Z0_t (stateArray_outS02ser[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S02reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS03ser[4]), .B0_t (stateArray_outS02ser[4]), .Z0_t (stateArray_S02reg_gff_1_SFF_4_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S02reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S02reg_gff_1_SFF_4_MUXInst_X), .Z0_t (stateArray_S02reg_gff_1_SFF_4_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S02reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (stateArray_S02reg_gff_1_SFF_4_MUXInst_Y), .B0_t (stateArray_outS03ser[4]), .Z0_t (stateArray_outS02ser[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S02reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS03ser[5]), .B0_t (stateArray_outS02ser[5]), .Z0_t (stateArray_S02reg_gff_1_SFF_5_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S02reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S02reg_gff_1_SFF_5_MUXInst_X), .Z0_t (stateArray_S02reg_gff_1_SFF_5_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S02reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (stateArray_S02reg_gff_1_SFF_5_MUXInst_Y), .B0_t (stateArray_outS03ser[5]), .Z0_t (stateArray_outS02ser[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S02reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS03ser[6]), .B0_t (stateArray_outS02ser[6]), .Z0_t (stateArray_S02reg_gff_1_SFF_6_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S02reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S02reg_gff_1_SFF_6_MUXInst_X), .Z0_t (stateArray_S02reg_gff_1_SFF_6_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S02reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (stateArray_S02reg_gff_1_SFF_6_MUXInst_Y), .B0_t (stateArray_outS03ser[6]), .Z0_t (stateArray_outS02ser[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S02reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS03ser[7]), .B0_t (stateArray_outS02ser[7]), .Z0_t (stateArray_S02reg_gff_1_SFF_7_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S02reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S02reg_gff_1_SFF_7_MUXInst_X), .Z0_t (stateArray_S02reg_gff_1_SFF_7_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S02reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (stateArray_S02reg_gff_1_SFF_7_MUXInst_Y), .B0_t (stateArray_outS03ser[7]), .Z0_t (stateArray_outS02ser[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S03reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS03ser[0]), .B0_t (stateArray_outS03ser[0]), .Z0_t (stateArray_S03reg_gff_1_SFF_0_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S03reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S03reg_gff_1_SFF_0_MUXInst_X), .Z0_t (stateArray_S03reg_gff_1_SFF_0_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S03reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (stateArray_S03reg_gff_1_SFF_0_MUXInst_Y), .B0_t (stateArray_inS03ser[0]), .Z0_t (stateArray_outS03ser[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S03reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS03ser[1]), .B0_t (stateArray_outS03ser[1]), .Z0_t (stateArray_S03reg_gff_1_SFF_1_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S03reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S03reg_gff_1_SFF_1_MUXInst_X), .Z0_t (stateArray_S03reg_gff_1_SFF_1_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S03reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (stateArray_S03reg_gff_1_SFF_1_MUXInst_Y), .B0_t (stateArray_inS03ser[1]), .Z0_t (stateArray_outS03ser[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S03reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS03ser[2]), .B0_t (stateArray_outS03ser[2]), .Z0_t (stateArray_S03reg_gff_1_SFF_2_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S03reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S03reg_gff_1_SFF_2_MUXInst_X), .Z0_t (stateArray_S03reg_gff_1_SFF_2_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S03reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (stateArray_S03reg_gff_1_SFF_2_MUXInst_Y), .B0_t (stateArray_inS03ser[2]), .Z0_t (stateArray_outS03ser[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S03reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS03ser[3]), .B0_t (stateArray_outS03ser[3]), .Z0_t (stateArray_S03reg_gff_1_SFF_3_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S03reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S03reg_gff_1_SFF_3_MUXInst_X), .Z0_t (stateArray_S03reg_gff_1_SFF_3_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S03reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (stateArray_S03reg_gff_1_SFF_3_MUXInst_Y), .B0_t (stateArray_inS03ser[3]), .Z0_t (stateArray_outS03ser[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S03reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS03ser[4]), .B0_t (stateArray_outS03ser[4]), .Z0_t (stateArray_S03reg_gff_1_SFF_4_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S03reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S03reg_gff_1_SFF_4_MUXInst_X), .Z0_t (stateArray_S03reg_gff_1_SFF_4_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S03reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (stateArray_S03reg_gff_1_SFF_4_MUXInst_Y), .B0_t (stateArray_inS03ser[4]), .Z0_t (stateArray_outS03ser[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S03reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS03ser[5]), .B0_t (stateArray_outS03ser[5]), .Z0_t (stateArray_S03reg_gff_1_SFF_5_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S03reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S03reg_gff_1_SFF_5_MUXInst_X), .Z0_t (stateArray_S03reg_gff_1_SFF_5_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S03reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (stateArray_S03reg_gff_1_SFF_5_MUXInst_Y), .B0_t (stateArray_inS03ser[5]), .Z0_t (stateArray_outS03ser[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S03reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS03ser[6]), .B0_t (stateArray_outS03ser[6]), .Z0_t (stateArray_S03reg_gff_1_SFF_6_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S03reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S03reg_gff_1_SFF_6_MUXInst_X), .Z0_t (stateArray_S03reg_gff_1_SFF_6_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S03reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (stateArray_S03reg_gff_1_SFF_6_MUXInst_Y), .B0_t (stateArray_inS03ser[6]), .Z0_t (stateArray_outS03ser[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S03reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS03ser[7]), .B0_t (stateArray_outS03ser[7]), .Z0_t (stateArray_S03reg_gff_1_SFF_7_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S03reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S03reg_gff_1_SFF_7_MUXInst_X), .Z0_t (stateArray_S03reg_gff_1_SFF_7_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S03reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (stateArray_S03reg_gff_1_SFF_7_MUXInst_Y), .B0_t (stateArray_inS03ser[7]), .Z0_t (stateArray_outS03ser[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S10reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS11ser[0]), .B0_t (stateArray_outS11ser[0]), .Z0_t (stateArray_S10reg_gff_1_SFF_0_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S10reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S10reg_gff_1_SFF_0_MUXInst_X), .Z0_t (stateArray_S10reg_gff_1_SFF_0_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S10reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (stateArray_S10reg_gff_1_SFF_0_MUXInst_Y), .B0_t (stateArray_outS11ser[0]), .Z0_t (MCin[16]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S10reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS11ser[1]), .B0_t (stateArray_outS11ser[1]), .Z0_t (stateArray_S10reg_gff_1_SFF_1_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S10reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S10reg_gff_1_SFF_1_MUXInst_X), .Z0_t (stateArray_S10reg_gff_1_SFF_1_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S10reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (stateArray_S10reg_gff_1_SFF_1_MUXInst_Y), .B0_t (stateArray_outS11ser[1]), .Z0_t (MixColumns_line1_S02[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S10reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS11ser[2]), .B0_t (stateArray_outS11ser[2]), .Z0_t (stateArray_S10reg_gff_1_SFF_2_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S10reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S10reg_gff_1_SFF_2_MUXInst_X), .Z0_t (stateArray_S10reg_gff_1_SFF_2_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S10reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (stateArray_S10reg_gff_1_SFF_2_MUXInst_Y), .B0_t (stateArray_outS11ser[2]), .Z0_t (MCin[18]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S10reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS11ser[3]), .B0_t (stateArray_outS11ser[3]), .Z0_t (stateArray_S10reg_gff_1_SFF_3_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S10reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S10reg_gff_1_SFF_3_MUXInst_X), .Z0_t (stateArray_S10reg_gff_1_SFF_3_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S10reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (stateArray_S10reg_gff_1_SFF_3_MUXInst_Y), .B0_t (stateArray_outS11ser[3]), .Z0_t (MCin[19]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S10reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS11ser[4]), .B0_t (stateArray_outS11ser[4]), .Z0_t (stateArray_S10reg_gff_1_SFF_4_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S10reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S10reg_gff_1_SFF_4_MUXInst_X), .Z0_t (stateArray_S10reg_gff_1_SFF_4_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S10reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (stateArray_S10reg_gff_1_SFF_4_MUXInst_Y), .B0_t (stateArray_outS11ser[4]), .Z0_t (MixColumns_line1_S02[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S10reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS11ser[5]), .B0_t (stateArray_outS11ser[5]), .Z0_t (stateArray_S10reg_gff_1_SFF_5_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S10reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S10reg_gff_1_SFF_5_MUXInst_X), .Z0_t (stateArray_S10reg_gff_1_SFF_5_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S10reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (stateArray_S10reg_gff_1_SFF_5_MUXInst_Y), .B0_t (stateArray_outS11ser[5]), .Z0_t (MixColumns_line1_S02[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S10reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS11ser[6]), .B0_t (stateArray_outS11ser[6]), .Z0_t (stateArray_S10reg_gff_1_SFF_6_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S10reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S10reg_gff_1_SFF_6_MUXInst_X), .Z0_t (stateArray_S10reg_gff_1_SFF_6_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S10reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (stateArray_S10reg_gff_1_SFF_6_MUXInst_Y), .B0_t (stateArray_outS11ser[6]), .Z0_t (MixColumns_line1_S02[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S10reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS11ser[7]), .B0_t (stateArray_outS11ser[7]), .Z0_t (stateArray_S10reg_gff_1_SFF_7_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S10reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S10reg_gff_1_SFF_7_MUXInst_X), .Z0_t (stateArray_S10reg_gff_1_SFF_7_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S10reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (stateArray_S10reg_gff_1_SFF_7_MUXInst_Y), .B0_t (stateArray_outS11ser[7]), .Z0_t (MixColumns_line1_S02[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S11reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS12ser[0]), .B0_t (stateArray_outS12ser[0]), .Z0_t (stateArray_S11reg_gff_1_SFF_0_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S11reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S11reg_gff_1_SFF_0_MUXInst_X), .Z0_t (stateArray_S11reg_gff_1_SFF_0_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S11reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (stateArray_S11reg_gff_1_SFF_0_MUXInst_Y), .B0_t (stateArray_outS12ser[0]), .Z0_t (stateArray_outS11ser[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S11reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS12ser[1]), .B0_t (stateArray_outS12ser[1]), .Z0_t (stateArray_S11reg_gff_1_SFF_1_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S11reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S11reg_gff_1_SFF_1_MUXInst_X), .Z0_t (stateArray_S11reg_gff_1_SFF_1_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S11reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (stateArray_S11reg_gff_1_SFF_1_MUXInst_Y), .B0_t (stateArray_outS12ser[1]), .Z0_t (stateArray_outS11ser[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S11reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS12ser[2]), .B0_t (stateArray_outS12ser[2]), .Z0_t (stateArray_S11reg_gff_1_SFF_2_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S11reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S11reg_gff_1_SFF_2_MUXInst_X), .Z0_t (stateArray_S11reg_gff_1_SFF_2_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S11reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (stateArray_S11reg_gff_1_SFF_2_MUXInst_Y), .B0_t (stateArray_outS12ser[2]), .Z0_t (stateArray_outS11ser[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S11reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS12ser[3]), .B0_t (stateArray_outS12ser[3]), .Z0_t (stateArray_S11reg_gff_1_SFF_3_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S11reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S11reg_gff_1_SFF_3_MUXInst_X), .Z0_t (stateArray_S11reg_gff_1_SFF_3_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S11reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (stateArray_S11reg_gff_1_SFF_3_MUXInst_Y), .B0_t (stateArray_outS12ser[3]), .Z0_t (stateArray_outS11ser[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S11reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS12ser[4]), .B0_t (stateArray_outS12ser[4]), .Z0_t (stateArray_S11reg_gff_1_SFF_4_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S11reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S11reg_gff_1_SFF_4_MUXInst_X), .Z0_t (stateArray_S11reg_gff_1_SFF_4_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S11reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (stateArray_S11reg_gff_1_SFF_4_MUXInst_Y), .B0_t (stateArray_outS12ser[4]), .Z0_t (stateArray_outS11ser[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S11reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS12ser[5]), .B0_t (stateArray_outS12ser[5]), .Z0_t (stateArray_S11reg_gff_1_SFF_5_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S11reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S11reg_gff_1_SFF_5_MUXInst_X), .Z0_t (stateArray_S11reg_gff_1_SFF_5_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S11reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (stateArray_S11reg_gff_1_SFF_5_MUXInst_Y), .B0_t (stateArray_outS12ser[5]), .Z0_t (stateArray_outS11ser[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S11reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS12ser[6]), .B0_t (stateArray_outS12ser[6]), .Z0_t (stateArray_S11reg_gff_1_SFF_6_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S11reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S11reg_gff_1_SFF_6_MUXInst_X), .Z0_t (stateArray_S11reg_gff_1_SFF_6_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S11reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (stateArray_S11reg_gff_1_SFF_6_MUXInst_Y), .B0_t (stateArray_outS12ser[6]), .Z0_t (stateArray_outS11ser[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S11reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS12ser[7]), .B0_t (stateArray_outS12ser[7]), .Z0_t (stateArray_S11reg_gff_1_SFF_7_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S11reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S11reg_gff_1_SFF_7_MUXInst_X), .Z0_t (stateArray_S11reg_gff_1_SFF_7_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S11reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (stateArray_S11reg_gff_1_SFF_7_MUXInst_Y), .B0_t (stateArray_outS12ser[7]), .Z0_t (stateArray_outS11ser[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S12reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS13ser[0]), .B0_t (stateArray_outS13ser[0]), .Z0_t (stateArray_S12reg_gff_1_SFF_0_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S12reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S12reg_gff_1_SFF_0_MUXInst_X), .Z0_t (stateArray_S12reg_gff_1_SFF_0_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S12reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (stateArray_S12reg_gff_1_SFF_0_MUXInst_Y), .B0_t (stateArray_outS13ser[0]), .Z0_t (stateArray_outS12ser[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S12reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS13ser[1]), .B0_t (stateArray_outS13ser[1]), .Z0_t (stateArray_S12reg_gff_1_SFF_1_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S12reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S12reg_gff_1_SFF_1_MUXInst_X), .Z0_t (stateArray_S12reg_gff_1_SFF_1_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S12reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (stateArray_S12reg_gff_1_SFF_1_MUXInst_Y), .B0_t (stateArray_outS13ser[1]), .Z0_t (stateArray_outS12ser[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S12reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS13ser[2]), .B0_t (stateArray_outS13ser[2]), .Z0_t (stateArray_S12reg_gff_1_SFF_2_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S12reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S12reg_gff_1_SFF_2_MUXInst_X), .Z0_t (stateArray_S12reg_gff_1_SFF_2_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S12reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (stateArray_S12reg_gff_1_SFF_2_MUXInst_Y), .B0_t (stateArray_outS13ser[2]), .Z0_t (stateArray_outS12ser[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S12reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS13ser[3]), .B0_t (stateArray_outS13ser[3]), .Z0_t (stateArray_S12reg_gff_1_SFF_3_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S12reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S12reg_gff_1_SFF_3_MUXInst_X), .Z0_t (stateArray_S12reg_gff_1_SFF_3_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S12reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (stateArray_S12reg_gff_1_SFF_3_MUXInst_Y), .B0_t (stateArray_outS13ser[3]), .Z0_t (stateArray_outS12ser[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S12reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS13ser[4]), .B0_t (stateArray_outS13ser[4]), .Z0_t (stateArray_S12reg_gff_1_SFF_4_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S12reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S12reg_gff_1_SFF_4_MUXInst_X), .Z0_t (stateArray_S12reg_gff_1_SFF_4_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S12reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (stateArray_S12reg_gff_1_SFF_4_MUXInst_Y), .B0_t (stateArray_outS13ser[4]), .Z0_t (stateArray_outS12ser[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S12reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS13ser[5]), .B0_t (stateArray_outS13ser[5]), .Z0_t (stateArray_S12reg_gff_1_SFF_5_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S12reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S12reg_gff_1_SFF_5_MUXInst_X), .Z0_t (stateArray_S12reg_gff_1_SFF_5_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S12reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (stateArray_S12reg_gff_1_SFF_5_MUXInst_Y), .B0_t (stateArray_outS13ser[5]), .Z0_t (stateArray_outS12ser[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S12reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS13ser[6]), .B0_t (stateArray_outS13ser[6]), .Z0_t (stateArray_S12reg_gff_1_SFF_6_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S12reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S12reg_gff_1_SFF_6_MUXInst_X), .Z0_t (stateArray_S12reg_gff_1_SFF_6_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S12reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (stateArray_S12reg_gff_1_SFF_6_MUXInst_Y), .B0_t (stateArray_outS13ser[6]), .Z0_t (stateArray_outS12ser[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S12reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS13ser[7]), .B0_t (stateArray_outS13ser[7]), .Z0_t (stateArray_S12reg_gff_1_SFF_7_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S12reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S12reg_gff_1_SFF_7_MUXInst_X), .Z0_t (stateArray_S12reg_gff_1_SFF_7_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S12reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (stateArray_S12reg_gff_1_SFF_7_MUXInst_Y), .B0_t (stateArray_outS13ser[7]), .Z0_t (stateArray_outS12ser[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S13reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS13ser[0]), .B0_t (MCin[16]), .Z0_t (stateArray_S13reg_gff_1_SFF_0_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S13reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S13reg_gff_1_SFF_0_MUXInst_X), .Z0_t (stateArray_S13reg_gff_1_SFF_0_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S13reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (stateArray_S13reg_gff_1_SFF_0_MUXInst_Y), .B0_t (stateArray_inS13ser[0]), .Z0_t (stateArray_outS13ser[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S13reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS13ser[1]), .B0_t (MixColumns_line1_S02[2]), .Z0_t (stateArray_S13reg_gff_1_SFF_1_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S13reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S13reg_gff_1_SFF_1_MUXInst_X), .Z0_t (stateArray_S13reg_gff_1_SFF_1_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S13reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (stateArray_S13reg_gff_1_SFF_1_MUXInst_Y), .B0_t (stateArray_inS13ser[1]), .Z0_t (stateArray_outS13ser[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S13reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS13ser[2]), .B0_t (MCin[18]), .Z0_t (stateArray_S13reg_gff_1_SFF_2_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S13reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S13reg_gff_1_SFF_2_MUXInst_X), .Z0_t (stateArray_S13reg_gff_1_SFF_2_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S13reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (stateArray_S13reg_gff_1_SFF_2_MUXInst_Y), .B0_t (stateArray_inS13ser[2]), .Z0_t (stateArray_outS13ser[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S13reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS13ser[3]), .B0_t (MCin[19]), .Z0_t (stateArray_S13reg_gff_1_SFF_3_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S13reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S13reg_gff_1_SFF_3_MUXInst_X), .Z0_t (stateArray_S13reg_gff_1_SFF_3_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S13reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (stateArray_S13reg_gff_1_SFF_3_MUXInst_Y), .B0_t (stateArray_inS13ser[3]), .Z0_t (stateArray_outS13ser[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S13reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS13ser[4]), .B0_t (MixColumns_line1_S02[5]), .Z0_t (stateArray_S13reg_gff_1_SFF_4_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S13reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S13reg_gff_1_SFF_4_MUXInst_X), .Z0_t (stateArray_S13reg_gff_1_SFF_4_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S13reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (stateArray_S13reg_gff_1_SFF_4_MUXInst_Y), .B0_t (stateArray_inS13ser[4]), .Z0_t (stateArray_outS13ser[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S13reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS13ser[5]), .B0_t (MixColumns_line1_S02[6]), .Z0_t (stateArray_S13reg_gff_1_SFF_5_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S13reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S13reg_gff_1_SFF_5_MUXInst_X), .Z0_t (stateArray_S13reg_gff_1_SFF_5_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S13reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (stateArray_S13reg_gff_1_SFF_5_MUXInst_Y), .B0_t (stateArray_inS13ser[5]), .Z0_t (stateArray_outS13ser[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S13reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS13ser[6]), .B0_t (MixColumns_line1_S02[7]), .Z0_t (stateArray_S13reg_gff_1_SFF_6_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S13reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S13reg_gff_1_SFF_6_MUXInst_X), .Z0_t (stateArray_S13reg_gff_1_SFF_6_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S13reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (stateArray_S13reg_gff_1_SFF_6_MUXInst_Y), .B0_t (stateArray_inS13ser[6]), .Z0_t (stateArray_outS13ser[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S13reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS13ser[7]), .B0_t (MixColumns_line1_S02[0]), .Z0_t (stateArray_S13reg_gff_1_SFF_7_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S13reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S13reg_gff_1_SFF_7_MUXInst_X), .Z0_t (stateArray_S13reg_gff_1_SFF_7_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S13reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (stateArray_S13reg_gff_1_SFF_7_MUXInst_Y), .B0_t (stateArray_inS13ser[7]), .Z0_t (stateArray_outS13ser[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S20reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS21ser[0]), .B0_t (stateArray_outS22ser[0]), .Z0_t (stateArray_S20reg_gff_1_SFF_0_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S20reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S20reg_gff_1_SFF_0_MUXInst_X), .Z0_t (stateArray_S20reg_gff_1_SFF_0_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S20reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (stateArray_S20reg_gff_1_SFF_0_MUXInst_Y), .B0_t (stateArray_outS21ser[0]), .Z0_t (MCin[8]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S20reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS21ser[1]), .B0_t (stateArray_outS22ser[1]), .Z0_t (stateArray_S20reg_gff_1_SFF_1_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S20reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S20reg_gff_1_SFF_1_MUXInst_X), .Z0_t (stateArray_S20reg_gff_1_SFF_1_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S20reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (stateArray_S20reg_gff_1_SFF_1_MUXInst_Y), .B0_t (stateArray_outS21ser[1]), .Z0_t (MixColumns_line2_S02[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S20reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS21ser[2]), .B0_t (stateArray_outS22ser[2]), .Z0_t (stateArray_S20reg_gff_1_SFF_2_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S20reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S20reg_gff_1_SFF_2_MUXInst_X), .Z0_t (stateArray_S20reg_gff_1_SFF_2_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S20reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (stateArray_S20reg_gff_1_SFF_2_MUXInst_Y), .B0_t (stateArray_outS21ser[2]), .Z0_t (MCin[10]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S20reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS21ser[3]), .B0_t (stateArray_outS22ser[3]), .Z0_t (stateArray_S20reg_gff_1_SFF_3_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S20reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S20reg_gff_1_SFF_3_MUXInst_X), .Z0_t (stateArray_S20reg_gff_1_SFF_3_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S20reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (stateArray_S20reg_gff_1_SFF_3_MUXInst_Y), .B0_t (stateArray_outS21ser[3]), .Z0_t (MCin[11]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S20reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS21ser[4]), .B0_t (stateArray_outS22ser[4]), .Z0_t (stateArray_S20reg_gff_1_SFF_4_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S20reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S20reg_gff_1_SFF_4_MUXInst_X), .Z0_t (stateArray_S20reg_gff_1_SFF_4_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S20reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (stateArray_S20reg_gff_1_SFF_4_MUXInst_Y), .B0_t (stateArray_outS21ser[4]), .Z0_t (MixColumns_line2_S02[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S20reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS21ser[5]), .B0_t (stateArray_outS22ser[5]), .Z0_t (stateArray_S20reg_gff_1_SFF_5_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S20reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S20reg_gff_1_SFF_5_MUXInst_X), .Z0_t (stateArray_S20reg_gff_1_SFF_5_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S20reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (stateArray_S20reg_gff_1_SFF_5_MUXInst_Y), .B0_t (stateArray_outS21ser[5]), .Z0_t (MixColumns_line2_S02[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S20reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS21ser[6]), .B0_t (stateArray_outS22ser[6]), .Z0_t (stateArray_S20reg_gff_1_SFF_6_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S20reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S20reg_gff_1_SFF_6_MUXInst_X), .Z0_t (stateArray_S20reg_gff_1_SFF_6_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S20reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (stateArray_S20reg_gff_1_SFF_6_MUXInst_Y), .B0_t (stateArray_outS21ser[6]), .Z0_t (MixColumns_line2_S02[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S20reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS21ser[7]), .B0_t (stateArray_outS22ser[7]), .Z0_t (stateArray_S20reg_gff_1_SFF_7_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S20reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S20reg_gff_1_SFF_7_MUXInst_X), .Z0_t (stateArray_S20reg_gff_1_SFF_7_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S20reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (stateArray_S20reg_gff_1_SFF_7_MUXInst_Y), .B0_t (stateArray_outS21ser[7]), .Z0_t (MixColumns_line2_S02[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S21reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS22ser[0]), .B0_t (stateArray_outS23ser[0]), .Z0_t (stateArray_S21reg_gff_1_SFF_0_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S21reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S21reg_gff_1_SFF_0_MUXInst_X), .Z0_t (stateArray_S21reg_gff_1_SFF_0_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S21reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (stateArray_S21reg_gff_1_SFF_0_MUXInst_Y), .B0_t (stateArray_outS22ser[0]), .Z0_t (stateArray_outS21ser[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S21reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS22ser[1]), .B0_t (stateArray_outS23ser[1]), .Z0_t (stateArray_S21reg_gff_1_SFF_1_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S21reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S21reg_gff_1_SFF_1_MUXInst_X), .Z0_t (stateArray_S21reg_gff_1_SFF_1_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S21reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (stateArray_S21reg_gff_1_SFF_1_MUXInst_Y), .B0_t (stateArray_outS22ser[1]), .Z0_t (stateArray_outS21ser[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S21reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS22ser[2]), .B0_t (stateArray_outS23ser[2]), .Z0_t (stateArray_S21reg_gff_1_SFF_2_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S21reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S21reg_gff_1_SFF_2_MUXInst_X), .Z0_t (stateArray_S21reg_gff_1_SFF_2_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S21reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (stateArray_S21reg_gff_1_SFF_2_MUXInst_Y), .B0_t (stateArray_outS22ser[2]), .Z0_t (stateArray_outS21ser[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S21reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS22ser[3]), .B0_t (stateArray_outS23ser[3]), .Z0_t (stateArray_S21reg_gff_1_SFF_3_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S21reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S21reg_gff_1_SFF_3_MUXInst_X), .Z0_t (stateArray_S21reg_gff_1_SFF_3_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S21reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (stateArray_S21reg_gff_1_SFF_3_MUXInst_Y), .B0_t (stateArray_outS22ser[3]), .Z0_t (stateArray_outS21ser[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S21reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS22ser[4]), .B0_t (stateArray_outS23ser[4]), .Z0_t (stateArray_S21reg_gff_1_SFF_4_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S21reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S21reg_gff_1_SFF_4_MUXInst_X), .Z0_t (stateArray_S21reg_gff_1_SFF_4_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S21reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (stateArray_S21reg_gff_1_SFF_4_MUXInst_Y), .B0_t (stateArray_outS22ser[4]), .Z0_t (stateArray_outS21ser[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S21reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS22ser[5]), .B0_t (stateArray_outS23ser[5]), .Z0_t (stateArray_S21reg_gff_1_SFF_5_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S21reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S21reg_gff_1_SFF_5_MUXInst_X), .Z0_t (stateArray_S21reg_gff_1_SFF_5_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S21reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (stateArray_S21reg_gff_1_SFF_5_MUXInst_Y), .B0_t (stateArray_outS22ser[5]), .Z0_t (stateArray_outS21ser[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S21reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS22ser[6]), .B0_t (stateArray_outS23ser[6]), .Z0_t (stateArray_S21reg_gff_1_SFF_6_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S21reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S21reg_gff_1_SFF_6_MUXInst_X), .Z0_t (stateArray_S21reg_gff_1_SFF_6_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S21reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (stateArray_S21reg_gff_1_SFF_6_MUXInst_Y), .B0_t (stateArray_outS22ser[6]), .Z0_t (stateArray_outS21ser[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S21reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS22ser[7]), .B0_t (stateArray_outS23ser[7]), .Z0_t (stateArray_S21reg_gff_1_SFF_7_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S21reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S21reg_gff_1_SFF_7_MUXInst_X), .Z0_t (stateArray_S21reg_gff_1_SFF_7_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S21reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (stateArray_S21reg_gff_1_SFF_7_MUXInst_Y), .B0_t (stateArray_outS22ser[7]), .Z0_t (stateArray_outS21ser[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S22reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS23ser[0]), .B0_t (MCin[8]), .Z0_t (stateArray_S22reg_gff_1_SFF_0_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S22reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S22reg_gff_1_SFF_0_MUXInst_X), .Z0_t (stateArray_S22reg_gff_1_SFF_0_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S22reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (stateArray_S22reg_gff_1_SFF_0_MUXInst_Y), .B0_t (stateArray_outS23ser[0]), .Z0_t (stateArray_outS22ser[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S22reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS23ser[1]), .B0_t (MixColumns_line2_S02[2]), .Z0_t (stateArray_S22reg_gff_1_SFF_1_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S22reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S22reg_gff_1_SFF_1_MUXInst_X), .Z0_t (stateArray_S22reg_gff_1_SFF_1_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S22reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (stateArray_S22reg_gff_1_SFF_1_MUXInst_Y), .B0_t (stateArray_outS23ser[1]), .Z0_t (stateArray_outS22ser[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S22reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS23ser[2]), .B0_t (MCin[10]), .Z0_t (stateArray_S22reg_gff_1_SFF_2_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S22reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S22reg_gff_1_SFF_2_MUXInst_X), .Z0_t (stateArray_S22reg_gff_1_SFF_2_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S22reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (stateArray_S22reg_gff_1_SFF_2_MUXInst_Y), .B0_t (stateArray_outS23ser[2]), .Z0_t (stateArray_outS22ser[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S22reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS23ser[3]), .B0_t (MCin[11]), .Z0_t (stateArray_S22reg_gff_1_SFF_3_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S22reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S22reg_gff_1_SFF_3_MUXInst_X), .Z0_t (stateArray_S22reg_gff_1_SFF_3_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S22reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (stateArray_S22reg_gff_1_SFF_3_MUXInst_Y), .B0_t (stateArray_outS23ser[3]), .Z0_t (stateArray_outS22ser[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S22reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS23ser[4]), .B0_t (MixColumns_line2_S02[5]), .Z0_t (stateArray_S22reg_gff_1_SFF_4_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S22reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S22reg_gff_1_SFF_4_MUXInst_X), .Z0_t (stateArray_S22reg_gff_1_SFF_4_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S22reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (stateArray_S22reg_gff_1_SFF_4_MUXInst_Y), .B0_t (stateArray_outS23ser[4]), .Z0_t (stateArray_outS22ser[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S22reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS23ser[5]), .B0_t (MixColumns_line2_S02[6]), .Z0_t (stateArray_S22reg_gff_1_SFF_5_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S22reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S22reg_gff_1_SFF_5_MUXInst_X), .Z0_t (stateArray_S22reg_gff_1_SFF_5_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S22reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (stateArray_S22reg_gff_1_SFF_5_MUXInst_Y), .B0_t (stateArray_outS23ser[5]), .Z0_t (stateArray_outS22ser[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S22reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS23ser[6]), .B0_t (MixColumns_line2_S02[7]), .Z0_t (stateArray_S22reg_gff_1_SFF_6_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S22reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S22reg_gff_1_SFF_6_MUXInst_X), .Z0_t (stateArray_S22reg_gff_1_SFF_6_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S22reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (stateArray_S22reg_gff_1_SFF_6_MUXInst_Y), .B0_t (stateArray_outS23ser[6]), .Z0_t (stateArray_outS22ser[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S22reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS23ser[7]), .B0_t (MixColumns_line2_S02[0]), .Z0_t (stateArray_S22reg_gff_1_SFF_7_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S22reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S22reg_gff_1_SFF_7_MUXInst_X), .Z0_t (stateArray_S22reg_gff_1_SFF_7_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S22reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (stateArray_S22reg_gff_1_SFF_7_MUXInst_Y), .B0_t (stateArray_outS23ser[7]), .Z0_t (stateArray_outS22ser[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S23reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS23ser[0]), .B0_t (stateArray_outS21ser[0]), .Z0_t (stateArray_S23reg_gff_1_SFF_0_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S23reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S23reg_gff_1_SFF_0_MUXInst_X), .Z0_t (stateArray_S23reg_gff_1_SFF_0_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S23reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (stateArray_S23reg_gff_1_SFF_0_MUXInst_Y), .B0_t (stateArray_inS23ser[0]), .Z0_t (stateArray_outS23ser[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S23reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS23ser[1]), .B0_t (stateArray_outS21ser[1]), .Z0_t (stateArray_S23reg_gff_1_SFF_1_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S23reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S23reg_gff_1_SFF_1_MUXInst_X), .Z0_t (stateArray_S23reg_gff_1_SFF_1_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S23reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (stateArray_S23reg_gff_1_SFF_1_MUXInst_Y), .B0_t (stateArray_inS23ser[1]), .Z0_t (stateArray_outS23ser[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S23reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS23ser[2]), .B0_t (stateArray_outS21ser[2]), .Z0_t (stateArray_S23reg_gff_1_SFF_2_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S23reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S23reg_gff_1_SFF_2_MUXInst_X), .Z0_t (stateArray_S23reg_gff_1_SFF_2_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S23reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (stateArray_S23reg_gff_1_SFF_2_MUXInst_Y), .B0_t (stateArray_inS23ser[2]), .Z0_t (stateArray_outS23ser[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S23reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS23ser[3]), .B0_t (stateArray_outS21ser[3]), .Z0_t (stateArray_S23reg_gff_1_SFF_3_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S23reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S23reg_gff_1_SFF_3_MUXInst_X), .Z0_t (stateArray_S23reg_gff_1_SFF_3_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S23reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (stateArray_S23reg_gff_1_SFF_3_MUXInst_Y), .B0_t (stateArray_inS23ser[3]), .Z0_t (stateArray_outS23ser[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S23reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS23ser[4]), .B0_t (stateArray_outS21ser[4]), .Z0_t (stateArray_S23reg_gff_1_SFF_4_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S23reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S23reg_gff_1_SFF_4_MUXInst_X), .Z0_t (stateArray_S23reg_gff_1_SFF_4_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S23reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (stateArray_S23reg_gff_1_SFF_4_MUXInst_Y), .B0_t (stateArray_inS23ser[4]), .Z0_t (stateArray_outS23ser[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S23reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS23ser[5]), .B0_t (stateArray_outS21ser[5]), .Z0_t (stateArray_S23reg_gff_1_SFF_5_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S23reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S23reg_gff_1_SFF_5_MUXInst_X), .Z0_t (stateArray_S23reg_gff_1_SFF_5_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S23reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (stateArray_S23reg_gff_1_SFF_5_MUXInst_Y), .B0_t (stateArray_inS23ser[5]), .Z0_t (stateArray_outS23ser[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S23reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS23ser[6]), .B0_t (stateArray_outS21ser[6]), .Z0_t (stateArray_S23reg_gff_1_SFF_6_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S23reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S23reg_gff_1_SFF_6_MUXInst_X), .Z0_t (stateArray_S23reg_gff_1_SFF_6_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S23reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (stateArray_S23reg_gff_1_SFF_6_MUXInst_Y), .B0_t (stateArray_inS23ser[6]), .Z0_t (stateArray_outS23ser[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S23reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS23ser[7]), .B0_t (stateArray_outS21ser[7]), .Z0_t (stateArray_S23reg_gff_1_SFF_7_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S23reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S23reg_gff_1_SFF_7_MUXInst_X), .Z0_t (stateArray_S23reg_gff_1_SFF_7_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S23reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (stateArray_S23reg_gff_1_SFF_7_MUXInst_Y), .B0_t (stateArray_inS23ser[7]), .Z0_t (stateArray_outS23ser[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S30reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS31ser[0]), .B0_t (stateArray_outS33ser[0]), .Z0_t (stateArray_S30reg_gff_1_SFF_0_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S30reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S30reg_gff_1_SFF_0_MUXInst_X), .Z0_t (stateArray_S30reg_gff_1_SFF_0_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S30reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (stateArray_S30reg_gff_1_SFF_0_MUXInst_Y), .B0_t (stateArray_outS31ser[0]), .Z0_t (MCin[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S30reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS31ser[1]), .B0_t (stateArray_outS33ser[1]), .Z0_t (stateArray_S30reg_gff_1_SFF_1_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S30reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S30reg_gff_1_SFF_1_MUXInst_X), .Z0_t (stateArray_S30reg_gff_1_SFF_1_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S30reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (stateArray_S30reg_gff_1_SFF_1_MUXInst_Y), .B0_t (stateArray_outS31ser[1]), .Z0_t (MixColumns_line3_S02[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S30reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS31ser[2]), .B0_t (stateArray_outS33ser[2]), .Z0_t (stateArray_S30reg_gff_1_SFF_2_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S30reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S30reg_gff_1_SFF_2_MUXInst_X), .Z0_t (stateArray_S30reg_gff_1_SFF_2_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S30reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (stateArray_S30reg_gff_1_SFF_2_MUXInst_Y), .B0_t (stateArray_outS31ser[2]), .Z0_t (MCin[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S30reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS31ser[3]), .B0_t (stateArray_outS33ser[3]), .Z0_t (stateArray_S30reg_gff_1_SFF_3_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S30reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S30reg_gff_1_SFF_3_MUXInst_X), .Z0_t (stateArray_S30reg_gff_1_SFF_3_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S30reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (stateArray_S30reg_gff_1_SFF_3_MUXInst_Y), .B0_t (stateArray_outS31ser[3]), .Z0_t (MCin[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S30reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS31ser[4]), .B0_t (stateArray_outS33ser[4]), .Z0_t (stateArray_S30reg_gff_1_SFF_4_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S30reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S30reg_gff_1_SFF_4_MUXInst_X), .Z0_t (stateArray_S30reg_gff_1_SFF_4_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S30reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (stateArray_S30reg_gff_1_SFF_4_MUXInst_Y), .B0_t (stateArray_outS31ser[4]), .Z0_t (MixColumns_line3_S02[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S30reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS31ser[5]), .B0_t (stateArray_outS33ser[5]), .Z0_t (stateArray_S30reg_gff_1_SFF_5_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S30reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S30reg_gff_1_SFF_5_MUXInst_X), .Z0_t (stateArray_S30reg_gff_1_SFF_5_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S30reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (stateArray_S30reg_gff_1_SFF_5_MUXInst_Y), .B0_t (stateArray_outS31ser[5]), .Z0_t (MixColumns_line3_S02[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S30reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS31ser[6]), .B0_t (stateArray_outS33ser[6]), .Z0_t (stateArray_S30reg_gff_1_SFF_6_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S30reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S30reg_gff_1_SFF_6_MUXInst_X), .Z0_t (stateArray_S30reg_gff_1_SFF_6_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S30reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (stateArray_S30reg_gff_1_SFF_6_MUXInst_Y), .B0_t (stateArray_outS31ser[6]), .Z0_t (MixColumns_line3_S02[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S30reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS31ser[7]), .B0_t (stateArray_outS33ser[7]), .Z0_t (stateArray_S30reg_gff_1_SFF_7_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S30reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S30reg_gff_1_SFF_7_MUXInst_X), .Z0_t (stateArray_S30reg_gff_1_SFF_7_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S30reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (stateArray_S30reg_gff_1_SFF_7_MUXInst_Y), .B0_t (stateArray_outS31ser[7]), .Z0_t (MixColumns_line3_S02[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S31reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS32ser[0]), .B0_t (MCin[0]), .Z0_t (stateArray_S31reg_gff_1_SFF_0_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S31reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S31reg_gff_1_SFF_0_MUXInst_X), .Z0_t (stateArray_S31reg_gff_1_SFF_0_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S31reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (stateArray_S31reg_gff_1_SFF_0_MUXInst_Y), .B0_t (stateArray_outS32ser[0]), .Z0_t (stateArray_outS31ser[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S31reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS32ser[1]), .B0_t (MixColumns_line3_S02[2]), .Z0_t (stateArray_S31reg_gff_1_SFF_1_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S31reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S31reg_gff_1_SFF_1_MUXInst_X), .Z0_t (stateArray_S31reg_gff_1_SFF_1_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S31reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (stateArray_S31reg_gff_1_SFF_1_MUXInst_Y), .B0_t (stateArray_outS32ser[1]), .Z0_t (stateArray_outS31ser[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S31reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS32ser[2]), .B0_t (MCin[2]), .Z0_t (stateArray_S31reg_gff_1_SFF_2_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S31reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S31reg_gff_1_SFF_2_MUXInst_X), .Z0_t (stateArray_S31reg_gff_1_SFF_2_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S31reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (stateArray_S31reg_gff_1_SFF_2_MUXInst_Y), .B0_t (stateArray_outS32ser[2]), .Z0_t (stateArray_outS31ser[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S31reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS32ser[3]), .B0_t (MCin[3]), .Z0_t (stateArray_S31reg_gff_1_SFF_3_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S31reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S31reg_gff_1_SFF_3_MUXInst_X), .Z0_t (stateArray_S31reg_gff_1_SFF_3_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S31reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (stateArray_S31reg_gff_1_SFF_3_MUXInst_Y), .B0_t (stateArray_outS32ser[3]), .Z0_t (stateArray_outS31ser[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S31reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS32ser[4]), .B0_t (MixColumns_line3_S02[5]), .Z0_t (stateArray_S31reg_gff_1_SFF_4_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S31reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S31reg_gff_1_SFF_4_MUXInst_X), .Z0_t (stateArray_S31reg_gff_1_SFF_4_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S31reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (stateArray_S31reg_gff_1_SFF_4_MUXInst_Y), .B0_t (stateArray_outS32ser[4]), .Z0_t (stateArray_outS31ser[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S31reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS32ser[5]), .B0_t (MixColumns_line3_S02[6]), .Z0_t (stateArray_S31reg_gff_1_SFF_5_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S31reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S31reg_gff_1_SFF_5_MUXInst_X), .Z0_t (stateArray_S31reg_gff_1_SFF_5_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S31reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (stateArray_S31reg_gff_1_SFF_5_MUXInst_Y), .B0_t (stateArray_outS32ser[5]), .Z0_t (stateArray_outS31ser[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S31reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS32ser[6]), .B0_t (MixColumns_line3_S02[7]), .Z0_t (stateArray_S31reg_gff_1_SFF_6_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S31reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S31reg_gff_1_SFF_6_MUXInst_X), .Z0_t (stateArray_S31reg_gff_1_SFF_6_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S31reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (stateArray_S31reg_gff_1_SFF_6_MUXInst_Y), .B0_t (stateArray_outS32ser[6]), .Z0_t (stateArray_outS31ser[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S31reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS32ser[7]), .B0_t (MixColumns_line3_S02[0]), .Z0_t (stateArray_S31reg_gff_1_SFF_7_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S31reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S31reg_gff_1_SFF_7_MUXInst_X), .Z0_t (stateArray_S31reg_gff_1_SFF_7_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S31reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (stateArray_S31reg_gff_1_SFF_7_MUXInst_Y), .B0_t (stateArray_outS32ser[7]), .Z0_t (stateArray_outS31ser[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S32reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS33ser[0]), .B0_t (stateArray_outS31ser[0]), .Z0_t (stateArray_S32reg_gff_1_SFF_0_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S32reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S32reg_gff_1_SFF_0_MUXInst_X), .Z0_t (stateArray_S32reg_gff_1_SFF_0_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S32reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (stateArray_S32reg_gff_1_SFF_0_MUXInst_Y), .B0_t (stateArray_outS33ser[0]), .Z0_t (stateArray_outS32ser[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S32reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS33ser[1]), .B0_t (stateArray_outS31ser[1]), .Z0_t (stateArray_S32reg_gff_1_SFF_1_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S32reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S32reg_gff_1_SFF_1_MUXInst_X), .Z0_t (stateArray_S32reg_gff_1_SFF_1_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S32reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (stateArray_S32reg_gff_1_SFF_1_MUXInst_Y), .B0_t (stateArray_outS33ser[1]), .Z0_t (stateArray_outS32ser[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S32reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS33ser[2]), .B0_t (stateArray_outS31ser[2]), .Z0_t (stateArray_S32reg_gff_1_SFF_2_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S32reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S32reg_gff_1_SFF_2_MUXInst_X), .Z0_t (stateArray_S32reg_gff_1_SFF_2_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S32reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (stateArray_S32reg_gff_1_SFF_2_MUXInst_Y), .B0_t (stateArray_outS33ser[2]), .Z0_t (stateArray_outS32ser[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S32reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS33ser[3]), .B0_t (stateArray_outS31ser[3]), .Z0_t (stateArray_S32reg_gff_1_SFF_3_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S32reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S32reg_gff_1_SFF_3_MUXInst_X), .Z0_t (stateArray_S32reg_gff_1_SFF_3_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S32reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (stateArray_S32reg_gff_1_SFF_3_MUXInst_Y), .B0_t (stateArray_outS33ser[3]), .Z0_t (stateArray_outS32ser[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S32reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS33ser[4]), .B0_t (stateArray_outS31ser[4]), .Z0_t (stateArray_S32reg_gff_1_SFF_4_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S32reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S32reg_gff_1_SFF_4_MUXInst_X), .Z0_t (stateArray_S32reg_gff_1_SFF_4_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S32reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (stateArray_S32reg_gff_1_SFF_4_MUXInst_Y), .B0_t (stateArray_outS33ser[4]), .Z0_t (stateArray_outS32ser[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S32reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS33ser[5]), .B0_t (stateArray_outS31ser[5]), .Z0_t (stateArray_S32reg_gff_1_SFF_5_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S32reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S32reg_gff_1_SFF_5_MUXInst_X), .Z0_t (stateArray_S32reg_gff_1_SFF_5_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S32reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (stateArray_S32reg_gff_1_SFF_5_MUXInst_Y), .B0_t (stateArray_outS33ser[5]), .Z0_t (stateArray_outS32ser[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S32reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS33ser[6]), .B0_t (stateArray_outS31ser[6]), .Z0_t (stateArray_S32reg_gff_1_SFF_6_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S32reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S32reg_gff_1_SFF_6_MUXInst_X), .Z0_t (stateArray_S32reg_gff_1_SFF_6_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S32reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (stateArray_S32reg_gff_1_SFF_6_MUXInst_Y), .B0_t (stateArray_outS33ser[6]), .Z0_t (stateArray_outS32ser[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S32reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS33ser[7]), .B0_t (stateArray_outS31ser[7]), .Z0_t (stateArray_S32reg_gff_1_SFF_7_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S32reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S32reg_gff_1_SFF_7_MUXInst_X), .Z0_t (stateArray_S32reg_gff_1_SFF_7_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S32reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (stateArray_S32reg_gff_1_SFF_7_MUXInst_Y), .B0_t (stateArray_outS33ser[7]), .Z0_t (stateArray_outS32ser[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S33reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS33ser[0]), .B0_t (stateArray_outS32ser[0]), .Z0_t (stateArray_S33reg_gff_1_SFF_0_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S33reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S33reg_gff_1_SFF_0_MUXInst_X), .Z0_t (stateArray_S33reg_gff_1_SFF_0_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S33reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (stateArray_S33reg_gff_1_SFF_0_MUXInst_Y), .B0_t (stateArray_inS33ser[0]), .Z0_t (stateArray_outS33ser[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S33reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS33ser[1]), .B0_t (stateArray_outS32ser[1]), .Z0_t (stateArray_S33reg_gff_1_SFF_1_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S33reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S33reg_gff_1_SFF_1_MUXInst_X), .Z0_t (stateArray_S33reg_gff_1_SFF_1_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S33reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (stateArray_S33reg_gff_1_SFF_1_MUXInst_Y), .B0_t (stateArray_inS33ser[1]), .Z0_t (stateArray_outS33ser[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S33reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS33ser[2]), .B0_t (stateArray_outS32ser[2]), .Z0_t (stateArray_S33reg_gff_1_SFF_2_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S33reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S33reg_gff_1_SFF_2_MUXInst_X), .Z0_t (stateArray_S33reg_gff_1_SFF_2_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S33reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (stateArray_S33reg_gff_1_SFF_2_MUXInst_Y), .B0_t (stateArray_inS33ser[2]), .Z0_t (stateArray_outS33ser[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S33reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS33ser[3]), .B0_t (stateArray_outS32ser[3]), .Z0_t (stateArray_S33reg_gff_1_SFF_3_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S33reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S33reg_gff_1_SFF_3_MUXInst_X), .Z0_t (stateArray_S33reg_gff_1_SFF_3_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S33reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (stateArray_S33reg_gff_1_SFF_3_MUXInst_Y), .B0_t (stateArray_inS33ser[3]), .Z0_t (stateArray_outS33ser[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S33reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS33ser[4]), .B0_t (stateArray_outS32ser[4]), .Z0_t (stateArray_S33reg_gff_1_SFF_4_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S33reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S33reg_gff_1_SFF_4_MUXInst_X), .Z0_t (stateArray_S33reg_gff_1_SFF_4_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S33reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (stateArray_S33reg_gff_1_SFF_4_MUXInst_Y), .B0_t (stateArray_inS33ser[4]), .Z0_t (stateArray_outS33ser[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S33reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS33ser[5]), .B0_t (stateArray_outS32ser[5]), .Z0_t (stateArray_S33reg_gff_1_SFF_5_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S33reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S33reg_gff_1_SFF_5_MUXInst_X), .Z0_t (stateArray_S33reg_gff_1_SFF_5_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S33reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (stateArray_S33reg_gff_1_SFF_5_MUXInst_Y), .B0_t (stateArray_inS33ser[5]), .Z0_t (stateArray_outS33ser[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S33reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS33ser[6]), .B0_t (stateArray_outS32ser[6]), .Z0_t (stateArray_S33reg_gff_1_SFF_6_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S33reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S33reg_gff_1_SFF_6_MUXInst_X), .Z0_t (stateArray_S33reg_gff_1_SFF_6_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S33reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (stateArray_S33reg_gff_1_SFF_6_MUXInst_Y), .B0_t (stateArray_inS33ser[6]), .Z0_t (stateArray_outS33ser[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S33reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS33ser[7]), .B0_t (stateArray_outS32ser[7]), .Z0_t (stateArray_S33reg_gff_1_SFF_7_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S33reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (ctrl_n4), .B0_t (stateArray_S33reg_gff_1_SFF_7_MUXInst_X), .Z0_t (stateArray_S33reg_gff_1_SFF_7_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S33reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (stateArray_S33reg_gff_1_SFF_7_MUXInst_Y), .B0_t (stateArray_inS33ser[7]), .Z0_t (stateArray_outS33ser[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_0_XOR1_U1 ( .A0_t (MCin[16]), .B0_t (StateInMC[24]), .Z0_t (stateArray_MUX_inS03ser_mux_inst_0_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_0_AND1_U1 ( .A0_t (stateArray_nReset_selMC), .B0_t (stateArray_MUX_inS03ser_mux_inst_0_X), .Z0_t (stateArray_MUX_inS03ser_mux_inst_0_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_0_XOR2_U1 ( .A0_t (stateArray_MUX_inS03ser_mux_inst_0_Y), .B0_t (MCin[16]), .Z0_t (stateArray_inS03ser[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_1_XOR1_U1 ( .A0_t (MixColumns_line1_S02[2]), .B0_t (StateInMC[25]), .Z0_t (stateArray_MUX_inS03ser_mux_inst_1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_1_AND1_U1 ( .A0_t (stateArray_nReset_selMC), .B0_t (stateArray_MUX_inS03ser_mux_inst_1_X), .Z0_t (stateArray_MUX_inS03ser_mux_inst_1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_1_XOR2_U1 ( .A0_t (stateArray_MUX_inS03ser_mux_inst_1_Y), .B0_t (MixColumns_line1_S02[2]), .Z0_t (stateArray_inS03ser[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_2_XOR1_U1 ( .A0_t (MCin[18]), .B0_t (StateInMC[26]), .Z0_t (stateArray_MUX_inS03ser_mux_inst_2_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_2_AND1_U1 ( .A0_t (stateArray_nReset_selMC), .B0_t (stateArray_MUX_inS03ser_mux_inst_2_X), .Z0_t (stateArray_MUX_inS03ser_mux_inst_2_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_2_XOR2_U1 ( .A0_t (stateArray_MUX_inS03ser_mux_inst_2_Y), .B0_t (MCin[18]), .Z0_t (stateArray_inS03ser[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_3_XOR1_U1 ( .A0_t (MCin[19]), .B0_t (StateInMC[27]), .Z0_t (stateArray_MUX_inS03ser_mux_inst_3_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_3_AND1_U1 ( .A0_t (stateArray_nReset_selMC), .B0_t (stateArray_MUX_inS03ser_mux_inst_3_X), .Z0_t (stateArray_MUX_inS03ser_mux_inst_3_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_3_XOR2_U1 ( .A0_t (stateArray_MUX_inS03ser_mux_inst_3_Y), .B0_t (MCin[19]), .Z0_t (stateArray_inS03ser[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_4_XOR1_U1 ( .A0_t (MixColumns_line1_S02[5]), .B0_t (StateInMC[28]), .Z0_t (stateArray_MUX_inS03ser_mux_inst_4_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_4_AND1_U1 ( .A0_t (stateArray_nReset_selMC), .B0_t (stateArray_MUX_inS03ser_mux_inst_4_X), .Z0_t (stateArray_MUX_inS03ser_mux_inst_4_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_4_XOR2_U1 ( .A0_t (stateArray_MUX_inS03ser_mux_inst_4_Y), .B0_t (MixColumns_line1_S02[5]), .Z0_t (stateArray_inS03ser[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_5_XOR1_U1 ( .A0_t (MixColumns_line1_S02[6]), .B0_t (StateInMC[29]), .Z0_t (stateArray_MUX_inS03ser_mux_inst_5_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_5_AND1_U1 ( .A0_t (stateArray_nReset_selMC), .B0_t (stateArray_MUX_inS03ser_mux_inst_5_X), .Z0_t (stateArray_MUX_inS03ser_mux_inst_5_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_5_XOR2_U1 ( .A0_t (stateArray_MUX_inS03ser_mux_inst_5_Y), .B0_t (MixColumns_line1_S02[6]), .Z0_t (stateArray_inS03ser[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_6_XOR1_U1 ( .A0_t (MixColumns_line1_S02[7]), .B0_t (StateInMC[30]), .Z0_t (stateArray_MUX_inS03ser_mux_inst_6_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_6_AND1_U1 ( .A0_t (stateArray_nReset_selMC), .B0_t (stateArray_MUX_inS03ser_mux_inst_6_X), .Z0_t (stateArray_MUX_inS03ser_mux_inst_6_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_6_XOR2_U1 ( .A0_t (stateArray_MUX_inS03ser_mux_inst_6_Y), .B0_t (MixColumns_line1_S02[7]), .Z0_t (stateArray_inS03ser[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_7_XOR1_U1 ( .A0_t (MixColumns_line1_S02[0]), .B0_t (StateInMC[31]), .Z0_t (stateArray_MUX_inS03ser_mux_inst_7_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_7_AND1_U1 ( .A0_t (stateArray_nReset_selMC), .B0_t (stateArray_MUX_inS03ser_mux_inst_7_X), .Z0_t (stateArray_MUX_inS03ser_mux_inst_7_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_7_XOR2_U1 ( .A0_t (stateArray_MUX_inS03ser_mux_inst_7_Y), .B0_t (MixColumns_line1_S02[0]), .Z0_t (stateArray_inS03ser[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_0_XOR1_U1 ( .A0_t (MCin[8]), .B0_t (StateInMC[16]), .Z0_t (stateArray_MUX_inS13ser_mux_inst_0_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_0_AND1_U1 ( .A0_t (stateArray_nReset_selMC), .B0_t (stateArray_MUX_inS13ser_mux_inst_0_X), .Z0_t (stateArray_MUX_inS13ser_mux_inst_0_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_0_XOR2_U1 ( .A0_t (stateArray_MUX_inS13ser_mux_inst_0_Y), .B0_t (MCin[8]), .Z0_t (stateArray_inS13ser[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_1_XOR1_U1 ( .A0_t (MixColumns_line2_S02[2]), .B0_t (StateInMC[17]), .Z0_t (stateArray_MUX_inS13ser_mux_inst_1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_1_AND1_U1 ( .A0_t (stateArray_nReset_selMC), .B0_t (stateArray_MUX_inS13ser_mux_inst_1_X), .Z0_t (stateArray_MUX_inS13ser_mux_inst_1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_1_XOR2_U1 ( .A0_t (stateArray_MUX_inS13ser_mux_inst_1_Y), .B0_t (MixColumns_line2_S02[2]), .Z0_t (stateArray_inS13ser[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_2_XOR1_U1 ( .A0_t (MCin[10]), .B0_t (StateInMC[18]), .Z0_t (stateArray_MUX_inS13ser_mux_inst_2_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_2_AND1_U1 ( .A0_t (stateArray_nReset_selMC), .B0_t (stateArray_MUX_inS13ser_mux_inst_2_X), .Z0_t (stateArray_MUX_inS13ser_mux_inst_2_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_2_XOR2_U1 ( .A0_t (stateArray_MUX_inS13ser_mux_inst_2_Y), .B0_t (MCin[10]), .Z0_t (stateArray_inS13ser[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_3_XOR1_U1 ( .A0_t (MCin[11]), .B0_t (StateInMC[19]), .Z0_t (stateArray_MUX_inS13ser_mux_inst_3_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_3_AND1_U1 ( .A0_t (stateArray_nReset_selMC), .B0_t (stateArray_MUX_inS13ser_mux_inst_3_X), .Z0_t (stateArray_MUX_inS13ser_mux_inst_3_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_3_XOR2_U1 ( .A0_t (stateArray_MUX_inS13ser_mux_inst_3_Y), .B0_t (MCin[11]), .Z0_t (stateArray_inS13ser[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_4_XOR1_U1 ( .A0_t (MixColumns_line2_S02[5]), .B0_t (StateInMC[20]), .Z0_t (stateArray_MUX_inS13ser_mux_inst_4_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_4_AND1_U1 ( .A0_t (stateArray_nReset_selMC), .B0_t (stateArray_MUX_inS13ser_mux_inst_4_X), .Z0_t (stateArray_MUX_inS13ser_mux_inst_4_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_4_XOR2_U1 ( .A0_t (stateArray_MUX_inS13ser_mux_inst_4_Y), .B0_t (MixColumns_line2_S02[5]), .Z0_t (stateArray_inS13ser[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_5_XOR1_U1 ( .A0_t (MixColumns_line2_S02[6]), .B0_t (StateInMC[21]), .Z0_t (stateArray_MUX_inS13ser_mux_inst_5_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_5_AND1_U1 ( .A0_t (stateArray_nReset_selMC), .B0_t (stateArray_MUX_inS13ser_mux_inst_5_X), .Z0_t (stateArray_MUX_inS13ser_mux_inst_5_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_5_XOR2_U1 ( .A0_t (stateArray_MUX_inS13ser_mux_inst_5_Y), .B0_t (MixColumns_line2_S02[6]), .Z0_t (stateArray_inS13ser[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_6_XOR1_U1 ( .A0_t (MixColumns_line2_S02[7]), .B0_t (StateInMC[22]), .Z0_t (stateArray_MUX_inS13ser_mux_inst_6_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_6_AND1_U1 ( .A0_t (stateArray_nReset_selMC), .B0_t (stateArray_MUX_inS13ser_mux_inst_6_X), .Z0_t (stateArray_MUX_inS13ser_mux_inst_6_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_6_XOR2_U1 ( .A0_t (stateArray_MUX_inS13ser_mux_inst_6_Y), .B0_t (MixColumns_line2_S02[7]), .Z0_t (stateArray_inS13ser[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_7_XOR1_U1 ( .A0_t (MixColumns_line2_S02[0]), .B0_t (StateInMC[23]), .Z0_t (stateArray_MUX_inS13ser_mux_inst_7_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_7_AND1_U1 ( .A0_t (stateArray_nReset_selMC), .B0_t (stateArray_MUX_inS13ser_mux_inst_7_X), .Z0_t (stateArray_MUX_inS13ser_mux_inst_7_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_7_XOR2_U1 ( .A0_t (stateArray_MUX_inS13ser_mux_inst_7_Y), .B0_t (MixColumns_line2_S02[0]), .Z0_t (stateArray_inS13ser[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_0_XOR1_U1 ( .A0_t (MCin[0]), .B0_t (StateInMC[8]), .Z0_t (stateArray_MUX_inS23ser_mux_inst_0_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_0_AND1_U1 ( .A0_t (stateArray_nReset_selMC), .B0_t (stateArray_MUX_inS23ser_mux_inst_0_X), .Z0_t (stateArray_MUX_inS23ser_mux_inst_0_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_0_XOR2_U1 ( .A0_t (stateArray_MUX_inS23ser_mux_inst_0_Y), .B0_t (MCin[0]), .Z0_t (stateArray_inS23ser[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_1_XOR1_U1 ( .A0_t (MixColumns_line3_S02[2]), .B0_t (StateInMC[9]), .Z0_t (stateArray_MUX_inS23ser_mux_inst_1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_1_AND1_U1 ( .A0_t (stateArray_nReset_selMC), .B0_t (stateArray_MUX_inS23ser_mux_inst_1_X), .Z0_t (stateArray_MUX_inS23ser_mux_inst_1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_1_XOR2_U1 ( .A0_t (stateArray_MUX_inS23ser_mux_inst_1_Y), .B0_t (MixColumns_line3_S02[2]), .Z0_t (stateArray_inS23ser[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_2_XOR1_U1 ( .A0_t (MCin[2]), .B0_t (StateInMC[10]), .Z0_t (stateArray_MUX_inS23ser_mux_inst_2_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_2_AND1_U1 ( .A0_t (stateArray_nReset_selMC), .B0_t (stateArray_MUX_inS23ser_mux_inst_2_X), .Z0_t (stateArray_MUX_inS23ser_mux_inst_2_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_2_XOR2_U1 ( .A0_t (stateArray_MUX_inS23ser_mux_inst_2_Y), .B0_t (MCin[2]), .Z0_t (stateArray_inS23ser[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_3_XOR1_U1 ( .A0_t (MCin[3]), .B0_t (StateInMC[11]), .Z0_t (stateArray_MUX_inS23ser_mux_inst_3_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_3_AND1_U1 ( .A0_t (stateArray_nReset_selMC), .B0_t (stateArray_MUX_inS23ser_mux_inst_3_X), .Z0_t (stateArray_MUX_inS23ser_mux_inst_3_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_3_XOR2_U1 ( .A0_t (stateArray_MUX_inS23ser_mux_inst_3_Y), .B0_t (MCin[3]), .Z0_t (stateArray_inS23ser[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_4_XOR1_U1 ( .A0_t (MixColumns_line3_S02[5]), .B0_t (StateInMC[12]), .Z0_t (stateArray_MUX_inS23ser_mux_inst_4_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_4_AND1_U1 ( .A0_t (stateArray_nReset_selMC), .B0_t (stateArray_MUX_inS23ser_mux_inst_4_X), .Z0_t (stateArray_MUX_inS23ser_mux_inst_4_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_4_XOR2_U1 ( .A0_t (stateArray_MUX_inS23ser_mux_inst_4_Y), .B0_t (MixColumns_line3_S02[5]), .Z0_t (stateArray_inS23ser[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_5_XOR1_U1 ( .A0_t (MixColumns_line3_S02[6]), .B0_t (StateInMC[13]), .Z0_t (stateArray_MUX_inS23ser_mux_inst_5_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_5_AND1_U1 ( .A0_t (stateArray_nReset_selMC), .B0_t (stateArray_MUX_inS23ser_mux_inst_5_X), .Z0_t (stateArray_MUX_inS23ser_mux_inst_5_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_5_XOR2_U1 ( .A0_t (stateArray_MUX_inS23ser_mux_inst_5_Y), .B0_t (MixColumns_line3_S02[6]), .Z0_t (stateArray_inS23ser[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_6_XOR1_U1 ( .A0_t (MixColumns_line3_S02[7]), .B0_t (StateInMC[14]), .Z0_t (stateArray_MUX_inS23ser_mux_inst_6_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_6_AND1_U1 ( .A0_t (stateArray_nReset_selMC), .B0_t (stateArray_MUX_inS23ser_mux_inst_6_X), .Z0_t (stateArray_MUX_inS23ser_mux_inst_6_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_6_XOR2_U1 ( .A0_t (stateArray_MUX_inS23ser_mux_inst_6_Y), .B0_t (MixColumns_line3_S02[7]), .Z0_t (stateArray_inS23ser[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_7_XOR1_U1 ( .A0_t (MixColumns_line3_S02[0]), .B0_t (StateInMC[15]), .Z0_t (stateArray_MUX_inS23ser_mux_inst_7_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_7_AND1_U1 ( .A0_t (stateArray_nReset_selMC), .B0_t (stateArray_MUX_inS23ser_mux_inst_7_X), .Z0_t (stateArray_MUX_inS23ser_mux_inst_7_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_7_XOR2_U1 ( .A0_t (stateArray_MUX_inS23ser_mux_inst_7_Y), .B0_t (MixColumns_line3_S02[0]), .Z0_t (stateArray_inS23ser[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_0_XOR1_U1 ( .A0_t (StateIn[0]), .B0_t (StateInMC[0]), .Z0_t (stateArray_MUX_input_MC_mux_inst_0_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_0_AND1_U1 ( .A0_t (selMC), .B0_t (stateArray_MUX_input_MC_mux_inst_0_X), .Z0_t (stateArray_MUX_input_MC_mux_inst_0_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_0_XOR2_U1 ( .A0_t (stateArray_MUX_input_MC_mux_inst_0_Y), .B0_t (StateIn[0]), .Z0_t (stateArray_input_MC[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_1_XOR1_U1 ( .A0_t (StateIn[1]), .B0_t (StateInMC[1]), .Z0_t (stateArray_MUX_input_MC_mux_inst_1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_1_AND1_U1 ( .A0_t (selMC), .B0_t (stateArray_MUX_input_MC_mux_inst_1_X), .Z0_t (stateArray_MUX_input_MC_mux_inst_1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_1_XOR2_U1 ( .A0_t (stateArray_MUX_input_MC_mux_inst_1_Y), .B0_t (StateIn[1]), .Z0_t (stateArray_input_MC[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_2_XOR1_U1 ( .A0_t (StateIn[2]), .B0_t (StateInMC[2]), .Z0_t (stateArray_MUX_input_MC_mux_inst_2_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_2_AND1_U1 ( .A0_t (selMC), .B0_t (stateArray_MUX_input_MC_mux_inst_2_X), .Z0_t (stateArray_MUX_input_MC_mux_inst_2_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_2_XOR2_U1 ( .A0_t (stateArray_MUX_input_MC_mux_inst_2_Y), .B0_t (StateIn[2]), .Z0_t (stateArray_input_MC[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_3_XOR1_U1 ( .A0_t (StateIn[3]), .B0_t (StateInMC[3]), .Z0_t (stateArray_MUX_input_MC_mux_inst_3_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_3_AND1_U1 ( .A0_t (selMC), .B0_t (stateArray_MUX_input_MC_mux_inst_3_X), .Z0_t (stateArray_MUX_input_MC_mux_inst_3_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_3_XOR2_U1 ( .A0_t (stateArray_MUX_input_MC_mux_inst_3_Y), .B0_t (StateIn[3]), .Z0_t (stateArray_input_MC[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_4_XOR1_U1 ( .A0_t (StateIn[4]), .B0_t (StateInMC[4]), .Z0_t (stateArray_MUX_input_MC_mux_inst_4_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_4_AND1_U1 ( .A0_t (selMC), .B0_t (stateArray_MUX_input_MC_mux_inst_4_X), .Z0_t (stateArray_MUX_input_MC_mux_inst_4_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_4_XOR2_U1 ( .A0_t (stateArray_MUX_input_MC_mux_inst_4_Y), .B0_t (StateIn[4]), .Z0_t (stateArray_input_MC[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_5_XOR1_U1 ( .A0_t (StateIn[5]), .B0_t (StateInMC[5]), .Z0_t (stateArray_MUX_input_MC_mux_inst_5_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_5_AND1_U1 ( .A0_t (selMC), .B0_t (stateArray_MUX_input_MC_mux_inst_5_X), .Z0_t (stateArray_MUX_input_MC_mux_inst_5_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_5_XOR2_U1 ( .A0_t (stateArray_MUX_input_MC_mux_inst_5_Y), .B0_t (StateIn[5]), .Z0_t (stateArray_input_MC[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_6_XOR1_U1 ( .A0_t (StateIn[6]), .B0_t (StateInMC[6]), .Z0_t (stateArray_MUX_input_MC_mux_inst_6_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_6_AND1_U1 ( .A0_t (selMC), .B0_t (stateArray_MUX_input_MC_mux_inst_6_X), .Z0_t (stateArray_MUX_input_MC_mux_inst_6_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_6_XOR2_U1 ( .A0_t (stateArray_MUX_input_MC_mux_inst_6_Y), .B0_t (StateIn[6]), .Z0_t (stateArray_input_MC[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_7_XOR1_U1 ( .A0_t (StateIn[7]), .B0_t (StateInMC[7]), .Z0_t (stateArray_MUX_input_MC_mux_inst_7_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_7_AND1_U1 ( .A0_t (selMC), .B0_t (stateArray_MUX_input_MC_mux_inst_7_X), .Z0_t (stateArray_MUX_input_MC_mux_inst_7_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_7_XOR2_U1 ( .A0_t (stateArray_MUX_input_MC_mux_inst_7_Y), .B0_t (StateIn[7]), .Z0_t (stateArray_input_MC[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_0_XOR1_U1 ( .A0_t (port_in[0]), .B0_t (stateArray_input_MC[0]), .Z0_t (stateArray_MUX_inS33ser_mux_inst_0_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_0_AND1_U1 ( .A0_t (start), .B0_t (stateArray_MUX_inS33ser_mux_inst_0_X), .Z0_t (stateArray_MUX_inS33ser_mux_inst_0_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_0_XOR2_U1 ( .A0_t (stateArray_MUX_inS33ser_mux_inst_0_Y), .B0_t (port_in[0]), .Z0_t (stateArray_inS33ser[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_1_XOR1_U1 ( .A0_t (port_in[1]), .B0_t (stateArray_input_MC[1]), .Z0_t (stateArray_MUX_inS33ser_mux_inst_1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_1_AND1_U1 ( .A0_t (start), .B0_t (stateArray_MUX_inS33ser_mux_inst_1_X), .Z0_t (stateArray_MUX_inS33ser_mux_inst_1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_1_XOR2_U1 ( .A0_t (stateArray_MUX_inS33ser_mux_inst_1_Y), .B0_t (port_in[1]), .Z0_t (stateArray_inS33ser[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_2_XOR1_U1 ( .A0_t (port_in[2]), .B0_t (stateArray_input_MC[2]), .Z0_t (stateArray_MUX_inS33ser_mux_inst_2_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_2_AND1_U1 ( .A0_t (start), .B0_t (stateArray_MUX_inS33ser_mux_inst_2_X), .Z0_t (stateArray_MUX_inS33ser_mux_inst_2_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_2_XOR2_U1 ( .A0_t (stateArray_MUX_inS33ser_mux_inst_2_Y), .B0_t (port_in[2]), .Z0_t (stateArray_inS33ser[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_3_XOR1_U1 ( .A0_t (port_in[3]), .B0_t (stateArray_input_MC[3]), .Z0_t (stateArray_MUX_inS33ser_mux_inst_3_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_3_AND1_U1 ( .A0_t (start), .B0_t (stateArray_MUX_inS33ser_mux_inst_3_X), .Z0_t (stateArray_MUX_inS33ser_mux_inst_3_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_3_XOR2_U1 ( .A0_t (stateArray_MUX_inS33ser_mux_inst_3_Y), .B0_t (port_in[3]), .Z0_t (stateArray_inS33ser[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_4_XOR1_U1 ( .A0_t (port_in[4]), .B0_t (stateArray_input_MC[4]), .Z0_t (stateArray_MUX_inS33ser_mux_inst_4_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_4_AND1_U1 ( .A0_t (start), .B0_t (stateArray_MUX_inS33ser_mux_inst_4_X), .Z0_t (stateArray_MUX_inS33ser_mux_inst_4_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_4_XOR2_U1 ( .A0_t (stateArray_MUX_inS33ser_mux_inst_4_Y), .B0_t (port_in[4]), .Z0_t (stateArray_inS33ser[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_5_XOR1_U1 ( .A0_t (port_in[5]), .B0_t (stateArray_input_MC[5]), .Z0_t (stateArray_MUX_inS33ser_mux_inst_5_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_5_AND1_U1 ( .A0_t (start), .B0_t (stateArray_MUX_inS33ser_mux_inst_5_X), .Z0_t (stateArray_MUX_inS33ser_mux_inst_5_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_5_XOR2_U1 ( .A0_t (stateArray_MUX_inS33ser_mux_inst_5_Y), .B0_t (port_in[5]), .Z0_t (stateArray_inS33ser[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_6_XOR1_U1 ( .A0_t (port_in[6]), .B0_t (stateArray_input_MC[6]), .Z0_t (stateArray_MUX_inS33ser_mux_inst_6_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_6_AND1_U1 ( .A0_t (start), .B0_t (stateArray_MUX_inS33ser_mux_inst_6_X), .Z0_t (stateArray_MUX_inS33ser_mux_inst_6_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_6_XOR2_U1 ( .A0_t (stateArray_MUX_inS33ser_mux_inst_6_Y), .B0_t (port_in[6]), .Z0_t (stateArray_inS33ser[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_7_XOR1_U1 ( .A0_t (port_in[7]), .B0_t (stateArray_input_MC[7]), .Z0_t (stateArray_MUX_inS33ser_mux_inst_7_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_7_AND1_U1 ( .A0_t (start), .B0_t (stateArray_MUX_inS33ser_mux_inst_7_X), .Z0_t (stateArray_MUX_inS33ser_mux_inst_7_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_7_XOR2_U1 ( .A0_t (stateArray_MUX_inS33ser_mux_inst_7_Y), .B0_t (port_in[7]), .Z0_t (stateArray_inS33ser[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_0_XOR1_U1 ( .A0_t (MCout[0]), .B0_t (MCin[0]), .Z0_t (MUX_StateInMC_mux_inst_0_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_0_AND1_U1 ( .A0_t (intFinal), .B0_t (MUX_StateInMC_mux_inst_0_X), .Z0_t (MUX_StateInMC_mux_inst_0_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_0_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_0_Y), .B0_t (MCout[0]), .Z0_t (StateInMC[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_1_XOR1_U1 ( .A0_t (MCout[1]), .B0_t (MixColumns_line3_S02[2]), .Z0_t (MUX_StateInMC_mux_inst_1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_1_AND1_U1 ( .A0_t (intFinal), .B0_t (MUX_StateInMC_mux_inst_1_X), .Z0_t (MUX_StateInMC_mux_inst_1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_1_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_1_Y), .B0_t (MCout[1]), .Z0_t (StateInMC[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_2_XOR1_U1 ( .A0_t (MCout[2]), .B0_t (MCin[2]), .Z0_t (MUX_StateInMC_mux_inst_2_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_2_AND1_U1 ( .A0_t (intFinal), .B0_t (MUX_StateInMC_mux_inst_2_X), .Z0_t (MUX_StateInMC_mux_inst_2_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_2_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_2_Y), .B0_t (MCout[2]), .Z0_t (StateInMC[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_3_XOR1_U1 ( .A0_t (MCout[3]), .B0_t (MCin[3]), .Z0_t (MUX_StateInMC_mux_inst_3_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_3_AND1_U1 ( .A0_t (intFinal), .B0_t (MUX_StateInMC_mux_inst_3_X), .Z0_t (MUX_StateInMC_mux_inst_3_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_3_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_3_Y), .B0_t (MCout[3]), .Z0_t (StateInMC[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_4_XOR1_U1 ( .A0_t (MCout[4]), .B0_t (MixColumns_line3_S02[5]), .Z0_t (MUX_StateInMC_mux_inst_4_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_4_AND1_U1 ( .A0_t (intFinal), .B0_t (MUX_StateInMC_mux_inst_4_X), .Z0_t (MUX_StateInMC_mux_inst_4_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_4_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_4_Y), .B0_t (MCout[4]), .Z0_t (StateInMC[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_5_XOR1_U1 ( .A0_t (MCout[5]), .B0_t (MixColumns_line3_S02[6]), .Z0_t (MUX_StateInMC_mux_inst_5_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_5_AND1_U1 ( .A0_t (intFinal), .B0_t (MUX_StateInMC_mux_inst_5_X), .Z0_t (MUX_StateInMC_mux_inst_5_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_5_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_5_Y), .B0_t (MCout[5]), .Z0_t (StateInMC[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_6_XOR1_U1 ( .A0_t (MCout[6]), .B0_t (MixColumns_line3_S02[7]), .Z0_t (MUX_StateInMC_mux_inst_6_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_6_AND1_U1 ( .A0_t (intFinal), .B0_t (MUX_StateInMC_mux_inst_6_X), .Z0_t (MUX_StateInMC_mux_inst_6_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_6_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_6_Y), .B0_t (MCout[6]), .Z0_t (StateInMC[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_7_XOR1_U1 ( .A0_t (MCout[7]), .B0_t (MixColumns_line3_S02[0]), .Z0_t (MUX_StateInMC_mux_inst_7_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_7_AND1_U1 ( .A0_t (intFinal), .B0_t (MUX_StateInMC_mux_inst_7_X), .Z0_t (MUX_StateInMC_mux_inst_7_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_7_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_7_Y), .B0_t (MCout[7]), .Z0_t (StateInMC[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_8_XOR1_U1 ( .A0_t (MCout[8]), .B0_t (MCin[8]), .Z0_t (MUX_StateInMC_mux_inst_8_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_8_AND1_U1 ( .A0_t (intFinal), .B0_t (MUX_StateInMC_mux_inst_8_X), .Z0_t (MUX_StateInMC_mux_inst_8_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_8_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_8_Y), .B0_t (MCout[8]), .Z0_t (StateInMC[8]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_9_XOR1_U1 ( .A0_t (MCout[9]), .B0_t (MixColumns_line2_S02[2]), .Z0_t (MUX_StateInMC_mux_inst_9_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_9_AND1_U1 ( .A0_t (intFinal), .B0_t (MUX_StateInMC_mux_inst_9_X), .Z0_t (MUX_StateInMC_mux_inst_9_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_9_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_9_Y), .B0_t (MCout[9]), .Z0_t (StateInMC[9]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_10_XOR1_U1 ( .A0_t (MCout[10]), .B0_t (MCin[10]), .Z0_t (MUX_StateInMC_mux_inst_10_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_10_AND1_U1 ( .A0_t (intFinal), .B0_t (MUX_StateInMC_mux_inst_10_X), .Z0_t (MUX_StateInMC_mux_inst_10_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_10_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_10_Y), .B0_t (MCout[10]), .Z0_t (StateInMC[10]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_11_XOR1_U1 ( .A0_t (MCout[11]), .B0_t (MCin[11]), .Z0_t (MUX_StateInMC_mux_inst_11_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_11_AND1_U1 ( .A0_t (intFinal), .B0_t (MUX_StateInMC_mux_inst_11_X), .Z0_t (MUX_StateInMC_mux_inst_11_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_11_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_11_Y), .B0_t (MCout[11]), .Z0_t (StateInMC[11]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_12_XOR1_U1 ( .A0_t (MCout[12]), .B0_t (MixColumns_line2_S02[5]), .Z0_t (MUX_StateInMC_mux_inst_12_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_12_AND1_U1 ( .A0_t (intFinal), .B0_t (MUX_StateInMC_mux_inst_12_X), .Z0_t (MUX_StateInMC_mux_inst_12_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_12_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_12_Y), .B0_t (MCout[12]), .Z0_t (StateInMC[12]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_13_XOR1_U1 ( .A0_t (MCout[13]), .B0_t (MixColumns_line2_S02[6]), .Z0_t (MUX_StateInMC_mux_inst_13_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_13_AND1_U1 ( .A0_t (intFinal), .B0_t (MUX_StateInMC_mux_inst_13_X), .Z0_t (MUX_StateInMC_mux_inst_13_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_13_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_13_Y), .B0_t (MCout[13]), .Z0_t (StateInMC[13]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_14_XOR1_U1 ( .A0_t (MCout[14]), .B0_t (MixColumns_line2_S02[7]), .Z0_t (MUX_StateInMC_mux_inst_14_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_14_AND1_U1 ( .A0_t (intFinal), .B0_t (MUX_StateInMC_mux_inst_14_X), .Z0_t (MUX_StateInMC_mux_inst_14_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_14_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_14_Y), .B0_t (MCout[14]), .Z0_t (StateInMC[14]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_15_XOR1_U1 ( .A0_t (MCout[15]), .B0_t (MixColumns_line2_S02[0]), .Z0_t (MUX_StateInMC_mux_inst_15_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_15_AND1_U1 ( .A0_t (intFinal), .B0_t (MUX_StateInMC_mux_inst_15_X), .Z0_t (MUX_StateInMC_mux_inst_15_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_15_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_15_Y), .B0_t (MCout[15]), .Z0_t (StateInMC[15]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_16_XOR1_U1 ( .A0_t (MCout[16]), .B0_t (MCin[16]), .Z0_t (MUX_StateInMC_mux_inst_16_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_16_AND1_U1 ( .A0_t (intFinal), .B0_t (MUX_StateInMC_mux_inst_16_X), .Z0_t (MUX_StateInMC_mux_inst_16_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_16_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_16_Y), .B0_t (MCout[16]), .Z0_t (StateInMC[16]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_17_XOR1_U1 ( .A0_t (MCout[17]), .B0_t (MixColumns_line1_S02[2]), .Z0_t (MUX_StateInMC_mux_inst_17_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_17_AND1_U1 ( .A0_t (intFinal), .B0_t (MUX_StateInMC_mux_inst_17_X), .Z0_t (MUX_StateInMC_mux_inst_17_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_17_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_17_Y), .B0_t (MCout[17]), .Z0_t (StateInMC[17]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_18_XOR1_U1 ( .A0_t (MCout[18]), .B0_t (MCin[18]), .Z0_t (MUX_StateInMC_mux_inst_18_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_18_AND1_U1 ( .A0_t (intFinal), .B0_t (MUX_StateInMC_mux_inst_18_X), .Z0_t (MUX_StateInMC_mux_inst_18_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_18_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_18_Y), .B0_t (MCout[18]), .Z0_t (StateInMC[18]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_19_XOR1_U1 ( .A0_t (MCout[19]), .B0_t (MCin[19]), .Z0_t (MUX_StateInMC_mux_inst_19_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_19_AND1_U1 ( .A0_t (intFinal), .B0_t (MUX_StateInMC_mux_inst_19_X), .Z0_t (MUX_StateInMC_mux_inst_19_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_19_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_19_Y), .B0_t (MCout[19]), .Z0_t (StateInMC[19]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_20_XOR1_U1 ( .A0_t (MCout[20]), .B0_t (MixColumns_line1_S02[5]), .Z0_t (MUX_StateInMC_mux_inst_20_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_20_AND1_U1 ( .A0_t (intFinal), .B0_t (MUX_StateInMC_mux_inst_20_X), .Z0_t (MUX_StateInMC_mux_inst_20_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_20_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_20_Y), .B0_t (MCout[20]), .Z0_t (StateInMC[20]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_21_XOR1_U1 ( .A0_t (MCout[21]), .B0_t (MixColumns_line1_S02[6]), .Z0_t (MUX_StateInMC_mux_inst_21_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_21_AND1_U1 ( .A0_t (intFinal), .B0_t (MUX_StateInMC_mux_inst_21_X), .Z0_t (MUX_StateInMC_mux_inst_21_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_21_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_21_Y), .B0_t (MCout[21]), .Z0_t (StateInMC[21]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_22_XOR1_U1 ( .A0_t (MCout[22]), .B0_t (MixColumns_line1_S02[7]), .Z0_t (MUX_StateInMC_mux_inst_22_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_22_AND1_U1 ( .A0_t (intFinal), .B0_t (MUX_StateInMC_mux_inst_22_X), .Z0_t (MUX_StateInMC_mux_inst_22_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_22_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_22_Y), .B0_t (MCout[22]), .Z0_t (StateInMC[22]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_23_XOR1_U1 ( .A0_t (MCout[23]), .B0_t (MixColumns_line1_S02[0]), .Z0_t (MUX_StateInMC_mux_inst_23_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_23_AND1_U1 ( .A0_t (intFinal), .B0_t (MUX_StateInMC_mux_inst_23_X), .Z0_t (MUX_StateInMC_mux_inst_23_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_23_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_23_Y), .B0_t (MCout[23]), .Z0_t (StateInMC[23]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_24_XOR1_U1 ( .A0_t (MCout[24]), .B0_t (port_out[0]), .Z0_t (MUX_StateInMC_mux_inst_24_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_24_AND1_U1 ( .A0_t (intFinal), .B0_t (MUX_StateInMC_mux_inst_24_X), .Z0_t (MUX_StateInMC_mux_inst_24_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_24_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_24_Y), .B0_t (MCout[24]), .Z0_t (StateInMC[24]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_25_XOR1_U1 ( .A0_t (MCout[25]), .B0_t (port_out[1]), .Z0_t (MUX_StateInMC_mux_inst_25_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_25_AND1_U1 ( .A0_t (intFinal), .B0_t (MUX_StateInMC_mux_inst_25_X), .Z0_t (MUX_StateInMC_mux_inst_25_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_25_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_25_Y), .B0_t (MCout[25]), .Z0_t (StateInMC[25]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_26_XOR1_U1 ( .A0_t (MCout[26]), .B0_t (port_out[2]), .Z0_t (MUX_StateInMC_mux_inst_26_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_26_AND1_U1 ( .A0_t (intFinal), .B0_t (MUX_StateInMC_mux_inst_26_X), .Z0_t (MUX_StateInMC_mux_inst_26_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_26_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_26_Y), .B0_t (MCout[26]), .Z0_t (StateInMC[26]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_27_XOR1_U1 ( .A0_t (MCout[27]), .B0_t (port_out[3]), .Z0_t (MUX_StateInMC_mux_inst_27_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_27_AND1_U1 ( .A0_t (intFinal), .B0_t (MUX_StateInMC_mux_inst_27_X), .Z0_t (MUX_StateInMC_mux_inst_27_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_27_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_27_Y), .B0_t (MCout[27]), .Z0_t (StateInMC[27]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_28_XOR1_U1 ( .A0_t (MCout[28]), .B0_t (port_out[4]), .Z0_t (MUX_StateInMC_mux_inst_28_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_28_AND1_U1 ( .A0_t (intFinal), .B0_t (MUX_StateInMC_mux_inst_28_X), .Z0_t (MUX_StateInMC_mux_inst_28_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_28_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_28_Y), .B0_t (MCout[28]), .Z0_t (StateInMC[28]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_29_XOR1_U1 ( .A0_t (MCout[29]), .B0_t (port_out[5]), .Z0_t (MUX_StateInMC_mux_inst_29_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_29_AND1_U1 ( .A0_t (intFinal), .B0_t (MUX_StateInMC_mux_inst_29_X), .Z0_t (MUX_StateInMC_mux_inst_29_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_29_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_29_Y), .B0_t (MCout[29]), .Z0_t (StateInMC[29]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_30_XOR1_U1 ( .A0_t (MCout[30]), .B0_t (port_out[6]), .Z0_t (MUX_StateInMC_mux_inst_30_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_30_AND1_U1 ( .A0_t (intFinal), .B0_t (MUX_StateInMC_mux_inst_30_X), .Z0_t (MUX_StateInMC_mux_inst_30_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_30_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_30_Y), .B0_t (MCout[30]), .Z0_t (StateInMC[30]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_31_XOR1_U1 ( .A0_t (MCout[31]), .B0_t (port_out[7]), .Z0_t (MUX_StateInMC_mux_inst_31_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_31_AND1_U1 ( .A0_t (intFinal), .B0_t (MUX_StateInMC_mux_inst_31_X), .Z0_t (MUX_StateInMC_mux_inst_31_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_31_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_31_Y), .B0_t (MCout[31]), .Z0_t (StateInMC[31]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_U32 ( .A0_t (KeyArray_outS01ser_7_), .B0_t (keyStateIn[7]), .Z0_t (KeyArray_outS01ser_XOR_00[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_U31 ( .A0_t (KeyArray_outS01ser_6_), .B0_t (keyStateIn[6]), .Z0_t (KeyArray_outS01ser_XOR_00[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_U30 ( .A0_t (KeyArray_outS01ser_5_), .B0_t (keyStateIn[5]), .Z0_t (KeyArray_outS01ser_XOR_00[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_U29 ( .A0_t (KeyArray_outS01ser_4_), .B0_t (keyStateIn[4]), .Z0_t (KeyArray_outS01ser_XOR_00[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_U28 ( .A0_t (KeyArray_outS01ser_3_), .B0_t (keyStateIn[3]), .Z0_t (KeyArray_outS01ser_XOR_00[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_U27 ( .A0_t (KeyArray_outS01ser_2_), .B0_t (keyStateIn[2]), .Z0_t (KeyArray_outS01ser_XOR_00[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_U26 ( .A0_t (KeyArray_outS01ser_1_), .B0_t (keyStateIn[1]), .Z0_t (KeyArray_outS01ser_XOR_00[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_U25 ( .A0_t (KeyArray_outS01ser_0_), .B0_t (keyStateIn[0]), .Z0_t (KeyArray_outS01ser_XOR_00[0]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) KeyArray_U24 ( .A0_t (start), .B0_t (intselXOR), .Z0_t (KeyArray_nReset_selXOR) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_U23 ( .A0_t (KeyArray_n32), .B0_t (keyStateIn[7]), .Z0_t (KeyArray_inS30par[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_U22 ( .A0_t (roundConstant[7]), .B0_t (SboxOut[7]), .Z0_t (KeyArray_n32) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_U21 ( .A0_t (KeyArray_n31), .B0_t (keyStateIn[6]), .Z0_t (KeyArray_inS30par[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_U20 ( .A0_t (roundConstant[6]), .B0_t (SboxOut[6]), .Z0_t (KeyArray_n31) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_U19 ( .A0_t (KeyArray_n30), .B0_t (keyStateIn[5]), .Z0_t (KeyArray_inS30par[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_U18 ( .A0_t (roundConstant[5]), .B0_t (SboxOut[5]), .Z0_t (KeyArray_n30) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_U17 ( .A0_t (KeyArray_n29), .B0_t (keyStateIn[4]), .Z0_t (KeyArray_inS30par[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_U16 ( .A0_t (roundConstant[4]), .B0_t (SboxOut[4]), .Z0_t (KeyArray_n29) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_U15 ( .A0_t (KeyArray_n28), .B0_t (keyStateIn[3]), .Z0_t (KeyArray_inS30par[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_U14 ( .A0_t (roundConstant[3]), .B0_t (SboxOut[3]), .Z0_t (KeyArray_n28) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_U13 ( .A0_t (KeyArray_n27), .B0_t (keyStateIn[2]), .Z0_t (KeyArray_inS30par[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_U12 ( .A0_t (roundConstant[2]), .B0_t (SboxOut[2]), .Z0_t (KeyArray_n27) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_U11 ( .A0_t (KeyArray_n26), .B0_t (keyStateIn[1]), .Z0_t (KeyArray_inS30par[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_U10 ( .A0_t (roundConstant[1]), .B0_t (SboxOut[1]), .Z0_t (KeyArray_n26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_U9 ( .A0_t (KeyArray_n25), .B0_t (keyStateIn[0]), .Z0_t (KeyArray_inS30par[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_U8 ( .A0_t (roundConstant[0]), .B0_t (SboxOut[0]), .Z0_t (KeyArray_n25) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S00reg_gff_1_SFF_0_U3 ( .A0_t (KeyArray_S00reg_gff_1_SFF_0_n2), .B0_t (KeyArray_S00reg_gff_1_SFF_0_n1), .Z0_t (keyStateIn[0]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_0_U2 ( .A0_t (enKS), .B0_t (keyStateIn[0]), .Z0_t (KeyArray_S00reg_gff_1_SFF_0_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_0_U1 ( .A0_t (KeyArray_S00reg_gff_1_SFF_0_QD), .B0_t (enKS), .Z0_t (KeyArray_S00reg_gff_1_SFF_0_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS00ser[0]), .B0_t (KeyArray_outS10ser[0]), .Z0_t (KeyArray_S00reg_gff_1_SFF_0_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S00reg_gff_1_SFF_0_MUXInst_X), .Z0_t (KeyArray_S00reg_gff_1_SFF_0_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S00reg_gff_1_SFF_0_MUXInst_Y), .B0_t (KeyArray_inS00ser[0]), .Z0_t (KeyArray_S00reg_gff_1_SFF_0_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S00reg_gff_1_SFF_1_U3 ( .A0_t (KeyArray_S00reg_gff_1_SFF_1_n2), .B0_t (KeyArray_S00reg_gff_1_SFF_1_n1), .Z0_t (keyStateIn[1]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_1_U2 ( .A0_t (enKS), .B0_t (keyStateIn[1]), .Z0_t (KeyArray_S00reg_gff_1_SFF_1_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_1_U1 ( .A0_t (KeyArray_S00reg_gff_1_SFF_1_QD), .B0_t (enKS), .Z0_t (KeyArray_S00reg_gff_1_SFF_1_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS00ser[1]), .B0_t (KeyArray_outS10ser[1]), .Z0_t (KeyArray_S00reg_gff_1_SFF_1_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S00reg_gff_1_SFF_1_MUXInst_X), .Z0_t (KeyArray_S00reg_gff_1_SFF_1_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S00reg_gff_1_SFF_1_MUXInst_Y), .B0_t (KeyArray_inS00ser[1]), .Z0_t (KeyArray_S00reg_gff_1_SFF_1_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S00reg_gff_1_SFF_2_U3 ( .A0_t (KeyArray_S00reg_gff_1_SFF_2_n2), .B0_t (KeyArray_S00reg_gff_1_SFF_2_n1), .Z0_t (keyStateIn[2]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_2_U2 ( .A0_t (enKS), .B0_t (keyStateIn[2]), .Z0_t (KeyArray_S00reg_gff_1_SFF_2_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_2_U1 ( .A0_t (KeyArray_S00reg_gff_1_SFF_2_QD), .B0_t (enKS), .Z0_t (KeyArray_S00reg_gff_1_SFF_2_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS00ser[2]), .B0_t (KeyArray_outS10ser[2]), .Z0_t (KeyArray_S00reg_gff_1_SFF_2_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S00reg_gff_1_SFF_2_MUXInst_X), .Z0_t (KeyArray_S00reg_gff_1_SFF_2_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S00reg_gff_1_SFF_2_MUXInst_Y), .B0_t (KeyArray_inS00ser[2]), .Z0_t (KeyArray_S00reg_gff_1_SFF_2_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S00reg_gff_1_SFF_3_U3 ( .A0_t (KeyArray_S00reg_gff_1_SFF_3_n2), .B0_t (KeyArray_S00reg_gff_1_SFF_3_n1), .Z0_t (keyStateIn[3]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_3_U2 ( .A0_t (enKS), .B0_t (keyStateIn[3]), .Z0_t (KeyArray_S00reg_gff_1_SFF_3_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_3_U1 ( .A0_t (KeyArray_S00reg_gff_1_SFF_3_QD), .B0_t (enKS), .Z0_t (KeyArray_S00reg_gff_1_SFF_3_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS00ser[3]), .B0_t (KeyArray_outS10ser[3]), .Z0_t (KeyArray_S00reg_gff_1_SFF_3_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S00reg_gff_1_SFF_3_MUXInst_X), .Z0_t (KeyArray_S00reg_gff_1_SFF_3_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S00reg_gff_1_SFF_3_MUXInst_Y), .B0_t (KeyArray_inS00ser[3]), .Z0_t (KeyArray_S00reg_gff_1_SFF_3_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S00reg_gff_1_SFF_4_U3 ( .A0_t (KeyArray_S00reg_gff_1_SFF_4_n2), .B0_t (KeyArray_S00reg_gff_1_SFF_4_n1), .Z0_t (keyStateIn[4]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_4_U2 ( .A0_t (enKS), .B0_t (keyStateIn[4]), .Z0_t (KeyArray_S00reg_gff_1_SFF_4_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_4_U1 ( .A0_t (KeyArray_S00reg_gff_1_SFF_4_QD), .B0_t (enKS), .Z0_t (KeyArray_S00reg_gff_1_SFF_4_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS00ser[4]), .B0_t (KeyArray_outS10ser[4]), .Z0_t (KeyArray_S00reg_gff_1_SFF_4_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S00reg_gff_1_SFF_4_MUXInst_X), .Z0_t (KeyArray_S00reg_gff_1_SFF_4_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S00reg_gff_1_SFF_4_MUXInst_Y), .B0_t (KeyArray_inS00ser[4]), .Z0_t (KeyArray_S00reg_gff_1_SFF_4_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S00reg_gff_1_SFF_5_U3 ( .A0_t (KeyArray_S00reg_gff_1_SFF_5_n2), .B0_t (KeyArray_S00reg_gff_1_SFF_5_n1), .Z0_t (keyStateIn[5]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_5_U2 ( .A0_t (enKS), .B0_t (keyStateIn[5]), .Z0_t (KeyArray_S00reg_gff_1_SFF_5_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_5_U1 ( .A0_t (KeyArray_S00reg_gff_1_SFF_5_QD), .B0_t (enKS), .Z0_t (KeyArray_S00reg_gff_1_SFF_5_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS00ser[5]), .B0_t (KeyArray_outS10ser[5]), .Z0_t (KeyArray_S00reg_gff_1_SFF_5_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S00reg_gff_1_SFF_5_MUXInst_X), .Z0_t (KeyArray_S00reg_gff_1_SFF_5_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S00reg_gff_1_SFF_5_MUXInst_Y), .B0_t (KeyArray_inS00ser[5]), .Z0_t (KeyArray_S00reg_gff_1_SFF_5_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S00reg_gff_1_SFF_6_U3 ( .A0_t (KeyArray_S00reg_gff_1_SFF_6_n2), .B0_t (KeyArray_S00reg_gff_1_SFF_6_n1), .Z0_t (keyStateIn[6]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_6_U2 ( .A0_t (enKS), .B0_t (keyStateIn[6]), .Z0_t (KeyArray_S00reg_gff_1_SFF_6_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_6_U1 ( .A0_t (KeyArray_S00reg_gff_1_SFF_6_QD), .B0_t (enKS), .Z0_t (KeyArray_S00reg_gff_1_SFF_6_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS00ser[6]), .B0_t (KeyArray_outS10ser[6]), .Z0_t (KeyArray_S00reg_gff_1_SFF_6_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S00reg_gff_1_SFF_6_MUXInst_X), .Z0_t (KeyArray_S00reg_gff_1_SFF_6_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S00reg_gff_1_SFF_6_MUXInst_Y), .B0_t (KeyArray_inS00ser[6]), .Z0_t (KeyArray_S00reg_gff_1_SFF_6_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S00reg_gff_1_SFF_7_U3 ( .A0_t (KeyArray_S00reg_gff_1_SFF_7_n2), .B0_t (KeyArray_S00reg_gff_1_SFF_7_n1), .Z0_t (keyStateIn[7]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_7_U2 ( .A0_t (enKS), .B0_t (keyStateIn[7]), .Z0_t (KeyArray_S00reg_gff_1_SFF_7_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_7_U1 ( .A0_t (KeyArray_S00reg_gff_1_SFF_7_QD), .B0_t (enKS), .Z0_t (KeyArray_S00reg_gff_1_SFF_7_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS00ser[7]), .B0_t (KeyArray_outS10ser[7]), .Z0_t (KeyArray_S00reg_gff_1_SFF_7_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S00reg_gff_1_SFF_7_MUXInst_X), .Z0_t (KeyArray_S00reg_gff_1_SFF_7_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S00reg_gff_1_SFF_7_MUXInst_Y), .B0_t (KeyArray_inS00ser[7]), .Z0_t (KeyArray_S00reg_gff_1_SFF_7_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S01reg_gff_1_SFF_0_U3 ( .A0_t (KeyArray_S01reg_gff_1_SFF_0_n2), .B0_t (KeyArray_S01reg_gff_1_SFF_0_n1), .Z0_t (KeyArray_outS01ser_0_) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_0_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS01ser_0_), .Z0_t (KeyArray_S01reg_gff_1_SFF_0_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_0_U1 ( .A0_t (KeyArray_S01reg_gff_1_SFF_0_QD), .B0_t (enKS), .Z0_t (KeyArray_S01reg_gff_1_SFF_0_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS02ser[0]), .B0_t (KeyArray_outS11ser[0]), .Z0_t (KeyArray_S01reg_gff_1_SFF_0_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S01reg_gff_1_SFF_0_MUXInst_X), .Z0_t (KeyArray_S01reg_gff_1_SFF_0_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S01reg_gff_1_SFF_0_MUXInst_Y), .B0_t (KeyArray_outS02ser[0]), .Z0_t (KeyArray_S01reg_gff_1_SFF_0_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S01reg_gff_1_SFF_1_U3 ( .A0_t (KeyArray_S01reg_gff_1_SFF_1_n2), .B0_t (KeyArray_S01reg_gff_1_SFF_1_n1), .Z0_t (KeyArray_outS01ser_1_) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_1_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS01ser_1_), .Z0_t (KeyArray_S01reg_gff_1_SFF_1_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_1_U1 ( .A0_t (KeyArray_S01reg_gff_1_SFF_1_QD), .B0_t (enKS), .Z0_t (KeyArray_S01reg_gff_1_SFF_1_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS02ser[1]), .B0_t (KeyArray_outS11ser[1]), .Z0_t (KeyArray_S01reg_gff_1_SFF_1_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S01reg_gff_1_SFF_1_MUXInst_X), .Z0_t (KeyArray_S01reg_gff_1_SFF_1_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S01reg_gff_1_SFF_1_MUXInst_Y), .B0_t (KeyArray_outS02ser[1]), .Z0_t (KeyArray_S01reg_gff_1_SFF_1_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S01reg_gff_1_SFF_2_U3 ( .A0_t (KeyArray_S01reg_gff_1_SFF_2_n2), .B0_t (KeyArray_S01reg_gff_1_SFF_2_n1), .Z0_t (KeyArray_outS01ser_2_) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_2_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS01ser_2_), .Z0_t (KeyArray_S01reg_gff_1_SFF_2_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_2_U1 ( .A0_t (KeyArray_S01reg_gff_1_SFF_2_QD), .B0_t (enKS), .Z0_t (KeyArray_S01reg_gff_1_SFF_2_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS02ser[2]), .B0_t (KeyArray_outS11ser[2]), .Z0_t (KeyArray_S01reg_gff_1_SFF_2_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S01reg_gff_1_SFF_2_MUXInst_X), .Z0_t (KeyArray_S01reg_gff_1_SFF_2_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S01reg_gff_1_SFF_2_MUXInst_Y), .B0_t (KeyArray_outS02ser[2]), .Z0_t (KeyArray_S01reg_gff_1_SFF_2_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S01reg_gff_1_SFF_3_U3 ( .A0_t (KeyArray_S01reg_gff_1_SFF_3_n2), .B0_t (KeyArray_S01reg_gff_1_SFF_3_n1), .Z0_t (KeyArray_outS01ser_3_) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_3_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS01ser_3_), .Z0_t (KeyArray_S01reg_gff_1_SFF_3_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_3_U1 ( .A0_t (KeyArray_S01reg_gff_1_SFF_3_QD), .B0_t (enKS), .Z0_t (KeyArray_S01reg_gff_1_SFF_3_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS02ser[3]), .B0_t (KeyArray_outS11ser[3]), .Z0_t (KeyArray_S01reg_gff_1_SFF_3_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S01reg_gff_1_SFF_3_MUXInst_X), .Z0_t (KeyArray_S01reg_gff_1_SFF_3_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S01reg_gff_1_SFF_3_MUXInst_Y), .B0_t (KeyArray_outS02ser[3]), .Z0_t (KeyArray_S01reg_gff_1_SFF_3_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S01reg_gff_1_SFF_4_U3 ( .A0_t (KeyArray_S01reg_gff_1_SFF_4_n2), .B0_t (KeyArray_S01reg_gff_1_SFF_4_n1), .Z0_t (KeyArray_outS01ser_4_) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_4_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS01ser_4_), .Z0_t (KeyArray_S01reg_gff_1_SFF_4_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_4_U1 ( .A0_t (KeyArray_S01reg_gff_1_SFF_4_QD), .B0_t (enKS), .Z0_t (KeyArray_S01reg_gff_1_SFF_4_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS02ser[4]), .B0_t (KeyArray_outS11ser[4]), .Z0_t (KeyArray_S01reg_gff_1_SFF_4_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S01reg_gff_1_SFF_4_MUXInst_X), .Z0_t (KeyArray_S01reg_gff_1_SFF_4_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S01reg_gff_1_SFF_4_MUXInst_Y), .B0_t (KeyArray_outS02ser[4]), .Z0_t (KeyArray_S01reg_gff_1_SFF_4_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S01reg_gff_1_SFF_5_U3 ( .A0_t (KeyArray_S01reg_gff_1_SFF_5_n2), .B0_t (KeyArray_S01reg_gff_1_SFF_5_n1), .Z0_t (KeyArray_outS01ser_5_) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_5_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS01ser_5_), .Z0_t (KeyArray_S01reg_gff_1_SFF_5_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_5_U1 ( .A0_t (KeyArray_S01reg_gff_1_SFF_5_QD), .B0_t (enKS), .Z0_t (KeyArray_S01reg_gff_1_SFF_5_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS02ser[5]), .B0_t (KeyArray_outS11ser[5]), .Z0_t (KeyArray_S01reg_gff_1_SFF_5_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S01reg_gff_1_SFF_5_MUXInst_X), .Z0_t (KeyArray_S01reg_gff_1_SFF_5_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S01reg_gff_1_SFF_5_MUXInst_Y), .B0_t (KeyArray_outS02ser[5]), .Z0_t (KeyArray_S01reg_gff_1_SFF_5_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S01reg_gff_1_SFF_6_U3 ( .A0_t (KeyArray_S01reg_gff_1_SFF_6_n2), .B0_t (KeyArray_S01reg_gff_1_SFF_6_n1), .Z0_t (KeyArray_outS01ser_6_) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_6_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS01ser_6_), .Z0_t (KeyArray_S01reg_gff_1_SFF_6_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_6_U1 ( .A0_t (KeyArray_S01reg_gff_1_SFF_6_QD), .B0_t (enKS), .Z0_t (KeyArray_S01reg_gff_1_SFF_6_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS02ser[6]), .B0_t (KeyArray_outS11ser[6]), .Z0_t (KeyArray_S01reg_gff_1_SFF_6_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S01reg_gff_1_SFF_6_MUXInst_X), .Z0_t (KeyArray_S01reg_gff_1_SFF_6_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S01reg_gff_1_SFF_6_MUXInst_Y), .B0_t (KeyArray_outS02ser[6]), .Z0_t (KeyArray_S01reg_gff_1_SFF_6_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S01reg_gff_1_SFF_7_U3 ( .A0_t (KeyArray_S01reg_gff_1_SFF_7_n2), .B0_t (KeyArray_S01reg_gff_1_SFF_7_n1), .Z0_t (KeyArray_outS01ser_7_) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_7_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS01ser_7_), .Z0_t (KeyArray_S01reg_gff_1_SFF_7_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_7_U1 ( .A0_t (KeyArray_S01reg_gff_1_SFF_7_QD), .B0_t (enKS), .Z0_t (KeyArray_S01reg_gff_1_SFF_7_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS02ser[7]), .B0_t (KeyArray_outS11ser[7]), .Z0_t (KeyArray_S01reg_gff_1_SFF_7_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S01reg_gff_1_SFF_7_MUXInst_X), .Z0_t (KeyArray_S01reg_gff_1_SFF_7_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S01reg_gff_1_SFF_7_MUXInst_Y), .B0_t (KeyArray_outS02ser[7]), .Z0_t (KeyArray_S01reg_gff_1_SFF_7_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S02reg_gff_1_SFF_0_U3 ( .A0_t (KeyArray_S02reg_gff_1_SFF_0_n2), .B0_t (KeyArray_S02reg_gff_1_SFF_0_n1), .Z0_t (KeyArray_outS02ser[0]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_0_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS02ser[0]), .Z0_t (KeyArray_S02reg_gff_1_SFF_0_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_0_U1 ( .A0_t (KeyArray_S02reg_gff_1_SFF_0_QD), .B0_t (enKS), .Z0_t (KeyArray_S02reg_gff_1_SFF_0_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS03ser[0]), .B0_t (KeyArray_outS12ser[0]), .Z0_t (KeyArray_S02reg_gff_1_SFF_0_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S02reg_gff_1_SFF_0_MUXInst_X), .Z0_t (KeyArray_S02reg_gff_1_SFF_0_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S02reg_gff_1_SFF_0_MUXInst_Y), .B0_t (KeyArray_outS03ser[0]), .Z0_t (KeyArray_S02reg_gff_1_SFF_0_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S02reg_gff_1_SFF_1_U3 ( .A0_t (KeyArray_S02reg_gff_1_SFF_1_n2), .B0_t (KeyArray_S02reg_gff_1_SFF_1_n1), .Z0_t (KeyArray_outS02ser[1]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_1_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS02ser[1]), .Z0_t (KeyArray_S02reg_gff_1_SFF_1_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_1_U1 ( .A0_t (KeyArray_S02reg_gff_1_SFF_1_QD), .B0_t (enKS), .Z0_t (KeyArray_S02reg_gff_1_SFF_1_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS03ser[1]), .B0_t (KeyArray_outS12ser[1]), .Z0_t (KeyArray_S02reg_gff_1_SFF_1_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S02reg_gff_1_SFF_1_MUXInst_X), .Z0_t (KeyArray_S02reg_gff_1_SFF_1_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S02reg_gff_1_SFF_1_MUXInst_Y), .B0_t (KeyArray_outS03ser[1]), .Z0_t (KeyArray_S02reg_gff_1_SFF_1_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S02reg_gff_1_SFF_2_U3 ( .A0_t (KeyArray_S02reg_gff_1_SFF_2_n2), .B0_t (KeyArray_S02reg_gff_1_SFF_2_n1), .Z0_t (KeyArray_outS02ser[2]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_2_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS02ser[2]), .Z0_t (KeyArray_S02reg_gff_1_SFF_2_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_2_U1 ( .A0_t (KeyArray_S02reg_gff_1_SFF_2_QD), .B0_t (enKS), .Z0_t (KeyArray_S02reg_gff_1_SFF_2_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS03ser[2]), .B0_t (KeyArray_outS12ser[2]), .Z0_t (KeyArray_S02reg_gff_1_SFF_2_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S02reg_gff_1_SFF_2_MUXInst_X), .Z0_t (KeyArray_S02reg_gff_1_SFF_2_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S02reg_gff_1_SFF_2_MUXInst_Y), .B0_t (KeyArray_outS03ser[2]), .Z0_t (KeyArray_S02reg_gff_1_SFF_2_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S02reg_gff_1_SFF_3_U3 ( .A0_t (KeyArray_S02reg_gff_1_SFF_3_n2), .B0_t (KeyArray_S02reg_gff_1_SFF_3_n1), .Z0_t (KeyArray_outS02ser[3]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_3_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS02ser[3]), .Z0_t (KeyArray_S02reg_gff_1_SFF_3_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_3_U1 ( .A0_t (KeyArray_S02reg_gff_1_SFF_3_QD), .B0_t (enKS), .Z0_t (KeyArray_S02reg_gff_1_SFF_3_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS03ser[3]), .B0_t (KeyArray_outS12ser[3]), .Z0_t (KeyArray_S02reg_gff_1_SFF_3_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S02reg_gff_1_SFF_3_MUXInst_X), .Z0_t (KeyArray_S02reg_gff_1_SFF_3_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S02reg_gff_1_SFF_3_MUXInst_Y), .B0_t (KeyArray_outS03ser[3]), .Z0_t (KeyArray_S02reg_gff_1_SFF_3_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S02reg_gff_1_SFF_4_U3 ( .A0_t (KeyArray_S02reg_gff_1_SFF_4_n2), .B0_t (KeyArray_S02reg_gff_1_SFF_4_n1), .Z0_t (KeyArray_outS02ser[4]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_4_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS02ser[4]), .Z0_t (KeyArray_S02reg_gff_1_SFF_4_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_4_U1 ( .A0_t (KeyArray_S02reg_gff_1_SFF_4_QD), .B0_t (enKS), .Z0_t (KeyArray_S02reg_gff_1_SFF_4_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS03ser[4]), .B0_t (KeyArray_outS12ser[4]), .Z0_t (KeyArray_S02reg_gff_1_SFF_4_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S02reg_gff_1_SFF_4_MUXInst_X), .Z0_t (KeyArray_S02reg_gff_1_SFF_4_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S02reg_gff_1_SFF_4_MUXInst_Y), .B0_t (KeyArray_outS03ser[4]), .Z0_t (KeyArray_S02reg_gff_1_SFF_4_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S02reg_gff_1_SFF_5_U3 ( .A0_t (KeyArray_S02reg_gff_1_SFF_5_n2), .B0_t (KeyArray_S02reg_gff_1_SFF_5_n1), .Z0_t (KeyArray_outS02ser[5]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_5_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS02ser[5]), .Z0_t (KeyArray_S02reg_gff_1_SFF_5_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_5_U1 ( .A0_t (KeyArray_S02reg_gff_1_SFF_5_QD), .B0_t (enKS), .Z0_t (KeyArray_S02reg_gff_1_SFF_5_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS03ser[5]), .B0_t (KeyArray_outS12ser[5]), .Z0_t (KeyArray_S02reg_gff_1_SFF_5_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S02reg_gff_1_SFF_5_MUXInst_X), .Z0_t (KeyArray_S02reg_gff_1_SFF_5_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S02reg_gff_1_SFF_5_MUXInst_Y), .B0_t (KeyArray_outS03ser[5]), .Z0_t (KeyArray_S02reg_gff_1_SFF_5_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S02reg_gff_1_SFF_6_U3 ( .A0_t (KeyArray_S02reg_gff_1_SFF_6_n2), .B0_t (KeyArray_S02reg_gff_1_SFF_6_n1), .Z0_t (KeyArray_outS02ser[6]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_6_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS02ser[6]), .Z0_t (KeyArray_S02reg_gff_1_SFF_6_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_6_U1 ( .A0_t (KeyArray_S02reg_gff_1_SFF_6_QD), .B0_t (enKS), .Z0_t (KeyArray_S02reg_gff_1_SFF_6_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS03ser[6]), .B0_t (KeyArray_outS12ser[6]), .Z0_t (KeyArray_S02reg_gff_1_SFF_6_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S02reg_gff_1_SFF_6_MUXInst_X), .Z0_t (KeyArray_S02reg_gff_1_SFF_6_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S02reg_gff_1_SFF_6_MUXInst_Y), .B0_t (KeyArray_outS03ser[6]), .Z0_t (KeyArray_S02reg_gff_1_SFF_6_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S02reg_gff_1_SFF_7_U3 ( .A0_t (KeyArray_S02reg_gff_1_SFF_7_n2), .B0_t (KeyArray_S02reg_gff_1_SFF_7_n1), .Z0_t (KeyArray_outS02ser[7]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_7_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS02ser[7]), .Z0_t (KeyArray_S02reg_gff_1_SFF_7_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_7_U1 ( .A0_t (KeyArray_S02reg_gff_1_SFF_7_QD), .B0_t (enKS), .Z0_t (KeyArray_S02reg_gff_1_SFF_7_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS03ser[7]), .B0_t (KeyArray_outS12ser[7]), .Z0_t (KeyArray_S02reg_gff_1_SFF_7_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S02reg_gff_1_SFF_7_MUXInst_X), .Z0_t (KeyArray_S02reg_gff_1_SFF_7_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S02reg_gff_1_SFF_7_MUXInst_Y), .B0_t (KeyArray_outS03ser[7]), .Z0_t (KeyArray_S02reg_gff_1_SFF_7_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S03reg_gff_1_SFF_0_U3 ( .A0_t (KeyArray_S03reg_gff_1_SFF_0_n2), .B0_t (KeyArray_S03reg_gff_1_SFF_0_n1), .Z0_t (KeyArray_outS03ser[0]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_0_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS03ser[0]), .Z0_t (KeyArray_S03reg_gff_1_SFF_0_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_0_U1 ( .A0_t (KeyArray_S03reg_gff_1_SFF_0_QD), .B0_t (enKS), .Z0_t (KeyArray_S03reg_gff_1_SFF_0_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS10ser[0]), .B0_t (keySBIn[0]), .Z0_t (KeyArray_S03reg_gff_1_SFF_0_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S03reg_gff_1_SFF_0_MUXInst_X), .Z0_t (KeyArray_S03reg_gff_1_SFF_0_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S03reg_gff_1_SFF_0_MUXInst_Y), .B0_t (KeyArray_outS10ser[0]), .Z0_t (KeyArray_S03reg_gff_1_SFF_0_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S03reg_gff_1_SFF_1_U3 ( .A0_t (KeyArray_S03reg_gff_1_SFF_1_n2), .B0_t (KeyArray_S03reg_gff_1_SFF_1_n1), .Z0_t (KeyArray_outS03ser[1]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_1_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS03ser[1]), .Z0_t (KeyArray_S03reg_gff_1_SFF_1_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_1_U1 ( .A0_t (KeyArray_S03reg_gff_1_SFF_1_QD), .B0_t (enKS), .Z0_t (KeyArray_S03reg_gff_1_SFF_1_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS10ser[1]), .B0_t (keySBIn[1]), .Z0_t (KeyArray_S03reg_gff_1_SFF_1_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S03reg_gff_1_SFF_1_MUXInst_X), .Z0_t (KeyArray_S03reg_gff_1_SFF_1_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S03reg_gff_1_SFF_1_MUXInst_Y), .B0_t (KeyArray_outS10ser[1]), .Z0_t (KeyArray_S03reg_gff_1_SFF_1_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S03reg_gff_1_SFF_2_U3 ( .A0_t (KeyArray_S03reg_gff_1_SFF_2_n2), .B0_t (KeyArray_S03reg_gff_1_SFF_2_n1), .Z0_t (KeyArray_outS03ser[2]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_2_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS03ser[2]), .Z0_t (KeyArray_S03reg_gff_1_SFF_2_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_2_U1 ( .A0_t (KeyArray_S03reg_gff_1_SFF_2_QD), .B0_t (enKS), .Z0_t (KeyArray_S03reg_gff_1_SFF_2_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS10ser[2]), .B0_t (keySBIn[2]), .Z0_t (KeyArray_S03reg_gff_1_SFF_2_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S03reg_gff_1_SFF_2_MUXInst_X), .Z0_t (KeyArray_S03reg_gff_1_SFF_2_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S03reg_gff_1_SFF_2_MUXInst_Y), .B0_t (KeyArray_outS10ser[2]), .Z0_t (KeyArray_S03reg_gff_1_SFF_2_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S03reg_gff_1_SFF_3_U3 ( .A0_t (KeyArray_S03reg_gff_1_SFF_3_n2), .B0_t (KeyArray_S03reg_gff_1_SFF_3_n1), .Z0_t (KeyArray_outS03ser[3]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_3_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS03ser[3]), .Z0_t (KeyArray_S03reg_gff_1_SFF_3_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_3_U1 ( .A0_t (KeyArray_S03reg_gff_1_SFF_3_QD), .B0_t (enKS), .Z0_t (KeyArray_S03reg_gff_1_SFF_3_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS10ser[3]), .B0_t (keySBIn[3]), .Z0_t (KeyArray_S03reg_gff_1_SFF_3_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S03reg_gff_1_SFF_3_MUXInst_X), .Z0_t (KeyArray_S03reg_gff_1_SFF_3_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S03reg_gff_1_SFF_3_MUXInst_Y), .B0_t (KeyArray_outS10ser[3]), .Z0_t (KeyArray_S03reg_gff_1_SFF_3_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S03reg_gff_1_SFF_4_U3 ( .A0_t (KeyArray_S03reg_gff_1_SFF_4_n2), .B0_t (KeyArray_S03reg_gff_1_SFF_4_n1), .Z0_t (KeyArray_outS03ser[4]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_4_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS03ser[4]), .Z0_t (KeyArray_S03reg_gff_1_SFF_4_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_4_U1 ( .A0_t (KeyArray_S03reg_gff_1_SFF_4_QD), .B0_t (enKS), .Z0_t (KeyArray_S03reg_gff_1_SFF_4_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS10ser[4]), .B0_t (keySBIn[4]), .Z0_t (KeyArray_S03reg_gff_1_SFF_4_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S03reg_gff_1_SFF_4_MUXInst_X), .Z0_t (KeyArray_S03reg_gff_1_SFF_4_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S03reg_gff_1_SFF_4_MUXInst_Y), .B0_t (KeyArray_outS10ser[4]), .Z0_t (KeyArray_S03reg_gff_1_SFF_4_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S03reg_gff_1_SFF_5_U3 ( .A0_t (KeyArray_S03reg_gff_1_SFF_5_n2), .B0_t (KeyArray_S03reg_gff_1_SFF_5_n1), .Z0_t (KeyArray_outS03ser[5]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_5_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS03ser[5]), .Z0_t (KeyArray_S03reg_gff_1_SFF_5_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_5_U1 ( .A0_t (KeyArray_S03reg_gff_1_SFF_5_QD), .B0_t (enKS), .Z0_t (KeyArray_S03reg_gff_1_SFF_5_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS10ser[5]), .B0_t (keySBIn[5]), .Z0_t (KeyArray_S03reg_gff_1_SFF_5_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S03reg_gff_1_SFF_5_MUXInst_X), .Z0_t (KeyArray_S03reg_gff_1_SFF_5_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S03reg_gff_1_SFF_5_MUXInst_Y), .B0_t (KeyArray_outS10ser[5]), .Z0_t (KeyArray_S03reg_gff_1_SFF_5_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S03reg_gff_1_SFF_6_U3 ( .A0_t (KeyArray_S03reg_gff_1_SFF_6_n2), .B0_t (KeyArray_S03reg_gff_1_SFF_6_n1), .Z0_t (KeyArray_outS03ser[6]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_6_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS03ser[6]), .Z0_t (KeyArray_S03reg_gff_1_SFF_6_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_6_U1 ( .A0_t (KeyArray_S03reg_gff_1_SFF_6_QD), .B0_t (enKS), .Z0_t (KeyArray_S03reg_gff_1_SFF_6_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS10ser[6]), .B0_t (keySBIn[6]), .Z0_t (KeyArray_S03reg_gff_1_SFF_6_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S03reg_gff_1_SFF_6_MUXInst_X), .Z0_t (KeyArray_S03reg_gff_1_SFF_6_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S03reg_gff_1_SFF_6_MUXInst_Y), .B0_t (KeyArray_outS10ser[6]), .Z0_t (KeyArray_S03reg_gff_1_SFF_6_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S03reg_gff_1_SFF_7_U3 ( .A0_t (KeyArray_S03reg_gff_1_SFF_7_n2), .B0_t (KeyArray_S03reg_gff_1_SFF_7_n1), .Z0_t (KeyArray_outS03ser[7]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_7_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS03ser[7]), .Z0_t (KeyArray_S03reg_gff_1_SFF_7_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_7_U1 ( .A0_t (KeyArray_S03reg_gff_1_SFF_7_QD), .B0_t (enKS), .Z0_t (KeyArray_S03reg_gff_1_SFF_7_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS10ser[7]), .B0_t (keySBIn[7]), .Z0_t (KeyArray_S03reg_gff_1_SFF_7_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S03reg_gff_1_SFF_7_MUXInst_X), .Z0_t (KeyArray_S03reg_gff_1_SFF_7_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S03reg_gff_1_SFF_7_MUXInst_Y), .B0_t (KeyArray_outS10ser[7]), .Z0_t (KeyArray_S03reg_gff_1_SFF_7_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S10reg_gff_1_SFF_0_U3 ( .A0_t (KeyArray_S10reg_gff_1_SFF_0_n2), .B0_t (KeyArray_S10reg_gff_1_SFF_0_n1), .Z0_t (KeyArray_outS10ser[0]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_0_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS10ser[0]), .Z0_t (KeyArray_S10reg_gff_1_SFF_0_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_0_U1 ( .A0_t (KeyArray_S10reg_gff_1_SFF_0_QD), .B0_t (enKS), .Z0_t (KeyArray_S10reg_gff_1_SFF_0_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS11ser[0]), .B0_t (KeyArray_outS20ser[0]), .Z0_t (KeyArray_S10reg_gff_1_SFF_0_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S10reg_gff_1_SFF_0_MUXInst_X), .Z0_t (KeyArray_S10reg_gff_1_SFF_0_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S10reg_gff_1_SFF_0_MUXInst_Y), .B0_t (KeyArray_outS11ser[0]), .Z0_t (KeyArray_S10reg_gff_1_SFF_0_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S10reg_gff_1_SFF_1_U3 ( .A0_t (KeyArray_S10reg_gff_1_SFF_1_n2), .B0_t (KeyArray_S10reg_gff_1_SFF_1_n1), .Z0_t (KeyArray_outS10ser[1]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_1_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS10ser[1]), .Z0_t (KeyArray_S10reg_gff_1_SFF_1_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_1_U1 ( .A0_t (KeyArray_S10reg_gff_1_SFF_1_QD), .B0_t (enKS), .Z0_t (KeyArray_S10reg_gff_1_SFF_1_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS11ser[1]), .B0_t (KeyArray_outS20ser[1]), .Z0_t (KeyArray_S10reg_gff_1_SFF_1_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S10reg_gff_1_SFF_1_MUXInst_X), .Z0_t (KeyArray_S10reg_gff_1_SFF_1_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S10reg_gff_1_SFF_1_MUXInst_Y), .B0_t (KeyArray_outS11ser[1]), .Z0_t (KeyArray_S10reg_gff_1_SFF_1_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S10reg_gff_1_SFF_2_U3 ( .A0_t (KeyArray_S10reg_gff_1_SFF_2_n2), .B0_t (KeyArray_S10reg_gff_1_SFF_2_n1), .Z0_t (KeyArray_outS10ser[2]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_2_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS10ser[2]), .Z0_t (KeyArray_S10reg_gff_1_SFF_2_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_2_U1 ( .A0_t (KeyArray_S10reg_gff_1_SFF_2_QD), .B0_t (enKS), .Z0_t (KeyArray_S10reg_gff_1_SFF_2_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS11ser[2]), .B0_t (KeyArray_outS20ser[2]), .Z0_t (KeyArray_S10reg_gff_1_SFF_2_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S10reg_gff_1_SFF_2_MUXInst_X), .Z0_t (KeyArray_S10reg_gff_1_SFF_2_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S10reg_gff_1_SFF_2_MUXInst_Y), .B0_t (KeyArray_outS11ser[2]), .Z0_t (KeyArray_S10reg_gff_1_SFF_2_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S10reg_gff_1_SFF_3_U3 ( .A0_t (KeyArray_S10reg_gff_1_SFF_3_n2), .B0_t (KeyArray_S10reg_gff_1_SFF_3_n1), .Z0_t (KeyArray_outS10ser[3]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_3_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS10ser[3]), .Z0_t (KeyArray_S10reg_gff_1_SFF_3_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_3_U1 ( .A0_t (KeyArray_S10reg_gff_1_SFF_3_QD), .B0_t (enKS), .Z0_t (KeyArray_S10reg_gff_1_SFF_3_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS11ser[3]), .B0_t (KeyArray_outS20ser[3]), .Z0_t (KeyArray_S10reg_gff_1_SFF_3_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S10reg_gff_1_SFF_3_MUXInst_X), .Z0_t (KeyArray_S10reg_gff_1_SFF_3_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S10reg_gff_1_SFF_3_MUXInst_Y), .B0_t (KeyArray_outS11ser[3]), .Z0_t (KeyArray_S10reg_gff_1_SFF_3_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S10reg_gff_1_SFF_4_U3 ( .A0_t (KeyArray_S10reg_gff_1_SFF_4_n2), .B0_t (KeyArray_S10reg_gff_1_SFF_4_n1), .Z0_t (KeyArray_outS10ser[4]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_4_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS10ser[4]), .Z0_t (KeyArray_S10reg_gff_1_SFF_4_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_4_U1 ( .A0_t (KeyArray_S10reg_gff_1_SFF_4_QD), .B0_t (enKS), .Z0_t (KeyArray_S10reg_gff_1_SFF_4_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS11ser[4]), .B0_t (KeyArray_outS20ser[4]), .Z0_t (KeyArray_S10reg_gff_1_SFF_4_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S10reg_gff_1_SFF_4_MUXInst_X), .Z0_t (KeyArray_S10reg_gff_1_SFF_4_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S10reg_gff_1_SFF_4_MUXInst_Y), .B0_t (KeyArray_outS11ser[4]), .Z0_t (KeyArray_S10reg_gff_1_SFF_4_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S10reg_gff_1_SFF_5_U3 ( .A0_t (KeyArray_S10reg_gff_1_SFF_5_n2), .B0_t (KeyArray_S10reg_gff_1_SFF_5_n1), .Z0_t (KeyArray_outS10ser[5]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_5_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS10ser[5]), .Z0_t (KeyArray_S10reg_gff_1_SFF_5_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_5_U1 ( .A0_t (KeyArray_S10reg_gff_1_SFF_5_QD), .B0_t (enKS), .Z0_t (KeyArray_S10reg_gff_1_SFF_5_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS11ser[5]), .B0_t (KeyArray_outS20ser[5]), .Z0_t (KeyArray_S10reg_gff_1_SFF_5_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S10reg_gff_1_SFF_5_MUXInst_X), .Z0_t (KeyArray_S10reg_gff_1_SFF_5_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S10reg_gff_1_SFF_5_MUXInst_Y), .B0_t (KeyArray_outS11ser[5]), .Z0_t (KeyArray_S10reg_gff_1_SFF_5_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S10reg_gff_1_SFF_6_U3 ( .A0_t (KeyArray_S10reg_gff_1_SFF_6_n2), .B0_t (KeyArray_S10reg_gff_1_SFF_6_n1), .Z0_t (KeyArray_outS10ser[6]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_6_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS10ser[6]), .Z0_t (KeyArray_S10reg_gff_1_SFF_6_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_6_U1 ( .A0_t (KeyArray_S10reg_gff_1_SFF_6_QD), .B0_t (enKS), .Z0_t (KeyArray_S10reg_gff_1_SFF_6_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS11ser[6]), .B0_t (KeyArray_outS20ser[6]), .Z0_t (KeyArray_S10reg_gff_1_SFF_6_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S10reg_gff_1_SFF_6_MUXInst_X), .Z0_t (KeyArray_S10reg_gff_1_SFF_6_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S10reg_gff_1_SFF_6_MUXInst_Y), .B0_t (KeyArray_outS11ser[6]), .Z0_t (KeyArray_S10reg_gff_1_SFF_6_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S10reg_gff_1_SFF_7_U3 ( .A0_t (KeyArray_S10reg_gff_1_SFF_7_n2), .B0_t (KeyArray_S10reg_gff_1_SFF_7_n1), .Z0_t (KeyArray_outS10ser[7]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_7_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS10ser[7]), .Z0_t (KeyArray_S10reg_gff_1_SFF_7_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_7_U1 ( .A0_t (KeyArray_S10reg_gff_1_SFF_7_QD), .B0_t (enKS), .Z0_t (KeyArray_S10reg_gff_1_SFF_7_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS11ser[7]), .B0_t (KeyArray_outS20ser[7]), .Z0_t (KeyArray_S10reg_gff_1_SFF_7_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S10reg_gff_1_SFF_7_MUXInst_X), .Z0_t (KeyArray_S10reg_gff_1_SFF_7_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S10reg_gff_1_SFF_7_MUXInst_Y), .B0_t (KeyArray_outS11ser[7]), .Z0_t (KeyArray_S10reg_gff_1_SFF_7_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S11reg_gff_1_SFF_0_U3 ( .A0_t (KeyArray_S11reg_gff_1_SFF_0_n2), .B0_t (KeyArray_S11reg_gff_1_SFF_0_n1), .Z0_t (KeyArray_outS11ser[0]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_0_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS11ser[0]), .Z0_t (KeyArray_S11reg_gff_1_SFF_0_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_0_U1 ( .A0_t (KeyArray_S11reg_gff_1_SFF_0_QD), .B0_t (enKS), .Z0_t (KeyArray_S11reg_gff_1_SFF_0_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS12ser[0]), .B0_t (KeyArray_outS21ser[0]), .Z0_t (KeyArray_S11reg_gff_1_SFF_0_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S11reg_gff_1_SFF_0_MUXInst_X), .Z0_t (KeyArray_S11reg_gff_1_SFF_0_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S11reg_gff_1_SFF_0_MUXInst_Y), .B0_t (KeyArray_outS12ser[0]), .Z0_t (KeyArray_S11reg_gff_1_SFF_0_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S11reg_gff_1_SFF_1_U3 ( .A0_t (KeyArray_S11reg_gff_1_SFF_1_n2), .B0_t (KeyArray_S11reg_gff_1_SFF_1_n1), .Z0_t (KeyArray_outS11ser[1]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_1_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS11ser[1]), .Z0_t (KeyArray_S11reg_gff_1_SFF_1_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_1_U1 ( .A0_t (KeyArray_S11reg_gff_1_SFF_1_QD), .B0_t (enKS), .Z0_t (KeyArray_S11reg_gff_1_SFF_1_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS12ser[1]), .B0_t (KeyArray_outS21ser[1]), .Z0_t (KeyArray_S11reg_gff_1_SFF_1_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S11reg_gff_1_SFF_1_MUXInst_X), .Z0_t (KeyArray_S11reg_gff_1_SFF_1_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S11reg_gff_1_SFF_1_MUXInst_Y), .B0_t (KeyArray_outS12ser[1]), .Z0_t (KeyArray_S11reg_gff_1_SFF_1_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S11reg_gff_1_SFF_2_U3 ( .A0_t (KeyArray_S11reg_gff_1_SFF_2_n2), .B0_t (KeyArray_S11reg_gff_1_SFF_2_n1), .Z0_t (KeyArray_outS11ser[2]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_2_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS11ser[2]), .Z0_t (KeyArray_S11reg_gff_1_SFF_2_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_2_U1 ( .A0_t (KeyArray_S11reg_gff_1_SFF_2_QD), .B0_t (enKS), .Z0_t (KeyArray_S11reg_gff_1_SFF_2_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS12ser[2]), .B0_t (KeyArray_outS21ser[2]), .Z0_t (KeyArray_S11reg_gff_1_SFF_2_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S11reg_gff_1_SFF_2_MUXInst_X), .Z0_t (KeyArray_S11reg_gff_1_SFF_2_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S11reg_gff_1_SFF_2_MUXInst_Y), .B0_t (KeyArray_outS12ser[2]), .Z0_t (KeyArray_S11reg_gff_1_SFF_2_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S11reg_gff_1_SFF_3_U3 ( .A0_t (KeyArray_S11reg_gff_1_SFF_3_n2), .B0_t (KeyArray_S11reg_gff_1_SFF_3_n1), .Z0_t (KeyArray_outS11ser[3]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_3_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS11ser[3]), .Z0_t (KeyArray_S11reg_gff_1_SFF_3_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_3_U1 ( .A0_t (KeyArray_S11reg_gff_1_SFF_3_QD), .B0_t (enKS), .Z0_t (KeyArray_S11reg_gff_1_SFF_3_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS12ser[3]), .B0_t (KeyArray_outS21ser[3]), .Z0_t (KeyArray_S11reg_gff_1_SFF_3_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S11reg_gff_1_SFF_3_MUXInst_X), .Z0_t (KeyArray_S11reg_gff_1_SFF_3_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S11reg_gff_1_SFF_3_MUXInst_Y), .B0_t (KeyArray_outS12ser[3]), .Z0_t (KeyArray_S11reg_gff_1_SFF_3_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S11reg_gff_1_SFF_4_U3 ( .A0_t (KeyArray_S11reg_gff_1_SFF_4_n2), .B0_t (KeyArray_S11reg_gff_1_SFF_4_n1), .Z0_t (KeyArray_outS11ser[4]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_4_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS11ser[4]), .Z0_t (KeyArray_S11reg_gff_1_SFF_4_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_4_U1 ( .A0_t (KeyArray_S11reg_gff_1_SFF_4_QD), .B0_t (enKS), .Z0_t (KeyArray_S11reg_gff_1_SFF_4_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS12ser[4]), .B0_t (KeyArray_outS21ser[4]), .Z0_t (KeyArray_S11reg_gff_1_SFF_4_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S11reg_gff_1_SFF_4_MUXInst_X), .Z0_t (KeyArray_S11reg_gff_1_SFF_4_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S11reg_gff_1_SFF_4_MUXInst_Y), .B0_t (KeyArray_outS12ser[4]), .Z0_t (KeyArray_S11reg_gff_1_SFF_4_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S11reg_gff_1_SFF_5_U3 ( .A0_t (KeyArray_S11reg_gff_1_SFF_5_n2), .B0_t (KeyArray_S11reg_gff_1_SFF_5_n1), .Z0_t (KeyArray_outS11ser[5]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_5_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS11ser[5]), .Z0_t (KeyArray_S11reg_gff_1_SFF_5_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_5_U1 ( .A0_t (KeyArray_S11reg_gff_1_SFF_5_QD), .B0_t (enKS), .Z0_t (KeyArray_S11reg_gff_1_SFF_5_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS12ser[5]), .B0_t (KeyArray_outS21ser[5]), .Z0_t (KeyArray_S11reg_gff_1_SFF_5_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S11reg_gff_1_SFF_5_MUXInst_X), .Z0_t (KeyArray_S11reg_gff_1_SFF_5_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S11reg_gff_1_SFF_5_MUXInst_Y), .B0_t (KeyArray_outS12ser[5]), .Z0_t (KeyArray_S11reg_gff_1_SFF_5_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S11reg_gff_1_SFF_6_U3 ( .A0_t (KeyArray_S11reg_gff_1_SFF_6_n2), .B0_t (KeyArray_S11reg_gff_1_SFF_6_n1), .Z0_t (KeyArray_outS11ser[6]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_6_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS11ser[6]), .Z0_t (KeyArray_S11reg_gff_1_SFF_6_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_6_U1 ( .A0_t (KeyArray_S11reg_gff_1_SFF_6_QD), .B0_t (enKS), .Z0_t (KeyArray_S11reg_gff_1_SFF_6_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS12ser[6]), .B0_t (KeyArray_outS21ser[6]), .Z0_t (KeyArray_S11reg_gff_1_SFF_6_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S11reg_gff_1_SFF_6_MUXInst_X), .Z0_t (KeyArray_S11reg_gff_1_SFF_6_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S11reg_gff_1_SFF_6_MUXInst_Y), .B0_t (KeyArray_outS12ser[6]), .Z0_t (KeyArray_S11reg_gff_1_SFF_6_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S11reg_gff_1_SFF_7_U3 ( .A0_t (KeyArray_S11reg_gff_1_SFF_7_n2), .B0_t (KeyArray_S11reg_gff_1_SFF_7_n1), .Z0_t (KeyArray_outS11ser[7]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_7_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS11ser[7]), .Z0_t (KeyArray_S11reg_gff_1_SFF_7_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_7_U1 ( .A0_t (KeyArray_S11reg_gff_1_SFF_7_QD), .B0_t (enKS), .Z0_t (KeyArray_S11reg_gff_1_SFF_7_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS12ser[7]), .B0_t (KeyArray_outS21ser[7]), .Z0_t (KeyArray_S11reg_gff_1_SFF_7_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S11reg_gff_1_SFF_7_MUXInst_X), .Z0_t (KeyArray_S11reg_gff_1_SFF_7_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S11reg_gff_1_SFF_7_MUXInst_Y), .B0_t (KeyArray_outS12ser[7]), .Z0_t (KeyArray_S11reg_gff_1_SFF_7_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S12reg_gff_1_SFF_0_U3 ( .A0_t (KeyArray_S12reg_gff_1_SFF_0_n2), .B0_t (KeyArray_S12reg_gff_1_SFF_0_n1), .Z0_t (KeyArray_outS12ser[0]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_0_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS12ser[0]), .Z0_t (KeyArray_S12reg_gff_1_SFF_0_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_0_U1 ( .A0_t (KeyArray_S12reg_gff_1_SFF_0_QD), .B0_t (enKS), .Z0_t (KeyArray_S12reg_gff_1_SFF_0_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (keySBIn[0]), .B0_t (KeyArray_outS22ser[0]), .Z0_t (KeyArray_S12reg_gff_1_SFF_0_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S12reg_gff_1_SFF_0_MUXInst_X), .Z0_t (KeyArray_S12reg_gff_1_SFF_0_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S12reg_gff_1_SFF_0_MUXInst_Y), .B0_t (keySBIn[0]), .Z0_t (KeyArray_S12reg_gff_1_SFF_0_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S12reg_gff_1_SFF_1_U3 ( .A0_t (KeyArray_S12reg_gff_1_SFF_1_n2), .B0_t (KeyArray_S12reg_gff_1_SFF_1_n1), .Z0_t (KeyArray_outS12ser[1]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_1_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS12ser[1]), .Z0_t (KeyArray_S12reg_gff_1_SFF_1_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_1_U1 ( .A0_t (KeyArray_S12reg_gff_1_SFF_1_QD), .B0_t (enKS), .Z0_t (KeyArray_S12reg_gff_1_SFF_1_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (keySBIn[1]), .B0_t (KeyArray_outS22ser[1]), .Z0_t (KeyArray_S12reg_gff_1_SFF_1_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S12reg_gff_1_SFF_1_MUXInst_X), .Z0_t (KeyArray_S12reg_gff_1_SFF_1_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S12reg_gff_1_SFF_1_MUXInst_Y), .B0_t (keySBIn[1]), .Z0_t (KeyArray_S12reg_gff_1_SFF_1_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S12reg_gff_1_SFF_2_U3 ( .A0_t (KeyArray_S12reg_gff_1_SFF_2_n2), .B0_t (KeyArray_S12reg_gff_1_SFF_2_n1), .Z0_t (KeyArray_outS12ser[2]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_2_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS12ser[2]), .Z0_t (KeyArray_S12reg_gff_1_SFF_2_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_2_U1 ( .A0_t (KeyArray_S12reg_gff_1_SFF_2_QD), .B0_t (enKS), .Z0_t (KeyArray_S12reg_gff_1_SFF_2_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (keySBIn[2]), .B0_t (KeyArray_outS22ser[2]), .Z0_t (KeyArray_S12reg_gff_1_SFF_2_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S12reg_gff_1_SFF_2_MUXInst_X), .Z0_t (KeyArray_S12reg_gff_1_SFF_2_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S12reg_gff_1_SFF_2_MUXInst_Y), .B0_t (keySBIn[2]), .Z0_t (KeyArray_S12reg_gff_1_SFF_2_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S12reg_gff_1_SFF_3_U3 ( .A0_t (KeyArray_S12reg_gff_1_SFF_3_n2), .B0_t (KeyArray_S12reg_gff_1_SFF_3_n1), .Z0_t (KeyArray_outS12ser[3]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_3_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS12ser[3]), .Z0_t (KeyArray_S12reg_gff_1_SFF_3_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_3_U1 ( .A0_t (KeyArray_S12reg_gff_1_SFF_3_QD), .B0_t (enKS), .Z0_t (KeyArray_S12reg_gff_1_SFF_3_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (keySBIn[3]), .B0_t (KeyArray_outS22ser[3]), .Z0_t (KeyArray_S12reg_gff_1_SFF_3_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S12reg_gff_1_SFF_3_MUXInst_X), .Z0_t (KeyArray_S12reg_gff_1_SFF_3_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S12reg_gff_1_SFF_3_MUXInst_Y), .B0_t (keySBIn[3]), .Z0_t (KeyArray_S12reg_gff_1_SFF_3_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S12reg_gff_1_SFF_4_U3 ( .A0_t (KeyArray_S12reg_gff_1_SFF_4_n2), .B0_t (KeyArray_S12reg_gff_1_SFF_4_n1), .Z0_t (KeyArray_outS12ser[4]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_4_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS12ser[4]), .Z0_t (KeyArray_S12reg_gff_1_SFF_4_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_4_U1 ( .A0_t (KeyArray_S12reg_gff_1_SFF_4_QD), .B0_t (enKS), .Z0_t (KeyArray_S12reg_gff_1_SFF_4_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (keySBIn[4]), .B0_t (KeyArray_outS22ser[4]), .Z0_t (KeyArray_S12reg_gff_1_SFF_4_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S12reg_gff_1_SFF_4_MUXInst_X), .Z0_t (KeyArray_S12reg_gff_1_SFF_4_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S12reg_gff_1_SFF_4_MUXInst_Y), .B0_t (keySBIn[4]), .Z0_t (KeyArray_S12reg_gff_1_SFF_4_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S12reg_gff_1_SFF_5_U3 ( .A0_t (KeyArray_S12reg_gff_1_SFF_5_n2), .B0_t (KeyArray_S12reg_gff_1_SFF_5_n1), .Z0_t (KeyArray_outS12ser[5]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_5_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS12ser[5]), .Z0_t (KeyArray_S12reg_gff_1_SFF_5_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_5_U1 ( .A0_t (KeyArray_S12reg_gff_1_SFF_5_QD), .B0_t (enKS), .Z0_t (KeyArray_S12reg_gff_1_SFF_5_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (keySBIn[5]), .B0_t (KeyArray_outS22ser[5]), .Z0_t (KeyArray_S12reg_gff_1_SFF_5_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S12reg_gff_1_SFF_5_MUXInst_X), .Z0_t (KeyArray_S12reg_gff_1_SFF_5_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S12reg_gff_1_SFF_5_MUXInst_Y), .B0_t (keySBIn[5]), .Z0_t (KeyArray_S12reg_gff_1_SFF_5_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S12reg_gff_1_SFF_6_U3 ( .A0_t (KeyArray_S12reg_gff_1_SFF_6_n2), .B0_t (KeyArray_S12reg_gff_1_SFF_6_n1), .Z0_t (KeyArray_outS12ser[6]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_6_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS12ser[6]), .Z0_t (KeyArray_S12reg_gff_1_SFF_6_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_6_U1 ( .A0_t (KeyArray_S12reg_gff_1_SFF_6_QD), .B0_t (enKS), .Z0_t (KeyArray_S12reg_gff_1_SFF_6_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (keySBIn[6]), .B0_t (KeyArray_outS22ser[6]), .Z0_t (KeyArray_S12reg_gff_1_SFF_6_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S12reg_gff_1_SFF_6_MUXInst_X), .Z0_t (KeyArray_S12reg_gff_1_SFF_6_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S12reg_gff_1_SFF_6_MUXInst_Y), .B0_t (keySBIn[6]), .Z0_t (KeyArray_S12reg_gff_1_SFF_6_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S12reg_gff_1_SFF_7_U3 ( .A0_t (KeyArray_S12reg_gff_1_SFF_7_n2), .B0_t (KeyArray_S12reg_gff_1_SFF_7_n1), .Z0_t (KeyArray_outS12ser[7]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_7_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS12ser[7]), .Z0_t (KeyArray_S12reg_gff_1_SFF_7_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_7_U1 ( .A0_t (KeyArray_S12reg_gff_1_SFF_7_QD), .B0_t (enKS), .Z0_t (KeyArray_S12reg_gff_1_SFF_7_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (keySBIn[7]), .B0_t (KeyArray_outS22ser[7]), .Z0_t (KeyArray_S12reg_gff_1_SFF_7_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S12reg_gff_1_SFF_7_MUXInst_X), .Z0_t (KeyArray_S12reg_gff_1_SFF_7_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S12reg_gff_1_SFF_7_MUXInst_Y), .B0_t (keySBIn[7]), .Z0_t (KeyArray_S12reg_gff_1_SFF_7_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S13reg_gff_1_SFF_0_U3 ( .A0_t (KeyArray_S13reg_gff_1_SFF_0_n2), .B0_t (KeyArray_S13reg_gff_1_SFF_0_n1), .Z0_t (keySBIn[0]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_0_U2 ( .A0_t (enKS), .B0_t (keySBIn[0]), .Z0_t (KeyArray_S13reg_gff_1_SFF_0_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_0_U1 ( .A0_t (KeyArray_S13reg_gff_1_SFF_0_QD), .B0_t (enKS), .Z0_t (KeyArray_S13reg_gff_1_SFF_0_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS20ser[0]), .B0_t (KeyArray_outS23ser[0]), .Z0_t (KeyArray_S13reg_gff_1_SFF_0_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S13reg_gff_1_SFF_0_MUXInst_X), .Z0_t (KeyArray_S13reg_gff_1_SFF_0_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S13reg_gff_1_SFF_0_MUXInst_Y), .B0_t (KeyArray_outS20ser[0]), .Z0_t (KeyArray_S13reg_gff_1_SFF_0_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S13reg_gff_1_SFF_1_U3 ( .A0_t (KeyArray_S13reg_gff_1_SFF_1_n2), .B0_t (KeyArray_S13reg_gff_1_SFF_1_n1), .Z0_t (keySBIn[1]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_1_U2 ( .A0_t (enKS), .B0_t (keySBIn[1]), .Z0_t (KeyArray_S13reg_gff_1_SFF_1_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_1_U1 ( .A0_t (KeyArray_S13reg_gff_1_SFF_1_QD), .B0_t (enKS), .Z0_t (KeyArray_S13reg_gff_1_SFF_1_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS20ser[1]), .B0_t (KeyArray_outS23ser[1]), .Z0_t (KeyArray_S13reg_gff_1_SFF_1_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S13reg_gff_1_SFF_1_MUXInst_X), .Z0_t (KeyArray_S13reg_gff_1_SFF_1_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S13reg_gff_1_SFF_1_MUXInst_Y), .B0_t (KeyArray_outS20ser[1]), .Z0_t (KeyArray_S13reg_gff_1_SFF_1_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S13reg_gff_1_SFF_2_U3 ( .A0_t (KeyArray_S13reg_gff_1_SFF_2_n2), .B0_t (KeyArray_S13reg_gff_1_SFF_2_n1), .Z0_t (keySBIn[2]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_2_U2 ( .A0_t (enKS), .B0_t (keySBIn[2]), .Z0_t (KeyArray_S13reg_gff_1_SFF_2_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_2_U1 ( .A0_t (KeyArray_S13reg_gff_1_SFF_2_QD), .B0_t (enKS), .Z0_t (KeyArray_S13reg_gff_1_SFF_2_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS20ser[2]), .B0_t (KeyArray_outS23ser[2]), .Z0_t (KeyArray_S13reg_gff_1_SFF_2_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S13reg_gff_1_SFF_2_MUXInst_X), .Z0_t (KeyArray_S13reg_gff_1_SFF_2_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S13reg_gff_1_SFF_2_MUXInst_Y), .B0_t (KeyArray_outS20ser[2]), .Z0_t (KeyArray_S13reg_gff_1_SFF_2_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S13reg_gff_1_SFF_3_U3 ( .A0_t (KeyArray_S13reg_gff_1_SFF_3_n2), .B0_t (KeyArray_S13reg_gff_1_SFF_3_n1), .Z0_t (keySBIn[3]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_3_U2 ( .A0_t (enKS), .B0_t (keySBIn[3]), .Z0_t (KeyArray_S13reg_gff_1_SFF_3_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_3_U1 ( .A0_t (KeyArray_S13reg_gff_1_SFF_3_QD), .B0_t (enKS), .Z0_t (KeyArray_S13reg_gff_1_SFF_3_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS20ser[3]), .B0_t (KeyArray_outS23ser[3]), .Z0_t (KeyArray_S13reg_gff_1_SFF_3_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S13reg_gff_1_SFF_3_MUXInst_X), .Z0_t (KeyArray_S13reg_gff_1_SFF_3_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S13reg_gff_1_SFF_3_MUXInst_Y), .B0_t (KeyArray_outS20ser[3]), .Z0_t (KeyArray_S13reg_gff_1_SFF_3_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S13reg_gff_1_SFF_4_U3 ( .A0_t (KeyArray_S13reg_gff_1_SFF_4_n2), .B0_t (KeyArray_S13reg_gff_1_SFF_4_n1), .Z0_t (keySBIn[4]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_4_U2 ( .A0_t (enKS), .B0_t (keySBIn[4]), .Z0_t (KeyArray_S13reg_gff_1_SFF_4_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_4_U1 ( .A0_t (KeyArray_S13reg_gff_1_SFF_4_QD), .B0_t (enKS), .Z0_t (KeyArray_S13reg_gff_1_SFF_4_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS20ser[4]), .B0_t (KeyArray_outS23ser[4]), .Z0_t (KeyArray_S13reg_gff_1_SFF_4_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S13reg_gff_1_SFF_4_MUXInst_X), .Z0_t (KeyArray_S13reg_gff_1_SFF_4_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S13reg_gff_1_SFF_4_MUXInst_Y), .B0_t (KeyArray_outS20ser[4]), .Z0_t (KeyArray_S13reg_gff_1_SFF_4_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S13reg_gff_1_SFF_5_U3 ( .A0_t (KeyArray_S13reg_gff_1_SFF_5_n2), .B0_t (KeyArray_S13reg_gff_1_SFF_5_n1), .Z0_t (keySBIn[5]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_5_U2 ( .A0_t (enKS), .B0_t (keySBIn[5]), .Z0_t (KeyArray_S13reg_gff_1_SFF_5_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_5_U1 ( .A0_t (KeyArray_S13reg_gff_1_SFF_5_QD), .B0_t (enKS), .Z0_t (KeyArray_S13reg_gff_1_SFF_5_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS20ser[5]), .B0_t (KeyArray_outS23ser[5]), .Z0_t (KeyArray_S13reg_gff_1_SFF_5_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S13reg_gff_1_SFF_5_MUXInst_X), .Z0_t (KeyArray_S13reg_gff_1_SFF_5_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S13reg_gff_1_SFF_5_MUXInst_Y), .B0_t (KeyArray_outS20ser[5]), .Z0_t (KeyArray_S13reg_gff_1_SFF_5_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S13reg_gff_1_SFF_6_U3 ( .A0_t (KeyArray_S13reg_gff_1_SFF_6_n2), .B0_t (KeyArray_S13reg_gff_1_SFF_6_n1), .Z0_t (keySBIn[6]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_6_U2 ( .A0_t (enKS), .B0_t (keySBIn[6]), .Z0_t (KeyArray_S13reg_gff_1_SFF_6_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_6_U1 ( .A0_t (KeyArray_S13reg_gff_1_SFF_6_QD), .B0_t (enKS), .Z0_t (KeyArray_S13reg_gff_1_SFF_6_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS20ser[6]), .B0_t (KeyArray_outS23ser[6]), .Z0_t (KeyArray_S13reg_gff_1_SFF_6_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S13reg_gff_1_SFF_6_MUXInst_X), .Z0_t (KeyArray_S13reg_gff_1_SFF_6_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S13reg_gff_1_SFF_6_MUXInst_Y), .B0_t (KeyArray_outS20ser[6]), .Z0_t (KeyArray_S13reg_gff_1_SFF_6_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S13reg_gff_1_SFF_7_U3 ( .A0_t (KeyArray_S13reg_gff_1_SFF_7_n2), .B0_t (KeyArray_S13reg_gff_1_SFF_7_n1), .Z0_t (keySBIn[7]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_7_U2 ( .A0_t (enKS), .B0_t (keySBIn[7]), .Z0_t (KeyArray_S13reg_gff_1_SFF_7_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_7_U1 ( .A0_t (KeyArray_S13reg_gff_1_SFF_7_QD), .B0_t (enKS), .Z0_t (KeyArray_S13reg_gff_1_SFF_7_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS20ser[7]), .B0_t (KeyArray_outS23ser[7]), .Z0_t (KeyArray_S13reg_gff_1_SFF_7_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S13reg_gff_1_SFF_7_MUXInst_X), .Z0_t (KeyArray_S13reg_gff_1_SFF_7_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S13reg_gff_1_SFF_7_MUXInst_Y), .B0_t (KeyArray_outS20ser[7]), .Z0_t (KeyArray_S13reg_gff_1_SFF_7_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S20reg_gff_1_SFF_0_U3 ( .A0_t (KeyArray_S20reg_gff_1_SFF_0_n2), .B0_t (KeyArray_S20reg_gff_1_SFF_0_n1), .Z0_t (KeyArray_outS20ser[0]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_0_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS20ser[0]), .Z0_t (KeyArray_S20reg_gff_1_SFF_0_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_0_U1 ( .A0_t (KeyArray_S20reg_gff_1_SFF_0_QD), .B0_t (enKS), .Z0_t (KeyArray_S20reg_gff_1_SFF_0_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS21ser[0]), .B0_t (KeyArray_outS30ser[0]), .Z0_t (KeyArray_S20reg_gff_1_SFF_0_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S20reg_gff_1_SFF_0_MUXInst_X), .Z0_t (KeyArray_S20reg_gff_1_SFF_0_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S20reg_gff_1_SFF_0_MUXInst_Y), .B0_t (KeyArray_outS21ser[0]), .Z0_t (KeyArray_S20reg_gff_1_SFF_0_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S20reg_gff_1_SFF_1_U3 ( .A0_t (KeyArray_S20reg_gff_1_SFF_1_n2), .B0_t (KeyArray_S20reg_gff_1_SFF_1_n1), .Z0_t (KeyArray_outS20ser[1]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_1_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS20ser[1]), .Z0_t (KeyArray_S20reg_gff_1_SFF_1_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_1_U1 ( .A0_t (KeyArray_S20reg_gff_1_SFF_1_QD), .B0_t (enKS), .Z0_t (KeyArray_S20reg_gff_1_SFF_1_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS21ser[1]), .B0_t (KeyArray_outS30ser[1]), .Z0_t (KeyArray_S20reg_gff_1_SFF_1_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S20reg_gff_1_SFF_1_MUXInst_X), .Z0_t (KeyArray_S20reg_gff_1_SFF_1_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S20reg_gff_1_SFF_1_MUXInst_Y), .B0_t (KeyArray_outS21ser[1]), .Z0_t (KeyArray_S20reg_gff_1_SFF_1_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S20reg_gff_1_SFF_2_U3 ( .A0_t (KeyArray_S20reg_gff_1_SFF_2_n2), .B0_t (KeyArray_S20reg_gff_1_SFF_2_n1), .Z0_t (KeyArray_outS20ser[2]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_2_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS20ser[2]), .Z0_t (KeyArray_S20reg_gff_1_SFF_2_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_2_U1 ( .A0_t (KeyArray_S20reg_gff_1_SFF_2_QD), .B0_t (enKS), .Z0_t (KeyArray_S20reg_gff_1_SFF_2_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS21ser[2]), .B0_t (KeyArray_outS30ser[2]), .Z0_t (KeyArray_S20reg_gff_1_SFF_2_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S20reg_gff_1_SFF_2_MUXInst_X), .Z0_t (KeyArray_S20reg_gff_1_SFF_2_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S20reg_gff_1_SFF_2_MUXInst_Y), .B0_t (KeyArray_outS21ser[2]), .Z0_t (KeyArray_S20reg_gff_1_SFF_2_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S20reg_gff_1_SFF_3_U3 ( .A0_t (KeyArray_S20reg_gff_1_SFF_3_n2), .B0_t (KeyArray_S20reg_gff_1_SFF_3_n1), .Z0_t (KeyArray_outS20ser[3]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_3_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS20ser[3]), .Z0_t (KeyArray_S20reg_gff_1_SFF_3_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_3_U1 ( .A0_t (KeyArray_S20reg_gff_1_SFF_3_QD), .B0_t (enKS), .Z0_t (KeyArray_S20reg_gff_1_SFF_3_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS21ser[3]), .B0_t (KeyArray_outS30ser[3]), .Z0_t (KeyArray_S20reg_gff_1_SFF_3_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S20reg_gff_1_SFF_3_MUXInst_X), .Z0_t (KeyArray_S20reg_gff_1_SFF_3_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S20reg_gff_1_SFF_3_MUXInst_Y), .B0_t (KeyArray_outS21ser[3]), .Z0_t (KeyArray_S20reg_gff_1_SFF_3_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S20reg_gff_1_SFF_4_U3 ( .A0_t (KeyArray_S20reg_gff_1_SFF_4_n2), .B0_t (KeyArray_S20reg_gff_1_SFF_4_n1), .Z0_t (KeyArray_outS20ser[4]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_4_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS20ser[4]), .Z0_t (KeyArray_S20reg_gff_1_SFF_4_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_4_U1 ( .A0_t (KeyArray_S20reg_gff_1_SFF_4_QD), .B0_t (enKS), .Z0_t (KeyArray_S20reg_gff_1_SFF_4_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS21ser[4]), .B0_t (KeyArray_outS30ser[4]), .Z0_t (KeyArray_S20reg_gff_1_SFF_4_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S20reg_gff_1_SFF_4_MUXInst_X), .Z0_t (KeyArray_S20reg_gff_1_SFF_4_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S20reg_gff_1_SFF_4_MUXInst_Y), .B0_t (KeyArray_outS21ser[4]), .Z0_t (KeyArray_S20reg_gff_1_SFF_4_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S20reg_gff_1_SFF_5_U3 ( .A0_t (KeyArray_S20reg_gff_1_SFF_5_n2), .B0_t (KeyArray_S20reg_gff_1_SFF_5_n1), .Z0_t (KeyArray_outS20ser[5]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_5_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS20ser[5]), .Z0_t (KeyArray_S20reg_gff_1_SFF_5_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_5_U1 ( .A0_t (KeyArray_S20reg_gff_1_SFF_5_QD), .B0_t (enKS), .Z0_t (KeyArray_S20reg_gff_1_SFF_5_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS21ser[5]), .B0_t (KeyArray_outS30ser[5]), .Z0_t (KeyArray_S20reg_gff_1_SFF_5_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S20reg_gff_1_SFF_5_MUXInst_X), .Z0_t (KeyArray_S20reg_gff_1_SFF_5_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S20reg_gff_1_SFF_5_MUXInst_Y), .B0_t (KeyArray_outS21ser[5]), .Z0_t (KeyArray_S20reg_gff_1_SFF_5_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S20reg_gff_1_SFF_6_U3 ( .A0_t (KeyArray_S20reg_gff_1_SFF_6_n2), .B0_t (KeyArray_S20reg_gff_1_SFF_6_n1), .Z0_t (KeyArray_outS20ser[6]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_6_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS20ser[6]), .Z0_t (KeyArray_S20reg_gff_1_SFF_6_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_6_U1 ( .A0_t (KeyArray_S20reg_gff_1_SFF_6_QD), .B0_t (enKS), .Z0_t (KeyArray_S20reg_gff_1_SFF_6_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS21ser[6]), .B0_t (KeyArray_outS30ser[6]), .Z0_t (KeyArray_S20reg_gff_1_SFF_6_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S20reg_gff_1_SFF_6_MUXInst_X), .Z0_t (KeyArray_S20reg_gff_1_SFF_6_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S20reg_gff_1_SFF_6_MUXInst_Y), .B0_t (KeyArray_outS21ser[6]), .Z0_t (KeyArray_S20reg_gff_1_SFF_6_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S20reg_gff_1_SFF_7_U3 ( .A0_t (KeyArray_S20reg_gff_1_SFF_7_n2), .B0_t (KeyArray_S20reg_gff_1_SFF_7_n1), .Z0_t (KeyArray_outS20ser[7]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_7_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS20ser[7]), .Z0_t (KeyArray_S20reg_gff_1_SFF_7_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_7_U1 ( .A0_t (KeyArray_S20reg_gff_1_SFF_7_QD), .B0_t (enKS), .Z0_t (KeyArray_S20reg_gff_1_SFF_7_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS21ser[7]), .B0_t (KeyArray_outS30ser[7]), .Z0_t (KeyArray_S20reg_gff_1_SFF_7_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S20reg_gff_1_SFF_7_MUXInst_X), .Z0_t (KeyArray_S20reg_gff_1_SFF_7_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S20reg_gff_1_SFF_7_MUXInst_Y), .B0_t (KeyArray_outS21ser[7]), .Z0_t (KeyArray_S20reg_gff_1_SFF_7_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S21reg_gff_1_SFF_0_U3 ( .A0_t (KeyArray_S21reg_gff_1_SFF_0_n2), .B0_t (KeyArray_S21reg_gff_1_SFF_0_n1), .Z0_t (KeyArray_outS21ser[0]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_0_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS21ser[0]), .Z0_t (KeyArray_S21reg_gff_1_SFF_0_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_0_U1 ( .A0_t (KeyArray_S21reg_gff_1_SFF_0_QD), .B0_t (enKS), .Z0_t (KeyArray_S21reg_gff_1_SFF_0_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS22ser[0]), .B0_t (KeyArray_outS31ser[0]), .Z0_t (KeyArray_S21reg_gff_1_SFF_0_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S21reg_gff_1_SFF_0_MUXInst_X), .Z0_t (KeyArray_S21reg_gff_1_SFF_0_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S21reg_gff_1_SFF_0_MUXInst_Y), .B0_t (KeyArray_outS22ser[0]), .Z0_t (KeyArray_S21reg_gff_1_SFF_0_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S21reg_gff_1_SFF_1_U3 ( .A0_t (KeyArray_S21reg_gff_1_SFF_1_n2), .B0_t (KeyArray_S21reg_gff_1_SFF_1_n1), .Z0_t (KeyArray_outS21ser[1]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_1_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS21ser[1]), .Z0_t (KeyArray_S21reg_gff_1_SFF_1_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_1_U1 ( .A0_t (KeyArray_S21reg_gff_1_SFF_1_QD), .B0_t (enKS), .Z0_t (KeyArray_S21reg_gff_1_SFF_1_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS22ser[1]), .B0_t (KeyArray_outS31ser[1]), .Z0_t (KeyArray_S21reg_gff_1_SFF_1_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S21reg_gff_1_SFF_1_MUXInst_X), .Z0_t (KeyArray_S21reg_gff_1_SFF_1_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S21reg_gff_1_SFF_1_MUXInst_Y), .B0_t (KeyArray_outS22ser[1]), .Z0_t (KeyArray_S21reg_gff_1_SFF_1_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S21reg_gff_1_SFF_2_U3 ( .A0_t (KeyArray_S21reg_gff_1_SFF_2_n2), .B0_t (KeyArray_S21reg_gff_1_SFF_2_n1), .Z0_t (KeyArray_outS21ser[2]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_2_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS21ser[2]), .Z0_t (KeyArray_S21reg_gff_1_SFF_2_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_2_U1 ( .A0_t (KeyArray_S21reg_gff_1_SFF_2_QD), .B0_t (enKS), .Z0_t (KeyArray_S21reg_gff_1_SFF_2_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS22ser[2]), .B0_t (KeyArray_outS31ser[2]), .Z0_t (KeyArray_S21reg_gff_1_SFF_2_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S21reg_gff_1_SFF_2_MUXInst_X), .Z0_t (KeyArray_S21reg_gff_1_SFF_2_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S21reg_gff_1_SFF_2_MUXInst_Y), .B0_t (KeyArray_outS22ser[2]), .Z0_t (KeyArray_S21reg_gff_1_SFF_2_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S21reg_gff_1_SFF_3_U3 ( .A0_t (KeyArray_S21reg_gff_1_SFF_3_n2), .B0_t (KeyArray_S21reg_gff_1_SFF_3_n1), .Z0_t (KeyArray_outS21ser[3]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_3_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS21ser[3]), .Z0_t (KeyArray_S21reg_gff_1_SFF_3_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_3_U1 ( .A0_t (KeyArray_S21reg_gff_1_SFF_3_QD), .B0_t (enKS), .Z0_t (KeyArray_S21reg_gff_1_SFF_3_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS22ser[3]), .B0_t (KeyArray_outS31ser[3]), .Z0_t (KeyArray_S21reg_gff_1_SFF_3_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S21reg_gff_1_SFF_3_MUXInst_X), .Z0_t (KeyArray_S21reg_gff_1_SFF_3_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S21reg_gff_1_SFF_3_MUXInst_Y), .B0_t (KeyArray_outS22ser[3]), .Z0_t (KeyArray_S21reg_gff_1_SFF_3_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S21reg_gff_1_SFF_4_U3 ( .A0_t (KeyArray_S21reg_gff_1_SFF_4_n2), .B0_t (KeyArray_S21reg_gff_1_SFF_4_n1), .Z0_t (KeyArray_outS21ser[4]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_4_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS21ser[4]), .Z0_t (KeyArray_S21reg_gff_1_SFF_4_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_4_U1 ( .A0_t (KeyArray_S21reg_gff_1_SFF_4_QD), .B0_t (enKS), .Z0_t (KeyArray_S21reg_gff_1_SFF_4_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS22ser[4]), .B0_t (KeyArray_outS31ser[4]), .Z0_t (KeyArray_S21reg_gff_1_SFF_4_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S21reg_gff_1_SFF_4_MUXInst_X), .Z0_t (KeyArray_S21reg_gff_1_SFF_4_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S21reg_gff_1_SFF_4_MUXInst_Y), .B0_t (KeyArray_outS22ser[4]), .Z0_t (KeyArray_S21reg_gff_1_SFF_4_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S21reg_gff_1_SFF_5_U3 ( .A0_t (KeyArray_S21reg_gff_1_SFF_5_n2), .B0_t (KeyArray_S21reg_gff_1_SFF_5_n1), .Z0_t (KeyArray_outS21ser[5]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_5_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS21ser[5]), .Z0_t (KeyArray_S21reg_gff_1_SFF_5_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_5_U1 ( .A0_t (KeyArray_S21reg_gff_1_SFF_5_QD), .B0_t (enKS), .Z0_t (KeyArray_S21reg_gff_1_SFF_5_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS22ser[5]), .B0_t (KeyArray_outS31ser[5]), .Z0_t (KeyArray_S21reg_gff_1_SFF_5_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S21reg_gff_1_SFF_5_MUXInst_X), .Z0_t (KeyArray_S21reg_gff_1_SFF_5_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S21reg_gff_1_SFF_5_MUXInst_Y), .B0_t (KeyArray_outS22ser[5]), .Z0_t (KeyArray_S21reg_gff_1_SFF_5_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S21reg_gff_1_SFF_6_U3 ( .A0_t (KeyArray_S21reg_gff_1_SFF_6_n2), .B0_t (KeyArray_S21reg_gff_1_SFF_6_n1), .Z0_t (KeyArray_outS21ser[6]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_6_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS21ser[6]), .Z0_t (KeyArray_S21reg_gff_1_SFF_6_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_6_U1 ( .A0_t (KeyArray_S21reg_gff_1_SFF_6_QD), .B0_t (enKS), .Z0_t (KeyArray_S21reg_gff_1_SFF_6_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS22ser[6]), .B0_t (KeyArray_outS31ser[6]), .Z0_t (KeyArray_S21reg_gff_1_SFF_6_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S21reg_gff_1_SFF_6_MUXInst_X), .Z0_t (KeyArray_S21reg_gff_1_SFF_6_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S21reg_gff_1_SFF_6_MUXInst_Y), .B0_t (KeyArray_outS22ser[6]), .Z0_t (KeyArray_S21reg_gff_1_SFF_6_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S21reg_gff_1_SFF_7_U3 ( .A0_t (KeyArray_S21reg_gff_1_SFF_7_n2), .B0_t (KeyArray_S21reg_gff_1_SFF_7_n1), .Z0_t (KeyArray_outS21ser[7]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_7_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS21ser[7]), .Z0_t (KeyArray_S21reg_gff_1_SFF_7_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_7_U1 ( .A0_t (KeyArray_S21reg_gff_1_SFF_7_QD), .B0_t (enKS), .Z0_t (KeyArray_S21reg_gff_1_SFF_7_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS22ser[7]), .B0_t (KeyArray_outS31ser[7]), .Z0_t (KeyArray_S21reg_gff_1_SFF_7_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S21reg_gff_1_SFF_7_MUXInst_X), .Z0_t (KeyArray_S21reg_gff_1_SFF_7_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S21reg_gff_1_SFF_7_MUXInst_Y), .B0_t (KeyArray_outS22ser[7]), .Z0_t (KeyArray_S21reg_gff_1_SFF_7_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S22reg_gff_1_SFF_0_U3 ( .A0_t (KeyArray_S22reg_gff_1_SFF_0_n2), .B0_t (KeyArray_S22reg_gff_1_SFF_0_n1), .Z0_t (KeyArray_outS22ser[0]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_0_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS22ser[0]), .Z0_t (KeyArray_S22reg_gff_1_SFF_0_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_0_U1 ( .A0_t (KeyArray_S22reg_gff_1_SFF_0_QD), .B0_t (enKS), .Z0_t (KeyArray_S22reg_gff_1_SFF_0_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS23ser[0]), .B0_t (KeyArray_outS32ser[0]), .Z0_t (KeyArray_S22reg_gff_1_SFF_0_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S22reg_gff_1_SFF_0_MUXInst_X), .Z0_t (KeyArray_S22reg_gff_1_SFF_0_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S22reg_gff_1_SFF_0_MUXInst_Y), .B0_t (KeyArray_outS23ser[0]), .Z0_t (KeyArray_S22reg_gff_1_SFF_0_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S22reg_gff_1_SFF_1_U3 ( .A0_t (KeyArray_S22reg_gff_1_SFF_1_n2), .B0_t (KeyArray_S22reg_gff_1_SFF_1_n1), .Z0_t (KeyArray_outS22ser[1]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_1_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS22ser[1]), .Z0_t (KeyArray_S22reg_gff_1_SFF_1_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_1_U1 ( .A0_t (KeyArray_S22reg_gff_1_SFF_1_QD), .B0_t (enKS), .Z0_t (KeyArray_S22reg_gff_1_SFF_1_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS23ser[1]), .B0_t (KeyArray_outS32ser[1]), .Z0_t (KeyArray_S22reg_gff_1_SFF_1_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S22reg_gff_1_SFF_1_MUXInst_X), .Z0_t (KeyArray_S22reg_gff_1_SFF_1_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S22reg_gff_1_SFF_1_MUXInst_Y), .B0_t (KeyArray_outS23ser[1]), .Z0_t (KeyArray_S22reg_gff_1_SFF_1_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S22reg_gff_1_SFF_2_U3 ( .A0_t (KeyArray_S22reg_gff_1_SFF_2_n2), .B0_t (KeyArray_S22reg_gff_1_SFF_2_n1), .Z0_t (KeyArray_outS22ser[2]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_2_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS22ser[2]), .Z0_t (KeyArray_S22reg_gff_1_SFF_2_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_2_U1 ( .A0_t (KeyArray_S22reg_gff_1_SFF_2_QD), .B0_t (enKS), .Z0_t (KeyArray_S22reg_gff_1_SFF_2_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS23ser[2]), .B0_t (KeyArray_outS32ser[2]), .Z0_t (KeyArray_S22reg_gff_1_SFF_2_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S22reg_gff_1_SFF_2_MUXInst_X), .Z0_t (KeyArray_S22reg_gff_1_SFF_2_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S22reg_gff_1_SFF_2_MUXInst_Y), .B0_t (KeyArray_outS23ser[2]), .Z0_t (KeyArray_S22reg_gff_1_SFF_2_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S22reg_gff_1_SFF_3_U3 ( .A0_t (KeyArray_S22reg_gff_1_SFF_3_n2), .B0_t (KeyArray_S22reg_gff_1_SFF_3_n1), .Z0_t (KeyArray_outS22ser[3]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_3_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS22ser[3]), .Z0_t (KeyArray_S22reg_gff_1_SFF_3_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_3_U1 ( .A0_t (KeyArray_S22reg_gff_1_SFF_3_QD), .B0_t (enKS), .Z0_t (KeyArray_S22reg_gff_1_SFF_3_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS23ser[3]), .B0_t (KeyArray_outS32ser[3]), .Z0_t (KeyArray_S22reg_gff_1_SFF_3_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S22reg_gff_1_SFF_3_MUXInst_X), .Z0_t (KeyArray_S22reg_gff_1_SFF_3_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S22reg_gff_1_SFF_3_MUXInst_Y), .B0_t (KeyArray_outS23ser[3]), .Z0_t (KeyArray_S22reg_gff_1_SFF_3_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S22reg_gff_1_SFF_4_U3 ( .A0_t (KeyArray_S22reg_gff_1_SFF_4_n2), .B0_t (KeyArray_S22reg_gff_1_SFF_4_n1), .Z0_t (KeyArray_outS22ser[4]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_4_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS22ser[4]), .Z0_t (KeyArray_S22reg_gff_1_SFF_4_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_4_U1 ( .A0_t (KeyArray_S22reg_gff_1_SFF_4_QD), .B0_t (enKS), .Z0_t (KeyArray_S22reg_gff_1_SFF_4_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS23ser[4]), .B0_t (KeyArray_outS32ser[4]), .Z0_t (KeyArray_S22reg_gff_1_SFF_4_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S22reg_gff_1_SFF_4_MUXInst_X), .Z0_t (KeyArray_S22reg_gff_1_SFF_4_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S22reg_gff_1_SFF_4_MUXInst_Y), .B0_t (KeyArray_outS23ser[4]), .Z0_t (KeyArray_S22reg_gff_1_SFF_4_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S22reg_gff_1_SFF_5_U3 ( .A0_t (KeyArray_S22reg_gff_1_SFF_5_n2), .B0_t (KeyArray_S22reg_gff_1_SFF_5_n1), .Z0_t (KeyArray_outS22ser[5]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_5_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS22ser[5]), .Z0_t (KeyArray_S22reg_gff_1_SFF_5_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_5_U1 ( .A0_t (KeyArray_S22reg_gff_1_SFF_5_QD), .B0_t (enKS), .Z0_t (KeyArray_S22reg_gff_1_SFF_5_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS23ser[5]), .B0_t (KeyArray_outS32ser[5]), .Z0_t (KeyArray_S22reg_gff_1_SFF_5_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S22reg_gff_1_SFF_5_MUXInst_X), .Z0_t (KeyArray_S22reg_gff_1_SFF_5_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S22reg_gff_1_SFF_5_MUXInst_Y), .B0_t (KeyArray_outS23ser[5]), .Z0_t (KeyArray_S22reg_gff_1_SFF_5_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S22reg_gff_1_SFF_6_U3 ( .A0_t (KeyArray_S22reg_gff_1_SFF_6_n2), .B0_t (KeyArray_S22reg_gff_1_SFF_6_n1), .Z0_t (KeyArray_outS22ser[6]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_6_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS22ser[6]), .Z0_t (KeyArray_S22reg_gff_1_SFF_6_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_6_U1 ( .A0_t (KeyArray_S22reg_gff_1_SFF_6_QD), .B0_t (enKS), .Z0_t (KeyArray_S22reg_gff_1_SFF_6_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS23ser[6]), .B0_t (KeyArray_outS32ser[6]), .Z0_t (KeyArray_S22reg_gff_1_SFF_6_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S22reg_gff_1_SFF_6_MUXInst_X), .Z0_t (KeyArray_S22reg_gff_1_SFF_6_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S22reg_gff_1_SFF_6_MUXInst_Y), .B0_t (KeyArray_outS23ser[6]), .Z0_t (KeyArray_S22reg_gff_1_SFF_6_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S22reg_gff_1_SFF_7_U3 ( .A0_t (KeyArray_S22reg_gff_1_SFF_7_n2), .B0_t (KeyArray_S22reg_gff_1_SFF_7_n1), .Z0_t (KeyArray_outS22ser[7]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_7_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS22ser[7]), .Z0_t (KeyArray_S22reg_gff_1_SFF_7_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_7_U1 ( .A0_t (KeyArray_S22reg_gff_1_SFF_7_QD), .B0_t (enKS), .Z0_t (KeyArray_S22reg_gff_1_SFF_7_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS23ser[7]), .B0_t (KeyArray_outS32ser[7]), .Z0_t (KeyArray_S22reg_gff_1_SFF_7_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S22reg_gff_1_SFF_7_MUXInst_X), .Z0_t (KeyArray_S22reg_gff_1_SFF_7_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S22reg_gff_1_SFF_7_MUXInst_Y), .B0_t (KeyArray_outS23ser[7]), .Z0_t (KeyArray_S22reg_gff_1_SFF_7_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S23reg_gff_1_SFF_0_U3 ( .A0_t (KeyArray_S23reg_gff_1_SFF_0_n2), .B0_t (KeyArray_S23reg_gff_1_SFF_0_n1), .Z0_t (KeyArray_outS23ser[0]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_0_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS23ser[0]), .Z0_t (KeyArray_S23reg_gff_1_SFF_0_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_0_U1 ( .A0_t (KeyArray_S23reg_gff_1_SFF_0_QD), .B0_t (enKS), .Z0_t (KeyArray_S23reg_gff_1_SFF_0_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS30ser[0]), .B0_t (KeyArray_outS33ser[0]), .Z0_t (KeyArray_S23reg_gff_1_SFF_0_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S23reg_gff_1_SFF_0_MUXInst_X), .Z0_t (KeyArray_S23reg_gff_1_SFF_0_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S23reg_gff_1_SFF_0_MUXInst_Y), .B0_t (KeyArray_outS30ser[0]), .Z0_t (KeyArray_S23reg_gff_1_SFF_0_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S23reg_gff_1_SFF_1_U3 ( .A0_t (KeyArray_S23reg_gff_1_SFF_1_n2), .B0_t (KeyArray_S23reg_gff_1_SFF_1_n1), .Z0_t (KeyArray_outS23ser[1]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_1_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS23ser[1]), .Z0_t (KeyArray_S23reg_gff_1_SFF_1_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_1_U1 ( .A0_t (KeyArray_S23reg_gff_1_SFF_1_QD), .B0_t (enKS), .Z0_t (KeyArray_S23reg_gff_1_SFF_1_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS30ser[1]), .B0_t (KeyArray_outS33ser[1]), .Z0_t (KeyArray_S23reg_gff_1_SFF_1_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S23reg_gff_1_SFF_1_MUXInst_X), .Z0_t (KeyArray_S23reg_gff_1_SFF_1_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S23reg_gff_1_SFF_1_MUXInst_Y), .B0_t (KeyArray_outS30ser[1]), .Z0_t (KeyArray_S23reg_gff_1_SFF_1_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S23reg_gff_1_SFF_2_U3 ( .A0_t (KeyArray_S23reg_gff_1_SFF_2_n2), .B0_t (KeyArray_S23reg_gff_1_SFF_2_n1), .Z0_t (KeyArray_outS23ser[2]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_2_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS23ser[2]), .Z0_t (KeyArray_S23reg_gff_1_SFF_2_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_2_U1 ( .A0_t (KeyArray_S23reg_gff_1_SFF_2_QD), .B0_t (enKS), .Z0_t (KeyArray_S23reg_gff_1_SFF_2_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS30ser[2]), .B0_t (KeyArray_outS33ser[2]), .Z0_t (KeyArray_S23reg_gff_1_SFF_2_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S23reg_gff_1_SFF_2_MUXInst_X), .Z0_t (KeyArray_S23reg_gff_1_SFF_2_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S23reg_gff_1_SFF_2_MUXInst_Y), .B0_t (KeyArray_outS30ser[2]), .Z0_t (KeyArray_S23reg_gff_1_SFF_2_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S23reg_gff_1_SFF_3_U3 ( .A0_t (KeyArray_S23reg_gff_1_SFF_3_n2), .B0_t (KeyArray_S23reg_gff_1_SFF_3_n1), .Z0_t (KeyArray_outS23ser[3]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_3_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS23ser[3]), .Z0_t (KeyArray_S23reg_gff_1_SFF_3_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_3_U1 ( .A0_t (KeyArray_S23reg_gff_1_SFF_3_QD), .B0_t (enKS), .Z0_t (KeyArray_S23reg_gff_1_SFF_3_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS30ser[3]), .B0_t (KeyArray_outS33ser[3]), .Z0_t (KeyArray_S23reg_gff_1_SFF_3_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S23reg_gff_1_SFF_3_MUXInst_X), .Z0_t (KeyArray_S23reg_gff_1_SFF_3_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S23reg_gff_1_SFF_3_MUXInst_Y), .B0_t (KeyArray_outS30ser[3]), .Z0_t (KeyArray_S23reg_gff_1_SFF_3_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S23reg_gff_1_SFF_4_U3 ( .A0_t (KeyArray_S23reg_gff_1_SFF_4_n2), .B0_t (KeyArray_S23reg_gff_1_SFF_4_n1), .Z0_t (KeyArray_outS23ser[4]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_4_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS23ser[4]), .Z0_t (KeyArray_S23reg_gff_1_SFF_4_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_4_U1 ( .A0_t (KeyArray_S23reg_gff_1_SFF_4_QD), .B0_t (enKS), .Z0_t (KeyArray_S23reg_gff_1_SFF_4_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS30ser[4]), .B0_t (KeyArray_outS33ser[4]), .Z0_t (KeyArray_S23reg_gff_1_SFF_4_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S23reg_gff_1_SFF_4_MUXInst_X), .Z0_t (KeyArray_S23reg_gff_1_SFF_4_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S23reg_gff_1_SFF_4_MUXInst_Y), .B0_t (KeyArray_outS30ser[4]), .Z0_t (KeyArray_S23reg_gff_1_SFF_4_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S23reg_gff_1_SFF_5_U3 ( .A0_t (KeyArray_S23reg_gff_1_SFF_5_n2), .B0_t (KeyArray_S23reg_gff_1_SFF_5_n1), .Z0_t (KeyArray_outS23ser[5]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_5_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS23ser[5]), .Z0_t (KeyArray_S23reg_gff_1_SFF_5_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_5_U1 ( .A0_t (KeyArray_S23reg_gff_1_SFF_5_QD), .B0_t (enKS), .Z0_t (KeyArray_S23reg_gff_1_SFF_5_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS30ser[5]), .B0_t (KeyArray_outS33ser[5]), .Z0_t (KeyArray_S23reg_gff_1_SFF_5_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S23reg_gff_1_SFF_5_MUXInst_X), .Z0_t (KeyArray_S23reg_gff_1_SFF_5_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S23reg_gff_1_SFF_5_MUXInst_Y), .B0_t (KeyArray_outS30ser[5]), .Z0_t (KeyArray_S23reg_gff_1_SFF_5_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S23reg_gff_1_SFF_6_U3 ( .A0_t (KeyArray_S23reg_gff_1_SFF_6_n2), .B0_t (KeyArray_S23reg_gff_1_SFF_6_n1), .Z0_t (KeyArray_outS23ser[6]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_6_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS23ser[6]), .Z0_t (KeyArray_S23reg_gff_1_SFF_6_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_6_U1 ( .A0_t (KeyArray_S23reg_gff_1_SFF_6_QD), .B0_t (enKS), .Z0_t (KeyArray_S23reg_gff_1_SFF_6_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS30ser[6]), .B0_t (KeyArray_outS33ser[6]), .Z0_t (KeyArray_S23reg_gff_1_SFF_6_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S23reg_gff_1_SFF_6_MUXInst_X), .Z0_t (KeyArray_S23reg_gff_1_SFF_6_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S23reg_gff_1_SFF_6_MUXInst_Y), .B0_t (KeyArray_outS30ser[6]), .Z0_t (KeyArray_S23reg_gff_1_SFF_6_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S23reg_gff_1_SFF_7_U3 ( .A0_t (KeyArray_S23reg_gff_1_SFF_7_n2), .B0_t (KeyArray_S23reg_gff_1_SFF_7_n1), .Z0_t (KeyArray_outS23ser[7]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_7_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS23ser[7]), .Z0_t (KeyArray_S23reg_gff_1_SFF_7_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_7_U1 ( .A0_t (KeyArray_S23reg_gff_1_SFF_7_QD), .B0_t (enKS), .Z0_t (KeyArray_S23reg_gff_1_SFF_7_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS30ser[7]), .B0_t (KeyArray_outS33ser[7]), .Z0_t (KeyArray_S23reg_gff_1_SFF_7_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S23reg_gff_1_SFF_7_MUXInst_X), .Z0_t (KeyArray_S23reg_gff_1_SFF_7_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S23reg_gff_1_SFF_7_MUXInst_Y), .B0_t (KeyArray_outS30ser[7]), .Z0_t (KeyArray_S23reg_gff_1_SFF_7_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S30reg_gff_1_SFF_0_U3 ( .A0_t (KeyArray_S30reg_gff_1_SFF_0_n2), .B0_t (KeyArray_S30reg_gff_1_SFF_0_n1), .Z0_t (KeyArray_outS30ser[0]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_0_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS30ser[0]), .Z0_t (KeyArray_S30reg_gff_1_SFF_0_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_0_U1 ( .A0_t (KeyArray_S30reg_gff_1_SFF_0_QD), .B0_t (enKS), .Z0_t (KeyArray_S30reg_gff_1_SFF_0_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS31ser[0]), .B0_t (KeyArray_inS30par[0]), .Z0_t (KeyArray_S30reg_gff_1_SFF_0_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S30reg_gff_1_SFF_0_MUXInst_X), .Z0_t (KeyArray_S30reg_gff_1_SFF_0_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S30reg_gff_1_SFF_0_MUXInst_Y), .B0_t (KeyArray_outS31ser[0]), .Z0_t (KeyArray_S30reg_gff_1_SFF_0_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S30reg_gff_1_SFF_1_U3 ( .A0_t (KeyArray_S30reg_gff_1_SFF_1_n2), .B0_t (KeyArray_S30reg_gff_1_SFF_1_n1), .Z0_t (KeyArray_outS30ser[1]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_1_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS30ser[1]), .Z0_t (KeyArray_S30reg_gff_1_SFF_1_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_1_U1 ( .A0_t (KeyArray_S30reg_gff_1_SFF_1_QD), .B0_t (enKS), .Z0_t (KeyArray_S30reg_gff_1_SFF_1_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS31ser[1]), .B0_t (KeyArray_inS30par[1]), .Z0_t (KeyArray_S30reg_gff_1_SFF_1_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S30reg_gff_1_SFF_1_MUXInst_X), .Z0_t (KeyArray_S30reg_gff_1_SFF_1_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S30reg_gff_1_SFF_1_MUXInst_Y), .B0_t (KeyArray_outS31ser[1]), .Z0_t (KeyArray_S30reg_gff_1_SFF_1_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S30reg_gff_1_SFF_2_U3 ( .A0_t (KeyArray_S30reg_gff_1_SFF_2_n2), .B0_t (KeyArray_S30reg_gff_1_SFF_2_n1), .Z0_t (KeyArray_outS30ser[2]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_2_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS30ser[2]), .Z0_t (KeyArray_S30reg_gff_1_SFF_2_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_2_U1 ( .A0_t (KeyArray_S30reg_gff_1_SFF_2_QD), .B0_t (enKS), .Z0_t (KeyArray_S30reg_gff_1_SFF_2_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS31ser[2]), .B0_t (KeyArray_inS30par[2]), .Z0_t (KeyArray_S30reg_gff_1_SFF_2_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S30reg_gff_1_SFF_2_MUXInst_X), .Z0_t (KeyArray_S30reg_gff_1_SFF_2_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S30reg_gff_1_SFF_2_MUXInst_Y), .B0_t (KeyArray_outS31ser[2]), .Z0_t (KeyArray_S30reg_gff_1_SFF_2_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S30reg_gff_1_SFF_3_U3 ( .A0_t (KeyArray_S30reg_gff_1_SFF_3_n2), .B0_t (KeyArray_S30reg_gff_1_SFF_3_n1), .Z0_t (KeyArray_outS30ser[3]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_3_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS30ser[3]), .Z0_t (KeyArray_S30reg_gff_1_SFF_3_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_3_U1 ( .A0_t (KeyArray_S30reg_gff_1_SFF_3_QD), .B0_t (enKS), .Z0_t (KeyArray_S30reg_gff_1_SFF_3_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS31ser[3]), .B0_t (KeyArray_inS30par[3]), .Z0_t (KeyArray_S30reg_gff_1_SFF_3_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S30reg_gff_1_SFF_3_MUXInst_X), .Z0_t (KeyArray_S30reg_gff_1_SFF_3_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S30reg_gff_1_SFF_3_MUXInst_Y), .B0_t (KeyArray_outS31ser[3]), .Z0_t (KeyArray_S30reg_gff_1_SFF_3_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S30reg_gff_1_SFF_4_U3 ( .A0_t (KeyArray_S30reg_gff_1_SFF_4_n2), .B0_t (KeyArray_S30reg_gff_1_SFF_4_n1), .Z0_t (KeyArray_outS30ser[4]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_4_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS30ser[4]), .Z0_t (KeyArray_S30reg_gff_1_SFF_4_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_4_U1 ( .A0_t (KeyArray_S30reg_gff_1_SFF_4_QD), .B0_t (enKS), .Z0_t (KeyArray_S30reg_gff_1_SFF_4_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS31ser[4]), .B0_t (KeyArray_inS30par[4]), .Z0_t (KeyArray_S30reg_gff_1_SFF_4_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S30reg_gff_1_SFF_4_MUXInst_X), .Z0_t (KeyArray_S30reg_gff_1_SFF_4_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S30reg_gff_1_SFF_4_MUXInst_Y), .B0_t (KeyArray_outS31ser[4]), .Z0_t (KeyArray_S30reg_gff_1_SFF_4_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S30reg_gff_1_SFF_5_U3 ( .A0_t (KeyArray_S30reg_gff_1_SFF_5_n2), .B0_t (KeyArray_S30reg_gff_1_SFF_5_n1), .Z0_t (KeyArray_outS30ser[5]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_5_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS30ser[5]), .Z0_t (KeyArray_S30reg_gff_1_SFF_5_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_5_U1 ( .A0_t (KeyArray_S30reg_gff_1_SFF_5_QD), .B0_t (enKS), .Z0_t (KeyArray_S30reg_gff_1_SFF_5_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS31ser[5]), .B0_t (KeyArray_inS30par[5]), .Z0_t (KeyArray_S30reg_gff_1_SFF_5_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S30reg_gff_1_SFF_5_MUXInst_X), .Z0_t (KeyArray_S30reg_gff_1_SFF_5_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S30reg_gff_1_SFF_5_MUXInst_Y), .B0_t (KeyArray_outS31ser[5]), .Z0_t (KeyArray_S30reg_gff_1_SFF_5_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S30reg_gff_1_SFF_6_U3 ( .A0_t (KeyArray_S30reg_gff_1_SFF_6_n2), .B0_t (KeyArray_S30reg_gff_1_SFF_6_n1), .Z0_t (KeyArray_outS30ser[6]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_6_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS30ser[6]), .Z0_t (KeyArray_S30reg_gff_1_SFF_6_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_6_U1 ( .A0_t (KeyArray_S30reg_gff_1_SFF_6_QD), .B0_t (enKS), .Z0_t (KeyArray_S30reg_gff_1_SFF_6_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS31ser[6]), .B0_t (KeyArray_inS30par[6]), .Z0_t (KeyArray_S30reg_gff_1_SFF_6_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S30reg_gff_1_SFF_6_MUXInst_X), .Z0_t (KeyArray_S30reg_gff_1_SFF_6_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S30reg_gff_1_SFF_6_MUXInst_Y), .B0_t (KeyArray_outS31ser[6]), .Z0_t (KeyArray_S30reg_gff_1_SFF_6_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S30reg_gff_1_SFF_7_U3 ( .A0_t (KeyArray_S30reg_gff_1_SFF_7_n2), .B0_t (KeyArray_S30reg_gff_1_SFF_7_n1), .Z0_t (KeyArray_outS30ser[7]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_7_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS30ser[7]), .Z0_t (KeyArray_S30reg_gff_1_SFF_7_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_7_U1 ( .A0_t (KeyArray_S30reg_gff_1_SFF_7_QD), .B0_t (enKS), .Z0_t (KeyArray_S30reg_gff_1_SFF_7_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS31ser[7]), .B0_t (KeyArray_inS30par[7]), .Z0_t (KeyArray_S30reg_gff_1_SFF_7_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S30reg_gff_1_SFF_7_MUXInst_X), .Z0_t (KeyArray_S30reg_gff_1_SFF_7_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S30reg_gff_1_SFF_7_MUXInst_Y), .B0_t (KeyArray_outS31ser[7]), .Z0_t (KeyArray_S30reg_gff_1_SFF_7_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S31reg_gff_1_SFF_0_U3 ( .A0_t (KeyArray_S31reg_gff_1_SFF_0_n2), .B0_t (KeyArray_S31reg_gff_1_SFF_0_n1), .Z0_t (KeyArray_outS31ser[0]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_0_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS31ser[0]), .Z0_t (KeyArray_S31reg_gff_1_SFF_0_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_0_U1 ( .A0_t (KeyArray_S31reg_gff_1_SFF_0_QD), .B0_t (enKS), .Z0_t (KeyArray_S31reg_gff_1_SFF_0_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS32ser[0]), .B0_t (KeyArray_outS01ser_0_), .Z0_t (KeyArray_S31reg_gff_1_SFF_0_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S31reg_gff_1_SFF_0_MUXInst_X), .Z0_t (KeyArray_S31reg_gff_1_SFF_0_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S31reg_gff_1_SFF_0_MUXInst_Y), .B0_t (KeyArray_outS32ser[0]), .Z0_t (KeyArray_S31reg_gff_1_SFF_0_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S31reg_gff_1_SFF_1_U3 ( .A0_t (KeyArray_S31reg_gff_1_SFF_1_n2), .B0_t (KeyArray_S31reg_gff_1_SFF_1_n1), .Z0_t (KeyArray_outS31ser[1]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_1_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS31ser[1]), .Z0_t (KeyArray_S31reg_gff_1_SFF_1_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_1_U1 ( .A0_t (KeyArray_S31reg_gff_1_SFF_1_QD), .B0_t (enKS), .Z0_t (KeyArray_S31reg_gff_1_SFF_1_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS32ser[1]), .B0_t (KeyArray_outS01ser_1_), .Z0_t (KeyArray_S31reg_gff_1_SFF_1_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S31reg_gff_1_SFF_1_MUXInst_X), .Z0_t (KeyArray_S31reg_gff_1_SFF_1_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S31reg_gff_1_SFF_1_MUXInst_Y), .B0_t (KeyArray_outS32ser[1]), .Z0_t (KeyArray_S31reg_gff_1_SFF_1_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S31reg_gff_1_SFF_2_U3 ( .A0_t (KeyArray_S31reg_gff_1_SFF_2_n2), .B0_t (KeyArray_S31reg_gff_1_SFF_2_n1), .Z0_t (KeyArray_outS31ser[2]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_2_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS31ser[2]), .Z0_t (KeyArray_S31reg_gff_1_SFF_2_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_2_U1 ( .A0_t (KeyArray_S31reg_gff_1_SFF_2_QD), .B0_t (enKS), .Z0_t (KeyArray_S31reg_gff_1_SFF_2_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS32ser[2]), .B0_t (KeyArray_outS01ser_2_), .Z0_t (KeyArray_S31reg_gff_1_SFF_2_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S31reg_gff_1_SFF_2_MUXInst_X), .Z0_t (KeyArray_S31reg_gff_1_SFF_2_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S31reg_gff_1_SFF_2_MUXInst_Y), .B0_t (KeyArray_outS32ser[2]), .Z0_t (KeyArray_S31reg_gff_1_SFF_2_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S31reg_gff_1_SFF_3_U3 ( .A0_t (KeyArray_S31reg_gff_1_SFF_3_n2), .B0_t (KeyArray_S31reg_gff_1_SFF_3_n1), .Z0_t (KeyArray_outS31ser[3]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_3_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS31ser[3]), .Z0_t (KeyArray_S31reg_gff_1_SFF_3_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_3_U1 ( .A0_t (KeyArray_S31reg_gff_1_SFF_3_QD), .B0_t (enKS), .Z0_t (KeyArray_S31reg_gff_1_SFF_3_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS32ser[3]), .B0_t (KeyArray_outS01ser_3_), .Z0_t (KeyArray_S31reg_gff_1_SFF_3_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S31reg_gff_1_SFF_3_MUXInst_X), .Z0_t (KeyArray_S31reg_gff_1_SFF_3_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S31reg_gff_1_SFF_3_MUXInst_Y), .B0_t (KeyArray_outS32ser[3]), .Z0_t (KeyArray_S31reg_gff_1_SFF_3_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S31reg_gff_1_SFF_4_U3 ( .A0_t (KeyArray_S31reg_gff_1_SFF_4_n2), .B0_t (KeyArray_S31reg_gff_1_SFF_4_n1), .Z0_t (KeyArray_outS31ser[4]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_4_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS31ser[4]), .Z0_t (KeyArray_S31reg_gff_1_SFF_4_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_4_U1 ( .A0_t (KeyArray_S31reg_gff_1_SFF_4_QD), .B0_t (enKS), .Z0_t (KeyArray_S31reg_gff_1_SFF_4_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS32ser[4]), .B0_t (KeyArray_outS01ser_4_), .Z0_t (KeyArray_S31reg_gff_1_SFF_4_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S31reg_gff_1_SFF_4_MUXInst_X), .Z0_t (KeyArray_S31reg_gff_1_SFF_4_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S31reg_gff_1_SFF_4_MUXInst_Y), .B0_t (KeyArray_outS32ser[4]), .Z0_t (KeyArray_S31reg_gff_1_SFF_4_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S31reg_gff_1_SFF_5_U3 ( .A0_t (KeyArray_S31reg_gff_1_SFF_5_n2), .B0_t (KeyArray_S31reg_gff_1_SFF_5_n1), .Z0_t (KeyArray_outS31ser[5]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_5_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS31ser[5]), .Z0_t (KeyArray_S31reg_gff_1_SFF_5_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_5_U1 ( .A0_t (KeyArray_S31reg_gff_1_SFF_5_QD), .B0_t (enKS), .Z0_t (KeyArray_S31reg_gff_1_SFF_5_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS32ser[5]), .B0_t (KeyArray_outS01ser_5_), .Z0_t (KeyArray_S31reg_gff_1_SFF_5_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S31reg_gff_1_SFF_5_MUXInst_X), .Z0_t (KeyArray_S31reg_gff_1_SFF_5_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S31reg_gff_1_SFF_5_MUXInst_Y), .B0_t (KeyArray_outS32ser[5]), .Z0_t (KeyArray_S31reg_gff_1_SFF_5_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S31reg_gff_1_SFF_6_U3 ( .A0_t (KeyArray_S31reg_gff_1_SFF_6_n2), .B0_t (KeyArray_S31reg_gff_1_SFF_6_n1), .Z0_t (KeyArray_outS31ser[6]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_6_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS31ser[6]), .Z0_t (KeyArray_S31reg_gff_1_SFF_6_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_6_U1 ( .A0_t (KeyArray_S31reg_gff_1_SFF_6_QD), .B0_t (enKS), .Z0_t (KeyArray_S31reg_gff_1_SFF_6_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS32ser[6]), .B0_t (KeyArray_outS01ser_6_), .Z0_t (KeyArray_S31reg_gff_1_SFF_6_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S31reg_gff_1_SFF_6_MUXInst_X), .Z0_t (KeyArray_S31reg_gff_1_SFF_6_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S31reg_gff_1_SFF_6_MUXInst_Y), .B0_t (KeyArray_outS32ser[6]), .Z0_t (KeyArray_S31reg_gff_1_SFF_6_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S31reg_gff_1_SFF_7_U3 ( .A0_t (KeyArray_S31reg_gff_1_SFF_7_n2), .B0_t (KeyArray_S31reg_gff_1_SFF_7_n1), .Z0_t (KeyArray_outS31ser[7]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_7_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS31ser[7]), .Z0_t (KeyArray_S31reg_gff_1_SFF_7_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_7_U1 ( .A0_t (KeyArray_S31reg_gff_1_SFF_7_QD), .B0_t (enKS), .Z0_t (KeyArray_S31reg_gff_1_SFF_7_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS32ser[7]), .B0_t (KeyArray_outS01ser_7_), .Z0_t (KeyArray_S31reg_gff_1_SFF_7_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S31reg_gff_1_SFF_7_MUXInst_X), .Z0_t (KeyArray_S31reg_gff_1_SFF_7_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S31reg_gff_1_SFF_7_MUXInst_Y), .B0_t (KeyArray_outS32ser[7]), .Z0_t (KeyArray_S31reg_gff_1_SFF_7_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S32reg_gff_1_SFF_0_U3 ( .A0_t (KeyArray_S32reg_gff_1_SFF_0_n2), .B0_t (KeyArray_S32reg_gff_1_SFF_0_n1), .Z0_t (KeyArray_outS32ser[0]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_0_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS32ser[0]), .Z0_t (KeyArray_S32reg_gff_1_SFF_0_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_0_U1 ( .A0_t (KeyArray_S32reg_gff_1_SFF_0_QD), .B0_t (enKS), .Z0_t (KeyArray_S32reg_gff_1_SFF_0_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS33ser[0]), .B0_t (KeyArray_outS02ser[0]), .Z0_t (KeyArray_S32reg_gff_1_SFF_0_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S32reg_gff_1_SFF_0_MUXInst_X), .Z0_t (KeyArray_S32reg_gff_1_SFF_0_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S32reg_gff_1_SFF_0_MUXInst_Y), .B0_t (KeyArray_outS33ser[0]), .Z0_t (KeyArray_S32reg_gff_1_SFF_0_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S32reg_gff_1_SFF_1_U3 ( .A0_t (KeyArray_S32reg_gff_1_SFF_1_n2), .B0_t (KeyArray_S32reg_gff_1_SFF_1_n1), .Z0_t (KeyArray_outS32ser[1]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_1_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS32ser[1]), .Z0_t (KeyArray_S32reg_gff_1_SFF_1_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_1_U1 ( .A0_t (KeyArray_S32reg_gff_1_SFF_1_QD), .B0_t (enKS), .Z0_t (KeyArray_S32reg_gff_1_SFF_1_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS33ser[1]), .B0_t (KeyArray_outS02ser[1]), .Z0_t (KeyArray_S32reg_gff_1_SFF_1_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S32reg_gff_1_SFF_1_MUXInst_X), .Z0_t (KeyArray_S32reg_gff_1_SFF_1_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S32reg_gff_1_SFF_1_MUXInst_Y), .B0_t (KeyArray_outS33ser[1]), .Z0_t (KeyArray_S32reg_gff_1_SFF_1_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S32reg_gff_1_SFF_2_U3 ( .A0_t (KeyArray_S32reg_gff_1_SFF_2_n2), .B0_t (KeyArray_S32reg_gff_1_SFF_2_n1), .Z0_t (KeyArray_outS32ser[2]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_2_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS32ser[2]), .Z0_t (KeyArray_S32reg_gff_1_SFF_2_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_2_U1 ( .A0_t (KeyArray_S32reg_gff_1_SFF_2_QD), .B0_t (enKS), .Z0_t (KeyArray_S32reg_gff_1_SFF_2_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS33ser[2]), .B0_t (KeyArray_outS02ser[2]), .Z0_t (KeyArray_S32reg_gff_1_SFF_2_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S32reg_gff_1_SFF_2_MUXInst_X), .Z0_t (KeyArray_S32reg_gff_1_SFF_2_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S32reg_gff_1_SFF_2_MUXInst_Y), .B0_t (KeyArray_outS33ser[2]), .Z0_t (KeyArray_S32reg_gff_1_SFF_2_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S32reg_gff_1_SFF_3_U3 ( .A0_t (KeyArray_S32reg_gff_1_SFF_3_n2), .B0_t (KeyArray_S32reg_gff_1_SFF_3_n1), .Z0_t (KeyArray_outS32ser[3]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_3_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS32ser[3]), .Z0_t (KeyArray_S32reg_gff_1_SFF_3_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_3_U1 ( .A0_t (KeyArray_S32reg_gff_1_SFF_3_QD), .B0_t (enKS), .Z0_t (KeyArray_S32reg_gff_1_SFF_3_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS33ser[3]), .B0_t (KeyArray_outS02ser[3]), .Z0_t (KeyArray_S32reg_gff_1_SFF_3_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S32reg_gff_1_SFF_3_MUXInst_X), .Z0_t (KeyArray_S32reg_gff_1_SFF_3_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S32reg_gff_1_SFF_3_MUXInst_Y), .B0_t (KeyArray_outS33ser[3]), .Z0_t (KeyArray_S32reg_gff_1_SFF_3_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S32reg_gff_1_SFF_4_U3 ( .A0_t (KeyArray_S32reg_gff_1_SFF_4_n2), .B0_t (KeyArray_S32reg_gff_1_SFF_4_n1), .Z0_t (KeyArray_outS32ser[4]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_4_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS32ser[4]), .Z0_t (KeyArray_S32reg_gff_1_SFF_4_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_4_U1 ( .A0_t (KeyArray_S32reg_gff_1_SFF_4_QD), .B0_t (enKS), .Z0_t (KeyArray_S32reg_gff_1_SFF_4_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS33ser[4]), .B0_t (KeyArray_outS02ser[4]), .Z0_t (KeyArray_S32reg_gff_1_SFF_4_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S32reg_gff_1_SFF_4_MUXInst_X), .Z0_t (KeyArray_S32reg_gff_1_SFF_4_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S32reg_gff_1_SFF_4_MUXInst_Y), .B0_t (KeyArray_outS33ser[4]), .Z0_t (KeyArray_S32reg_gff_1_SFF_4_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S32reg_gff_1_SFF_5_U3 ( .A0_t (KeyArray_S32reg_gff_1_SFF_5_n2), .B0_t (KeyArray_S32reg_gff_1_SFF_5_n1), .Z0_t (KeyArray_outS32ser[5]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_5_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS32ser[5]), .Z0_t (KeyArray_S32reg_gff_1_SFF_5_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_5_U1 ( .A0_t (KeyArray_S32reg_gff_1_SFF_5_QD), .B0_t (enKS), .Z0_t (KeyArray_S32reg_gff_1_SFF_5_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS33ser[5]), .B0_t (KeyArray_outS02ser[5]), .Z0_t (KeyArray_S32reg_gff_1_SFF_5_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S32reg_gff_1_SFF_5_MUXInst_X), .Z0_t (KeyArray_S32reg_gff_1_SFF_5_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S32reg_gff_1_SFF_5_MUXInst_Y), .B0_t (KeyArray_outS33ser[5]), .Z0_t (KeyArray_S32reg_gff_1_SFF_5_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S32reg_gff_1_SFF_6_U3 ( .A0_t (KeyArray_S32reg_gff_1_SFF_6_n2), .B0_t (KeyArray_S32reg_gff_1_SFF_6_n1), .Z0_t (KeyArray_outS32ser[6]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_6_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS32ser[6]), .Z0_t (KeyArray_S32reg_gff_1_SFF_6_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_6_U1 ( .A0_t (KeyArray_S32reg_gff_1_SFF_6_QD), .B0_t (enKS), .Z0_t (KeyArray_S32reg_gff_1_SFF_6_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS33ser[6]), .B0_t (KeyArray_outS02ser[6]), .Z0_t (KeyArray_S32reg_gff_1_SFF_6_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S32reg_gff_1_SFF_6_MUXInst_X), .Z0_t (KeyArray_S32reg_gff_1_SFF_6_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S32reg_gff_1_SFF_6_MUXInst_Y), .B0_t (KeyArray_outS33ser[6]), .Z0_t (KeyArray_S32reg_gff_1_SFF_6_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S32reg_gff_1_SFF_7_U3 ( .A0_t (KeyArray_S32reg_gff_1_SFF_7_n2), .B0_t (KeyArray_S32reg_gff_1_SFF_7_n1), .Z0_t (KeyArray_outS32ser[7]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_7_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS32ser[7]), .Z0_t (KeyArray_S32reg_gff_1_SFF_7_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_7_U1 ( .A0_t (KeyArray_S32reg_gff_1_SFF_7_QD), .B0_t (enKS), .Z0_t (KeyArray_S32reg_gff_1_SFF_7_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS33ser[7]), .B0_t (KeyArray_outS02ser[7]), .Z0_t (KeyArray_S32reg_gff_1_SFF_7_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S32reg_gff_1_SFF_7_MUXInst_X), .Z0_t (KeyArray_S32reg_gff_1_SFF_7_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S32reg_gff_1_SFF_7_MUXInst_Y), .B0_t (KeyArray_outS33ser[7]), .Z0_t (KeyArray_S32reg_gff_1_SFF_7_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S33reg_gff_1_SFF_0_U3 ( .A0_t (KeyArray_S33reg_gff_1_SFF_0_n2), .B0_t (KeyArray_S33reg_gff_1_SFF_0_n1), .Z0_t (KeyArray_outS33ser[0]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_0_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS33ser[0]), .Z0_t (KeyArray_S33reg_gff_1_SFF_0_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_0_U1 ( .A0_t (KeyArray_S33reg_gff_1_SFF_0_QD), .B0_t (enKS), .Z0_t (KeyArray_S33reg_gff_1_SFF_0_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS33ser[0]), .B0_t (KeyArray_outS03ser[0]), .Z0_t (KeyArray_S33reg_gff_1_SFF_0_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S33reg_gff_1_SFF_0_MUXInst_X), .Z0_t (KeyArray_S33reg_gff_1_SFF_0_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S33reg_gff_1_SFF_0_MUXInst_Y), .B0_t (KeyArray_inS33ser[0]), .Z0_t (KeyArray_S33reg_gff_1_SFF_0_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S33reg_gff_1_SFF_1_U3 ( .A0_t (KeyArray_S33reg_gff_1_SFF_1_n2), .B0_t (KeyArray_S33reg_gff_1_SFF_1_n1), .Z0_t (KeyArray_outS33ser[1]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_1_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS33ser[1]), .Z0_t (KeyArray_S33reg_gff_1_SFF_1_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_1_U1 ( .A0_t (KeyArray_S33reg_gff_1_SFF_1_QD), .B0_t (enKS), .Z0_t (KeyArray_S33reg_gff_1_SFF_1_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS33ser[1]), .B0_t (KeyArray_outS03ser[1]), .Z0_t (KeyArray_S33reg_gff_1_SFF_1_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S33reg_gff_1_SFF_1_MUXInst_X), .Z0_t (KeyArray_S33reg_gff_1_SFF_1_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S33reg_gff_1_SFF_1_MUXInst_Y), .B0_t (KeyArray_inS33ser[1]), .Z0_t (KeyArray_S33reg_gff_1_SFF_1_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S33reg_gff_1_SFF_2_U3 ( .A0_t (KeyArray_S33reg_gff_1_SFF_2_n2), .B0_t (KeyArray_S33reg_gff_1_SFF_2_n1), .Z0_t (KeyArray_outS33ser[2]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_2_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS33ser[2]), .Z0_t (KeyArray_S33reg_gff_1_SFF_2_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_2_U1 ( .A0_t (KeyArray_S33reg_gff_1_SFF_2_QD), .B0_t (enKS), .Z0_t (KeyArray_S33reg_gff_1_SFF_2_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS33ser[2]), .B0_t (KeyArray_outS03ser[2]), .Z0_t (KeyArray_S33reg_gff_1_SFF_2_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S33reg_gff_1_SFF_2_MUXInst_X), .Z0_t (KeyArray_S33reg_gff_1_SFF_2_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S33reg_gff_1_SFF_2_MUXInst_Y), .B0_t (KeyArray_inS33ser[2]), .Z0_t (KeyArray_S33reg_gff_1_SFF_2_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S33reg_gff_1_SFF_3_U3 ( .A0_t (KeyArray_S33reg_gff_1_SFF_3_n2), .B0_t (KeyArray_S33reg_gff_1_SFF_3_n1), .Z0_t (KeyArray_outS33ser[3]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_3_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS33ser[3]), .Z0_t (KeyArray_S33reg_gff_1_SFF_3_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_3_U1 ( .A0_t (KeyArray_S33reg_gff_1_SFF_3_QD), .B0_t (enKS), .Z0_t (KeyArray_S33reg_gff_1_SFF_3_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS33ser[3]), .B0_t (KeyArray_outS03ser[3]), .Z0_t (KeyArray_S33reg_gff_1_SFF_3_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S33reg_gff_1_SFF_3_MUXInst_X), .Z0_t (KeyArray_S33reg_gff_1_SFF_3_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S33reg_gff_1_SFF_3_MUXInst_Y), .B0_t (KeyArray_inS33ser[3]), .Z0_t (KeyArray_S33reg_gff_1_SFF_3_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S33reg_gff_1_SFF_4_U3 ( .A0_t (KeyArray_S33reg_gff_1_SFF_4_n2), .B0_t (KeyArray_S33reg_gff_1_SFF_4_n1), .Z0_t (KeyArray_outS33ser[4]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_4_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS33ser[4]), .Z0_t (KeyArray_S33reg_gff_1_SFF_4_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_4_U1 ( .A0_t (KeyArray_S33reg_gff_1_SFF_4_QD), .B0_t (enKS), .Z0_t (KeyArray_S33reg_gff_1_SFF_4_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS33ser[4]), .B0_t (KeyArray_outS03ser[4]), .Z0_t (KeyArray_S33reg_gff_1_SFF_4_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S33reg_gff_1_SFF_4_MUXInst_X), .Z0_t (KeyArray_S33reg_gff_1_SFF_4_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S33reg_gff_1_SFF_4_MUXInst_Y), .B0_t (KeyArray_inS33ser[4]), .Z0_t (KeyArray_S33reg_gff_1_SFF_4_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S33reg_gff_1_SFF_5_U3 ( .A0_t (KeyArray_S33reg_gff_1_SFF_5_n2), .B0_t (KeyArray_S33reg_gff_1_SFF_5_n1), .Z0_t (KeyArray_outS33ser[5]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_5_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS33ser[5]), .Z0_t (KeyArray_S33reg_gff_1_SFF_5_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_5_U1 ( .A0_t (KeyArray_S33reg_gff_1_SFF_5_QD), .B0_t (enKS), .Z0_t (KeyArray_S33reg_gff_1_SFF_5_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS33ser[5]), .B0_t (KeyArray_outS03ser[5]), .Z0_t (KeyArray_S33reg_gff_1_SFF_5_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S33reg_gff_1_SFF_5_MUXInst_X), .Z0_t (KeyArray_S33reg_gff_1_SFF_5_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S33reg_gff_1_SFF_5_MUXInst_Y), .B0_t (KeyArray_inS33ser[5]), .Z0_t (KeyArray_S33reg_gff_1_SFF_5_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S33reg_gff_1_SFF_6_U3 ( .A0_t (KeyArray_S33reg_gff_1_SFF_6_n2), .B0_t (KeyArray_S33reg_gff_1_SFF_6_n1), .Z0_t (KeyArray_outS33ser[6]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_6_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS33ser[6]), .Z0_t (KeyArray_S33reg_gff_1_SFF_6_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_6_U1 ( .A0_t (KeyArray_S33reg_gff_1_SFF_6_QD), .B0_t (enKS), .Z0_t (KeyArray_S33reg_gff_1_SFF_6_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS33ser[6]), .B0_t (KeyArray_outS03ser[6]), .Z0_t (KeyArray_S33reg_gff_1_SFF_6_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S33reg_gff_1_SFF_6_MUXInst_X), .Z0_t (KeyArray_S33reg_gff_1_SFF_6_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S33reg_gff_1_SFF_6_MUXInst_Y), .B0_t (KeyArray_inS33ser[6]), .Z0_t (KeyArray_S33reg_gff_1_SFF_6_QD) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S33reg_gff_1_SFF_7_U3 ( .A0_t (KeyArray_S33reg_gff_1_SFF_7_n2), .B0_t (KeyArray_S33reg_gff_1_SFF_7_n1), .Z0_t (KeyArray_outS33ser[7]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_7_U2 ( .A0_t (enKS), .B0_t (KeyArray_outS33ser[7]), .Z0_t (KeyArray_S33reg_gff_1_SFF_7_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_7_U1 ( .A0_t (KeyArray_S33reg_gff_1_SFF_7_QD), .B0_t (enKS), .Z0_t (KeyArray_S33reg_gff_1_SFF_7_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS33ser[7]), .B0_t (KeyArray_outS03ser[7]), .Z0_t (KeyArray_S33reg_gff_1_SFF_7_MUXInst_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (selMC), .B0_t (KeyArray_S33reg_gff_1_SFF_7_MUXInst_X), .Z0_t (KeyArray_S33reg_gff_1_SFF_7_MUXInst_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S33reg_gff_1_SFF_7_MUXInst_Y), .B0_t (KeyArray_inS33ser[7]), .Z0_t (KeyArray_S33reg_gff_1_SFF_7_QD) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_0_XOR1_U1 ( .A0_t (KeyArray_outS01ser_0_), .B0_t (KeyArray_outS01ser_XOR_00[0]), .Z0_t (KeyArray_MUX_inS00ser_mux_inst_0_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_0_AND1_U1 ( .A0_t (KeyArray_nReset_selXOR), .B0_t (KeyArray_MUX_inS00ser_mux_inst_0_X), .Z0_t (KeyArray_MUX_inS00ser_mux_inst_0_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_0_XOR2_U1 ( .A0_t (KeyArray_MUX_inS00ser_mux_inst_0_Y), .B0_t (KeyArray_outS01ser_0_), .Z0_t (KeyArray_inS00ser[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_1_XOR1_U1 ( .A0_t (KeyArray_outS01ser_1_), .B0_t (KeyArray_outS01ser_XOR_00[1]), .Z0_t (KeyArray_MUX_inS00ser_mux_inst_1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_1_AND1_U1 ( .A0_t (KeyArray_nReset_selXOR), .B0_t (KeyArray_MUX_inS00ser_mux_inst_1_X), .Z0_t (KeyArray_MUX_inS00ser_mux_inst_1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_1_XOR2_U1 ( .A0_t (KeyArray_MUX_inS00ser_mux_inst_1_Y), .B0_t (KeyArray_outS01ser_1_), .Z0_t (KeyArray_inS00ser[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_2_XOR1_U1 ( .A0_t (KeyArray_outS01ser_2_), .B0_t (KeyArray_outS01ser_XOR_00[2]), .Z0_t (KeyArray_MUX_inS00ser_mux_inst_2_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_2_AND1_U1 ( .A0_t (KeyArray_nReset_selXOR), .B0_t (KeyArray_MUX_inS00ser_mux_inst_2_X), .Z0_t (KeyArray_MUX_inS00ser_mux_inst_2_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_2_XOR2_U1 ( .A0_t (KeyArray_MUX_inS00ser_mux_inst_2_Y), .B0_t (KeyArray_outS01ser_2_), .Z0_t (KeyArray_inS00ser[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_3_XOR1_U1 ( .A0_t (KeyArray_outS01ser_3_), .B0_t (KeyArray_outS01ser_XOR_00[3]), .Z0_t (KeyArray_MUX_inS00ser_mux_inst_3_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_3_AND1_U1 ( .A0_t (KeyArray_nReset_selXOR), .B0_t (KeyArray_MUX_inS00ser_mux_inst_3_X), .Z0_t (KeyArray_MUX_inS00ser_mux_inst_3_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_3_XOR2_U1 ( .A0_t (KeyArray_MUX_inS00ser_mux_inst_3_Y), .B0_t (KeyArray_outS01ser_3_), .Z0_t (KeyArray_inS00ser[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_4_XOR1_U1 ( .A0_t (KeyArray_outS01ser_4_), .B0_t (KeyArray_outS01ser_XOR_00[4]), .Z0_t (KeyArray_MUX_inS00ser_mux_inst_4_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_4_AND1_U1 ( .A0_t (KeyArray_nReset_selXOR), .B0_t (KeyArray_MUX_inS00ser_mux_inst_4_X), .Z0_t (KeyArray_MUX_inS00ser_mux_inst_4_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_4_XOR2_U1 ( .A0_t (KeyArray_MUX_inS00ser_mux_inst_4_Y), .B0_t (KeyArray_outS01ser_4_), .Z0_t (KeyArray_inS00ser[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_5_XOR1_U1 ( .A0_t (KeyArray_outS01ser_5_), .B0_t (KeyArray_outS01ser_XOR_00[5]), .Z0_t (KeyArray_MUX_inS00ser_mux_inst_5_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_5_AND1_U1 ( .A0_t (KeyArray_nReset_selXOR), .B0_t (KeyArray_MUX_inS00ser_mux_inst_5_X), .Z0_t (KeyArray_MUX_inS00ser_mux_inst_5_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_5_XOR2_U1 ( .A0_t (KeyArray_MUX_inS00ser_mux_inst_5_Y), .B0_t (KeyArray_outS01ser_5_), .Z0_t (KeyArray_inS00ser[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_6_XOR1_U1 ( .A0_t (KeyArray_outS01ser_6_), .B0_t (KeyArray_outS01ser_XOR_00[6]), .Z0_t (KeyArray_MUX_inS00ser_mux_inst_6_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_6_AND1_U1 ( .A0_t (KeyArray_nReset_selXOR), .B0_t (KeyArray_MUX_inS00ser_mux_inst_6_X), .Z0_t (KeyArray_MUX_inS00ser_mux_inst_6_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_6_XOR2_U1 ( .A0_t (KeyArray_MUX_inS00ser_mux_inst_6_Y), .B0_t (KeyArray_outS01ser_6_), .Z0_t (KeyArray_inS00ser[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_7_XOR1_U1 ( .A0_t (KeyArray_outS01ser_7_), .B0_t (KeyArray_outS01ser_XOR_00[7]), .Z0_t (KeyArray_MUX_inS00ser_mux_inst_7_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_7_AND1_U1 ( .A0_t (KeyArray_nReset_selXOR), .B0_t (KeyArray_MUX_inS00ser_mux_inst_7_X), .Z0_t (KeyArray_MUX_inS00ser_mux_inst_7_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_7_XOR2_U1 ( .A0_t (KeyArray_MUX_inS00ser_mux_inst_7_Y), .B0_t (KeyArray_outS01ser_7_), .Z0_t (KeyArray_inS00ser[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_0_XOR1_U1 ( .A0_t (port_out[0]), .B0_t (keyStateIn[0]), .Z0_t (KeyArray_MUX_inS33ser_mux_inst_0_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_0_AND1_U1 ( .A0_t (start), .B0_t (KeyArray_MUX_inS33ser_mux_inst_0_X), .Z0_t (KeyArray_MUX_inS33ser_mux_inst_0_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_0_XOR2_U1 ( .A0_t (KeyArray_MUX_inS33ser_mux_inst_0_Y), .B0_t (port_out[0]), .Z0_t (KeyArray_inS33ser[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_1_XOR1_U1 ( .A0_t (port_out[1]), .B0_t (keyStateIn[1]), .Z0_t (KeyArray_MUX_inS33ser_mux_inst_1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_1_AND1_U1 ( .A0_t (start), .B0_t (KeyArray_MUX_inS33ser_mux_inst_1_X), .Z0_t (KeyArray_MUX_inS33ser_mux_inst_1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_1_XOR2_U1 ( .A0_t (KeyArray_MUX_inS33ser_mux_inst_1_Y), .B0_t (port_out[1]), .Z0_t (KeyArray_inS33ser[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_2_XOR1_U1 ( .A0_t (port_out[2]), .B0_t (keyStateIn[2]), .Z0_t (KeyArray_MUX_inS33ser_mux_inst_2_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_2_AND1_U1 ( .A0_t (start), .B0_t (KeyArray_MUX_inS33ser_mux_inst_2_X), .Z0_t (KeyArray_MUX_inS33ser_mux_inst_2_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_2_XOR2_U1 ( .A0_t (KeyArray_MUX_inS33ser_mux_inst_2_Y), .B0_t (port_out[2]), .Z0_t (KeyArray_inS33ser[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_3_XOR1_U1 ( .A0_t (port_out[3]), .B0_t (keyStateIn[3]), .Z0_t (KeyArray_MUX_inS33ser_mux_inst_3_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_3_AND1_U1 ( .A0_t (start), .B0_t (KeyArray_MUX_inS33ser_mux_inst_3_X), .Z0_t (KeyArray_MUX_inS33ser_mux_inst_3_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_3_XOR2_U1 ( .A0_t (KeyArray_MUX_inS33ser_mux_inst_3_Y), .B0_t (port_out[3]), .Z0_t (KeyArray_inS33ser[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_4_XOR1_U1 ( .A0_t (port_out[4]), .B0_t (keyStateIn[4]), .Z0_t (KeyArray_MUX_inS33ser_mux_inst_4_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_4_AND1_U1 ( .A0_t (start), .B0_t (KeyArray_MUX_inS33ser_mux_inst_4_X), .Z0_t (KeyArray_MUX_inS33ser_mux_inst_4_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_4_XOR2_U1 ( .A0_t (KeyArray_MUX_inS33ser_mux_inst_4_Y), .B0_t (port_out[4]), .Z0_t (KeyArray_inS33ser[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_5_XOR1_U1 ( .A0_t (port_out[5]), .B0_t (keyStateIn[5]), .Z0_t (KeyArray_MUX_inS33ser_mux_inst_5_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_5_AND1_U1 ( .A0_t (start), .B0_t (KeyArray_MUX_inS33ser_mux_inst_5_X), .Z0_t (KeyArray_MUX_inS33ser_mux_inst_5_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_5_XOR2_U1 ( .A0_t (KeyArray_MUX_inS33ser_mux_inst_5_Y), .B0_t (port_out[5]), .Z0_t (KeyArray_inS33ser[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_6_XOR1_U1 ( .A0_t (port_out[6]), .B0_t (keyStateIn[6]), .Z0_t (KeyArray_MUX_inS33ser_mux_inst_6_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_6_AND1_U1 ( .A0_t (start), .B0_t (KeyArray_MUX_inS33ser_mux_inst_6_X), .Z0_t (KeyArray_MUX_inS33ser_mux_inst_6_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_6_XOR2_U1 ( .A0_t (KeyArray_MUX_inS33ser_mux_inst_6_Y), .B0_t (port_out[6]), .Z0_t (KeyArray_inS33ser[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_7_XOR1_U1 ( .A0_t (port_out[7]), .B0_t (keyStateIn[7]), .Z0_t (KeyArray_MUX_inS33ser_mux_inst_7_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_7_AND1_U1 ( .A0_t (start), .B0_t (KeyArray_MUX_inS33ser_mux_inst_7_X), .Z0_t (KeyArray_MUX_inS33ser_mux_inst_7_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_7_XOR2_U1 ( .A0_t (KeyArray_MUX_inS33ser_mux_inst_7_Y), .B0_t (port_out[7]), .Z0_t (KeyArray_inS33ser[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line0_U24 ( .A0_t (MixColumns_line0_n16), .B0_t (MixColumns_line0_n15), .Z0_t (MCout[31]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line0_U23 ( .A0_t (MixColumns_line2_S02[0]), .B0_t (MixColumns_line3_S02[0]), .Z0_t (MixColumns_line0_n15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_U22 ( .A0_t (port_out[6]), .B0_t (MixColumns_line0_S13[7]), .Z0_t (MixColumns_line0_n16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line0_U21 ( .A0_t (MixColumns_line0_n14), .B0_t (MixColumns_line0_n13), .Z0_t (MCout[30]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line0_U20 ( .A0_t (MixColumns_line2_S02[7]), .B0_t (MixColumns_line3_S02[7]), .Z0_t (MixColumns_line0_n13) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_U19 ( .A0_t (port_out[5]), .B0_t (MixColumns_line0_S13[6]), .Z0_t (MixColumns_line0_n14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line0_U18 ( .A0_t (MixColumns_line0_n12), .B0_t (MixColumns_line0_n11), .Z0_t (MCout[29]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line0_U17 ( .A0_t (MixColumns_line2_S02[6]), .B0_t (MixColumns_line3_S02[6]), .Z0_t (MixColumns_line0_n11) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_U16 ( .A0_t (port_out[4]), .B0_t (MixColumns_line0_S13[5]), .Z0_t (MixColumns_line0_n12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line0_U15 ( .A0_t (MixColumns_line0_n10), .B0_t (MixColumns_line0_n9), .Z0_t (MCout[28]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line0_U14 ( .A0_t (MixColumns_line2_S02[5]), .B0_t (MixColumns_line3_S02[5]), .Z0_t (MixColumns_line0_n9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_U13 ( .A0_t (MixColumns_line0_S02[4]), .B0_t (MixColumns_line0_S13[4]), .Z0_t (MixColumns_line0_n10) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line0_U12 ( .A0_t (MixColumns_line0_n8), .B0_t (MixColumns_line0_n7), .Z0_t (MCout[27]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line0_U11 ( .A0_t (MCin[11]), .B0_t (MCin[3]), .Z0_t (MixColumns_line0_n7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_U10 ( .A0_t (MixColumns_line0_S02[3]), .B0_t (MixColumns_line0_S13[3]), .Z0_t (MixColumns_line0_n8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line0_U9 ( .A0_t (MixColumns_line0_n6), .B0_t (MixColumns_line0_n5), .Z0_t (MCout[26]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line0_U8 ( .A0_t (MCin[10]), .B0_t (MCin[2]), .Z0_t (MixColumns_line0_n5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_U7 ( .A0_t (port_out[1]), .B0_t (MixColumns_line0_S13[2]), .Z0_t (MixColumns_line0_n6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line0_U6 ( .A0_t (MixColumns_line0_n4), .B0_t (MixColumns_line0_n3), .Z0_t (MCout[25]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line0_U5 ( .A0_t (MixColumns_line3_S02[2]), .B0_t (MixColumns_line2_S02[2]), .Z0_t (MixColumns_line0_n3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_U4 ( .A0_t (MixColumns_line0_S02[1]), .B0_t (MixColumns_line0_S13[1]), .Z0_t (MixColumns_line0_n4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line0_U3 ( .A0_t (MixColumns_line0_n2), .B0_t (MixColumns_line0_n1), .Z0_t (MCout[24]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line0_U2 ( .A0_t (MCin[0]), .B0_t (MCin[8]), .Z0_t (MixColumns_line0_n1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_U1 ( .A0_t (port_out[7]), .B0_t (MixColumns_line0_S13[0]), .Z0_t (MixColumns_line0_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_timesTWO_U3 ( .A0_t (port_out[7]), .B0_t (port_out[3]), .Z0_t (MixColumns_line0_S02[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_timesTWO_U2 ( .A0_t (port_out[7]), .B0_t (port_out[2]), .Z0_t (MixColumns_line0_S02[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_timesTWO_U1 ( .A0_t (port_out[7]), .B0_t (port_out[0]), .Z0_t (MixColumns_line0_S02[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_timesTHREE_U8 ( .A0_t (MixColumns_line1_S02[0]), .B0_t (MixColumns_line1_S02[7]), .Z0_t (MixColumns_line0_S13[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_timesTHREE_U7 ( .A0_t (MixColumns_line1_S02[7]), .B0_t (MixColumns_line1_S02[6]), .Z0_t (MixColumns_line0_S13[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_timesTHREE_U6 ( .A0_t (MixColumns_line1_S02[6]), .B0_t (MixColumns_line1_S02[5]), .Z0_t (MixColumns_line0_S13[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_timesTHREE_U5 ( .A0_t (MixColumns_line1_S02[5]), .B0_t (MixColumns_line0_timesTHREE_input2[4]), .Z0_t (MixColumns_line0_S13[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_timesTHREE_U4 ( .A0_t (MCin[19]), .B0_t (MixColumns_line0_timesTHREE_input2[3]), .Z0_t (MixColumns_line0_S13[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_timesTHREE_U3 ( .A0_t (MCin[18]), .B0_t (MixColumns_line1_S02[2]), .Z0_t (MixColumns_line0_S13[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_timesTHREE_U2 ( .A0_t (MixColumns_line1_S02[2]), .B0_t (MixColumns_line0_timesTHREE_input2[1]), .Z0_t (MixColumns_line0_S13[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_timesTHREE_U1 ( .A0_t (MCin[16]), .B0_t (MixColumns_line1_S02[0]), .Z0_t (MixColumns_line0_S13[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_timesTHREE_timesTWO_U3 ( .A0_t (MixColumns_line1_S02[0]), .B0_t (MCin[19]), .Z0_t (MixColumns_line0_timesTHREE_input2[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_timesTHREE_timesTWO_U2 ( .A0_t (MixColumns_line1_S02[0]), .B0_t (MCin[18]), .Z0_t (MixColumns_line0_timesTHREE_input2[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_timesTHREE_timesTWO_U1 ( .A0_t (MixColumns_line1_S02[0]), .B0_t (MCin[16]), .Z0_t (MixColumns_line0_timesTHREE_input2[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line1_U24 ( .A0_t (MixColumns_line1_n16), .B0_t (MixColumns_line1_n15), .Z0_t (MCout[23]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line1_U23 ( .A0_t (MixColumns_line3_S02[0]), .B0_t (port_out[7]), .Z0_t (MixColumns_line1_n15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_U22 ( .A0_t (MixColumns_line1_S02[7]), .B0_t (MixColumns_line1_S13[7]), .Z0_t (MixColumns_line1_n16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line1_U21 ( .A0_t (MixColumns_line1_n14), .B0_t (MixColumns_line1_n13), .Z0_t (MCout[22]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line1_U20 ( .A0_t (MixColumns_line3_S02[7]), .B0_t (port_out[6]), .Z0_t (MixColumns_line1_n13) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_U19 ( .A0_t (MixColumns_line1_S02[6]), .B0_t (MixColumns_line1_S13[6]), .Z0_t (MixColumns_line1_n14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line1_U18 ( .A0_t (MixColumns_line1_n12), .B0_t (MixColumns_line1_n11), .Z0_t (MCout[21]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line1_U17 ( .A0_t (MixColumns_line3_S02[6]), .B0_t (port_out[5]), .Z0_t (MixColumns_line1_n11) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_U16 ( .A0_t (MixColumns_line1_S02[5]), .B0_t (MixColumns_line1_S13[5]), .Z0_t (MixColumns_line1_n12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line1_U15 ( .A0_t (MixColumns_line1_n10), .B0_t (MixColumns_line1_n9), .Z0_t (MCout[20]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line1_U14 ( .A0_t (MixColumns_line3_S02[5]), .B0_t (port_out[4]), .Z0_t (MixColumns_line1_n9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_U13 ( .A0_t (MixColumns_line1_S02[4]), .B0_t (MixColumns_line1_S13[4]), .Z0_t (MixColumns_line1_n10) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line1_U12 ( .A0_t (MixColumns_line1_n8), .B0_t (MixColumns_line1_n7), .Z0_t (MCout[19]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line1_U11 ( .A0_t (MCin[3]), .B0_t (port_out[3]), .Z0_t (MixColumns_line1_n7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_U10 ( .A0_t (MixColumns_line1_S02[3]), .B0_t (MixColumns_line1_S13[3]), .Z0_t (MixColumns_line1_n8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line1_U9 ( .A0_t (MixColumns_line1_n6), .B0_t (MixColumns_line1_n5), .Z0_t (MCout[18]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line1_U8 ( .A0_t (MCin[2]), .B0_t (port_out[2]), .Z0_t (MixColumns_line1_n5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_U7 ( .A0_t (MixColumns_line1_S02[2]), .B0_t (MixColumns_line1_S13[2]), .Z0_t (MixColumns_line1_n6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line1_U6 ( .A0_t (MixColumns_line1_n4), .B0_t (MixColumns_line1_n3), .Z0_t (MCout[17]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line1_U5 ( .A0_t (port_out[1]), .B0_t (MixColumns_line3_S02[2]), .Z0_t (MixColumns_line1_n3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_U4 ( .A0_t (MixColumns_line1_S02[1]), .B0_t (MixColumns_line1_S13[1]), .Z0_t (MixColumns_line1_n4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line1_U3 ( .A0_t (MixColumns_line1_n2), .B0_t (MixColumns_line1_n1), .Z0_t (MCout[16]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line1_U2 ( .A0_t (port_out[0]), .B0_t (MCin[0]), .Z0_t (MixColumns_line1_n1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_U1 ( .A0_t (MixColumns_line1_S02[0]), .B0_t (MixColumns_line1_S13[0]), .Z0_t (MixColumns_line1_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_timesTWO_U3 ( .A0_t (MixColumns_line1_S02[0]), .B0_t (MCin[19]), .Z0_t (MixColumns_line1_S02[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_timesTWO_U2 ( .A0_t (MixColumns_line1_S02[0]), .B0_t (MCin[18]), .Z0_t (MixColumns_line1_S02[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_timesTWO_U1 ( .A0_t (MixColumns_line1_S02[0]), .B0_t (MCin[16]), .Z0_t (MixColumns_line1_S02[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_timesTHREE_U8 ( .A0_t (MixColumns_line2_S02[0]), .B0_t (MixColumns_line2_S02[7]), .Z0_t (MixColumns_line1_S13[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_timesTHREE_U7 ( .A0_t (MixColumns_line2_S02[7]), .B0_t (MixColumns_line2_S02[6]), .Z0_t (MixColumns_line1_S13[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_timesTHREE_U6 ( .A0_t (MixColumns_line2_S02[6]), .B0_t (MixColumns_line2_S02[5]), .Z0_t (MixColumns_line1_S13[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_timesTHREE_U5 ( .A0_t (MixColumns_line2_S02[5]), .B0_t (MixColumns_line1_timesTHREE_input2[4]), .Z0_t (MixColumns_line1_S13[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_timesTHREE_U4 ( .A0_t (MCin[11]), .B0_t (MixColumns_line1_timesTHREE_input2[3]), .Z0_t (MixColumns_line1_S13[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_timesTHREE_U3 ( .A0_t (MCin[10]), .B0_t (MixColumns_line2_S02[2]), .Z0_t (MixColumns_line1_S13[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_timesTHREE_U2 ( .A0_t (MixColumns_line2_S02[2]), .B0_t (MixColumns_line1_timesTHREE_input2[1]), .Z0_t (MixColumns_line1_S13[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_timesTHREE_U1 ( .A0_t (MCin[8]), .B0_t (MixColumns_line2_S02[0]), .Z0_t (MixColumns_line1_S13[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_timesTHREE_timesTWO_U3 ( .A0_t (MixColumns_line2_S02[0]), .B0_t (MCin[11]), .Z0_t (MixColumns_line1_timesTHREE_input2[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_timesTHREE_timesTWO_U2 ( .A0_t (MixColumns_line2_S02[0]), .B0_t (MCin[10]), .Z0_t (MixColumns_line1_timesTHREE_input2[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_timesTHREE_timesTWO_U1 ( .A0_t (MixColumns_line2_S02[0]), .B0_t (MCin[8]), .Z0_t (MixColumns_line1_timesTHREE_input2[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line2_U24 ( .A0_t (MixColumns_line2_n16), .B0_t (MixColumns_line2_n15), .Z0_t (MCout[15]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line2_U23 ( .A0_t (port_out[7]), .B0_t (MixColumns_line1_S02[0]), .Z0_t (MixColumns_line2_n15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_U22 ( .A0_t (MixColumns_line2_S02[7]), .B0_t (MixColumns_line2_S13[7]), .Z0_t (MixColumns_line2_n16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line2_U21 ( .A0_t (MixColumns_line2_n14), .B0_t (MixColumns_line2_n13), .Z0_t (MCout[14]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line2_U20 ( .A0_t (port_out[6]), .B0_t (MixColumns_line1_S02[7]), .Z0_t (MixColumns_line2_n13) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_U19 ( .A0_t (MixColumns_line2_S02[6]), .B0_t (MixColumns_line2_S13[6]), .Z0_t (MixColumns_line2_n14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line2_U18 ( .A0_t (MixColumns_line2_n12), .B0_t (MixColumns_line2_n11), .Z0_t (MCout[13]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line2_U17 ( .A0_t (port_out[5]), .B0_t (MixColumns_line1_S02[6]), .Z0_t (MixColumns_line2_n11) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_U16 ( .A0_t (MixColumns_line2_S02[5]), .B0_t (MixColumns_line2_S13[5]), .Z0_t (MixColumns_line2_n12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line2_U15 ( .A0_t (MixColumns_line2_n10), .B0_t (MixColumns_line2_n9), .Z0_t (MCout[12]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line2_U14 ( .A0_t (port_out[4]), .B0_t (MixColumns_line1_S02[5]), .Z0_t (MixColumns_line2_n9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_U13 ( .A0_t (MixColumns_line2_S02[4]), .B0_t (MixColumns_line2_S13[4]), .Z0_t (MixColumns_line2_n10) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line2_U12 ( .A0_t (MixColumns_line2_n8), .B0_t (MixColumns_line2_n7), .Z0_t (MCout[11]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line2_U11 ( .A0_t (port_out[3]), .B0_t (MCin[19]), .Z0_t (MixColumns_line2_n7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_U10 ( .A0_t (MixColumns_line2_S02[3]), .B0_t (MixColumns_line2_S13[3]), .Z0_t (MixColumns_line2_n8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line2_U9 ( .A0_t (MixColumns_line2_n6), .B0_t (MixColumns_line2_n5), .Z0_t (MCout[10]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line2_U8 ( .A0_t (port_out[2]), .B0_t (MCin[18]), .Z0_t (MixColumns_line2_n5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_U7 ( .A0_t (MixColumns_line2_S02[2]), .B0_t (MixColumns_line2_S13[2]), .Z0_t (MixColumns_line2_n6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line2_U6 ( .A0_t (MixColumns_line2_n4), .B0_t (MixColumns_line2_n3), .Z0_t (MCout[9]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line2_U5 ( .A0_t (MixColumns_line1_S02[2]), .B0_t (port_out[1]), .Z0_t (MixColumns_line2_n3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_U4 ( .A0_t (MixColumns_line2_S02[1]), .B0_t (MixColumns_line2_S13[1]), .Z0_t (MixColumns_line2_n4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line2_U3 ( .A0_t (MixColumns_line2_n2), .B0_t (MixColumns_line2_n1), .Z0_t (MCout[8]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line2_U2 ( .A0_t (MCin[16]), .B0_t (port_out[0]), .Z0_t (MixColumns_line2_n1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_U1 ( .A0_t (MixColumns_line2_S02[0]), .B0_t (MixColumns_line2_S13[0]), .Z0_t (MixColumns_line2_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_timesTWO_U3 ( .A0_t (MixColumns_line2_S02[0]), .B0_t (MCin[11]), .Z0_t (MixColumns_line2_S02[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_timesTWO_U2 ( .A0_t (MixColumns_line2_S02[0]), .B0_t (MCin[10]), .Z0_t (MixColumns_line2_S02[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_timesTWO_U1 ( .A0_t (MixColumns_line2_S02[0]), .B0_t (MCin[8]), .Z0_t (MixColumns_line2_S02[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_timesTHREE_U8 ( .A0_t (MixColumns_line3_S02[0]), .B0_t (MixColumns_line3_S02[7]), .Z0_t (MixColumns_line2_S13[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_timesTHREE_U7 ( .A0_t (MixColumns_line3_S02[7]), .B0_t (MixColumns_line3_S02[6]), .Z0_t (MixColumns_line2_S13[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_timesTHREE_U6 ( .A0_t (MixColumns_line3_S02[6]), .B0_t (MixColumns_line3_S02[5]), .Z0_t (MixColumns_line2_S13[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_timesTHREE_U5 ( .A0_t (MixColumns_line3_S02[5]), .B0_t (MixColumns_line2_timesTHREE_input2[4]), .Z0_t (MixColumns_line2_S13[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_timesTHREE_U4 ( .A0_t (MCin[3]), .B0_t (MixColumns_line2_timesTHREE_input2[3]), .Z0_t (MixColumns_line2_S13[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_timesTHREE_U3 ( .A0_t (MCin[2]), .B0_t (MixColumns_line3_S02[2]), .Z0_t (MixColumns_line2_S13[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_timesTHREE_U2 ( .A0_t (MixColumns_line3_S02[2]), .B0_t (MixColumns_line2_timesTHREE_input2[1]), .Z0_t (MixColumns_line2_S13[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_timesTHREE_U1 ( .A0_t (MCin[0]), .B0_t (MixColumns_line3_S02[0]), .Z0_t (MixColumns_line2_S13[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_timesTHREE_timesTWO_U3 ( .A0_t (MixColumns_line3_S02[0]), .B0_t (MCin[3]), .Z0_t (MixColumns_line2_timesTHREE_input2[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_timesTHREE_timesTWO_U2 ( .A0_t (MixColumns_line3_S02[0]), .B0_t (MCin[2]), .Z0_t (MixColumns_line2_timesTHREE_input2[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_timesTHREE_timesTWO_U1 ( .A0_t (MixColumns_line3_S02[0]), .B0_t (MCin[0]), .Z0_t (MixColumns_line2_timesTHREE_input2[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line3_U24 ( .A0_t (MixColumns_line3_n16), .B0_t (MixColumns_line3_n15), .Z0_t (MCout[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line3_U23 ( .A0_t (MixColumns_line1_S02[0]), .B0_t (MixColumns_line2_S02[0]), .Z0_t (MixColumns_line3_n15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_U22 ( .A0_t (MixColumns_line3_S02[7]), .B0_t (MixColumns_line3_S13[7]), .Z0_t (MixColumns_line3_n16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line3_U21 ( .A0_t (MixColumns_line3_n14), .B0_t (MixColumns_line3_n13), .Z0_t (MCout[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line3_U20 ( .A0_t (MixColumns_line1_S02[7]), .B0_t (MixColumns_line2_S02[7]), .Z0_t (MixColumns_line3_n13) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_U19 ( .A0_t (MixColumns_line3_S02[6]), .B0_t (MixColumns_line3_S13[6]), .Z0_t (MixColumns_line3_n14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line3_U18 ( .A0_t (MixColumns_line3_n12), .B0_t (MixColumns_line3_n11), .Z0_t (MCout[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line3_U17 ( .A0_t (MixColumns_line1_S02[6]), .B0_t (MixColumns_line2_S02[6]), .Z0_t (MixColumns_line3_n11) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_U16 ( .A0_t (MixColumns_line3_S02[5]), .B0_t (MixColumns_line3_S13[5]), .Z0_t (MixColumns_line3_n12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line3_U15 ( .A0_t (MixColumns_line3_n10), .B0_t (MixColumns_line3_n9), .Z0_t (MCout[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line3_U14 ( .A0_t (MixColumns_line1_S02[5]), .B0_t (MixColumns_line2_S02[5]), .Z0_t (MixColumns_line3_n9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_U13 ( .A0_t (MixColumns_line3_S02[4]), .B0_t (MixColumns_line3_S13[4]), .Z0_t (MixColumns_line3_n10) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line3_U12 ( .A0_t (MixColumns_line3_n8), .B0_t (MixColumns_line3_n7), .Z0_t (MCout[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line3_U11 ( .A0_t (MCin[19]), .B0_t (MCin[11]), .Z0_t (MixColumns_line3_n7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_U10 ( .A0_t (MixColumns_line3_S02[3]), .B0_t (MixColumns_line3_S13[3]), .Z0_t (MixColumns_line3_n8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line3_U9 ( .A0_t (MixColumns_line3_n6), .B0_t (MixColumns_line3_n5), .Z0_t (MCout[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line3_U8 ( .A0_t (MCin[18]), .B0_t (MCin[10]), .Z0_t (MixColumns_line3_n5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_U7 ( .A0_t (MixColumns_line3_S02[2]), .B0_t (MixColumns_line3_S13[2]), .Z0_t (MixColumns_line3_n6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line3_U6 ( .A0_t (MixColumns_line3_n4), .B0_t (MixColumns_line3_n3), .Z0_t (MCout[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line3_U5 ( .A0_t (MixColumns_line2_S02[2]), .B0_t (MixColumns_line1_S02[2]), .Z0_t (MixColumns_line3_n3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_U4 ( .A0_t (MixColumns_line3_S02[1]), .B0_t (MixColumns_line3_S13[1]), .Z0_t (MixColumns_line3_n4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line3_U3 ( .A0_t (MixColumns_line3_n2), .B0_t (MixColumns_line3_n1), .Z0_t (MCout[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line3_U2 ( .A0_t (MCin[8]), .B0_t (MCin[16]), .Z0_t (MixColumns_line3_n1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_U1 ( .A0_t (MixColumns_line3_S02[0]), .B0_t (MixColumns_line3_S13[0]), .Z0_t (MixColumns_line3_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_timesTWO_U3 ( .A0_t (MixColumns_line3_S02[0]), .B0_t (MCin[3]), .Z0_t (MixColumns_line3_S02[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_timesTWO_U2 ( .A0_t (MixColumns_line3_S02[0]), .B0_t (MCin[2]), .Z0_t (MixColumns_line3_S02[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_timesTWO_U1 ( .A0_t (MixColumns_line3_S02[0]), .B0_t (MCin[0]), .Z0_t (MixColumns_line3_S02[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_timesTHREE_U8 ( .A0_t (port_out[7]), .B0_t (port_out[6]), .Z0_t (MixColumns_line3_S13[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_timesTHREE_U7 ( .A0_t (port_out[6]), .B0_t (port_out[5]), .Z0_t (MixColumns_line3_S13[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_timesTHREE_U6 ( .A0_t (port_out[5]), .B0_t (port_out[4]), .Z0_t (MixColumns_line3_S13[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_timesTHREE_U5 ( .A0_t (port_out[4]), .B0_t (MixColumns_line3_timesTHREE_input2_4_), .Z0_t (MixColumns_line3_S13[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_timesTHREE_U4 ( .A0_t (port_out[3]), .B0_t (MixColumns_line3_timesTHREE_input2_3_), .Z0_t (MixColumns_line3_S13[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_timesTHREE_U3 ( .A0_t (port_out[2]), .B0_t (port_out[1]), .Z0_t (MixColumns_line3_S13[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_timesTHREE_U2 ( .A0_t (port_out[1]), .B0_t (MixColumns_line3_timesTHREE_input2_1_), .Z0_t (MixColumns_line3_S13[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_timesTHREE_U1 ( .A0_t (port_out[0]), .B0_t (port_out[7]), .Z0_t (MixColumns_line3_S13[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_timesTHREE_timesTWO_U3 ( .A0_t (port_out[7]), .B0_t (port_out[3]), .Z0_t (MixColumns_line3_timesTHREE_input2_4_) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_timesTHREE_timesTWO_U2 ( .A0_t (port_out[7]), .B0_t (port_out[2]), .Z0_t (MixColumns_line3_timesTHREE_input2_3_) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_timesTHREE_timesTWO_U1 ( .A0_t (port_out[7]), .B0_t (port_out[0]), .Z0_t (MixColumns_line3_timesTHREE_input2_1_) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U53 ( .A0_t (calcRCon_s_current_state_7_), .B0_t (enRCon), .Z0_t (roundConstant[7]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U52 ( .A0_t (calcRCon_s_current_state_6_), .B0_t (enRCon), .Z0_t (roundConstant[6]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U51 ( .A0_t (calcRCon_s_current_state_5_), .B0_t (enRCon), .Z0_t (roundConstant[5]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U50 ( .A0_t (calcRCon_s_current_state_4_), .B0_t (enRCon), .Z0_t (roundConstant[4]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U49 ( .A0_t (calcRCon_s_current_state_3_), .B0_t (enRCon), .Z0_t (roundConstant[3]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U48 ( .A0_t (calcRCon_s_current_state_2_), .B0_t (enRCon), .Z0_t (roundConstant[2]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U47 ( .A0_t (calcRCon_s_current_state_1_), .B0_t (enRCon), .Z0_t (roundConstant[1]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U46 ( .A0_t (calcRCon_s_current_state_0_), .B0_t (enRCon), .Z0_t (roundConstant[0]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) calcRCon_U44 ( .A0_t (calcRCon_n42), .B0_t (calcRCon_n41), .Z0_t (notFirst) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U43 ( .A0_t (calcRCon_n40), .B0_t (calcRCon_n39), .Z0_t (calcRCon_n41) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) calcRCon_U42 ( .A0_t (calcRCon_s_current_state_6_), .B0_t (calcRCon_s_current_state_5_), .Z0_t (calcRCon_n39) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) calcRCon_U41 ( .A0_t (calcRCon_s_current_state_3_), .B0_t (calcRCon_s_current_state_7_), .Z0_t (calcRCon_n40) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U40 ( .A0_t (calcRCon_n38), .B0_t (calcRCon_n37), .Z0_t (calcRCon_n42) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) calcRCon_U39 ( .A0_t (calcRCon_s_current_state_2_), .B0_t (calcRCon_s_current_state_0_), .Z0_t (calcRCon_n37) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) calcRCon_U38 ( .A0_t (calcRCon_s_current_state_1_), .B0_t (calcRCon_s_current_state_4_), .Z0_t (calcRCon_n38) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1), .NL(1'b1)) calcRCon_U37 ( .A0_t (calcRCon_n36), .B0_t (calcRCon_n35), .Z0_t (calcRCon_s_current_state_0_) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) calcRCon_U36 ( .A0_t (calcRCon_n34), .B0_t (calcRCon_s_current_state_0_), .Z0_t (calcRCon_n35) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U35 ( .A0_t (start), .B0_t (calcRCon_n33), .Z0_t (calcRCon_n36) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U34 ( .A0_t (calcRCon_n34), .B0_t (calcRCon_s_current_state_7_), .Z0_t (calcRCon_n33) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1), .NL(1'b1)) calcRCon_U33 ( .A0_t (calcRCon_n32), .B0_t (calcRCon_n31), .Z0_t (calcRCon_s_current_state_1_) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) calcRCon_U32 ( .A0_t (calcRCon_n34), .B0_t (calcRCon_s_current_state_1_), .Z0_t (calcRCon_n31) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) calcRCon_U31 ( .A0_t (calcRCon_n30), .B0_t (calcRCon_n29), .Z0_t (calcRCon_n32) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) calcRCon_U30 ( .A0_t (calcRCon_s_current_state_0_), .B0_t (calcRCon_s_current_state_7_), .Z0_t (calcRCon_n30) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b1), .NL(1'b1)) calcRCon_U29 ( .A0_t (start), .B0_t (calcRCon_n28), .Z0_t (calcRCon_s_current_state_2_) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U28 ( .A0_t (calcRCon_n27), .B0_t (calcRCon_n26), .Z0_t (calcRCon_n28) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U27 ( .A0_t (ctrl_n4), .B0_t (calcRCon_s_current_state_2_), .Z0_t (calcRCon_n26) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U26 ( .A0_t (calcRCon_n34), .B0_t (calcRCon_s_current_state_1_), .Z0_t (calcRCon_n27) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1), .NL(1'b1)) calcRCon_U25 ( .A0_t (calcRCon_n25), .B0_t (calcRCon_n24), .Z0_t (calcRCon_s_current_state_3_) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) calcRCon_U24 ( .A0_t (calcRCon_n34), .B0_t (calcRCon_s_current_state_3_), .Z0_t (calcRCon_n24) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U23 ( .A0_t (calcRCon_n23), .B0_t (start), .Z0_t (calcRCon_n25) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U22 ( .A0_t (calcRCon_n34), .B0_t (calcRCon_n22), .Z0_t (calcRCon_n23) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) calcRCon_U21 ( .A0_t (calcRCon_s_current_state_2_), .B0_t (calcRCon_s_current_state_7_), .Z0_t (calcRCon_n22) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1), .NL(1'b1)) calcRCon_U20 ( .A0_t (calcRCon_n21), .B0_t (calcRCon_n20), .Z0_t (calcRCon_s_current_state_4_) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) calcRCon_U19 ( .A0_t (calcRCon_n34), .B0_t (calcRCon_s_current_state_4_), .Z0_t (calcRCon_n20) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) calcRCon_U18 ( .A0_t (calcRCon_n19), .B0_t (calcRCon_n29), .Z0_t (calcRCon_n21) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) calcRCon_U17 ( .A0_t (calcRCon_s_current_state_3_), .B0_t (calcRCon_s_current_state_7_), .Z0_t (calcRCon_n19) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1), .NL(1'b1)) calcRCon_U16 ( .A0_t (calcRCon_n18), .B0_t (calcRCon_n17), .Z0_t (calcRCon_s_current_state_5_) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) calcRCon_U15 ( .A0_t (calcRCon_s_current_state_5_), .B0_t (calcRCon_n34), .Z0_t (calcRCon_n17) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) calcRCon_U14 ( .A0_t (calcRCon_s_current_state_4_), .B0_t (calcRCon_n29), .Z0_t (calcRCon_n18) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1), .NL(1'b1)) calcRCon_U13 ( .A0_t (calcRCon_n16), .B0_t (calcRCon_n15), .Z0_t (calcRCon_s_current_state_6_) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) calcRCon_U12 ( .A0_t (calcRCon_s_current_state_6_), .B0_t (calcRCon_n34), .Z0_t (calcRCon_n15) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) calcRCon_U11 ( .A0_t (calcRCon_s_current_state_5_), .B0_t (calcRCon_n29), .Z0_t (calcRCon_n16) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U10 ( .A0_t (calcRCon_n34), .B0_t (start), .Z0_t (calcRCon_n29) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b1), .NL(1'b1)) calcRCon_U9 ( .A0_t (start), .B0_t (calcRCon_n14), .Z0_t (calcRCon_s_current_state_7_) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U8 ( .A0_t (calcRCon_n13), .B0_t (calcRCon_n9), .Z0_t (calcRCon_n14) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U7 ( .A0_t (ctrl_n4), .B0_t (calcRCon_s_current_state_7_), .Z0_t (calcRCon_n9) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U6 ( .A0_t (calcRCon_n34), .B0_t (calcRCon_s_current_state_6_), .Z0_t (calcRCon_n13) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) calcRCon_U5 ( .A0_t (calcRCon_s_current_state_5_), .B0_t (calcRCon_s_current_state_4_), .Z0_t (calcRCon_n7) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) calcRCon_U4 ( .A0_t (calcRCon_s_current_state_1_), .B0_t (calcRCon_s_current_state_2_), .Z0_t (calcRCon_n8) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U2 ( .A0_t (ctrl_n4), .B0_t (start), .Z0_t (calcRCon_n34) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U1 ( .A0_t (calcRCon_n8), .B0_t (calcRCon_n7), .Z0_t (intFinal) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_0_XOR1_U1 ( .A0_t (StateOutXORroundKey[0]), .B0_t (keySBIn[0]), .Z0_t (MUX_SboxIn_mux_inst_0_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_0_AND1_U1 ( .A0_t (selMC), .B0_t (MUX_SboxIn_mux_inst_0_X), .Z0_t (MUX_SboxIn_mux_inst_0_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_0_XOR2_U1 ( .A0_t (MUX_SboxIn_mux_inst_0_Y), .B0_t (StateOutXORroundKey[0]), .Z0_t (SboxIn[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_1_XOR1_U1 ( .A0_t (StateOutXORroundKey[1]), .B0_t (keySBIn[1]), .Z0_t (MUX_SboxIn_mux_inst_1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_1_AND1_U1 ( .A0_t (selMC), .B0_t (MUX_SboxIn_mux_inst_1_X), .Z0_t (MUX_SboxIn_mux_inst_1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_1_XOR2_U1 ( .A0_t (MUX_SboxIn_mux_inst_1_Y), .B0_t (StateOutXORroundKey[1]), .Z0_t (SboxIn[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_2_XOR1_U1 ( .A0_t (StateOutXORroundKey[2]), .B0_t (keySBIn[2]), .Z0_t (MUX_SboxIn_mux_inst_2_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_2_AND1_U1 ( .A0_t (selMC), .B0_t (MUX_SboxIn_mux_inst_2_X), .Z0_t (MUX_SboxIn_mux_inst_2_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_2_XOR2_U1 ( .A0_t (MUX_SboxIn_mux_inst_2_Y), .B0_t (StateOutXORroundKey[2]), .Z0_t (SboxIn[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_3_XOR1_U1 ( .A0_t (StateOutXORroundKey[3]), .B0_t (keySBIn[3]), .Z0_t (MUX_SboxIn_mux_inst_3_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_3_AND1_U1 ( .A0_t (selMC), .B0_t (MUX_SboxIn_mux_inst_3_X), .Z0_t (MUX_SboxIn_mux_inst_3_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_3_XOR2_U1 ( .A0_t (MUX_SboxIn_mux_inst_3_Y), .B0_t (StateOutXORroundKey[3]), .Z0_t (SboxIn[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_4_XOR1_U1 ( .A0_t (StateOutXORroundKey[4]), .B0_t (keySBIn[4]), .Z0_t (MUX_SboxIn_mux_inst_4_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_4_AND1_U1 ( .A0_t (selMC), .B0_t (MUX_SboxIn_mux_inst_4_X), .Z0_t (MUX_SboxIn_mux_inst_4_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_4_XOR2_U1 ( .A0_t (MUX_SboxIn_mux_inst_4_Y), .B0_t (StateOutXORroundKey[4]), .Z0_t (SboxIn[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_5_XOR1_U1 ( .A0_t (StateOutXORroundKey[5]), .B0_t (keySBIn[5]), .Z0_t (MUX_SboxIn_mux_inst_5_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_5_AND1_U1 ( .A0_t (selMC), .B0_t (MUX_SboxIn_mux_inst_5_X), .Z0_t (MUX_SboxIn_mux_inst_5_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_5_XOR2_U1 ( .A0_t (MUX_SboxIn_mux_inst_5_Y), .B0_t (StateOutXORroundKey[5]), .Z0_t (SboxIn[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_6_XOR1_U1 ( .A0_t (StateOutXORroundKey[6]), .B0_t (keySBIn[6]), .Z0_t (MUX_SboxIn_mux_inst_6_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_6_AND1_U1 ( .A0_t (selMC), .B0_t (MUX_SboxIn_mux_inst_6_X), .Z0_t (MUX_SboxIn_mux_inst_6_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_6_XOR2_U1 ( .A0_t (MUX_SboxIn_mux_inst_6_Y), .B0_t (StateOutXORroundKey[6]), .Z0_t (SboxIn[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_7_XOR1_U1 ( .A0_t (StateOutXORroundKey[7]), .B0_t (keySBIn[7]), .Z0_t (MUX_SboxIn_mux_inst_7_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_7_AND1_U1 ( .A0_t (selMC), .B0_t (MUX_SboxIn_mux_inst_7_X), .Z0_t (MUX_SboxIn_mux_inst_7_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_7_XOR2_U1 ( .A0_t (MUX_SboxIn_mux_inst_7_Y), .B0_t (StateOutXORroundKey[7]), .Z0_t (SboxIn[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T1_U1 ( .A0_t (SboxIn[7]), .B0_t (SboxIn[4]), .Z0_t (Inst_bSbox_T1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T2_U1 ( .A0_t (SboxIn[7]), .B0_t (SboxIn[2]), .Z0_t (Inst_bSbox_T2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T3_U1 ( .A0_t (SboxIn[7]), .B0_t (SboxIn[1]), .Z0_t (Inst_bSbox_T3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T4_U1 ( .A0_t (SboxIn[4]), .B0_t (SboxIn[2]), .Z0_t (Inst_bSbox_T4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T5_U1 ( .A0_t (SboxIn[3]), .B0_t (SboxIn[1]), .Z0_t (Inst_bSbox_T5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T6_U1 ( .A0_t (Inst_bSbox_T1), .B0_t (Inst_bSbox_T5), .Z0_t (Inst_bSbox_T6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T7_U1 ( .A0_t (SboxIn[6]), .B0_t (SboxIn[5]), .Z0_t (Inst_bSbox_T7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T8_U1 ( .A0_t (SboxIn[0]), .B0_t (Inst_bSbox_T6), .Z0_t (Inst_bSbox_T8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T9_U1 ( .A0_t (SboxIn[0]), .B0_t (Inst_bSbox_T7), .Z0_t (Inst_bSbox_T9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T10_U1 ( .A0_t (Inst_bSbox_T6), .B0_t (Inst_bSbox_T7), .Z0_t (Inst_bSbox_T10) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T11_U1 ( .A0_t (SboxIn[6]), .B0_t (SboxIn[2]), .Z0_t (Inst_bSbox_T11) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T12_U1 ( .A0_t (SboxIn[5]), .B0_t (SboxIn[2]), .Z0_t (Inst_bSbox_T12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T13_U1 ( .A0_t (Inst_bSbox_T3), .B0_t (Inst_bSbox_T4), .Z0_t (Inst_bSbox_T13) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T14_U1 ( .A0_t (Inst_bSbox_T6), .B0_t (Inst_bSbox_T11), .Z0_t (Inst_bSbox_T14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T15_U1 ( .A0_t (Inst_bSbox_T5), .B0_t (Inst_bSbox_T11), .Z0_t (Inst_bSbox_T15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T16_U1 ( .A0_t (Inst_bSbox_T5), .B0_t (Inst_bSbox_T12), .Z0_t (Inst_bSbox_T16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T17_U1 ( .A0_t (Inst_bSbox_T9), .B0_t (Inst_bSbox_T16), .Z0_t (Inst_bSbox_T17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T18_U1 ( .A0_t (SboxIn[4]), .B0_t (SboxIn[0]), .Z0_t (Inst_bSbox_T18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T19_U1 ( .A0_t (Inst_bSbox_T7), .B0_t (Inst_bSbox_T18), .Z0_t (Inst_bSbox_T19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T20_U1 ( .A0_t (Inst_bSbox_T1), .B0_t (Inst_bSbox_T19), .Z0_t (Inst_bSbox_T20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T21_U1 ( .A0_t (SboxIn[1]), .B0_t (SboxIn[0]), .Z0_t (Inst_bSbox_T21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T22_U1 ( .A0_t (Inst_bSbox_T7), .B0_t (Inst_bSbox_T21), .Z0_t (Inst_bSbox_T22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T23_U1 ( .A0_t (Inst_bSbox_T2), .B0_t (Inst_bSbox_T22), .Z0_t (Inst_bSbox_T23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T24_U1 ( .A0_t (Inst_bSbox_T2), .B0_t (Inst_bSbox_T10), .Z0_t (Inst_bSbox_T24) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T25_U1 ( .A0_t (Inst_bSbox_T20), .B0_t (Inst_bSbox_T17), .Z0_t (Inst_bSbox_T25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T26_U1 ( .A0_t (Inst_bSbox_T3), .B0_t (Inst_bSbox_T16), .Z0_t (Inst_bSbox_T26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T27_U1 ( .A0_t (Inst_bSbox_T1), .B0_t (Inst_bSbox_T12), .Z0_t (Inst_bSbox_T27) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M1_U1 ( .A0_t (Inst_bSbox_T13), .B0_t (Inst_bSbox_T6), .Z0_t (Inst_bSbox_M1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M2_U1 ( .A0_t (Inst_bSbox_T23), .B0_t (Inst_bSbox_T8), .Z0_t (Inst_bSbox_M2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M3_U1 ( .A0_t (Inst_bSbox_T14), .B0_t (Inst_bSbox_M1), .Z0_t (Inst_bSbox_M3) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M4_U1 ( .A0_t (Inst_bSbox_T19), .B0_t (SboxIn[0]), .Z0_t (Inst_bSbox_M4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M5_U1 ( .A0_t (Inst_bSbox_M4), .B0_t (Inst_bSbox_M1), .Z0_t (Inst_bSbox_M5) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M6_U1 ( .A0_t (Inst_bSbox_T3), .B0_t (Inst_bSbox_T16), .Z0_t (Inst_bSbox_M6) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M7_U1 ( .A0_t (Inst_bSbox_T22), .B0_t (Inst_bSbox_T9), .Z0_t (Inst_bSbox_M7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M8_U1 ( .A0_t (Inst_bSbox_T26), .B0_t (Inst_bSbox_M6), .Z0_t (Inst_bSbox_M8) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M9_U1 ( .A0_t (Inst_bSbox_T20), .B0_t (Inst_bSbox_T17), .Z0_t (Inst_bSbox_M9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M10_U1 ( .A0_t (Inst_bSbox_M9), .B0_t (Inst_bSbox_M6), .Z0_t (Inst_bSbox_M10) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M11_U1 ( .A0_t (Inst_bSbox_T1), .B0_t (Inst_bSbox_T15), .Z0_t (Inst_bSbox_M11) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M12_U1 ( .A0_t (Inst_bSbox_T4), .B0_t (Inst_bSbox_T27), .Z0_t (Inst_bSbox_M12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M13_U1 ( .A0_t (Inst_bSbox_M12), .B0_t (Inst_bSbox_M11), .Z0_t (Inst_bSbox_M13) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M14_U1 ( .A0_t (Inst_bSbox_T2), .B0_t (Inst_bSbox_T10), .Z0_t (Inst_bSbox_M14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M15_U1 ( .A0_t (Inst_bSbox_M14), .B0_t (Inst_bSbox_M11), .Z0_t (Inst_bSbox_M15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M16_U1 ( .A0_t (Inst_bSbox_M3), .B0_t (Inst_bSbox_M2), .Z0_t (Inst_bSbox_M16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M17_U1 ( .A0_t (Inst_bSbox_M5), .B0_t (Inst_bSbox_T24), .Z0_t (Inst_bSbox_M17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M18_U1 ( .A0_t (Inst_bSbox_M8), .B0_t (Inst_bSbox_M7), .Z0_t (Inst_bSbox_M18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M19_U1 ( .A0_t (Inst_bSbox_M10), .B0_t (Inst_bSbox_M15), .Z0_t (Inst_bSbox_M19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M20_U1 ( .A0_t (Inst_bSbox_M16), .B0_t (Inst_bSbox_M13), .Z0_t (Inst_bSbox_M20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M21_U1 ( .A0_t (Inst_bSbox_M17), .B0_t (Inst_bSbox_M15), .Z0_t (Inst_bSbox_M21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M22_U1 ( .A0_t (Inst_bSbox_M18), .B0_t (Inst_bSbox_M13), .Z0_t (Inst_bSbox_M22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M23_U1 ( .A0_t (Inst_bSbox_M19), .B0_t (Inst_bSbox_T25), .Z0_t (Inst_bSbox_M23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M24_U1 ( .A0_t (Inst_bSbox_M22), .B0_t (Inst_bSbox_M23), .Z0_t (Inst_bSbox_M24) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M25_U1 ( .A0_t (Inst_bSbox_M22), .B0_t (Inst_bSbox_M20), .Z0_t (Inst_bSbox_M25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M26_U1 ( .A0_t (Inst_bSbox_M21), .B0_t (Inst_bSbox_M25), .Z0_t (Inst_bSbox_M26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M27_U1 ( .A0_t (Inst_bSbox_M20), .B0_t (Inst_bSbox_M21), .Z0_t (Inst_bSbox_M27) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M28_U1 ( .A0_t (Inst_bSbox_M23), .B0_t (Inst_bSbox_M25), .Z0_t (Inst_bSbox_M28) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M29_U1 ( .A0_t (Inst_bSbox_M28), .B0_t (Inst_bSbox_M27), .Z0_t (Inst_bSbox_M29) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M30_U1 ( .A0_t (Inst_bSbox_M26), .B0_t (Inst_bSbox_M24), .Z0_t (Inst_bSbox_M30) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M31_U1 ( .A0_t (Inst_bSbox_M20), .B0_t (Inst_bSbox_M23), .Z0_t (Inst_bSbox_M31) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M32_U1 ( .A0_t (Inst_bSbox_M27), .B0_t (Inst_bSbox_M31), .Z0_t (Inst_bSbox_M32) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M33_U1 ( .A0_t (Inst_bSbox_M27), .B0_t (Inst_bSbox_M25), .Z0_t (Inst_bSbox_M33) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M34_U1 ( .A0_t (Inst_bSbox_M21), .B0_t (Inst_bSbox_M22), .Z0_t (Inst_bSbox_M34) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M35_U1 ( .A0_t (Inst_bSbox_M24), .B0_t (Inst_bSbox_M34), .Z0_t (Inst_bSbox_M35) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M36_U1 ( .A0_t (Inst_bSbox_M24), .B0_t (Inst_bSbox_M25), .Z0_t (Inst_bSbox_M36) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M37_U1 ( .A0_t (Inst_bSbox_M21), .B0_t (Inst_bSbox_M29), .Z0_t (Inst_bSbox_M37) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M38_U1 ( .A0_t (Inst_bSbox_M32), .B0_t (Inst_bSbox_M33), .Z0_t (Inst_bSbox_M38) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M39_U1 ( .A0_t (Inst_bSbox_M23), .B0_t (Inst_bSbox_M30), .Z0_t (Inst_bSbox_M39) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M40_U1 ( .A0_t (Inst_bSbox_M35), .B0_t (Inst_bSbox_M36), .Z0_t (Inst_bSbox_M40) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M41_U1 ( .A0_t (Inst_bSbox_M38), .B0_t (Inst_bSbox_M40), .Z0_t (Inst_bSbox_M41) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M42_U1 ( .A0_t (Inst_bSbox_M37), .B0_t (Inst_bSbox_M39), .Z0_t (Inst_bSbox_M42) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M43_U1 ( .A0_t (Inst_bSbox_M37), .B0_t (Inst_bSbox_M38), .Z0_t (Inst_bSbox_M43) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M44_U1 ( .A0_t (Inst_bSbox_M39), .B0_t (Inst_bSbox_M40), .Z0_t (Inst_bSbox_M44) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M45_U1 ( .A0_t (Inst_bSbox_M42), .B0_t (Inst_bSbox_M41), .Z0_t (Inst_bSbox_M45) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M46_U1 ( .A0_t (Inst_bSbox_M44), .B0_t (Inst_bSbox_T6), .Z0_t (Inst_bSbox_M46) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M47_U1 ( .A0_t (Inst_bSbox_M40), .B0_t (Inst_bSbox_T8), .Z0_t (Inst_bSbox_M47) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M48_U1 ( .A0_t (Inst_bSbox_M39), .B0_t (SboxIn[0]), .Z0_t (Inst_bSbox_M48) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M49_U1 ( .A0_t (Inst_bSbox_M43), .B0_t (Inst_bSbox_T16), .Z0_t (Inst_bSbox_M49) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M50_U1 ( .A0_t (Inst_bSbox_M38), .B0_t (Inst_bSbox_T9), .Z0_t (Inst_bSbox_M50) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M51_U1 ( .A0_t (Inst_bSbox_M37), .B0_t (Inst_bSbox_T17), .Z0_t (Inst_bSbox_M51) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M52_U1 ( .A0_t (Inst_bSbox_M42), .B0_t (Inst_bSbox_T15), .Z0_t (Inst_bSbox_M52) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M53_U1 ( .A0_t (Inst_bSbox_M45), .B0_t (Inst_bSbox_T27), .Z0_t (Inst_bSbox_M53) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M54_U1 ( .A0_t (Inst_bSbox_M41), .B0_t (Inst_bSbox_T10), .Z0_t (Inst_bSbox_M54) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M55_U1 ( .A0_t (Inst_bSbox_M44), .B0_t (Inst_bSbox_T13), .Z0_t (Inst_bSbox_M55) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M56_U1 ( .A0_t (Inst_bSbox_M40), .B0_t (Inst_bSbox_T23), .Z0_t (Inst_bSbox_M56) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M57_U1 ( .A0_t (Inst_bSbox_M39), .B0_t (Inst_bSbox_T19), .Z0_t (Inst_bSbox_M57) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M58_U1 ( .A0_t (Inst_bSbox_M43), .B0_t (Inst_bSbox_T3), .Z0_t (Inst_bSbox_M58) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M59_U1 ( .A0_t (Inst_bSbox_M38), .B0_t (Inst_bSbox_T22), .Z0_t (Inst_bSbox_M59) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M60_U1 ( .A0_t (Inst_bSbox_M37), .B0_t (Inst_bSbox_T20), .Z0_t (Inst_bSbox_M60) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M61_U1 ( .A0_t (Inst_bSbox_M42), .B0_t (Inst_bSbox_T1), .Z0_t (Inst_bSbox_M61) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M62_U1 ( .A0_t (Inst_bSbox_M45), .B0_t (Inst_bSbox_T4), .Z0_t (Inst_bSbox_M62) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M63_U1 ( .A0_t (Inst_bSbox_M41), .B0_t (Inst_bSbox_T2), .Z0_t (Inst_bSbox_M63) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L0_U1 ( .A0_t (Inst_bSbox_M61), .B0_t (Inst_bSbox_M62), .Z0_t (Inst_bSbox_L0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L1_U1 ( .A0_t (Inst_bSbox_M50), .B0_t (Inst_bSbox_M56), .Z0_t (Inst_bSbox_L1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L2_U1 ( .A0_t (Inst_bSbox_M46), .B0_t (Inst_bSbox_M48), .Z0_t (Inst_bSbox_L2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L3_U1 ( .A0_t (Inst_bSbox_M47), .B0_t (Inst_bSbox_M55), .Z0_t (Inst_bSbox_L3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L4_U1 ( .A0_t (Inst_bSbox_M54), .B0_t (Inst_bSbox_M58), .Z0_t (Inst_bSbox_L4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L5_U1 ( .A0_t (Inst_bSbox_M49), .B0_t (Inst_bSbox_M61), .Z0_t (Inst_bSbox_L5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L6_U1 ( .A0_t (Inst_bSbox_M62), .B0_t (Inst_bSbox_L5), .Z0_t (Inst_bSbox_L6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L7_U1 ( .A0_t (Inst_bSbox_M46), .B0_t (Inst_bSbox_L3), .Z0_t (Inst_bSbox_L7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L8_U1 ( .A0_t (Inst_bSbox_M51), .B0_t (Inst_bSbox_M59), .Z0_t (Inst_bSbox_L8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L9_U1 ( .A0_t (Inst_bSbox_M52), .B0_t (Inst_bSbox_M53), .Z0_t (Inst_bSbox_L9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L10_U1 ( .A0_t (Inst_bSbox_M53), .B0_t (Inst_bSbox_L4), .Z0_t (Inst_bSbox_L10) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L11_U1 ( .A0_t (Inst_bSbox_M60), .B0_t (Inst_bSbox_L2), .Z0_t (Inst_bSbox_L11) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L12_U1 ( .A0_t (Inst_bSbox_M48), .B0_t (Inst_bSbox_M51), .Z0_t (Inst_bSbox_L12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L13_U1 ( .A0_t (Inst_bSbox_M50), .B0_t (Inst_bSbox_L0), .Z0_t (Inst_bSbox_L13) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L14_U1 ( .A0_t (Inst_bSbox_M52), .B0_t (Inst_bSbox_M61), .Z0_t (Inst_bSbox_L14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L15_U1 ( .A0_t (Inst_bSbox_M55), .B0_t (Inst_bSbox_L1), .Z0_t (Inst_bSbox_L15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L16_U1 ( .A0_t (Inst_bSbox_M56), .B0_t (Inst_bSbox_L0), .Z0_t (Inst_bSbox_L16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L17_U1 ( .A0_t (Inst_bSbox_M57), .B0_t (Inst_bSbox_L1), .Z0_t (Inst_bSbox_L17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L18_U1 ( .A0_t (Inst_bSbox_M58), .B0_t (Inst_bSbox_L8), .Z0_t (Inst_bSbox_L18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L19_U1 ( .A0_t (Inst_bSbox_M63), .B0_t (Inst_bSbox_L4), .Z0_t (Inst_bSbox_L19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L20_U1 ( .A0_t (Inst_bSbox_L0), .B0_t (Inst_bSbox_L1), .Z0_t (Inst_bSbox_L20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L21_U1 ( .A0_t (Inst_bSbox_L1), .B0_t (Inst_bSbox_L7), .Z0_t (Inst_bSbox_L21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L22_U1 ( .A0_t (Inst_bSbox_L3), .B0_t (Inst_bSbox_L12), .Z0_t (Inst_bSbox_L22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L23_U1 ( .A0_t (Inst_bSbox_L18), .B0_t (Inst_bSbox_L2), .Z0_t (Inst_bSbox_L23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L24_U1 ( .A0_t (Inst_bSbox_L15), .B0_t (Inst_bSbox_L9), .Z0_t (Inst_bSbox_L24) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L25_U1 ( .A0_t (Inst_bSbox_L6), .B0_t (Inst_bSbox_L10), .Z0_t (Inst_bSbox_L25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L26_U1 ( .A0_t (Inst_bSbox_L7), .B0_t (Inst_bSbox_L9), .Z0_t (Inst_bSbox_L26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L27_U1 ( .A0_t (Inst_bSbox_L8), .B0_t (Inst_bSbox_L10), .Z0_t (Inst_bSbox_L27) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L28_U1 ( .A0_t (Inst_bSbox_L11), .B0_t (Inst_bSbox_L14), .Z0_t (Inst_bSbox_L28) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L29_U1 ( .A0_t (Inst_bSbox_L11), .B0_t (Inst_bSbox_L17), .Z0_t (Inst_bSbox_L29) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_S0_U1 ( .A0_t (Inst_bSbox_L6), .B0_t (Inst_bSbox_L24), .Z0_t (SboxOut[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Inst_bSbox_XOR_S1_U1 ( .A0_t (Inst_bSbox_L16), .B0_t (Inst_bSbox_L26), .Z0_t (SboxOut[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Inst_bSbox_XOR_S2_U1 ( .A0_t (Inst_bSbox_L19), .B0_t (Inst_bSbox_L28), .Z0_t (SboxOut[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_S3_U1 ( .A0_t (Inst_bSbox_L6), .B0_t (Inst_bSbox_L21), .Z0_t (SboxOut[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_S4_U1 ( .A0_t (Inst_bSbox_L20), .B0_t (Inst_bSbox_L22), .Z0_t (SboxOut[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_S5_U1 ( .A0_t (Inst_bSbox_L25), .B0_t (Inst_bSbox_L29), .Z0_t (SboxOut[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Inst_bSbox_XOR_S6_U1 ( .A0_t (Inst_bSbox_L13), .B0_t (Inst_bSbox_L27), .Z0_t (SboxOut[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Inst_bSbox_XOR_S7_U1 ( .A0_t (Inst_bSbox_L6), .B0_t (Inst_bSbox_L23), .Z0_t (SboxOut[0]) ) ;

    /* register cells */
endmodule
