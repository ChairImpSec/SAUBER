
module AES ( clk, start, port_in, port_out, done );
  input [7:0] port_in;
  output [7:0] port_out;
  input clk, start;
  output done;
  wire   selMC, selSR, selXOR, enRCon, intFinal, enKS, intselXOR, notFirst, n2,
         ctrl_n24, ctrl_n19, ctrl_n18, ctrl_n17, ctrl_n14, ctrl_n13, ctrl_n12,
         ctrl_n11, ctrl_n10, ctrl_n9, ctrl_n7, ctrl_n6, ctrl_n4,
         ctrl_finalStep, ctrl_n2, ctrl_n15, ctrl_n20, ctrl_n16, ctrl_n5,
         ctrl_n21, ctrl_seq4Out_1_, ctrl_seq4In_1_, ctrl_nRstSeq4, ctrl_n22,
         ctrl_seq6Out_4_, ctrl_seq6In_1_, ctrl_seq6In_2_, ctrl_seq6In_3_,
         ctrl_seq6In_4_, ctrl_n23, ctrl_seq6_SFF_0_n2, ctrl_seq6_SFF_0_n1,
         ctrl_seq6_SFF_0_n3, ctrl_seq6_SFF_0_n5, ctrl_seq6_SFF_0_QD,
         ctrl_seq6_SFF_0_MUXInst_Y, ctrl_seq6_SFF_0_MUXInst_X,
         ctrl_seq6_SFF_1_n2, ctrl_seq6_SFF_1_n1, ctrl_seq6_SFF_1_n10,
         ctrl_seq6_SFF_1_n5, ctrl_seq6_SFF_1_QD, ctrl_seq6_SFF_1_MUXInst_Y,
         ctrl_seq6_SFF_1_MUXInst_X, ctrl_seq6_SFF_2_n2, ctrl_seq6_SFF_2_n1,
         ctrl_seq6_SFF_2_n10, ctrl_seq6_SFF_2_n5, ctrl_seq6_SFF_2_QD,
         ctrl_seq6_SFF_2_MUXInst_Y, ctrl_seq6_SFF_2_MUXInst_X,
         ctrl_seq6_SFF_3_n2, ctrl_seq6_SFF_3_n1, ctrl_seq6_SFF_3_n10,
         ctrl_seq6_SFF_3_n5, ctrl_seq6_SFF_3_QD, ctrl_seq6_SFF_3_MUXInst_Y,
         ctrl_seq6_SFF_3_MUXInst_X, ctrl_seq6_SFF_4_n2, ctrl_seq6_SFF_4_n1,
         ctrl_seq6_SFF_4_n10, ctrl_seq6_SFF_4_n5, ctrl_seq6_SFF_4_QD,
         ctrl_seq6_SFF_4_MUXInst_Y, ctrl_seq6_SFF_4_MUXInst_X,
         ctrl_seq4_SFF_0_n2, ctrl_seq4_SFF_0_n1, ctrl_seq4_SFF_0_n10,
         ctrl_seq4_SFF_0_n5, ctrl_seq4_SFF_0_QD, ctrl_seq4_SFF_0_MUXInst_Y,
         ctrl_seq4_SFF_0_MUXInst_X, ctrl_seq4_SFF_1_n2, ctrl_seq4_SFF_1_n1,
         ctrl_seq4_SFF_1_n10, ctrl_seq4_SFF_1_n5, ctrl_seq4_SFF_1_QD,
         ctrl_seq4_SFF_1_MUXInst_Y, ctrl_seq4_SFF_1_MUXInst_X,
         MUX_StateIn_mux_inst_0_Y, MUX_StateIn_mux_inst_0_X,
         MUX_StateIn_mux_inst_1_Y, MUX_StateIn_mux_inst_1_X,
         MUX_StateIn_mux_inst_2_Y, MUX_StateIn_mux_inst_2_X,
         MUX_StateIn_mux_inst_3_Y, MUX_StateIn_mux_inst_3_X,
         MUX_StateIn_mux_inst_4_Y, MUX_StateIn_mux_inst_4_X,
         MUX_StateIn_mux_inst_5_Y, MUX_StateIn_mux_inst_5_X,
         MUX_StateIn_mux_inst_6_Y, MUX_StateIn_mux_inst_6_X,
         MUX_StateIn_mux_inst_7_Y, MUX_StateIn_mux_inst_7_X, stateArray_n8,
         stateArray_n7, stateArray_n6, stateArray_nReset_selMC,
         stateArray_S00reg_gff_1_SFF_0_QD,
         stateArray_S00reg_gff_1_SFF_0_MUXInst_Y,
         stateArray_S00reg_gff_1_SFF_0_MUXInst_X,
         stateArray_S00reg_gff_1_SFF_0_Q_reg_QN,
         stateArray_S00reg_gff_1_SFF_1_QD,
         stateArray_S00reg_gff_1_SFF_1_MUXInst_Y,
         stateArray_S00reg_gff_1_SFF_1_MUXInst_X,
         stateArray_S00reg_gff_1_SFF_1_Q_reg_QN,
         stateArray_S00reg_gff_1_SFF_2_QD,
         stateArray_S00reg_gff_1_SFF_2_MUXInst_Y,
         stateArray_S00reg_gff_1_SFF_2_MUXInst_X,
         stateArray_S00reg_gff_1_SFF_2_Q_reg_QN,
         stateArray_S00reg_gff_1_SFF_3_QD,
         stateArray_S00reg_gff_1_SFF_3_MUXInst_Y,
         stateArray_S00reg_gff_1_SFF_3_MUXInst_X,
         stateArray_S00reg_gff_1_SFF_3_Q_reg_QN,
         stateArray_S00reg_gff_1_SFF_4_QD,
         stateArray_S00reg_gff_1_SFF_4_MUXInst_Y,
         stateArray_S00reg_gff_1_SFF_4_MUXInst_X,
         stateArray_S00reg_gff_1_SFF_4_Q_reg_QN,
         stateArray_S00reg_gff_1_SFF_5_QD,
         stateArray_S00reg_gff_1_SFF_5_MUXInst_Y,
         stateArray_S00reg_gff_1_SFF_5_MUXInst_X,
         stateArray_S00reg_gff_1_SFF_5_Q_reg_QN,
         stateArray_S00reg_gff_1_SFF_6_QD,
         stateArray_S00reg_gff_1_SFF_6_MUXInst_Y,
         stateArray_S00reg_gff_1_SFF_6_MUXInst_X,
         stateArray_S00reg_gff_1_SFF_6_Q_reg_QN,
         stateArray_S00reg_gff_1_SFF_7_QD,
         stateArray_S00reg_gff_1_SFF_7_MUXInst_Y,
         stateArray_S00reg_gff_1_SFF_7_MUXInst_X,
         stateArray_S00reg_gff_1_SFF_7_Q_reg_QN,
         stateArray_S01reg_gff_1_SFF_0_QD,
         stateArray_S01reg_gff_1_SFF_0_MUXInst_Y,
         stateArray_S01reg_gff_1_SFF_0_MUXInst_X,
         stateArray_S01reg_gff_1_SFF_0_Q_reg_QN,
         stateArray_S01reg_gff_1_SFF_1_QD,
         stateArray_S01reg_gff_1_SFF_1_MUXInst_Y,
         stateArray_S01reg_gff_1_SFF_1_MUXInst_X,
         stateArray_S01reg_gff_1_SFF_1_Q_reg_QN,
         stateArray_S01reg_gff_1_SFF_2_QD,
         stateArray_S01reg_gff_1_SFF_2_MUXInst_Y,
         stateArray_S01reg_gff_1_SFF_2_MUXInst_X,
         stateArray_S01reg_gff_1_SFF_2_Q_reg_QN,
         stateArray_S01reg_gff_1_SFF_3_QD,
         stateArray_S01reg_gff_1_SFF_3_MUXInst_Y,
         stateArray_S01reg_gff_1_SFF_3_MUXInst_X,
         stateArray_S01reg_gff_1_SFF_3_Q_reg_QN,
         stateArray_S01reg_gff_1_SFF_4_QD,
         stateArray_S01reg_gff_1_SFF_4_MUXInst_Y,
         stateArray_S01reg_gff_1_SFF_4_MUXInst_X,
         stateArray_S01reg_gff_1_SFF_4_Q_reg_QN,
         stateArray_S01reg_gff_1_SFF_5_QD,
         stateArray_S01reg_gff_1_SFF_5_MUXInst_Y,
         stateArray_S01reg_gff_1_SFF_5_MUXInst_X,
         stateArray_S01reg_gff_1_SFF_5_Q_reg_QN,
         stateArray_S01reg_gff_1_SFF_6_QD,
         stateArray_S01reg_gff_1_SFF_6_MUXInst_Y,
         stateArray_S01reg_gff_1_SFF_6_MUXInst_X,
         stateArray_S01reg_gff_1_SFF_6_Q_reg_QN,
         stateArray_S01reg_gff_1_SFF_7_QD,
         stateArray_S01reg_gff_1_SFF_7_MUXInst_Y,
         stateArray_S01reg_gff_1_SFF_7_MUXInst_X,
         stateArray_S01reg_gff_1_SFF_7_Q_reg_QN,
         stateArray_S02reg_gff_1_SFF_0_QD,
         stateArray_S02reg_gff_1_SFF_0_MUXInst_Y,
         stateArray_S02reg_gff_1_SFF_0_MUXInst_X,
         stateArray_S02reg_gff_1_SFF_0_Q_reg_QN,
         stateArray_S02reg_gff_1_SFF_1_QD,
         stateArray_S02reg_gff_1_SFF_1_MUXInst_Y,
         stateArray_S02reg_gff_1_SFF_1_MUXInst_X,
         stateArray_S02reg_gff_1_SFF_1_Q_reg_QN,
         stateArray_S02reg_gff_1_SFF_2_QD,
         stateArray_S02reg_gff_1_SFF_2_MUXInst_Y,
         stateArray_S02reg_gff_1_SFF_2_MUXInst_X,
         stateArray_S02reg_gff_1_SFF_2_Q_reg_QN,
         stateArray_S02reg_gff_1_SFF_3_QD,
         stateArray_S02reg_gff_1_SFF_3_MUXInst_Y,
         stateArray_S02reg_gff_1_SFF_3_MUXInst_X,
         stateArray_S02reg_gff_1_SFF_3_Q_reg_QN,
         stateArray_S02reg_gff_1_SFF_4_QD,
         stateArray_S02reg_gff_1_SFF_4_MUXInst_Y,
         stateArray_S02reg_gff_1_SFF_4_MUXInst_X,
         stateArray_S02reg_gff_1_SFF_4_Q_reg_QN,
         stateArray_S02reg_gff_1_SFF_5_QD,
         stateArray_S02reg_gff_1_SFF_5_MUXInst_Y,
         stateArray_S02reg_gff_1_SFF_5_MUXInst_X,
         stateArray_S02reg_gff_1_SFF_5_Q_reg_QN,
         stateArray_S02reg_gff_1_SFF_6_QD,
         stateArray_S02reg_gff_1_SFF_6_MUXInst_Y,
         stateArray_S02reg_gff_1_SFF_6_MUXInst_X,
         stateArray_S02reg_gff_1_SFF_6_Q_reg_QN,
         stateArray_S02reg_gff_1_SFF_7_QD,
         stateArray_S02reg_gff_1_SFF_7_MUXInst_Y,
         stateArray_S02reg_gff_1_SFF_7_MUXInst_X,
         stateArray_S02reg_gff_1_SFF_7_Q_reg_QN,
         stateArray_S03reg_gff_1_SFF_0_QD,
         stateArray_S03reg_gff_1_SFF_0_MUXInst_Y,
         stateArray_S03reg_gff_1_SFF_0_MUXInst_X,
         stateArray_S03reg_gff_1_SFF_0_Q_reg_QN,
         stateArray_S03reg_gff_1_SFF_1_QD,
         stateArray_S03reg_gff_1_SFF_1_MUXInst_Y,
         stateArray_S03reg_gff_1_SFF_1_MUXInst_X,
         stateArray_S03reg_gff_1_SFF_1_Q_reg_QN,
         stateArray_S03reg_gff_1_SFF_2_QD,
         stateArray_S03reg_gff_1_SFF_2_MUXInst_Y,
         stateArray_S03reg_gff_1_SFF_2_MUXInst_X,
         stateArray_S03reg_gff_1_SFF_2_Q_reg_QN,
         stateArray_S03reg_gff_1_SFF_3_QD,
         stateArray_S03reg_gff_1_SFF_3_MUXInst_Y,
         stateArray_S03reg_gff_1_SFF_3_MUXInst_X,
         stateArray_S03reg_gff_1_SFF_3_Q_reg_QN,
         stateArray_S03reg_gff_1_SFF_4_QD,
         stateArray_S03reg_gff_1_SFF_4_MUXInst_Y,
         stateArray_S03reg_gff_1_SFF_4_MUXInst_X,
         stateArray_S03reg_gff_1_SFF_4_Q_reg_QN,
         stateArray_S03reg_gff_1_SFF_5_QD,
         stateArray_S03reg_gff_1_SFF_5_MUXInst_Y,
         stateArray_S03reg_gff_1_SFF_5_MUXInst_X,
         stateArray_S03reg_gff_1_SFF_5_Q_reg_QN,
         stateArray_S03reg_gff_1_SFF_6_QD,
         stateArray_S03reg_gff_1_SFF_6_MUXInst_Y,
         stateArray_S03reg_gff_1_SFF_6_MUXInst_X,
         stateArray_S03reg_gff_1_SFF_6_Q_reg_QN,
         stateArray_S03reg_gff_1_SFF_7_QD,
         stateArray_S03reg_gff_1_SFF_7_MUXInst_Y,
         stateArray_S03reg_gff_1_SFF_7_MUXInst_X,
         stateArray_S03reg_gff_1_SFF_7_Q_reg_QN,
         stateArray_S10reg_gff_1_SFF_0_QD,
         stateArray_S10reg_gff_1_SFF_0_MUXInst_Y,
         stateArray_S10reg_gff_1_SFF_0_MUXInst_X,
         stateArray_S10reg_gff_1_SFF_0_Q_reg_QN,
         stateArray_S10reg_gff_1_SFF_1_QD,
         stateArray_S10reg_gff_1_SFF_1_MUXInst_Y,
         stateArray_S10reg_gff_1_SFF_1_MUXInst_X,
         stateArray_S10reg_gff_1_SFF_1_Q_reg_QN,
         stateArray_S10reg_gff_1_SFF_2_QD,
         stateArray_S10reg_gff_1_SFF_2_MUXInst_Y,
         stateArray_S10reg_gff_1_SFF_2_MUXInst_X,
         stateArray_S10reg_gff_1_SFF_2_Q_reg_QN,
         stateArray_S10reg_gff_1_SFF_3_QD,
         stateArray_S10reg_gff_1_SFF_3_MUXInst_Y,
         stateArray_S10reg_gff_1_SFF_3_MUXInst_X,
         stateArray_S10reg_gff_1_SFF_3_Q_reg_QN,
         stateArray_S10reg_gff_1_SFF_4_QD,
         stateArray_S10reg_gff_1_SFF_4_MUXInst_Y,
         stateArray_S10reg_gff_1_SFF_4_MUXInst_X,
         stateArray_S10reg_gff_1_SFF_4_Q_reg_QN,
         stateArray_S10reg_gff_1_SFF_5_QD,
         stateArray_S10reg_gff_1_SFF_5_MUXInst_Y,
         stateArray_S10reg_gff_1_SFF_5_MUXInst_X,
         stateArray_S10reg_gff_1_SFF_5_Q_reg_QN,
         stateArray_S10reg_gff_1_SFF_6_QD,
         stateArray_S10reg_gff_1_SFF_6_MUXInst_Y,
         stateArray_S10reg_gff_1_SFF_6_MUXInst_X,
         stateArray_S10reg_gff_1_SFF_6_Q_reg_QN,
         stateArray_S10reg_gff_1_SFF_7_QD,
         stateArray_S10reg_gff_1_SFF_7_MUXInst_Y,
         stateArray_S10reg_gff_1_SFF_7_MUXInst_X,
         stateArray_S10reg_gff_1_SFF_7_Q_reg_QN,
         stateArray_S11reg_gff_1_SFF_0_QD,
         stateArray_S11reg_gff_1_SFF_0_MUXInst_Y,
         stateArray_S11reg_gff_1_SFF_0_MUXInst_X,
         stateArray_S11reg_gff_1_SFF_0_Q_reg_QN,
         stateArray_S11reg_gff_1_SFF_1_QD,
         stateArray_S11reg_gff_1_SFF_1_MUXInst_Y,
         stateArray_S11reg_gff_1_SFF_1_MUXInst_X,
         stateArray_S11reg_gff_1_SFF_1_Q_reg_QN,
         stateArray_S11reg_gff_1_SFF_2_QD,
         stateArray_S11reg_gff_1_SFF_2_MUXInst_Y,
         stateArray_S11reg_gff_1_SFF_2_MUXInst_X,
         stateArray_S11reg_gff_1_SFF_2_Q_reg_QN,
         stateArray_S11reg_gff_1_SFF_3_QD,
         stateArray_S11reg_gff_1_SFF_3_MUXInst_Y,
         stateArray_S11reg_gff_1_SFF_3_MUXInst_X,
         stateArray_S11reg_gff_1_SFF_3_Q_reg_QN,
         stateArray_S11reg_gff_1_SFF_4_QD,
         stateArray_S11reg_gff_1_SFF_4_MUXInst_Y,
         stateArray_S11reg_gff_1_SFF_4_MUXInst_X,
         stateArray_S11reg_gff_1_SFF_4_Q_reg_QN,
         stateArray_S11reg_gff_1_SFF_5_QD,
         stateArray_S11reg_gff_1_SFF_5_MUXInst_Y,
         stateArray_S11reg_gff_1_SFF_5_MUXInst_X,
         stateArray_S11reg_gff_1_SFF_5_Q_reg_QN,
         stateArray_S11reg_gff_1_SFF_6_QD,
         stateArray_S11reg_gff_1_SFF_6_MUXInst_Y,
         stateArray_S11reg_gff_1_SFF_6_MUXInst_X,
         stateArray_S11reg_gff_1_SFF_6_Q_reg_QN,
         stateArray_S11reg_gff_1_SFF_7_QD,
         stateArray_S11reg_gff_1_SFF_7_MUXInst_Y,
         stateArray_S11reg_gff_1_SFF_7_MUXInst_X,
         stateArray_S11reg_gff_1_SFF_7_Q_reg_QN,
         stateArray_S12reg_gff_1_SFF_0_QD,
         stateArray_S12reg_gff_1_SFF_0_MUXInst_Y,
         stateArray_S12reg_gff_1_SFF_0_MUXInst_X,
         stateArray_S12reg_gff_1_SFF_0_Q_reg_QN,
         stateArray_S12reg_gff_1_SFF_1_QD,
         stateArray_S12reg_gff_1_SFF_1_MUXInst_Y,
         stateArray_S12reg_gff_1_SFF_1_MUXInst_X,
         stateArray_S12reg_gff_1_SFF_1_Q_reg_QN,
         stateArray_S12reg_gff_1_SFF_2_QD,
         stateArray_S12reg_gff_1_SFF_2_MUXInst_Y,
         stateArray_S12reg_gff_1_SFF_2_MUXInst_X,
         stateArray_S12reg_gff_1_SFF_2_Q_reg_QN,
         stateArray_S12reg_gff_1_SFF_3_QD,
         stateArray_S12reg_gff_1_SFF_3_MUXInst_Y,
         stateArray_S12reg_gff_1_SFF_3_MUXInst_X,
         stateArray_S12reg_gff_1_SFF_3_Q_reg_QN,
         stateArray_S12reg_gff_1_SFF_4_QD,
         stateArray_S12reg_gff_1_SFF_4_MUXInst_Y,
         stateArray_S12reg_gff_1_SFF_4_MUXInst_X,
         stateArray_S12reg_gff_1_SFF_4_Q_reg_QN,
         stateArray_S12reg_gff_1_SFF_5_QD,
         stateArray_S12reg_gff_1_SFF_5_MUXInst_Y,
         stateArray_S12reg_gff_1_SFF_5_MUXInst_X,
         stateArray_S12reg_gff_1_SFF_5_Q_reg_QN,
         stateArray_S12reg_gff_1_SFF_6_QD,
         stateArray_S12reg_gff_1_SFF_6_MUXInst_Y,
         stateArray_S12reg_gff_1_SFF_6_MUXInst_X,
         stateArray_S12reg_gff_1_SFF_6_Q_reg_QN,
         stateArray_S12reg_gff_1_SFF_7_QD,
         stateArray_S12reg_gff_1_SFF_7_MUXInst_Y,
         stateArray_S12reg_gff_1_SFF_7_MUXInst_X,
         stateArray_S12reg_gff_1_SFF_7_Q_reg_QN,
         stateArray_S13reg_gff_1_SFF_0_QD,
         stateArray_S13reg_gff_1_SFF_0_MUXInst_Y,
         stateArray_S13reg_gff_1_SFF_0_MUXInst_X,
         stateArray_S13reg_gff_1_SFF_0_Q_reg_QN,
         stateArray_S13reg_gff_1_SFF_1_QD,
         stateArray_S13reg_gff_1_SFF_1_MUXInst_Y,
         stateArray_S13reg_gff_1_SFF_1_MUXInst_X,
         stateArray_S13reg_gff_1_SFF_1_Q_reg_QN,
         stateArray_S13reg_gff_1_SFF_2_QD,
         stateArray_S13reg_gff_1_SFF_2_MUXInst_Y,
         stateArray_S13reg_gff_1_SFF_2_MUXInst_X,
         stateArray_S13reg_gff_1_SFF_2_Q_reg_QN,
         stateArray_S13reg_gff_1_SFF_3_QD,
         stateArray_S13reg_gff_1_SFF_3_MUXInst_Y,
         stateArray_S13reg_gff_1_SFF_3_MUXInst_X,
         stateArray_S13reg_gff_1_SFF_3_Q_reg_QN,
         stateArray_S13reg_gff_1_SFF_4_QD,
         stateArray_S13reg_gff_1_SFF_4_MUXInst_Y,
         stateArray_S13reg_gff_1_SFF_4_MUXInst_X,
         stateArray_S13reg_gff_1_SFF_4_Q_reg_QN,
         stateArray_S13reg_gff_1_SFF_5_QD,
         stateArray_S13reg_gff_1_SFF_5_MUXInst_Y,
         stateArray_S13reg_gff_1_SFF_5_MUXInst_X,
         stateArray_S13reg_gff_1_SFF_5_Q_reg_QN,
         stateArray_S13reg_gff_1_SFF_6_QD,
         stateArray_S13reg_gff_1_SFF_6_MUXInst_Y,
         stateArray_S13reg_gff_1_SFF_6_MUXInst_X,
         stateArray_S13reg_gff_1_SFF_6_Q_reg_QN,
         stateArray_S13reg_gff_1_SFF_7_QD,
         stateArray_S13reg_gff_1_SFF_7_MUXInst_Y,
         stateArray_S13reg_gff_1_SFF_7_MUXInst_X,
         stateArray_S13reg_gff_1_SFF_7_Q_reg_QN,
         stateArray_S20reg_gff_1_SFF_0_QD,
         stateArray_S20reg_gff_1_SFF_0_MUXInst_Y,
         stateArray_S20reg_gff_1_SFF_0_MUXInst_X,
         stateArray_S20reg_gff_1_SFF_0_Q_reg_QN,
         stateArray_S20reg_gff_1_SFF_1_QD,
         stateArray_S20reg_gff_1_SFF_1_MUXInst_Y,
         stateArray_S20reg_gff_1_SFF_1_MUXInst_X,
         stateArray_S20reg_gff_1_SFF_1_Q_reg_QN,
         stateArray_S20reg_gff_1_SFF_2_QD,
         stateArray_S20reg_gff_1_SFF_2_MUXInst_Y,
         stateArray_S20reg_gff_1_SFF_2_MUXInst_X,
         stateArray_S20reg_gff_1_SFF_2_Q_reg_QN,
         stateArray_S20reg_gff_1_SFF_3_QD,
         stateArray_S20reg_gff_1_SFF_3_MUXInst_Y,
         stateArray_S20reg_gff_1_SFF_3_MUXInst_X,
         stateArray_S20reg_gff_1_SFF_3_Q_reg_QN,
         stateArray_S20reg_gff_1_SFF_4_QD,
         stateArray_S20reg_gff_1_SFF_4_MUXInst_Y,
         stateArray_S20reg_gff_1_SFF_4_MUXInst_X,
         stateArray_S20reg_gff_1_SFF_4_Q_reg_QN,
         stateArray_S20reg_gff_1_SFF_5_QD,
         stateArray_S20reg_gff_1_SFF_5_MUXInst_Y,
         stateArray_S20reg_gff_1_SFF_5_MUXInst_X,
         stateArray_S20reg_gff_1_SFF_5_Q_reg_QN,
         stateArray_S20reg_gff_1_SFF_6_QD,
         stateArray_S20reg_gff_1_SFF_6_MUXInst_Y,
         stateArray_S20reg_gff_1_SFF_6_MUXInst_X,
         stateArray_S20reg_gff_1_SFF_6_Q_reg_QN,
         stateArray_S20reg_gff_1_SFF_7_QD,
         stateArray_S20reg_gff_1_SFF_7_MUXInst_Y,
         stateArray_S20reg_gff_1_SFF_7_MUXInst_X,
         stateArray_S20reg_gff_1_SFF_7_Q_reg_QN,
         stateArray_S21reg_gff_1_SFF_0_QD,
         stateArray_S21reg_gff_1_SFF_0_MUXInst_Y,
         stateArray_S21reg_gff_1_SFF_0_MUXInst_X,
         stateArray_S21reg_gff_1_SFF_0_Q_reg_QN,
         stateArray_S21reg_gff_1_SFF_1_QD,
         stateArray_S21reg_gff_1_SFF_1_MUXInst_Y,
         stateArray_S21reg_gff_1_SFF_1_MUXInst_X,
         stateArray_S21reg_gff_1_SFF_1_Q_reg_QN,
         stateArray_S21reg_gff_1_SFF_2_QD,
         stateArray_S21reg_gff_1_SFF_2_MUXInst_Y,
         stateArray_S21reg_gff_1_SFF_2_MUXInst_X,
         stateArray_S21reg_gff_1_SFF_2_Q_reg_QN,
         stateArray_S21reg_gff_1_SFF_3_QD,
         stateArray_S21reg_gff_1_SFF_3_MUXInst_Y,
         stateArray_S21reg_gff_1_SFF_3_MUXInst_X,
         stateArray_S21reg_gff_1_SFF_3_Q_reg_QN,
         stateArray_S21reg_gff_1_SFF_4_QD,
         stateArray_S21reg_gff_1_SFF_4_MUXInst_Y,
         stateArray_S21reg_gff_1_SFF_4_MUXInst_X,
         stateArray_S21reg_gff_1_SFF_4_Q_reg_QN,
         stateArray_S21reg_gff_1_SFF_5_QD,
         stateArray_S21reg_gff_1_SFF_5_MUXInst_Y,
         stateArray_S21reg_gff_1_SFF_5_MUXInst_X,
         stateArray_S21reg_gff_1_SFF_5_Q_reg_QN,
         stateArray_S21reg_gff_1_SFF_6_QD,
         stateArray_S21reg_gff_1_SFF_6_MUXInst_Y,
         stateArray_S21reg_gff_1_SFF_6_MUXInst_X,
         stateArray_S21reg_gff_1_SFF_6_Q_reg_QN,
         stateArray_S21reg_gff_1_SFF_7_QD,
         stateArray_S21reg_gff_1_SFF_7_MUXInst_Y,
         stateArray_S21reg_gff_1_SFF_7_MUXInst_X,
         stateArray_S21reg_gff_1_SFF_7_Q_reg_QN,
         stateArray_S22reg_gff_1_SFF_0_QD,
         stateArray_S22reg_gff_1_SFF_0_MUXInst_Y,
         stateArray_S22reg_gff_1_SFF_0_MUXInst_X,
         stateArray_S22reg_gff_1_SFF_0_Q_reg_QN,
         stateArray_S22reg_gff_1_SFF_1_QD,
         stateArray_S22reg_gff_1_SFF_1_MUXInst_Y,
         stateArray_S22reg_gff_1_SFF_1_MUXInst_X,
         stateArray_S22reg_gff_1_SFF_1_Q_reg_QN,
         stateArray_S22reg_gff_1_SFF_2_QD,
         stateArray_S22reg_gff_1_SFF_2_MUXInst_Y,
         stateArray_S22reg_gff_1_SFF_2_MUXInst_X,
         stateArray_S22reg_gff_1_SFF_2_Q_reg_QN,
         stateArray_S22reg_gff_1_SFF_3_QD,
         stateArray_S22reg_gff_1_SFF_3_MUXInst_Y,
         stateArray_S22reg_gff_1_SFF_3_MUXInst_X,
         stateArray_S22reg_gff_1_SFF_3_Q_reg_QN,
         stateArray_S22reg_gff_1_SFF_4_QD,
         stateArray_S22reg_gff_1_SFF_4_MUXInst_Y,
         stateArray_S22reg_gff_1_SFF_4_MUXInst_X,
         stateArray_S22reg_gff_1_SFF_4_Q_reg_QN,
         stateArray_S22reg_gff_1_SFF_5_QD,
         stateArray_S22reg_gff_1_SFF_5_MUXInst_Y,
         stateArray_S22reg_gff_1_SFF_5_MUXInst_X,
         stateArray_S22reg_gff_1_SFF_5_Q_reg_QN,
         stateArray_S22reg_gff_1_SFF_6_QD,
         stateArray_S22reg_gff_1_SFF_6_MUXInst_Y,
         stateArray_S22reg_gff_1_SFF_6_MUXInst_X,
         stateArray_S22reg_gff_1_SFF_6_Q_reg_QN,
         stateArray_S22reg_gff_1_SFF_7_QD,
         stateArray_S22reg_gff_1_SFF_7_MUXInst_Y,
         stateArray_S22reg_gff_1_SFF_7_MUXInst_X,
         stateArray_S22reg_gff_1_SFF_7_Q_reg_QN,
         stateArray_S23reg_gff_1_SFF_0_QD,
         stateArray_S23reg_gff_1_SFF_0_MUXInst_Y,
         stateArray_S23reg_gff_1_SFF_0_MUXInst_X,
         stateArray_S23reg_gff_1_SFF_0_Q_reg_QN,
         stateArray_S23reg_gff_1_SFF_1_QD,
         stateArray_S23reg_gff_1_SFF_1_MUXInst_Y,
         stateArray_S23reg_gff_1_SFF_1_MUXInst_X,
         stateArray_S23reg_gff_1_SFF_1_Q_reg_QN,
         stateArray_S23reg_gff_1_SFF_2_QD,
         stateArray_S23reg_gff_1_SFF_2_MUXInst_Y,
         stateArray_S23reg_gff_1_SFF_2_MUXInst_X,
         stateArray_S23reg_gff_1_SFF_2_Q_reg_QN,
         stateArray_S23reg_gff_1_SFF_3_QD,
         stateArray_S23reg_gff_1_SFF_3_MUXInst_Y,
         stateArray_S23reg_gff_1_SFF_3_MUXInst_X,
         stateArray_S23reg_gff_1_SFF_3_Q_reg_QN,
         stateArray_S23reg_gff_1_SFF_4_QD,
         stateArray_S23reg_gff_1_SFF_4_MUXInst_Y,
         stateArray_S23reg_gff_1_SFF_4_MUXInst_X,
         stateArray_S23reg_gff_1_SFF_4_Q_reg_QN,
         stateArray_S23reg_gff_1_SFF_5_QD,
         stateArray_S23reg_gff_1_SFF_5_MUXInst_Y,
         stateArray_S23reg_gff_1_SFF_5_MUXInst_X,
         stateArray_S23reg_gff_1_SFF_5_Q_reg_QN,
         stateArray_S23reg_gff_1_SFF_6_QD,
         stateArray_S23reg_gff_1_SFF_6_MUXInst_Y,
         stateArray_S23reg_gff_1_SFF_6_MUXInst_X,
         stateArray_S23reg_gff_1_SFF_6_Q_reg_QN,
         stateArray_S23reg_gff_1_SFF_7_QD,
         stateArray_S23reg_gff_1_SFF_7_MUXInst_Y,
         stateArray_S23reg_gff_1_SFF_7_MUXInst_X,
         stateArray_S23reg_gff_1_SFF_7_Q_reg_QN,
         stateArray_S30reg_gff_1_SFF_0_QD,
         stateArray_S30reg_gff_1_SFF_0_MUXInst_Y,
         stateArray_S30reg_gff_1_SFF_0_MUXInst_X,
         stateArray_S30reg_gff_1_SFF_0_Q_reg_QN,
         stateArray_S30reg_gff_1_SFF_1_QD,
         stateArray_S30reg_gff_1_SFF_1_MUXInst_Y,
         stateArray_S30reg_gff_1_SFF_1_MUXInst_X,
         stateArray_S30reg_gff_1_SFF_1_Q_reg_QN,
         stateArray_S30reg_gff_1_SFF_2_QD,
         stateArray_S30reg_gff_1_SFF_2_MUXInst_Y,
         stateArray_S30reg_gff_1_SFF_2_MUXInst_X,
         stateArray_S30reg_gff_1_SFF_2_Q_reg_QN,
         stateArray_S30reg_gff_1_SFF_3_QD,
         stateArray_S30reg_gff_1_SFF_3_MUXInst_Y,
         stateArray_S30reg_gff_1_SFF_3_MUXInst_X,
         stateArray_S30reg_gff_1_SFF_3_Q_reg_QN,
         stateArray_S30reg_gff_1_SFF_4_QD,
         stateArray_S30reg_gff_1_SFF_4_MUXInst_Y,
         stateArray_S30reg_gff_1_SFF_4_MUXInst_X,
         stateArray_S30reg_gff_1_SFF_4_Q_reg_QN,
         stateArray_S30reg_gff_1_SFF_5_QD,
         stateArray_S30reg_gff_1_SFF_5_MUXInst_Y,
         stateArray_S30reg_gff_1_SFF_5_MUXInst_X,
         stateArray_S30reg_gff_1_SFF_5_Q_reg_QN,
         stateArray_S30reg_gff_1_SFF_6_QD,
         stateArray_S30reg_gff_1_SFF_6_MUXInst_Y,
         stateArray_S30reg_gff_1_SFF_6_MUXInst_X,
         stateArray_S30reg_gff_1_SFF_6_Q_reg_QN,
         stateArray_S30reg_gff_1_SFF_7_QD,
         stateArray_S30reg_gff_1_SFF_7_MUXInst_Y,
         stateArray_S30reg_gff_1_SFF_7_MUXInst_X,
         stateArray_S30reg_gff_1_SFF_7_Q_reg_QN,
         stateArray_S31reg_gff_1_SFF_0_QD,
         stateArray_S31reg_gff_1_SFF_0_MUXInst_Y,
         stateArray_S31reg_gff_1_SFF_0_MUXInst_X,
         stateArray_S31reg_gff_1_SFF_0_Q_reg_QN,
         stateArray_S31reg_gff_1_SFF_1_QD,
         stateArray_S31reg_gff_1_SFF_1_MUXInst_Y,
         stateArray_S31reg_gff_1_SFF_1_MUXInst_X,
         stateArray_S31reg_gff_1_SFF_1_Q_reg_QN,
         stateArray_S31reg_gff_1_SFF_2_QD,
         stateArray_S31reg_gff_1_SFF_2_MUXInst_Y,
         stateArray_S31reg_gff_1_SFF_2_MUXInst_X,
         stateArray_S31reg_gff_1_SFF_2_Q_reg_QN,
         stateArray_S31reg_gff_1_SFF_3_QD,
         stateArray_S31reg_gff_1_SFF_3_MUXInst_Y,
         stateArray_S31reg_gff_1_SFF_3_MUXInst_X,
         stateArray_S31reg_gff_1_SFF_3_Q_reg_QN,
         stateArray_S31reg_gff_1_SFF_4_QD,
         stateArray_S31reg_gff_1_SFF_4_MUXInst_Y,
         stateArray_S31reg_gff_1_SFF_4_MUXInst_X,
         stateArray_S31reg_gff_1_SFF_4_Q_reg_QN,
         stateArray_S31reg_gff_1_SFF_5_QD,
         stateArray_S31reg_gff_1_SFF_5_MUXInst_Y,
         stateArray_S31reg_gff_1_SFF_5_MUXInst_X,
         stateArray_S31reg_gff_1_SFF_5_Q_reg_QN,
         stateArray_S31reg_gff_1_SFF_6_QD,
         stateArray_S31reg_gff_1_SFF_6_MUXInst_Y,
         stateArray_S31reg_gff_1_SFF_6_MUXInst_X,
         stateArray_S31reg_gff_1_SFF_6_Q_reg_QN,
         stateArray_S31reg_gff_1_SFF_7_QD,
         stateArray_S31reg_gff_1_SFF_7_MUXInst_Y,
         stateArray_S31reg_gff_1_SFF_7_MUXInst_X,
         stateArray_S31reg_gff_1_SFF_7_Q_reg_QN,
         stateArray_S32reg_gff_1_SFF_0_QD,
         stateArray_S32reg_gff_1_SFF_0_MUXInst_Y,
         stateArray_S32reg_gff_1_SFF_0_MUXInst_X,
         stateArray_S32reg_gff_1_SFF_0_Q_reg_QN,
         stateArray_S32reg_gff_1_SFF_1_QD,
         stateArray_S32reg_gff_1_SFF_1_MUXInst_Y,
         stateArray_S32reg_gff_1_SFF_1_MUXInst_X,
         stateArray_S32reg_gff_1_SFF_1_Q_reg_QN,
         stateArray_S32reg_gff_1_SFF_2_QD,
         stateArray_S32reg_gff_1_SFF_2_MUXInst_Y,
         stateArray_S32reg_gff_1_SFF_2_MUXInst_X,
         stateArray_S32reg_gff_1_SFF_2_Q_reg_QN,
         stateArray_S32reg_gff_1_SFF_3_QD,
         stateArray_S32reg_gff_1_SFF_3_MUXInst_Y,
         stateArray_S32reg_gff_1_SFF_3_MUXInst_X,
         stateArray_S32reg_gff_1_SFF_3_Q_reg_QN,
         stateArray_S32reg_gff_1_SFF_4_QD,
         stateArray_S32reg_gff_1_SFF_4_MUXInst_Y,
         stateArray_S32reg_gff_1_SFF_4_MUXInst_X,
         stateArray_S32reg_gff_1_SFF_4_Q_reg_QN,
         stateArray_S32reg_gff_1_SFF_5_QD,
         stateArray_S32reg_gff_1_SFF_5_MUXInst_Y,
         stateArray_S32reg_gff_1_SFF_5_MUXInst_X,
         stateArray_S32reg_gff_1_SFF_5_Q_reg_QN,
         stateArray_S32reg_gff_1_SFF_6_QD,
         stateArray_S32reg_gff_1_SFF_6_MUXInst_Y,
         stateArray_S32reg_gff_1_SFF_6_MUXInst_X,
         stateArray_S32reg_gff_1_SFF_6_Q_reg_QN,
         stateArray_S32reg_gff_1_SFF_7_QD,
         stateArray_S32reg_gff_1_SFF_7_MUXInst_Y,
         stateArray_S32reg_gff_1_SFF_7_MUXInst_X,
         stateArray_S32reg_gff_1_SFF_7_Q_reg_QN,
         stateArray_S33reg_gff_1_SFF_0_QD,
         stateArray_S33reg_gff_1_SFF_0_MUXInst_Y,
         stateArray_S33reg_gff_1_SFF_0_MUXInst_X,
         stateArray_S33reg_gff_1_SFF_0_Q_reg_QN,
         stateArray_S33reg_gff_1_SFF_1_QD,
         stateArray_S33reg_gff_1_SFF_1_MUXInst_Y,
         stateArray_S33reg_gff_1_SFF_1_MUXInst_X,
         stateArray_S33reg_gff_1_SFF_1_Q_reg_QN,
         stateArray_S33reg_gff_1_SFF_2_QD,
         stateArray_S33reg_gff_1_SFF_2_MUXInst_Y,
         stateArray_S33reg_gff_1_SFF_2_MUXInst_X,
         stateArray_S33reg_gff_1_SFF_2_Q_reg_QN,
         stateArray_S33reg_gff_1_SFF_3_QD,
         stateArray_S33reg_gff_1_SFF_3_MUXInst_Y,
         stateArray_S33reg_gff_1_SFF_3_MUXInst_X,
         stateArray_S33reg_gff_1_SFF_3_Q_reg_QN,
         stateArray_S33reg_gff_1_SFF_4_QD,
         stateArray_S33reg_gff_1_SFF_4_MUXInst_Y,
         stateArray_S33reg_gff_1_SFF_4_MUXInst_X,
         stateArray_S33reg_gff_1_SFF_4_Q_reg_QN,
         stateArray_S33reg_gff_1_SFF_5_QD,
         stateArray_S33reg_gff_1_SFF_5_MUXInst_Y,
         stateArray_S33reg_gff_1_SFF_5_MUXInst_X,
         stateArray_S33reg_gff_1_SFF_5_Q_reg_QN,
         stateArray_S33reg_gff_1_SFF_6_QD,
         stateArray_S33reg_gff_1_SFF_6_MUXInst_Y,
         stateArray_S33reg_gff_1_SFF_6_MUXInst_X,
         stateArray_S33reg_gff_1_SFF_6_Q_reg_QN,
         stateArray_S33reg_gff_1_SFF_7_QD,
         stateArray_S33reg_gff_1_SFF_7_MUXInst_Y,
         stateArray_S33reg_gff_1_SFF_7_MUXInst_X,
         stateArray_S33reg_gff_1_SFF_7_Q_reg_QN,
         stateArray_MUX_inS03ser_mux_inst_0_Y,
         stateArray_MUX_inS03ser_mux_inst_0_X,
         stateArray_MUX_inS03ser_mux_inst_1_Y,
         stateArray_MUX_inS03ser_mux_inst_1_X,
         stateArray_MUX_inS03ser_mux_inst_2_Y,
         stateArray_MUX_inS03ser_mux_inst_2_X,
         stateArray_MUX_inS03ser_mux_inst_3_Y,
         stateArray_MUX_inS03ser_mux_inst_3_X,
         stateArray_MUX_inS03ser_mux_inst_4_Y,
         stateArray_MUX_inS03ser_mux_inst_4_X,
         stateArray_MUX_inS03ser_mux_inst_5_Y,
         stateArray_MUX_inS03ser_mux_inst_5_X,
         stateArray_MUX_inS03ser_mux_inst_6_Y,
         stateArray_MUX_inS03ser_mux_inst_6_X,
         stateArray_MUX_inS03ser_mux_inst_7_Y,
         stateArray_MUX_inS03ser_mux_inst_7_X,
         stateArray_MUX_inS13ser_mux_inst_0_Y,
         stateArray_MUX_inS13ser_mux_inst_0_X,
         stateArray_MUX_inS13ser_mux_inst_1_Y,
         stateArray_MUX_inS13ser_mux_inst_1_X,
         stateArray_MUX_inS13ser_mux_inst_2_Y,
         stateArray_MUX_inS13ser_mux_inst_2_X,
         stateArray_MUX_inS13ser_mux_inst_3_Y,
         stateArray_MUX_inS13ser_mux_inst_3_X,
         stateArray_MUX_inS13ser_mux_inst_4_Y,
         stateArray_MUX_inS13ser_mux_inst_4_X,
         stateArray_MUX_inS13ser_mux_inst_5_Y,
         stateArray_MUX_inS13ser_mux_inst_5_X,
         stateArray_MUX_inS13ser_mux_inst_6_Y,
         stateArray_MUX_inS13ser_mux_inst_6_X,
         stateArray_MUX_inS13ser_mux_inst_7_Y,
         stateArray_MUX_inS13ser_mux_inst_7_X,
         stateArray_MUX_inS23ser_mux_inst_0_Y,
         stateArray_MUX_inS23ser_mux_inst_0_X,
         stateArray_MUX_inS23ser_mux_inst_1_Y,
         stateArray_MUX_inS23ser_mux_inst_1_X,
         stateArray_MUX_inS23ser_mux_inst_2_Y,
         stateArray_MUX_inS23ser_mux_inst_2_X,
         stateArray_MUX_inS23ser_mux_inst_3_Y,
         stateArray_MUX_inS23ser_mux_inst_3_X,
         stateArray_MUX_inS23ser_mux_inst_4_Y,
         stateArray_MUX_inS23ser_mux_inst_4_X,
         stateArray_MUX_inS23ser_mux_inst_5_Y,
         stateArray_MUX_inS23ser_mux_inst_5_X,
         stateArray_MUX_inS23ser_mux_inst_6_Y,
         stateArray_MUX_inS23ser_mux_inst_6_X,
         stateArray_MUX_inS23ser_mux_inst_7_Y,
         stateArray_MUX_inS23ser_mux_inst_7_X,
         stateArray_MUX_input_MC_mux_inst_0_Y,
         stateArray_MUX_input_MC_mux_inst_0_X,
         stateArray_MUX_input_MC_mux_inst_1_Y,
         stateArray_MUX_input_MC_mux_inst_1_X,
         stateArray_MUX_input_MC_mux_inst_2_Y,
         stateArray_MUX_input_MC_mux_inst_2_X,
         stateArray_MUX_input_MC_mux_inst_3_Y,
         stateArray_MUX_input_MC_mux_inst_3_X,
         stateArray_MUX_input_MC_mux_inst_4_Y,
         stateArray_MUX_input_MC_mux_inst_4_X,
         stateArray_MUX_input_MC_mux_inst_5_Y,
         stateArray_MUX_input_MC_mux_inst_5_X,
         stateArray_MUX_input_MC_mux_inst_6_Y,
         stateArray_MUX_input_MC_mux_inst_6_X,
         stateArray_MUX_input_MC_mux_inst_7_Y,
         stateArray_MUX_input_MC_mux_inst_7_X,
         stateArray_MUX_inS33ser_mux_inst_0_Y,
         stateArray_MUX_inS33ser_mux_inst_0_X,
         stateArray_MUX_inS33ser_mux_inst_1_Y,
         stateArray_MUX_inS33ser_mux_inst_1_X,
         stateArray_MUX_inS33ser_mux_inst_2_Y,
         stateArray_MUX_inS33ser_mux_inst_2_X,
         stateArray_MUX_inS33ser_mux_inst_3_Y,
         stateArray_MUX_inS33ser_mux_inst_3_X,
         stateArray_MUX_inS33ser_mux_inst_4_Y,
         stateArray_MUX_inS33ser_mux_inst_4_X,
         stateArray_MUX_inS33ser_mux_inst_5_Y,
         stateArray_MUX_inS33ser_mux_inst_5_X,
         stateArray_MUX_inS33ser_mux_inst_6_Y,
         stateArray_MUX_inS33ser_mux_inst_6_X,
         stateArray_MUX_inS33ser_mux_inst_7_Y,
         stateArray_MUX_inS33ser_mux_inst_7_X, MUX_StateInMC_n4,
         MUX_StateInMC_n3, MUX_StateInMC_mux_inst_0_Y,
         MUX_StateInMC_mux_inst_0_X, MUX_StateInMC_mux_inst_1_Y,
         MUX_StateInMC_mux_inst_1_X, MUX_StateInMC_mux_inst_2_Y,
         MUX_StateInMC_mux_inst_2_X, MUX_StateInMC_mux_inst_3_Y,
         MUX_StateInMC_mux_inst_3_X, MUX_StateInMC_mux_inst_4_Y,
         MUX_StateInMC_mux_inst_4_X, MUX_StateInMC_mux_inst_5_Y,
         MUX_StateInMC_mux_inst_5_X, MUX_StateInMC_mux_inst_6_Y,
         MUX_StateInMC_mux_inst_6_X, MUX_StateInMC_mux_inst_7_Y,
         MUX_StateInMC_mux_inst_7_X, MUX_StateInMC_mux_inst_8_Y,
         MUX_StateInMC_mux_inst_8_X, MUX_StateInMC_mux_inst_9_Y,
         MUX_StateInMC_mux_inst_9_X, MUX_StateInMC_mux_inst_10_Y,
         MUX_StateInMC_mux_inst_10_X, MUX_StateInMC_mux_inst_11_Y,
         MUX_StateInMC_mux_inst_11_X, MUX_StateInMC_mux_inst_12_Y,
         MUX_StateInMC_mux_inst_12_X, MUX_StateInMC_mux_inst_13_Y,
         MUX_StateInMC_mux_inst_13_X, MUX_StateInMC_mux_inst_14_Y,
         MUX_StateInMC_mux_inst_14_X, MUX_StateInMC_mux_inst_15_Y,
         MUX_StateInMC_mux_inst_15_X, MUX_StateInMC_mux_inst_16_Y,
         MUX_StateInMC_mux_inst_16_X, MUX_StateInMC_mux_inst_17_Y,
         MUX_StateInMC_mux_inst_17_X, MUX_StateInMC_mux_inst_18_Y,
         MUX_StateInMC_mux_inst_18_X, MUX_StateInMC_mux_inst_19_Y,
         MUX_StateInMC_mux_inst_19_X, MUX_StateInMC_mux_inst_20_Y,
         MUX_StateInMC_mux_inst_20_X, MUX_StateInMC_mux_inst_21_Y,
         MUX_StateInMC_mux_inst_21_X, MUX_StateInMC_mux_inst_22_Y,
         MUX_StateInMC_mux_inst_22_X, MUX_StateInMC_mux_inst_23_Y,
         MUX_StateInMC_mux_inst_23_X, MUX_StateInMC_mux_inst_24_Y,
         MUX_StateInMC_mux_inst_24_X, MUX_StateInMC_mux_inst_25_Y,
         MUX_StateInMC_mux_inst_25_X, MUX_StateInMC_mux_inst_26_Y,
         MUX_StateInMC_mux_inst_26_X, MUX_StateInMC_mux_inst_27_Y,
         MUX_StateInMC_mux_inst_27_X, MUX_StateInMC_mux_inst_28_Y,
         MUX_StateInMC_mux_inst_28_X, MUX_StateInMC_mux_inst_29_Y,
         MUX_StateInMC_mux_inst_29_X, MUX_StateInMC_mux_inst_30_Y,
         MUX_StateInMC_mux_inst_30_X, MUX_StateInMC_mux_inst_31_Y,
         MUX_StateInMC_mux_inst_31_X, KeyArray_n32, KeyArray_n31, KeyArray_n30,
         KeyArray_n29, KeyArray_n28, KeyArray_n27, KeyArray_n26, KeyArray_n25,
         KeyArray_n24, KeyArray_n23, KeyArray_n22, KeyArray_n21, KeyArray_n20,
         KeyArray_n19, KeyArray_n18, KeyArray_nReset_selXOR,
         KeyArray_outS01ser_0_, KeyArray_outS01ser_1_, KeyArray_outS01ser_2_,
         KeyArray_outS01ser_3_, KeyArray_outS01ser_4_, KeyArray_outS01ser_5_,
         KeyArray_outS01ser_6_, KeyArray_outS01ser_7_,
         KeyArray_S00reg_gff_1_SFF_0_n2, KeyArray_S00reg_gff_1_SFF_0_n1,
         KeyArray_S00reg_gff_1_SFF_0_n3, KeyArray_S00reg_gff_1_SFF_0_n6,
         KeyArray_S00reg_gff_1_SFF_0_QD, KeyArray_S00reg_gff_1_SFF_0_MUXInst_Y,
         KeyArray_S00reg_gff_1_SFF_0_MUXInst_X, KeyArray_S00reg_gff_1_SFF_1_n2,
         KeyArray_S00reg_gff_1_SFF_1_n1, KeyArray_S00reg_gff_1_SFF_1_n11,
         KeyArray_S00reg_gff_1_SFF_1_n6, KeyArray_S00reg_gff_1_SFF_1_QD,
         KeyArray_S00reg_gff_1_SFF_1_MUXInst_Y,
         KeyArray_S00reg_gff_1_SFF_1_MUXInst_X, KeyArray_S00reg_gff_1_SFF_2_n2,
         KeyArray_S00reg_gff_1_SFF_2_n1, KeyArray_S00reg_gff_1_SFF_2_n11,
         KeyArray_S00reg_gff_1_SFF_2_n6, KeyArray_S00reg_gff_1_SFF_2_QD,
         KeyArray_S00reg_gff_1_SFF_2_MUXInst_Y,
         KeyArray_S00reg_gff_1_SFF_2_MUXInst_X, KeyArray_S00reg_gff_1_SFF_3_n2,
         KeyArray_S00reg_gff_1_SFF_3_n1, KeyArray_S00reg_gff_1_SFF_3_n11,
         KeyArray_S00reg_gff_1_SFF_3_n6, KeyArray_S00reg_gff_1_SFF_3_QD,
         KeyArray_S00reg_gff_1_SFF_3_MUXInst_Y,
         KeyArray_S00reg_gff_1_SFF_3_MUXInst_X, KeyArray_S00reg_gff_1_SFF_4_n2,
         KeyArray_S00reg_gff_1_SFF_4_n1, KeyArray_S00reg_gff_1_SFF_4_n11,
         KeyArray_S00reg_gff_1_SFF_4_n6, KeyArray_S00reg_gff_1_SFF_4_QD,
         KeyArray_S00reg_gff_1_SFF_4_MUXInst_Y,
         KeyArray_S00reg_gff_1_SFF_4_MUXInst_X, KeyArray_S00reg_gff_1_SFF_5_n2,
         KeyArray_S00reg_gff_1_SFF_5_n1, KeyArray_S00reg_gff_1_SFF_5_n11,
         KeyArray_S00reg_gff_1_SFF_5_n6, KeyArray_S00reg_gff_1_SFF_5_QD,
         KeyArray_S00reg_gff_1_SFF_5_MUXInst_Y,
         KeyArray_S00reg_gff_1_SFF_5_MUXInst_X, KeyArray_S00reg_gff_1_SFF_6_n2,
         KeyArray_S00reg_gff_1_SFF_6_n1, KeyArray_S00reg_gff_1_SFF_6_n11,
         KeyArray_S00reg_gff_1_SFF_6_n6, KeyArray_S00reg_gff_1_SFF_6_QD,
         KeyArray_S00reg_gff_1_SFF_6_MUXInst_Y,
         KeyArray_S00reg_gff_1_SFF_6_MUXInst_X, KeyArray_S00reg_gff_1_SFF_7_n2,
         KeyArray_S00reg_gff_1_SFF_7_n1, KeyArray_S00reg_gff_1_SFF_7_n11,
         KeyArray_S00reg_gff_1_SFF_7_n6, KeyArray_S00reg_gff_1_SFF_7_QD,
         KeyArray_S00reg_gff_1_SFF_7_MUXInst_Y,
         KeyArray_S00reg_gff_1_SFF_7_MUXInst_X, KeyArray_S01reg_gff_1_SFF_0_n2,
         KeyArray_S01reg_gff_1_SFF_0_n1, KeyArray_S01reg_gff_1_SFF_0_n11,
         KeyArray_S01reg_gff_1_SFF_0_n6, KeyArray_S01reg_gff_1_SFF_0_QD,
         KeyArray_S01reg_gff_1_SFF_0_MUXInst_Y,
         KeyArray_S01reg_gff_1_SFF_0_MUXInst_X, KeyArray_S01reg_gff_1_SFF_1_n2,
         KeyArray_S01reg_gff_1_SFF_1_n1, KeyArray_S01reg_gff_1_SFF_1_n11,
         KeyArray_S01reg_gff_1_SFF_1_n6, KeyArray_S01reg_gff_1_SFF_1_QD,
         KeyArray_S01reg_gff_1_SFF_1_MUXInst_Y,
         KeyArray_S01reg_gff_1_SFF_1_MUXInst_X, KeyArray_S01reg_gff_1_SFF_2_n2,
         KeyArray_S01reg_gff_1_SFF_2_n1, KeyArray_S01reg_gff_1_SFF_2_n11,
         KeyArray_S01reg_gff_1_SFF_2_n6, KeyArray_S01reg_gff_1_SFF_2_QD,
         KeyArray_S01reg_gff_1_SFF_2_MUXInst_Y,
         KeyArray_S01reg_gff_1_SFF_2_MUXInst_X, KeyArray_S01reg_gff_1_SFF_3_n2,
         KeyArray_S01reg_gff_1_SFF_3_n1, KeyArray_S01reg_gff_1_SFF_3_n11,
         KeyArray_S01reg_gff_1_SFF_3_n6, KeyArray_S01reg_gff_1_SFF_3_QD,
         KeyArray_S01reg_gff_1_SFF_3_MUXInst_Y,
         KeyArray_S01reg_gff_1_SFF_3_MUXInst_X, KeyArray_S01reg_gff_1_SFF_4_n2,
         KeyArray_S01reg_gff_1_SFF_4_n1, KeyArray_S01reg_gff_1_SFF_4_n11,
         KeyArray_S01reg_gff_1_SFF_4_n6, KeyArray_S01reg_gff_1_SFF_4_QD,
         KeyArray_S01reg_gff_1_SFF_4_MUXInst_Y,
         KeyArray_S01reg_gff_1_SFF_4_MUXInst_X, KeyArray_S01reg_gff_1_SFF_5_n2,
         KeyArray_S01reg_gff_1_SFF_5_n1, KeyArray_S01reg_gff_1_SFF_5_n11,
         KeyArray_S01reg_gff_1_SFF_5_n6, KeyArray_S01reg_gff_1_SFF_5_QD,
         KeyArray_S01reg_gff_1_SFF_5_MUXInst_Y,
         KeyArray_S01reg_gff_1_SFF_5_MUXInst_X, KeyArray_S01reg_gff_1_SFF_6_n2,
         KeyArray_S01reg_gff_1_SFF_6_n1, KeyArray_S01reg_gff_1_SFF_6_n11,
         KeyArray_S01reg_gff_1_SFF_6_n6, KeyArray_S01reg_gff_1_SFF_6_QD,
         KeyArray_S01reg_gff_1_SFF_6_MUXInst_Y,
         KeyArray_S01reg_gff_1_SFF_6_MUXInst_X, KeyArray_S01reg_gff_1_SFF_7_n2,
         KeyArray_S01reg_gff_1_SFF_7_n1, KeyArray_S01reg_gff_1_SFF_7_n11,
         KeyArray_S01reg_gff_1_SFF_7_n6, KeyArray_S01reg_gff_1_SFF_7_QD,
         KeyArray_S01reg_gff_1_SFF_7_MUXInst_Y,
         KeyArray_S01reg_gff_1_SFF_7_MUXInst_X, KeyArray_S02reg_gff_1_SFF_0_n2,
         KeyArray_S02reg_gff_1_SFF_0_n1, KeyArray_S02reg_gff_1_SFF_0_n11,
         KeyArray_S02reg_gff_1_SFF_0_n6, KeyArray_S02reg_gff_1_SFF_0_QD,
         KeyArray_S02reg_gff_1_SFF_0_MUXInst_Y,
         KeyArray_S02reg_gff_1_SFF_0_MUXInst_X, KeyArray_S02reg_gff_1_SFF_1_n2,
         KeyArray_S02reg_gff_1_SFF_1_n1, KeyArray_S02reg_gff_1_SFF_1_n11,
         KeyArray_S02reg_gff_1_SFF_1_n6, KeyArray_S02reg_gff_1_SFF_1_QD,
         KeyArray_S02reg_gff_1_SFF_1_MUXInst_Y,
         KeyArray_S02reg_gff_1_SFF_1_MUXInst_X, KeyArray_S02reg_gff_1_SFF_2_n2,
         KeyArray_S02reg_gff_1_SFF_2_n1, KeyArray_S02reg_gff_1_SFF_2_n11,
         KeyArray_S02reg_gff_1_SFF_2_n6, KeyArray_S02reg_gff_1_SFF_2_QD,
         KeyArray_S02reg_gff_1_SFF_2_MUXInst_Y,
         KeyArray_S02reg_gff_1_SFF_2_MUXInst_X, KeyArray_S02reg_gff_1_SFF_3_n2,
         KeyArray_S02reg_gff_1_SFF_3_n1, KeyArray_S02reg_gff_1_SFF_3_n11,
         KeyArray_S02reg_gff_1_SFF_3_n6, KeyArray_S02reg_gff_1_SFF_3_QD,
         KeyArray_S02reg_gff_1_SFF_3_MUXInst_Y,
         KeyArray_S02reg_gff_1_SFF_3_MUXInst_X, KeyArray_S02reg_gff_1_SFF_4_n2,
         KeyArray_S02reg_gff_1_SFF_4_n1, KeyArray_S02reg_gff_1_SFF_4_n11,
         KeyArray_S02reg_gff_1_SFF_4_n6, KeyArray_S02reg_gff_1_SFF_4_QD,
         KeyArray_S02reg_gff_1_SFF_4_MUXInst_Y,
         KeyArray_S02reg_gff_1_SFF_4_MUXInst_X, KeyArray_S02reg_gff_1_SFF_5_n2,
         KeyArray_S02reg_gff_1_SFF_5_n1, KeyArray_S02reg_gff_1_SFF_5_n11,
         KeyArray_S02reg_gff_1_SFF_5_n6, KeyArray_S02reg_gff_1_SFF_5_QD,
         KeyArray_S02reg_gff_1_SFF_5_MUXInst_Y,
         KeyArray_S02reg_gff_1_SFF_5_MUXInst_X, KeyArray_S02reg_gff_1_SFF_6_n2,
         KeyArray_S02reg_gff_1_SFF_6_n1, KeyArray_S02reg_gff_1_SFF_6_n11,
         KeyArray_S02reg_gff_1_SFF_6_n6, KeyArray_S02reg_gff_1_SFF_6_QD,
         KeyArray_S02reg_gff_1_SFF_6_MUXInst_Y,
         KeyArray_S02reg_gff_1_SFF_6_MUXInst_X, KeyArray_S02reg_gff_1_SFF_7_n2,
         KeyArray_S02reg_gff_1_SFF_7_n1, KeyArray_S02reg_gff_1_SFF_7_n11,
         KeyArray_S02reg_gff_1_SFF_7_n6, KeyArray_S02reg_gff_1_SFF_7_QD,
         KeyArray_S02reg_gff_1_SFF_7_MUXInst_Y,
         KeyArray_S02reg_gff_1_SFF_7_MUXInst_X, KeyArray_S03reg_gff_1_SFF_0_n2,
         KeyArray_S03reg_gff_1_SFF_0_n1, KeyArray_S03reg_gff_1_SFF_0_n11,
         KeyArray_S03reg_gff_1_SFF_0_n6, KeyArray_S03reg_gff_1_SFF_0_QD,
         KeyArray_S03reg_gff_1_SFF_0_MUXInst_Y,
         KeyArray_S03reg_gff_1_SFF_0_MUXInst_X, KeyArray_S03reg_gff_1_SFF_1_n2,
         KeyArray_S03reg_gff_1_SFF_1_n1, KeyArray_S03reg_gff_1_SFF_1_n11,
         KeyArray_S03reg_gff_1_SFF_1_n6, KeyArray_S03reg_gff_1_SFF_1_QD,
         KeyArray_S03reg_gff_1_SFF_1_MUXInst_Y,
         KeyArray_S03reg_gff_1_SFF_1_MUXInst_X, KeyArray_S03reg_gff_1_SFF_2_n2,
         KeyArray_S03reg_gff_1_SFF_2_n1, KeyArray_S03reg_gff_1_SFF_2_n11,
         KeyArray_S03reg_gff_1_SFF_2_n6, KeyArray_S03reg_gff_1_SFF_2_QD,
         KeyArray_S03reg_gff_1_SFF_2_MUXInst_Y,
         KeyArray_S03reg_gff_1_SFF_2_MUXInst_X, KeyArray_S03reg_gff_1_SFF_3_n2,
         KeyArray_S03reg_gff_1_SFF_3_n1, KeyArray_S03reg_gff_1_SFF_3_n11,
         KeyArray_S03reg_gff_1_SFF_3_n6, KeyArray_S03reg_gff_1_SFF_3_QD,
         KeyArray_S03reg_gff_1_SFF_3_MUXInst_Y,
         KeyArray_S03reg_gff_1_SFF_3_MUXInst_X, KeyArray_S03reg_gff_1_SFF_4_n2,
         KeyArray_S03reg_gff_1_SFF_4_n1, KeyArray_S03reg_gff_1_SFF_4_n11,
         KeyArray_S03reg_gff_1_SFF_4_n6, KeyArray_S03reg_gff_1_SFF_4_QD,
         KeyArray_S03reg_gff_1_SFF_4_MUXInst_Y,
         KeyArray_S03reg_gff_1_SFF_4_MUXInst_X, KeyArray_S03reg_gff_1_SFF_5_n2,
         KeyArray_S03reg_gff_1_SFF_5_n1, KeyArray_S03reg_gff_1_SFF_5_n3,
         KeyArray_S03reg_gff_1_SFF_5_n5, KeyArray_S03reg_gff_1_SFF_5_QD,
         KeyArray_S03reg_gff_1_SFF_5_MUXInst_Y,
         KeyArray_S03reg_gff_1_SFF_5_MUXInst_X, KeyArray_S03reg_gff_1_SFF_6_n2,
         KeyArray_S03reg_gff_1_SFF_6_n1, KeyArray_S03reg_gff_1_SFF_6_n10,
         KeyArray_S03reg_gff_1_SFF_6_n5, KeyArray_S03reg_gff_1_SFF_6_QD,
         KeyArray_S03reg_gff_1_SFF_6_MUXInst_Y,
         KeyArray_S03reg_gff_1_SFF_6_MUXInst_X, KeyArray_S03reg_gff_1_SFF_7_n2,
         KeyArray_S03reg_gff_1_SFF_7_n1, KeyArray_S03reg_gff_1_SFF_7_n10,
         KeyArray_S03reg_gff_1_SFF_7_n5, KeyArray_S03reg_gff_1_SFF_7_QD,
         KeyArray_S03reg_gff_1_SFF_7_MUXInst_Y,
         KeyArray_S03reg_gff_1_SFF_7_MUXInst_X, KeyArray_S10reg_gff_1_SFF_0_n2,
         KeyArray_S10reg_gff_1_SFF_0_n1, KeyArray_S10reg_gff_1_SFF_0_n10,
         KeyArray_S10reg_gff_1_SFF_0_n5, KeyArray_S10reg_gff_1_SFF_0_QD,
         KeyArray_S10reg_gff_1_SFF_0_MUXInst_Y,
         KeyArray_S10reg_gff_1_SFF_0_MUXInst_X, KeyArray_S10reg_gff_1_SFF_1_n2,
         KeyArray_S10reg_gff_1_SFF_1_n1, KeyArray_S10reg_gff_1_SFF_1_n10,
         KeyArray_S10reg_gff_1_SFF_1_n5, KeyArray_S10reg_gff_1_SFF_1_QD,
         KeyArray_S10reg_gff_1_SFF_1_MUXInst_Y,
         KeyArray_S10reg_gff_1_SFF_1_MUXInst_X, KeyArray_S10reg_gff_1_SFF_2_n2,
         KeyArray_S10reg_gff_1_SFF_2_n1, KeyArray_S10reg_gff_1_SFF_2_n10,
         KeyArray_S10reg_gff_1_SFF_2_n5, KeyArray_S10reg_gff_1_SFF_2_QD,
         KeyArray_S10reg_gff_1_SFF_2_MUXInst_Y,
         KeyArray_S10reg_gff_1_SFF_2_MUXInst_X, KeyArray_S10reg_gff_1_SFF_3_n2,
         KeyArray_S10reg_gff_1_SFF_3_n1, KeyArray_S10reg_gff_1_SFF_3_n10,
         KeyArray_S10reg_gff_1_SFF_3_n5, KeyArray_S10reg_gff_1_SFF_3_QD,
         KeyArray_S10reg_gff_1_SFF_3_MUXInst_Y,
         KeyArray_S10reg_gff_1_SFF_3_MUXInst_X, KeyArray_S10reg_gff_1_SFF_4_n2,
         KeyArray_S10reg_gff_1_SFF_4_n1, KeyArray_S10reg_gff_1_SFF_4_n10,
         KeyArray_S10reg_gff_1_SFF_4_n5, KeyArray_S10reg_gff_1_SFF_4_QD,
         KeyArray_S10reg_gff_1_SFF_4_MUXInst_Y,
         KeyArray_S10reg_gff_1_SFF_4_MUXInst_X, KeyArray_S10reg_gff_1_SFF_5_n2,
         KeyArray_S10reg_gff_1_SFF_5_n1, KeyArray_S10reg_gff_1_SFF_5_n10,
         KeyArray_S10reg_gff_1_SFF_5_n5, KeyArray_S10reg_gff_1_SFF_5_QD,
         KeyArray_S10reg_gff_1_SFF_5_MUXInst_Y,
         KeyArray_S10reg_gff_1_SFF_5_MUXInst_X, KeyArray_S10reg_gff_1_SFF_6_n2,
         KeyArray_S10reg_gff_1_SFF_6_n1, KeyArray_S10reg_gff_1_SFF_6_n10,
         KeyArray_S10reg_gff_1_SFF_6_n5, KeyArray_S10reg_gff_1_SFF_6_QD,
         KeyArray_S10reg_gff_1_SFF_6_MUXInst_Y,
         KeyArray_S10reg_gff_1_SFF_6_MUXInst_X, KeyArray_S10reg_gff_1_SFF_7_n2,
         KeyArray_S10reg_gff_1_SFF_7_n1, KeyArray_S10reg_gff_1_SFF_7_n10,
         KeyArray_S10reg_gff_1_SFF_7_n5, KeyArray_S10reg_gff_1_SFF_7_QD,
         KeyArray_S10reg_gff_1_SFF_7_MUXInst_Y,
         KeyArray_S10reg_gff_1_SFF_7_MUXInst_X, KeyArray_S11reg_gff_1_SFF_0_n2,
         KeyArray_S11reg_gff_1_SFF_0_n1, KeyArray_S11reg_gff_1_SFF_0_n11,
         KeyArray_S11reg_gff_1_SFF_0_n6, KeyArray_S11reg_gff_1_SFF_0_QD,
         KeyArray_S11reg_gff_1_SFF_0_MUXInst_Y,
         KeyArray_S11reg_gff_1_SFF_0_MUXInst_X, KeyArray_S11reg_gff_1_SFF_1_n2,
         KeyArray_S11reg_gff_1_SFF_1_n1, KeyArray_S11reg_gff_1_SFF_1_n11,
         KeyArray_S11reg_gff_1_SFF_1_n6, KeyArray_S11reg_gff_1_SFF_1_QD,
         KeyArray_S11reg_gff_1_SFF_1_MUXInst_Y,
         KeyArray_S11reg_gff_1_SFF_1_MUXInst_X, KeyArray_S11reg_gff_1_SFF_2_n2,
         KeyArray_S11reg_gff_1_SFF_2_n1, KeyArray_S11reg_gff_1_SFF_2_n11,
         KeyArray_S11reg_gff_1_SFF_2_n6, KeyArray_S11reg_gff_1_SFF_2_QD,
         KeyArray_S11reg_gff_1_SFF_2_MUXInst_Y,
         KeyArray_S11reg_gff_1_SFF_2_MUXInst_X, KeyArray_S11reg_gff_1_SFF_3_n2,
         KeyArray_S11reg_gff_1_SFF_3_n1, KeyArray_S11reg_gff_1_SFF_3_n11,
         KeyArray_S11reg_gff_1_SFF_3_n6, KeyArray_S11reg_gff_1_SFF_3_QD,
         KeyArray_S11reg_gff_1_SFF_3_MUXInst_Y,
         KeyArray_S11reg_gff_1_SFF_3_MUXInst_X, KeyArray_S11reg_gff_1_SFF_4_n2,
         KeyArray_S11reg_gff_1_SFF_4_n1, KeyArray_S11reg_gff_1_SFF_4_n11,
         KeyArray_S11reg_gff_1_SFF_4_n6, KeyArray_S11reg_gff_1_SFF_4_QD,
         KeyArray_S11reg_gff_1_SFF_4_MUXInst_Y,
         KeyArray_S11reg_gff_1_SFF_4_MUXInst_X, KeyArray_S11reg_gff_1_SFF_5_n2,
         KeyArray_S11reg_gff_1_SFF_5_n1, KeyArray_S11reg_gff_1_SFF_5_n11,
         KeyArray_S11reg_gff_1_SFF_5_n6, KeyArray_S11reg_gff_1_SFF_5_QD,
         KeyArray_S11reg_gff_1_SFF_5_MUXInst_Y,
         KeyArray_S11reg_gff_1_SFF_5_MUXInst_X, KeyArray_S11reg_gff_1_SFF_6_n2,
         KeyArray_S11reg_gff_1_SFF_6_n1, KeyArray_S11reg_gff_1_SFF_6_n11,
         KeyArray_S11reg_gff_1_SFF_6_n6, KeyArray_S11reg_gff_1_SFF_6_QD,
         KeyArray_S11reg_gff_1_SFF_6_MUXInst_Y,
         KeyArray_S11reg_gff_1_SFF_6_MUXInst_X, KeyArray_S11reg_gff_1_SFF_7_n2,
         KeyArray_S11reg_gff_1_SFF_7_n1, KeyArray_S11reg_gff_1_SFF_7_n11,
         KeyArray_S11reg_gff_1_SFF_7_n6, KeyArray_S11reg_gff_1_SFF_7_QD,
         KeyArray_S11reg_gff_1_SFF_7_MUXInst_Y,
         KeyArray_S11reg_gff_1_SFF_7_MUXInst_X, KeyArray_S12reg_gff_1_SFF_0_n2,
         KeyArray_S12reg_gff_1_SFF_0_n1, KeyArray_S12reg_gff_1_SFF_0_n11,
         KeyArray_S12reg_gff_1_SFF_0_n6, KeyArray_S12reg_gff_1_SFF_0_QD,
         KeyArray_S12reg_gff_1_SFF_0_MUXInst_Y,
         KeyArray_S12reg_gff_1_SFF_0_MUXInst_X, KeyArray_S12reg_gff_1_SFF_1_n2,
         KeyArray_S12reg_gff_1_SFF_1_n1, KeyArray_S12reg_gff_1_SFF_1_n11,
         KeyArray_S12reg_gff_1_SFF_1_n6, KeyArray_S12reg_gff_1_SFF_1_QD,
         KeyArray_S12reg_gff_1_SFF_1_MUXInst_Y,
         KeyArray_S12reg_gff_1_SFF_1_MUXInst_X, KeyArray_S12reg_gff_1_SFF_2_n2,
         KeyArray_S12reg_gff_1_SFF_2_n1, KeyArray_S12reg_gff_1_SFF_2_n11,
         KeyArray_S12reg_gff_1_SFF_2_n6, KeyArray_S12reg_gff_1_SFF_2_QD,
         KeyArray_S12reg_gff_1_SFF_2_MUXInst_Y,
         KeyArray_S12reg_gff_1_SFF_2_MUXInst_X, KeyArray_S12reg_gff_1_SFF_3_n2,
         KeyArray_S12reg_gff_1_SFF_3_n1, KeyArray_S12reg_gff_1_SFF_3_n11,
         KeyArray_S12reg_gff_1_SFF_3_n6, KeyArray_S12reg_gff_1_SFF_3_QD,
         KeyArray_S12reg_gff_1_SFF_3_MUXInst_Y,
         KeyArray_S12reg_gff_1_SFF_3_MUXInst_X, KeyArray_S12reg_gff_1_SFF_4_n2,
         KeyArray_S12reg_gff_1_SFF_4_n1, KeyArray_S12reg_gff_1_SFF_4_n11,
         KeyArray_S12reg_gff_1_SFF_4_n6, KeyArray_S12reg_gff_1_SFF_4_QD,
         KeyArray_S12reg_gff_1_SFF_4_MUXInst_Y,
         KeyArray_S12reg_gff_1_SFF_4_MUXInst_X, KeyArray_S12reg_gff_1_SFF_5_n2,
         KeyArray_S12reg_gff_1_SFF_5_n1, KeyArray_S12reg_gff_1_SFF_5_n11,
         KeyArray_S12reg_gff_1_SFF_5_n6, KeyArray_S12reg_gff_1_SFF_5_QD,
         KeyArray_S12reg_gff_1_SFF_5_MUXInst_Y,
         KeyArray_S12reg_gff_1_SFF_5_MUXInst_X, KeyArray_S12reg_gff_1_SFF_6_n2,
         KeyArray_S12reg_gff_1_SFF_6_n1, KeyArray_S12reg_gff_1_SFF_6_n11,
         KeyArray_S12reg_gff_1_SFF_6_n6, KeyArray_S12reg_gff_1_SFF_6_QD,
         KeyArray_S12reg_gff_1_SFF_6_MUXInst_Y,
         KeyArray_S12reg_gff_1_SFF_6_MUXInst_X, KeyArray_S12reg_gff_1_SFF_7_n2,
         KeyArray_S12reg_gff_1_SFF_7_n1, KeyArray_S12reg_gff_1_SFF_7_n11,
         KeyArray_S12reg_gff_1_SFF_7_n6, KeyArray_S12reg_gff_1_SFF_7_QD,
         KeyArray_S12reg_gff_1_SFF_7_MUXInst_Y,
         KeyArray_S12reg_gff_1_SFF_7_MUXInst_X, KeyArray_S13reg_gff_1_SFF_0_n2,
         KeyArray_S13reg_gff_1_SFF_0_n1, KeyArray_S13reg_gff_1_SFF_0_n11,
         KeyArray_S13reg_gff_1_SFF_0_n6, KeyArray_S13reg_gff_1_SFF_0_QD,
         KeyArray_S13reg_gff_1_SFF_0_MUXInst_Y,
         KeyArray_S13reg_gff_1_SFF_0_MUXInst_X, KeyArray_S13reg_gff_1_SFF_1_n2,
         KeyArray_S13reg_gff_1_SFF_1_n1, KeyArray_S13reg_gff_1_SFF_1_n11,
         KeyArray_S13reg_gff_1_SFF_1_n6, KeyArray_S13reg_gff_1_SFF_1_QD,
         KeyArray_S13reg_gff_1_SFF_1_MUXInst_Y,
         KeyArray_S13reg_gff_1_SFF_1_MUXInst_X, KeyArray_S13reg_gff_1_SFF_2_n2,
         KeyArray_S13reg_gff_1_SFF_2_n1, KeyArray_S13reg_gff_1_SFF_2_n11,
         KeyArray_S13reg_gff_1_SFF_2_n6, KeyArray_S13reg_gff_1_SFF_2_QD,
         KeyArray_S13reg_gff_1_SFF_2_MUXInst_Y,
         KeyArray_S13reg_gff_1_SFF_2_MUXInst_X, KeyArray_S13reg_gff_1_SFF_3_n2,
         KeyArray_S13reg_gff_1_SFF_3_n1, KeyArray_S13reg_gff_1_SFF_3_n11,
         KeyArray_S13reg_gff_1_SFF_3_n6, KeyArray_S13reg_gff_1_SFF_3_QD,
         KeyArray_S13reg_gff_1_SFF_3_MUXInst_Y,
         KeyArray_S13reg_gff_1_SFF_3_MUXInst_X, KeyArray_S13reg_gff_1_SFF_4_n2,
         KeyArray_S13reg_gff_1_SFF_4_n1, KeyArray_S13reg_gff_1_SFF_4_n11,
         KeyArray_S13reg_gff_1_SFF_4_n6, KeyArray_S13reg_gff_1_SFF_4_QD,
         KeyArray_S13reg_gff_1_SFF_4_MUXInst_Y,
         KeyArray_S13reg_gff_1_SFF_4_MUXInst_X, KeyArray_S13reg_gff_1_SFF_5_n2,
         KeyArray_S13reg_gff_1_SFF_5_n1, KeyArray_S13reg_gff_1_SFF_5_n10,
         KeyArray_S13reg_gff_1_SFF_5_n5, KeyArray_S13reg_gff_1_SFF_5_QD,
         KeyArray_S13reg_gff_1_SFF_5_MUXInst_Y,
         KeyArray_S13reg_gff_1_SFF_5_MUXInst_X, KeyArray_S13reg_gff_1_SFF_6_n2,
         KeyArray_S13reg_gff_1_SFF_6_n1, KeyArray_S13reg_gff_1_SFF_6_n10,
         KeyArray_S13reg_gff_1_SFF_6_n5, KeyArray_S13reg_gff_1_SFF_6_QD,
         KeyArray_S13reg_gff_1_SFF_6_MUXInst_Y,
         KeyArray_S13reg_gff_1_SFF_6_MUXInst_X, KeyArray_S13reg_gff_1_SFF_7_n2,
         KeyArray_S13reg_gff_1_SFF_7_n1, KeyArray_S13reg_gff_1_SFF_7_n10,
         KeyArray_S13reg_gff_1_SFF_7_n5, KeyArray_S13reg_gff_1_SFF_7_QD,
         KeyArray_S13reg_gff_1_SFF_7_MUXInst_Y,
         KeyArray_S13reg_gff_1_SFF_7_MUXInst_X, KeyArray_S20reg_gff_1_SFF_0_n2,
         KeyArray_S20reg_gff_1_SFF_0_n1, KeyArray_S20reg_gff_1_SFF_0_n10,
         KeyArray_S20reg_gff_1_SFF_0_n5, KeyArray_S20reg_gff_1_SFF_0_QD,
         KeyArray_S20reg_gff_1_SFF_0_MUXInst_Y,
         KeyArray_S20reg_gff_1_SFF_0_MUXInst_X, KeyArray_S20reg_gff_1_SFF_1_n2,
         KeyArray_S20reg_gff_1_SFF_1_n1, KeyArray_S20reg_gff_1_SFF_1_n10,
         KeyArray_S20reg_gff_1_SFF_1_n5, KeyArray_S20reg_gff_1_SFF_1_QD,
         KeyArray_S20reg_gff_1_SFF_1_MUXInst_Y,
         KeyArray_S20reg_gff_1_SFF_1_MUXInst_X, KeyArray_S20reg_gff_1_SFF_2_n2,
         KeyArray_S20reg_gff_1_SFF_2_n1, KeyArray_S20reg_gff_1_SFF_2_n10,
         KeyArray_S20reg_gff_1_SFF_2_n5, KeyArray_S20reg_gff_1_SFF_2_QD,
         KeyArray_S20reg_gff_1_SFF_2_MUXInst_Y,
         KeyArray_S20reg_gff_1_SFF_2_MUXInst_X, KeyArray_S20reg_gff_1_SFF_3_n2,
         KeyArray_S20reg_gff_1_SFF_3_n1, KeyArray_S20reg_gff_1_SFF_3_n10,
         KeyArray_S20reg_gff_1_SFF_3_n5, KeyArray_S20reg_gff_1_SFF_3_QD,
         KeyArray_S20reg_gff_1_SFF_3_MUXInst_Y,
         KeyArray_S20reg_gff_1_SFF_3_MUXInst_X, KeyArray_S20reg_gff_1_SFF_4_n2,
         KeyArray_S20reg_gff_1_SFF_4_n1, KeyArray_S20reg_gff_1_SFF_4_n10,
         KeyArray_S20reg_gff_1_SFF_4_n5, KeyArray_S20reg_gff_1_SFF_4_QD,
         KeyArray_S20reg_gff_1_SFF_4_MUXInst_Y,
         KeyArray_S20reg_gff_1_SFF_4_MUXInst_X, KeyArray_S20reg_gff_1_SFF_5_n2,
         KeyArray_S20reg_gff_1_SFF_5_n1, KeyArray_S20reg_gff_1_SFF_5_n10,
         KeyArray_S20reg_gff_1_SFF_5_n5, KeyArray_S20reg_gff_1_SFF_5_QD,
         KeyArray_S20reg_gff_1_SFF_5_MUXInst_Y,
         KeyArray_S20reg_gff_1_SFF_5_MUXInst_X, KeyArray_S20reg_gff_1_SFF_6_n2,
         KeyArray_S20reg_gff_1_SFF_6_n1, KeyArray_S20reg_gff_1_SFF_6_n10,
         KeyArray_S20reg_gff_1_SFF_6_n5, KeyArray_S20reg_gff_1_SFF_6_QD,
         KeyArray_S20reg_gff_1_SFF_6_MUXInst_Y,
         KeyArray_S20reg_gff_1_SFF_6_MUXInst_X, KeyArray_S20reg_gff_1_SFF_7_n2,
         KeyArray_S20reg_gff_1_SFF_7_n1, KeyArray_S20reg_gff_1_SFF_7_n10,
         KeyArray_S20reg_gff_1_SFF_7_n5, KeyArray_S20reg_gff_1_SFF_7_QD,
         KeyArray_S20reg_gff_1_SFF_7_MUXInst_Y,
         KeyArray_S20reg_gff_1_SFF_7_MUXInst_X, KeyArray_S21reg_gff_1_SFF_0_n2,
         KeyArray_S21reg_gff_1_SFF_0_n1, KeyArray_S21reg_gff_1_SFF_0_n11,
         KeyArray_S21reg_gff_1_SFF_0_n6, KeyArray_S21reg_gff_1_SFF_0_QD,
         KeyArray_S21reg_gff_1_SFF_0_MUXInst_Y,
         KeyArray_S21reg_gff_1_SFF_0_MUXInst_X, KeyArray_S21reg_gff_1_SFF_1_n2,
         KeyArray_S21reg_gff_1_SFF_1_n1, KeyArray_S21reg_gff_1_SFF_1_n11,
         KeyArray_S21reg_gff_1_SFF_1_n6, KeyArray_S21reg_gff_1_SFF_1_QD,
         KeyArray_S21reg_gff_1_SFF_1_MUXInst_Y,
         KeyArray_S21reg_gff_1_SFF_1_MUXInst_X, KeyArray_S21reg_gff_1_SFF_2_n2,
         KeyArray_S21reg_gff_1_SFF_2_n1, KeyArray_S21reg_gff_1_SFF_2_n11,
         KeyArray_S21reg_gff_1_SFF_2_n6, KeyArray_S21reg_gff_1_SFF_2_QD,
         KeyArray_S21reg_gff_1_SFF_2_MUXInst_Y,
         KeyArray_S21reg_gff_1_SFF_2_MUXInst_X, KeyArray_S21reg_gff_1_SFF_3_n2,
         KeyArray_S21reg_gff_1_SFF_3_n1, KeyArray_S21reg_gff_1_SFF_3_n11,
         KeyArray_S21reg_gff_1_SFF_3_n6, KeyArray_S21reg_gff_1_SFF_3_QD,
         KeyArray_S21reg_gff_1_SFF_3_MUXInst_Y,
         KeyArray_S21reg_gff_1_SFF_3_MUXInst_X, KeyArray_S21reg_gff_1_SFF_4_n2,
         KeyArray_S21reg_gff_1_SFF_4_n1, KeyArray_S21reg_gff_1_SFF_4_n11,
         KeyArray_S21reg_gff_1_SFF_4_n6, KeyArray_S21reg_gff_1_SFF_4_QD,
         KeyArray_S21reg_gff_1_SFF_4_MUXInst_Y,
         KeyArray_S21reg_gff_1_SFF_4_MUXInst_X, KeyArray_S21reg_gff_1_SFF_5_n2,
         KeyArray_S21reg_gff_1_SFF_5_n1, KeyArray_S21reg_gff_1_SFF_5_n11,
         KeyArray_S21reg_gff_1_SFF_5_n6, KeyArray_S21reg_gff_1_SFF_5_QD,
         KeyArray_S21reg_gff_1_SFF_5_MUXInst_Y,
         KeyArray_S21reg_gff_1_SFF_5_MUXInst_X, KeyArray_S21reg_gff_1_SFF_6_n2,
         KeyArray_S21reg_gff_1_SFF_6_n1, KeyArray_S21reg_gff_1_SFF_6_n11,
         KeyArray_S21reg_gff_1_SFF_6_n6, KeyArray_S21reg_gff_1_SFF_6_QD,
         KeyArray_S21reg_gff_1_SFF_6_MUXInst_Y,
         KeyArray_S21reg_gff_1_SFF_6_MUXInst_X, KeyArray_S21reg_gff_1_SFF_7_n2,
         KeyArray_S21reg_gff_1_SFF_7_n1, KeyArray_S21reg_gff_1_SFF_7_n11,
         KeyArray_S21reg_gff_1_SFF_7_n6, KeyArray_S21reg_gff_1_SFF_7_QD,
         KeyArray_S21reg_gff_1_SFF_7_MUXInst_Y,
         KeyArray_S21reg_gff_1_SFF_7_MUXInst_X, KeyArray_S22reg_gff_1_SFF_0_n2,
         KeyArray_S22reg_gff_1_SFF_0_n1, KeyArray_S22reg_gff_1_SFF_0_n11,
         KeyArray_S22reg_gff_1_SFF_0_n6, KeyArray_S22reg_gff_1_SFF_0_QD,
         KeyArray_S22reg_gff_1_SFF_0_MUXInst_Y,
         KeyArray_S22reg_gff_1_SFF_0_MUXInst_X, KeyArray_S22reg_gff_1_SFF_1_n2,
         KeyArray_S22reg_gff_1_SFF_1_n1, KeyArray_S22reg_gff_1_SFF_1_n11,
         KeyArray_S22reg_gff_1_SFF_1_n6, KeyArray_S22reg_gff_1_SFF_1_QD,
         KeyArray_S22reg_gff_1_SFF_1_MUXInst_Y,
         KeyArray_S22reg_gff_1_SFF_1_MUXInst_X, KeyArray_S22reg_gff_1_SFF_2_n2,
         KeyArray_S22reg_gff_1_SFF_2_n1, KeyArray_S22reg_gff_1_SFF_2_n11,
         KeyArray_S22reg_gff_1_SFF_2_n6, KeyArray_S22reg_gff_1_SFF_2_QD,
         KeyArray_S22reg_gff_1_SFF_2_MUXInst_Y,
         KeyArray_S22reg_gff_1_SFF_2_MUXInst_X, KeyArray_S22reg_gff_1_SFF_3_n2,
         KeyArray_S22reg_gff_1_SFF_3_n1, KeyArray_S22reg_gff_1_SFF_3_n11,
         KeyArray_S22reg_gff_1_SFF_3_n6, KeyArray_S22reg_gff_1_SFF_3_QD,
         KeyArray_S22reg_gff_1_SFF_3_MUXInst_Y,
         KeyArray_S22reg_gff_1_SFF_3_MUXInst_X, KeyArray_S22reg_gff_1_SFF_4_n2,
         KeyArray_S22reg_gff_1_SFF_4_n1, KeyArray_S22reg_gff_1_SFF_4_n11,
         KeyArray_S22reg_gff_1_SFF_4_n6, KeyArray_S22reg_gff_1_SFF_4_QD,
         KeyArray_S22reg_gff_1_SFF_4_MUXInst_Y,
         KeyArray_S22reg_gff_1_SFF_4_MUXInst_X, KeyArray_S22reg_gff_1_SFF_5_n2,
         KeyArray_S22reg_gff_1_SFF_5_n1, KeyArray_S22reg_gff_1_SFF_5_n11,
         KeyArray_S22reg_gff_1_SFF_5_n6, KeyArray_S22reg_gff_1_SFF_5_QD,
         KeyArray_S22reg_gff_1_SFF_5_MUXInst_Y,
         KeyArray_S22reg_gff_1_SFF_5_MUXInst_X, KeyArray_S22reg_gff_1_SFF_6_n2,
         KeyArray_S22reg_gff_1_SFF_6_n1, KeyArray_S22reg_gff_1_SFF_6_n11,
         KeyArray_S22reg_gff_1_SFF_6_n6, KeyArray_S22reg_gff_1_SFF_6_QD,
         KeyArray_S22reg_gff_1_SFF_6_MUXInst_Y,
         KeyArray_S22reg_gff_1_SFF_6_MUXInst_X, KeyArray_S22reg_gff_1_SFF_7_n2,
         KeyArray_S22reg_gff_1_SFF_7_n1, KeyArray_S22reg_gff_1_SFF_7_n11,
         KeyArray_S22reg_gff_1_SFF_7_n6, KeyArray_S22reg_gff_1_SFF_7_QD,
         KeyArray_S22reg_gff_1_SFF_7_MUXInst_Y,
         KeyArray_S22reg_gff_1_SFF_7_MUXInst_X, KeyArray_S23reg_gff_1_SFF_0_n2,
         KeyArray_S23reg_gff_1_SFF_0_n1, KeyArray_S23reg_gff_1_SFF_0_n11,
         KeyArray_S23reg_gff_1_SFF_0_n6, KeyArray_S23reg_gff_1_SFF_0_QD,
         KeyArray_S23reg_gff_1_SFF_0_MUXInst_Y,
         KeyArray_S23reg_gff_1_SFF_0_MUXInst_X, KeyArray_S23reg_gff_1_SFF_1_n2,
         KeyArray_S23reg_gff_1_SFF_1_n1, KeyArray_S23reg_gff_1_SFF_1_n11,
         KeyArray_S23reg_gff_1_SFF_1_n6, KeyArray_S23reg_gff_1_SFF_1_QD,
         KeyArray_S23reg_gff_1_SFF_1_MUXInst_Y,
         KeyArray_S23reg_gff_1_SFF_1_MUXInst_X, KeyArray_S23reg_gff_1_SFF_2_n2,
         KeyArray_S23reg_gff_1_SFF_2_n1, KeyArray_S23reg_gff_1_SFF_2_n11,
         KeyArray_S23reg_gff_1_SFF_2_n6, KeyArray_S23reg_gff_1_SFF_2_QD,
         KeyArray_S23reg_gff_1_SFF_2_MUXInst_Y,
         KeyArray_S23reg_gff_1_SFF_2_MUXInst_X, KeyArray_S23reg_gff_1_SFF_3_n2,
         KeyArray_S23reg_gff_1_SFF_3_n1, KeyArray_S23reg_gff_1_SFF_3_n11,
         KeyArray_S23reg_gff_1_SFF_3_n6, KeyArray_S23reg_gff_1_SFF_3_QD,
         KeyArray_S23reg_gff_1_SFF_3_MUXInst_Y,
         KeyArray_S23reg_gff_1_SFF_3_MUXInst_X, KeyArray_S23reg_gff_1_SFF_4_n2,
         KeyArray_S23reg_gff_1_SFF_4_n1, KeyArray_S23reg_gff_1_SFF_4_n11,
         KeyArray_S23reg_gff_1_SFF_4_n6, KeyArray_S23reg_gff_1_SFF_4_QD,
         KeyArray_S23reg_gff_1_SFF_4_MUXInst_Y,
         KeyArray_S23reg_gff_1_SFF_4_MUXInst_X, KeyArray_S23reg_gff_1_SFF_5_n2,
         KeyArray_S23reg_gff_1_SFF_5_n1, KeyArray_S23reg_gff_1_SFF_5_n10,
         KeyArray_S23reg_gff_1_SFF_5_n5, KeyArray_S23reg_gff_1_SFF_5_QD,
         KeyArray_S23reg_gff_1_SFF_5_MUXInst_Y,
         KeyArray_S23reg_gff_1_SFF_5_MUXInst_X, KeyArray_S23reg_gff_1_SFF_6_n2,
         KeyArray_S23reg_gff_1_SFF_6_n1, KeyArray_S23reg_gff_1_SFF_6_n10,
         KeyArray_S23reg_gff_1_SFF_6_n5, KeyArray_S23reg_gff_1_SFF_6_QD,
         KeyArray_S23reg_gff_1_SFF_6_MUXInst_Y,
         KeyArray_S23reg_gff_1_SFF_6_MUXInst_X, KeyArray_S23reg_gff_1_SFF_7_n2,
         KeyArray_S23reg_gff_1_SFF_7_n1, KeyArray_S23reg_gff_1_SFF_7_n10,
         KeyArray_S23reg_gff_1_SFF_7_n5, KeyArray_S23reg_gff_1_SFF_7_QD,
         KeyArray_S23reg_gff_1_SFF_7_MUXInst_Y,
         KeyArray_S23reg_gff_1_SFF_7_MUXInst_X, KeyArray_S30reg_gff_1_SFF_0_n2,
         KeyArray_S30reg_gff_1_SFF_0_n1, KeyArray_S30reg_gff_1_SFF_0_n10,
         KeyArray_S30reg_gff_1_SFF_0_n5, KeyArray_S30reg_gff_1_SFF_0_QD,
         KeyArray_S30reg_gff_1_SFF_0_MUXInst_Y,
         KeyArray_S30reg_gff_1_SFF_0_MUXInst_X, KeyArray_S30reg_gff_1_SFF_1_n2,
         KeyArray_S30reg_gff_1_SFF_1_n1, KeyArray_S30reg_gff_1_SFF_1_n10,
         KeyArray_S30reg_gff_1_SFF_1_n5, KeyArray_S30reg_gff_1_SFF_1_QD,
         KeyArray_S30reg_gff_1_SFF_1_MUXInst_Y,
         KeyArray_S30reg_gff_1_SFF_1_MUXInst_X, KeyArray_S30reg_gff_1_SFF_2_n2,
         KeyArray_S30reg_gff_1_SFF_2_n1, KeyArray_S30reg_gff_1_SFF_2_n10,
         KeyArray_S30reg_gff_1_SFF_2_n5, KeyArray_S30reg_gff_1_SFF_2_QD,
         KeyArray_S30reg_gff_1_SFF_2_MUXInst_Y,
         KeyArray_S30reg_gff_1_SFF_2_MUXInst_X, KeyArray_S30reg_gff_1_SFF_3_n2,
         KeyArray_S30reg_gff_1_SFF_3_n1, KeyArray_S30reg_gff_1_SFF_3_n10,
         KeyArray_S30reg_gff_1_SFF_3_n5, KeyArray_S30reg_gff_1_SFF_3_QD,
         KeyArray_S30reg_gff_1_SFF_3_MUXInst_Y,
         KeyArray_S30reg_gff_1_SFF_3_MUXInst_X, KeyArray_S30reg_gff_1_SFF_4_n2,
         KeyArray_S30reg_gff_1_SFF_4_n1, KeyArray_S30reg_gff_1_SFF_4_n10,
         KeyArray_S30reg_gff_1_SFF_4_n5, KeyArray_S30reg_gff_1_SFF_4_QD,
         KeyArray_S30reg_gff_1_SFF_4_MUXInst_Y,
         KeyArray_S30reg_gff_1_SFF_4_MUXInst_X, KeyArray_S30reg_gff_1_SFF_5_n2,
         KeyArray_S30reg_gff_1_SFF_5_n1, KeyArray_S30reg_gff_1_SFF_5_n10,
         KeyArray_S30reg_gff_1_SFF_5_n5, KeyArray_S30reg_gff_1_SFF_5_QD,
         KeyArray_S30reg_gff_1_SFF_5_MUXInst_Y,
         KeyArray_S30reg_gff_1_SFF_5_MUXInst_X, KeyArray_S30reg_gff_1_SFF_6_n2,
         KeyArray_S30reg_gff_1_SFF_6_n1, KeyArray_S30reg_gff_1_SFF_6_n10,
         KeyArray_S30reg_gff_1_SFF_6_n5, KeyArray_S30reg_gff_1_SFF_6_QD,
         KeyArray_S30reg_gff_1_SFF_6_MUXInst_Y,
         KeyArray_S30reg_gff_1_SFF_6_MUXInst_X, KeyArray_S30reg_gff_1_SFF_7_n2,
         KeyArray_S30reg_gff_1_SFF_7_n1, KeyArray_S30reg_gff_1_SFF_7_n10,
         KeyArray_S30reg_gff_1_SFF_7_n5, KeyArray_S30reg_gff_1_SFF_7_QD,
         KeyArray_S30reg_gff_1_SFF_7_MUXInst_Y,
         KeyArray_S30reg_gff_1_SFF_7_MUXInst_X, KeyArray_S31reg_gff_1_SFF_0_n2,
         KeyArray_S31reg_gff_1_SFF_0_n1, KeyArray_S31reg_gff_1_SFF_0_n11,
         KeyArray_S31reg_gff_1_SFF_0_n6, KeyArray_S31reg_gff_1_SFF_0_QD,
         KeyArray_S31reg_gff_1_SFF_0_MUXInst_Y,
         KeyArray_S31reg_gff_1_SFF_0_MUXInst_X, KeyArray_S31reg_gff_1_SFF_1_n2,
         KeyArray_S31reg_gff_1_SFF_1_n1, KeyArray_S31reg_gff_1_SFF_1_n11,
         KeyArray_S31reg_gff_1_SFF_1_n6, KeyArray_S31reg_gff_1_SFF_1_QD,
         KeyArray_S31reg_gff_1_SFF_1_MUXInst_Y,
         KeyArray_S31reg_gff_1_SFF_1_MUXInst_X, KeyArray_S31reg_gff_1_SFF_2_n2,
         KeyArray_S31reg_gff_1_SFF_2_n1, KeyArray_S31reg_gff_1_SFF_2_n11,
         KeyArray_S31reg_gff_1_SFF_2_n6, KeyArray_S31reg_gff_1_SFF_2_QD,
         KeyArray_S31reg_gff_1_SFF_2_MUXInst_Y,
         KeyArray_S31reg_gff_1_SFF_2_MUXInst_X, KeyArray_S31reg_gff_1_SFF_3_n2,
         KeyArray_S31reg_gff_1_SFF_3_n1, KeyArray_S31reg_gff_1_SFF_3_n11,
         KeyArray_S31reg_gff_1_SFF_3_n6, KeyArray_S31reg_gff_1_SFF_3_QD,
         KeyArray_S31reg_gff_1_SFF_3_MUXInst_Y,
         KeyArray_S31reg_gff_1_SFF_3_MUXInst_X, KeyArray_S31reg_gff_1_SFF_4_n2,
         KeyArray_S31reg_gff_1_SFF_4_n1, KeyArray_S31reg_gff_1_SFF_4_n11,
         KeyArray_S31reg_gff_1_SFF_4_n6, KeyArray_S31reg_gff_1_SFF_4_QD,
         KeyArray_S31reg_gff_1_SFF_4_MUXInst_Y,
         KeyArray_S31reg_gff_1_SFF_4_MUXInst_X, KeyArray_S31reg_gff_1_SFF_5_n2,
         KeyArray_S31reg_gff_1_SFF_5_n1, KeyArray_S31reg_gff_1_SFF_5_n11,
         KeyArray_S31reg_gff_1_SFF_5_n6, KeyArray_S31reg_gff_1_SFF_5_QD,
         KeyArray_S31reg_gff_1_SFF_5_MUXInst_Y,
         KeyArray_S31reg_gff_1_SFF_5_MUXInst_X, KeyArray_S31reg_gff_1_SFF_6_n2,
         KeyArray_S31reg_gff_1_SFF_6_n1, KeyArray_S31reg_gff_1_SFF_6_n11,
         KeyArray_S31reg_gff_1_SFF_6_n6, KeyArray_S31reg_gff_1_SFF_6_QD,
         KeyArray_S31reg_gff_1_SFF_6_MUXInst_Y,
         KeyArray_S31reg_gff_1_SFF_6_MUXInst_X, KeyArray_S31reg_gff_1_SFF_7_n2,
         KeyArray_S31reg_gff_1_SFF_7_n1, KeyArray_S31reg_gff_1_SFF_7_n11,
         KeyArray_S31reg_gff_1_SFF_7_n6, KeyArray_S31reg_gff_1_SFF_7_QD,
         KeyArray_S31reg_gff_1_SFF_7_MUXInst_Y,
         KeyArray_S31reg_gff_1_SFF_7_MUXInst_X, KeyArray_S32reg_gff_1_SFF_0_n2,
         KeyArray_S32reg_gff_1_SFF_0_n1, KeyArray_S32reg_gff_1_SFF_0_n11,
         KeyArray_S32reg_gff_1_SFF_0_n6, KeyArray_S32reg_gff_1_SFF_0_QD,
         KeyArray_S32reg_gff_1_SFF_0_MUXInst_Y,
         KeyArray_S32reg_gff_1_SFF_0_MUXInst_X, KeyArray_S32reg_gff_1_SFF_1_n2,
         KeyArray_S32reg_gff_1_SFF_1_n1, KeyArray_S32reg_gff_1_SFF_1_n11,
         KeyArray_S32reg_gff_1_SFF_1_n6, KeyArray_S32reg_gff_1_SFF_1_QD,
         KeyArray_S32reg_gff_1_SFF_1_MUXInst_Y,
         KeyArray_S32reg_gff_1_SFF_1_MUXInst_X, KeyArray_S32reg_gff_1_SFF_2_n2,
         KeyArray_S32reg_gff_1_SFF_2_n1, KeyArray_S32reg_gff_1_SFF_2_n11,
         KeyArray_S32reg_gff_1_SFF_2_n6, KeyArray_S32reg_gff_1_SFF_2_QD,
         KeyArray_S32reg_gff_1_SFF_2_MUXInst_Y,
         KeyArray_S32reg_gff_1_SFF_2_MUXInst_X, KeyArray_S32reg_gff_1_SFF_3_n2,
         KeyArray_S32reg_gff_1_SFF_3_n1, KeyArray_S32reg_gff_1_SFF_3_n11,
         KeyArray_S32reg_gff_1_SFF_3_n6, KeyArray_S32reg_gff_1_SFF_3_QD,
         KeyArray_S32reg_gff_1_SFF_3_MUXInst_Y,
         KeyArray_S32reg_gff_1_SFF_3_MUXInst_X, KeyArray_S32reg_gff_1_SFF_4_n2,
         KeyArray_S32reg_gff_1_SFF_4_n1, KeyArray_S32reg_gff_1_SFF_4_n11,
         KeyArray_S32reg_gff_1_SFF_4_n6, KeyArray_S32reg_gff_1_SFF_4_QD,
         KeyArray_S32reg_gff_1_SFF_4_MUXInst_Y,
         KeyArray_S32reg_gff_1_SFF_4_MUXInst_X, KeyArray_S32reg_gff_1_SFF_5_n2,
         KeyArray_S32reg_gff_1_SFF_5_n1, KeyArray_S32reg_gff_1_SFF_5_n10,
         KeyArray_S32reg_gff_1_SFF_5_n5, KeyArray_S32reg_gff_1_SFF_5_QD,
         KeyArray_S32reg_gff_1_SFF_5_MUXInst_Y,
         KeyArray_S32reg_gff_1_SFF_5_MUXInst_X, KeyArray_S32reg_gff_1_SFF_6_n2,
         KeyArray_S32reg_gff_1_SFF_6_n1, KeyArray_S32reg_gff_1_SFF_6_n10,
         KeyArray_S32reg_gff_1_SFF_6_n5, KeyArray_S32reg_gff_1_SFF_6_QD,
         KeyArray_S32reg_gff_1_SFF_6_MUXInst_Y,
         KeyArray_S32reg_gff_1_SFF_6_MUXInst_X, KeyArray_S32reg_gff_1_SFF_7_n2,
         KeyArray_S32reg_gff_1_SFF_7_n1, KeyArray_S32reg_gff_1_SFF_7_n10,
         KeyArray_S32reg_gff_1_SFF_7_n5, KeyArray_S32reg_gff_1_SFF_7_QD,
         KeyArray_S32reg_gff_1_SFF_7_MUXInst_Y,
         KeyArray_S32reg_gff_1_SFF_7_MUXInst_X, KeyArray_S33reg_gff_1_SFF_0_n2,
         KeyArray_S33reg_gff_1_SFF_0_n1, KeyArray_S33reg_gff_1_SFF_0_n10,
         KeyArray_S33reg_gff_1_SFF_0_n5, KeyArray_S33reg_gff_1_SFF_0_QD,
         KeyArray_S33reg_gff_1_SFF_0_MUXInst_Y,
         KeyArray_S33reg_gff_1_SFF_0_MUXInst_X, KeyArray_S33reg_gff_1_SFF_1_n2,
         KeyArray_S33reg_gff_1_SFF_1_n1, KeyArray_S33reg_gff_1_SFF_1_n10,
         KeyArray_S33reg_gff_1_SFF_1_n5, KeyArray_S33reg_gff_1_SFF_1_QD,
         KeyArray_S33reg_gff_1_SFF_1_MUXInst_Y,
         KeyArray_S33reg_gff_1_SFF_1_MUXInst_X, KeyArray_S33reg_gff_1_SFF_2_n2,
         KeyArray_S33reg_gff_1_SFF_2_n1, KeyArray_S33reg_gff_1_SFF_2_n10,
         KeyArray_S33reg_gff_1_SFF_2_n5, KeyArray_S33reg_gff_1_SFF_2_QD,
         KeyArray_S33reg_gff_1_SFF_2_MUXInst_Y,
         KeyArray_S33reg_gff_1_SFF_2_MUXInst_X, KeyArray_S33reg_gff_1_SFF_3_n2,
         KeyArray_S33reg_gff_1_SFF_3_n1, KeyArray_S33reg_gff_1_SFF_3_n10,
         KeyArray_S33reg_gff_1_SFF_3_n5, KeyArray_S33reg_gff_1_SFF_3_QD,
         KeyArray_S33reg_gff_1_SFF_3_MUXInst_Y,
         KeyArray_S33reg_gff_1_SFF_3_MUXInst_X, KeyArray_S33reg_gff_1_SFF_4_n2,
         KeyArray_S33reg_gff_1_SFF_4_n1, KeyArray_S33reg_gff_1_SFF_4_n10,
         KeyArray_S33reg_gff_1_SFF_4_n5, KeyArray_S33reg_gff_1_SFF_4_QD,
         KeyArray_S33reg_gff_1_SFF_4_MUXInst_Y,
         KeyArray_S33reg_gff_1_SFF_4_MUXInst_X, KeyArray_S33reg_gff_1_SFF_5_n2,
         KeyArray_S33reg_gff_1_SFF_5_n1, KeyArray_S33reg_gff_1_SFF_5_n10,
         KeyArray_S33reg_gff_1_SFF_5_n5, KeyArray_S33reg_gff_1_SFF_5_QD,
         KeyArray_S33reg_gff_1_SFF_5_MUXInst_Y,
         KeyArray_S33reg_gff_1_SFF_5_MUXInst_X, KeyArray_S33reg_gff_1_SFF_6_n2,
         KeyArray_S33reg_gff_1_SFF_6_n1, KeyArray_S33reg_gff_1_SFF_6_n10,
         KeyArray_S33reg_gff_1_SFF_6_n5, KeyArray_S33reg_gff_1_SFF_6_QD,
         KeyArray_S33reg_gff_1_SFF_6_MUXInst_Y,
         KeyArray_S33reg_gff_1_SFF_6_MUXInst_X, KeyArray_S33reg_gff_1_SFF_7_n2,
         KeyArray_S33reg_gff_1_SFF_7_n1, KeyArray_S33reg_gff_1_SFF_7_n10,
         KeyArray_S33reg_gff_1_SFF_7_n5, KeyArray_S33reg_gff_1_SFF_7_QD,
         KeyArray_S33reg_gff_1_SFF_7_MUXInst_Y,
         KeyArray_S33reg_gff_1_SFF_7_MUXInst_X,
         KeyArray_MUX_inS00ser_mux_inst_0_Y,
         KeyArray_MUX_inS00ser_mux_inst_0_X,
         KeyArray_MUX_inS00ser_mux_inst_1_Y,
         KeyArray_MUX_inS00ser_mux_inst_1_X,
         KeyArray_MUX_inS00ser_mux_inst_2_Y,
         KeyArray_MUX_inS00ser_mux_inst_2_X,
         KeyArray_MUX_inS00ser_mux_inst_3_Y,
         KeyArray_MUX_inS00ser_mux_inst_3_X,
         KeyArray_MUX_inS00ser_mux_inst_4_Y,
         KeyArray_MUX_inS00ser_mux_inst_4_X,
         KeyArray_MUX_inS00ser_mux_inst_5_Y,
         KeyArray_MUX_inS00ser_mux_inst_5_X,
         KeyArray_MUX_inS00ser_mux_inst_6_Y,
         KeyArray_MUX_inS00ser_mux_inst_6_X,
         KeyArray_MUX_inS00ser_mux_inst_7_Y,
         KeyArray_MUX_inS00ser_mux_inst_7_X,
         KeyArray_MUX_inS33ser_mux_inst_0_Y,
         KeyArray_MUX_inS33ser_mux_inst_0_X,
         KeyArray_MUX_inS33ser_mux_inst_1_Y,
         KeyArray_MUX_inS33ser_mux_inst_1_X,
         KeyArray_MUX_inS33ser_mux_inst_2_Y,
         KeyArray_MUX_inS33ser_mux_inst_2_X,
         KeyArray_MUX_inS33ser_mux_inst_3_Y,
         KeyArray_MUX_inS33ser_mux_inst_3_X,
         KeyArray_MUX_inS33ser_mux_inst_4_Y,
         KeyArray_MUX_inS33ser_mux_inst_4_X,
         KeyArray_MUX_inS33ser_mux_inst_5_Y,
         KeyArray_MUX_inS33ser_mux_inst_5_X,
         KeyArray_MUX_inS33ser_mux_inst_6_Y,
         KeyArray_MUX_inS33ser_mux_inst_6_X,
         KeyArray_MUX_inS33ser_mux_inst_7_Y,
         KeyArray_MUX_inS33ser_mux_inst_7_X, MixColumns_line0_n16,
         MixColumns_line0_n15, MixColumns_line0_n14, MixColumns_line0_n13,
         MixColumns_line0_n12, MixColumns_line0_n11, MixColumns_line0_n10,
         MixColumns_line0_n9, MixColumns_line0_n8, MixColumns_line0_n7,
         MixColumns_line0_n6, MixColumns_line0_n5, MixColumns_line0_n4,
         MixColumns_line0_n3, MixColumns_line0_n2, MixColumns_line0_n1,
         MixColumns_line1_n16, MixColumns_line1_n15, MixColumns_line1_n14,
         MixColumns_line1_n13, MixColumns_line1_n12, MixColumns_line1_n11,
         MixColumns_line1_n10, MixColumns_line1_n9, MixColumns_line1_n8,
         MixColumns_line1_n7, MixColumns_line1_n6, MixColumns_line1_n5,
         MixColumns_line1_n4, MixColumns_line1_n3, MixColumns_line1_n2,
         MixColumns_line1_n1, MixColumns_line2_n16, MixColumns_line2_n15,
         MixColumns_line2_n14, MixColumns_line2_n13, MixColumns_line2_n12,
         MixColumns_line2_n11, MixColumns_line2_n10, MixColumns_line2_n9,
         MixColumns_line2_n8, MixColumns_line2_n7, MixColumns_line2_n6,
         MixColumns_line2_n5, MixColumns_line2_n4, MixColumns_line2_n3,
         MixColumns_line2_n2, MixColumns_line2_n1, MixColumns_line3_n16,
         MixColumns_line3_n15, MixColumns_line3_n14, MixColumns_line3_n13,
         MixColumns_line3_n12, MixColumns_line3_n11, MixColumns_line3_n10,
         MixColumns_line3_n9, MixColumns_line3_n8, MixColumns_line3_n7,
         MixColumns_line3_n6, MixColumns_line3_n5, MixColumns_line3_n4,
         MixColumns_line3_n3, MixColumns_line3_n2, MixColumns_line3_n1,
         MixColumns_line3_timesTHREE_input2_1_,
         MixColumns_line3_timesTHREE_input2_3_,
         MixColumns_line3_timesTHREE_input2_4_, calcRCon_n43, calcRCon_n42,
         calcRCon_n41, calcRCon_n40, calcRCon_n39, calcRCon_n38, calcRCon_n37,
         calcRCon_n36, calcRCon_n35, calcRCon_n34, calcRCon_n33, calcRCon_n32,
         calcRCon_n31, calcRCon_n30, calcRCon_n29, calcRCon_n28, calcRCon_n27,
         calcRCon_n26, calcRCon_n25, calcRCon_n24, calcRCon_n23, calcRCon_n22,
         calcRCon_n21, calcRCon_n20, calcRCon_n19, calcRCon_n18, calcRCon_n17,
         calcRCon_n16, calcRCon_n15, calcRCon_n14, calcRCon_n13, calcRCon_n9,
         calcRCon_n8, calcRCon_n7, calcRCon_n6, calcRCon_n4, calcRCon_n3,
         calcRCon_n2, calcRCon_n1, calcRCon_n10, calcRCon_n44, calcRCon_n45,
         calcRCon_n46, calcRCon_n47, calcRCon_n48, calcRCon_n11, calcRCon_n49,
         calcRCon_n50, calcRCon_n12, calcRCon_s_current_state_0_,
         calcRCon_s_current_state_1_, calcRCon_s_current_state_2_,
         calcRCon_s_current_state_3_, calcRCon_s_current_state_4_,
         calcRCon_s_current_state_5_, calcRCon_s_current_state_6_,
         calcRCon_s_current_state_7_, calcRCon_n51,
         calcRCon_s_current_state_reg_3__QN, MUX_SboxIn_mux_inst_0_Y,
         MUX_SboxIn_mux_inst_0_X, MUX_SboxIn_mux_inst_1_Y,
         MUX_SboxIn_mux_inst_1_X, MUX_SboxIn_mux_inst_2_Y,
         MUX_SboxIn_mux_inst_2_X, MUX_SboxIn_mux_inst_3_Y,
         MUX_SboxIn_mux_inst_3_X, MUX_SboxIn_mux_inst_4_Y,
         MUX_SboxIn_mux_inst_4_X, MUX_SboxIn_mux_inst_5_Y,
         MUX_SboxIn_mux_inst_5_X, MUX_SboxIn_mux_inst_6_Y,
         MUX_SboxIn_mux_inst_6_X, MUX_SboxIn_mux_inst_7_Y,
         MUX_SboxIn_mux_inst_7_X, Inst_bSbox_L29, Inst_bSbox_L28,
         Inst_bSbox_L27, Inst_bSbox_L26, Inst_bSbox_L25, Inst_bSbox_L24,
         Inst_bSbox_L23, Inst_bSbox_L22, Inst_bSbox_L21, Inst_bSbox_L20,
         Inst_bSbox_L19, Inst_bSbox_L18, Inst_bSbox_L17, Inst_bSbox_L16,
         Inst_bSbox_L15, Inst_bSbox_L14, Inst_bSbox_L13, Inst_bSbox_L12,
         Inst_bSbox_L11, Inst_bSbox_L10, Inst_bSbox_L9, Inst_bSbox_L8,
         Inst_bSbox_L7, Inst_bSbox_L6, Inst_bSbox_L5, Inst_bSbox_L4,
         Inst_bSbox_L3, Inst_bSbox_L2, Inst_bSbox_L1, Inst_bSbox_L0,
         Inst_bSbox_M63, Inst_bSbox_M62, Inst_bSbox_M61, Inst_bSbox_M60,
         Inst_bSbox_M59, Inst_bSbox_M58, Inst_bSbox_M57, Inst_bSbox_M56,
         Inst_bSbox_M55, Inst_bSbox_M54, Inst_bSbox_M53, Inst_bSbox_M52,
         Inst_bSbox_M51, Inst_bSbox_M50, Inst_bSbox_M49, Inst_bSbox_M48,
         Inst_bSbox_M47, Inst_bSbox_M46, Inst_bSbox_M45, Inst_bSbox_M44,
         Inst_bSbox_M43, Inst_bSbox_M42, Inst_bSbox_M41, Inst_bSbox_M40,
         Inst_bSbox_M39, Inst_bSbox_M38, Inst_bSbox_M37, Inst_bSbox_M36,
         Inst_bSbox_M35, Inst_bSbox_M34, Inst_bSbox_M33, Inst_bSbox_M32,
         Inst_bSbox_M31, Inst_bSbox_M30, Inst_bSbox_M29, Inst_bSbox_M28,
         Inst_bSbox_M27, Inst_bSbox_M26, Inst_bSbox_M25, Inst_bSbox_M24,
         Inst_bSbox_M23, Inst_bSbox_M22, Inst_bSbox_M21, Inst_bSbox_M20,
         Inst_bSbox_M19, Inst_bSbox_M18, Inst_bSbox_M17, Inst_bSbox_M16,
         Inst_bSbox_M15, Inst_bSbox_M14, Inst_bSbox_M13, Inst_bSbox_M12,
         Inst_bSbox_M11, Inst_bSbox_M10, Inst_bSbox_M9, Inst_bSbox_M8,
         Inst_bSbox_M7, Inst_bSbox_M6, Inst_bSbox_M5, Inst_bSbox_M4,
         Inst_bSbox_M3, Inst_bSbox_M2, Inst_bSbox_M1, Inst_bSbox_T27,
         Inst_bSbox_T26, Inst_bSbox_T25, Inst_bSbox_T24, Inst_bSbox_T23,
         Inst_bSbox_T22, Inst_bSbox_T21, Inst_bSbox_T20, Inst_bSbox_T19,
         Inst_bSbox_T18, Inst_bSbox_T17, Inst_bSbox_T16, Inst_bSbox_T15,
         Inst_bSbox_T14, Inst_bSbox_T13, Inst_bSbox_T12, Inst_bSbox_T11,
         Inst_bSbox_T10, Inst_bSbox_T9, Inst_bSbox_T8, Inst_bSbox_T7,
         Inst_bSbox_T6, Inst_bSbox_T5, Inst_bSbox_T4, Inst_bSbox_T3,
         Inst_bSbox_T2, Inst_bSbox_T1;
  wire   [7:0] SboxOut;
  wire   [7:0] StateOutXORroundKey;
  wire   [7:0] StateIn;
  wire   [31:0] StateInMC;
  wire   [19:0] MCin;
  wire   [31:0] MCout;
  wire   [7:0] keyStateIn;
  wire   [7:0] roundConstant;
  wire   [7:0] keySBIn;
  wire   [7:0] SboxIn;
  wire   [7:0] stateArray_input_MC;
  wire   [7:0] stateArray_inS33ser;
  wire   [7:0] stateArray_outS33ser;
  wire   [7:0] stateArray_outS32ser;
  wire   [7:0] stateArray_outS31ser;
  wire   [7:0] stateArray_inS23ser;
  wire   [7:0] stateArray_outS23ser;
  wire   [7:0] stateArray_outS22ser;
  wire   [7:0] stateArray_outS21ser;
  wire   [7:0] stateArray_inS13ser;
  wire   [7:0] stateArray_outS13ser;
  wire   [7:0] stateArray_outS12ser;
  wire   [7:0] stateArray_outS11ser;
  wire   [7:0] stateArray_inS03ser;
  wire   [7:0] stateArray_outS03ser;
  wire   [7:0] stateArray_outS02ser;
  wire   [7:0] stateArray_outS01ser;
  wire   [7:0] KeyArray_outS01ser_XOR_00;
  wire   [7:0] KeyArray_inS33ser;
  wire   [7:0] KeyArray_outS33ser;
  wire   [7:0] KeyArray_outS32ser;
  wire   [7:0] KeyArray_inS30par;
  wire   [7:0] KeyArray_outS31ser;
  wire   [7:0] KeyArray_outS30ser;
  wire   [7:0] KeyArray_outS23ser;
  wire   [7:0] KeyArray_outS22ser;
  wire   [7:0] KeyArray_outS21ser;
  wire   [7:0] KeyArray_outS20ser;
  wire   [7:0] KeyArray_outS12ser;
  wire   [7:0] KeyArray_outS11ser;
  wire   [7:0] KeyArray_outS10ser;
  wire   [7:0] KeyArray_outS03ser;
  wire   [7:0] KeyArray_outS02ser;
  wire   [7:0] KeyArray_inS00ser;
  wire   [7:0] MixColumns_line0_S13;
  wire   [4:1] MixColumns_line0_S02;
  wire   [4:1] MixColumns_line0_timesTHREE_input2;
  wire   [7:0] MixColumns_line1_S13;
  wire   [7:0] MixColumns_line1_S02;
  wire   [4:1] MixColumns_line1_timesTHREE_input2;
  wire   [7:0] MixColumns_line2_S13;
  wire   [7:0] MixColumns_line2_S02;
  wire   [4:1] MixColumns_line2_timesTHREE_input2;
  wire   [7:0] MixColumns_line3_S13;
  wire   [7:0] MixColumns_line3_S02;

  NAND2_X1 U23 ( .A1(selSR), .A2(n2), .ZN(enKS) );
  INV_X1 U24 ( .A(start), .ZN(n2) );
  XOR2_X1 U25 ( .A(keyStateIn[0]), .B(port_out[0]), .Z(StateOutXORroundKey[0])
         );
  XOR2_X1 U26 ( .A(keyStateIn[1]), .B(port_out[1]), .Z(StateOutXORroundKey[1])
         );
  XOR2_X1 U27 ( .A(keyStateIn[2]), .B(port_out[2]), .Z(StateOutXORroundKey[2])
         );
  XOR2_X1 U28 ( .A(keyStateIn[3]), .B(port_out[3]), .Z(StateOutXORroundKey[3])
         );
  XOR2_X1 U29 ( .A(keyStateIn[4]), .B(port_out[4]), .Z(StateOutXORroundKey[4])
         );
  XOR2_X1 U30 ( .A(keyStateIn[5]), .B(port_out[5]), .Z(StateOutXORroundKey[5])
         );
  XOR2_X1 U31 ( .A(keyStateIn[6]), .B(port_out[6]), .Z(StateOutXORroundKey[6])
         );
  XOR2_X1 U32 ( .A(keyStateIn[7]), .B(port_out[7]), .Z(StateOutXORroundKey[7])
         );
  AND2_X1 U33 ( .A1(notFirst), .A2(selXOR), .ZN(intselXOR) );
  INV_X1 ctrl_U26 ( .A(ctrl_seq4Out_1_), .ZN(ctrl_n2) );
  NOR2_X1 ctrl_U25 ( .A1(ctrl_n24), .A2(ctrl_n7), .ZN(ctrl_nRstSeq4) );
  XNOR2_X1 ctrl_U24 ( .A(ctrl_seq6Out_4_), .B(ctrl_seq6In_1_), .ZN(ctrl_n22)
         );
  NAND2_X1 ctrl_U23 ( .A1(ctrl_n4), .A2(ctrl_n19), .ZN(ctrl_n21) );
  NAND2_X1 ctrl_U22 ( .A1(selXOR), .A2(ctrl_n5), .ZN(ctrl_n19) );
  NOR2_X1 ctrl_U21 ( .A1(ctrl_n7), .A2(ctrl_n18), .ZN(selXOR) );
  NOR2_X1 ctrl_U20 ( .A1(ctrl_seq4Out_1_), .A2(ctrl_seq4In_1_), .ZN(ctrl_n18)
         );
  OR2_X1 ctrl_U19 ( .A1(selSR), .A2(ctrl_n17), .ZN(ctrl_n20) );
  NOR2_X1 ctrl_U18 ( .A1(ctrl_n15), .A2(ctrl_n23), .ZN(ctrl_n17) );
  NAND2_X1 ctrl_U17 ( .A1(ctrl_n6), .A2(ctrl_n24), .ZN(ctrl_n14) );
  NOR2_X1 ctrl_U16 ( .A1(ctrl_seq4Out_1_), .A2(ctrl_n12), .ZN(ctrl_finalStep)
         );
  NAND2_X1 ctrl_U15 ( .A1(ctrl_n24), .A2(ctrl_seq4In_1_), .ZN(ctrl_n12) );
  NAND2_X1 ctrl_U14 ( .A1(ctrl_n10), .A2(ctrl_n9), .ZN(ctrl_n11) );
  NOR2_X1 ctrl_U13 ( .A1(ctrl_seq6In_3_), .A2(ctrl_seq6Out_4_), .ZN(ctrl_n9)
         );
  NOR2_X1 ctrl_U12 ( .A1(ctrl_seq6In_1_), .A2(ctrl_seq6In_4_), .ZN(ctrl_n10)
         );
  INV_X1 ctrl_U11 ( .A(n2), .ZN(ctrl_n7) );
  INV_X1 ctrl_U10 ( .A(ctrl_n7), .ZN(ctrl_n6) );
  NOR2_X1 ctrl_U9 ( .A1(ctrl_seq6In_2_), .A2(ctrl_n11), .ZN(ctrl_n24) );
  NAND2_X1 ctrl_U8 ( .A1(ctrl_n6), .A2(ctrl_n13), .ZN(ctrl_n23) );
  INV_X1 ctrl_U7 ( .A(ctrl_n23), .ZN(done) );
  AND2_X1 ctrl_U6 ( .A1(ctrl_finalStep), .A2(intFinal), .ZN(ctrl_n13) );
  OR2_X1 ctrl_U5 ( .A1(done), .A2(ctrl_n14), .ZN(ctrl_n4) );
  INV_X1 ctrl_U4 ( .A(ctrl_n4), .ZN(selSR) );
  NOR2_X2 ctrl_U3 ( .A1(ctrl_n16), .A2(ctrl_n7), .ZN(selMC) );
  NAND2_X1 ctrl_seq6_SFF_0_U3 ( .A1(ctrl_seq6_SFF_0_n2), .A2(
        ctrl_seq6_SFF_0_n1), .ZN(ctrl_seq6_SFF_0_n5) );
  OR2_X1 ctrl_seq6_SFF_0_U2 ( .A1(ctrl_n23), .A2(ctrl_seq6_SFF_0_n3), .ZN(
        ctrl_seq6_SFF_0_n1) );
  NAND2_X1 ctrl_seq6_SFF_0_U1 ( .A1(ctrl_seq6_SFF_0_QD), .A2(ctrl_n23), .ZN(
        ctrl_seq6_SFF_0_n2) );
  XOR2_X1 ctrl_seq6_SFF_0_MUXInst_XOR1_U1 ( .A(1'b1), .B(ctrl_n22), .Z(
        ctrl_seq6_SFF_0_MUXInst_X) );
  AND2_X1 ctrl_seq6_SFF_0_MUXInst_AND1_U1 ( .A1(ctrl_n6), .A2(
        ctrl_seq6_SFF_0_MUXInst_X), .ZN(ctrl_seq6_SFF_0_MUXInst_Y) );
  XOR2_X1 ctrl_seq6_SFF_0_MUXInst_XOR2_U1 ( .A(ctrl_seq6_SFF_0_MUXInst_Y), .B(
        1'b1), .Z(ctrl_seq6_SFF_0_QD) );
  INV_X1 ctrl_seq6_SFF_0_Q_reg_U1 ( .A(ctrl_seq6In_1_), .ZN(ctrl_seq6_SFF_0_n3) );
  DFF_X1 ctrl_seq6_SFF_0_Q_reg_FF_FF ( .D(ctrl_seq6_SFF_0_n5), .CK(clk), .Q(
        ctrl_seq6In_1_), .QN() );
  NAND2_X1 ctrl_seq6_SFF_1_U3 ( .A1(ctrl_seq6_SFF_1_n2), .A2(
        ctrl_seq6_SFF_1_n1), .ZN(ctrl_seq6_SFF_1_n5) );
  OR2_X1 ctrl_seq6_SFF_1_U2 ( .A1(ctrl_n23), .A2(ctrl_seq6_SFF_1_n10), .ZN(
        ctrl_seq6_SFF_1_n1) );
  NAND2_X1 ctrl_seq6_SFF_1_U1 ( .A1(ctrl_seq6_SFF_1_QD), .A2(ctrl_n23), .ZN(
        ctrl_seq6_SFF_1_n2) );
  XOR2_X1 ctrl_seq6_SFF_1_MUXInst_XOR1_U1 ( .A(1'b0), .B(ctrl_seq6In_1_), .Z(
        ctrl_seq6_SFF_1_MUXInst_X) );
  AND2_X1 ctrl_seq6_SFF_1_MUXInst_AND1_U1 ( .A1(ctrl_n6), .A2(
        ctrl_seq6_SFF_1_MUXInst_X), .ZN(ctrl_seq6_SFF_1_MUXInst_Y) );
  XOR2_X1 ctrl_seq6_SFF_1_MUXInst_XOR2_U1 ( .A(ctrl_seq6_SFF_1_MUXInst_Y), .B(
        1'b0), .Z(ctrl_seq6_SFF_1_QD) );
  INV_X1 ctrl_seq6_SFF_1_Q_reg_U1 ( .A(ctrl_seq6In_2_), .ZN(
        ctrl_seq6_SFF_1_n10) );
  DFF_X1 ctrl_seq6_SFF_1_Q_reg_FF_FF ( .D(ctrl_seq6_SFF_1_n5), .CK(clk), .Q(
        ctrl_seq6In_2_), .QN() );
  NAND2_X1 ctrl_seq6_SFF_2_U3 ( .A1(ctrl_seq6_SFF_2_n2), .A2(
        ctrl_seq6_SFF_2_n1), .ZN(ctrl_seq6_SFF_2_n5) );
  OR2_X1 ctrl_seq6_SFF_2_U2 ( .A1(ctrl_n23), .A2(ctrl_seq6_SFF_2_n10), .ZN(
        ctrl_seq6_SFF_2_n1) );
  NAND2_X1 ctrl_seq6_SFF_2_U1 ( .A1(ctrl_seq6_SFF_2_QD), .A2(ctrl_n23), .ZN(
        ctrl_seq6_SFF_2_n2) );
  XOR2_X1 ctrl_seq6_SFF_2_MUXInst_XOR1_U1 ( .A(1'b1), .B(ctrl_seq6In_2_), .Z(
        ctrl_seq6_SFF_2_MUXInst_X) );
  AND2_X1 ctrl_seq6_SFF_2_MUXInst_AND1_U1 ( .A1(ctrl_n6), .A2(
        ctrl_seq6_SFF_2_MUXInst_X), .ZN(ctrl_seq6_SFF_2_MUXInst_Y) );
  XOR2_X1 ctrl_seq6_SFF_2_MUXInst_XOR2_U1 ( .A(ctrl_seq6_SFF_2_MUXInst_Y), .B(
        1'b1), .Z(ctrl_seq6_SFF_2_QD) );
  INV_X1 ctrl_seq6_SFF_2_Q_reg_U1 ( .A(ctrl_seq6In_3_), .ZN(
        ctrl_seq6_SFF_2_n10) );
  DFF_X1 ctrl_seq6_SFF_2_Q_reg_FF_FF ( .D(ctrl_seq6_SFF_2_n5), .CK(clk), .Q(
        ctrl_seq6In_3_), .QN() );
  NAND2_X1 ctrl_seq6_SFF_3_U3 ( .A1(ctrl_seq6_SFF_3_n2), .A2(
        ctrl_seq6_SFF_3_n1), .ZN(ctrl_seq6_SFF_3_n5) );
  OR2_X1 ctrl_seq6_SFF_3_U2 ( .A1(ctrl_n23), .A2(ctrl_seq6_SFF_3_n10), .ZN(
        ctrl_seq6_SFF_3_n1) );
  NAND2_X1 ctrl_seq6_SFF_3_U1 ( .A1(ctrl_seq6_SFF_3_QD), .A2(ctrl_n23), .ZN(
        ctrl_seq6_SFF_3_n2) );
  XOR2_X1 ctrl_seq6_SFF_3_MUXInst_XOR1_U1 ( .A(1'b0), .B(ctrl_seq6In_3_), .Z(
        ctrl_seq6_SFF_3_MUXInst_X) );
  AND2_X1 ctrl_seq6_SFF_3_MUXInst_AND1_U1 ( .A1(ctrl_n6), .A2(
        ctrl_seq6_SFF_3_MUXInst_X), .ZN(ctrl_seq6_SFF_3_MUXInst_Y) );
  XOR2_X1 ctrl_seq6_SFF_3_MUXInst_XOR2_U1 ( .A(ctrl_seq6_SFF_3_MUXInst_Y), .B(
        1'b0), .Z(ctrl_seq6_SFF_3_QD) );
  INV_X1 ctrl_seq6_SFF_3_Q_reg_U1 ( .A(ctrl_seq6In_4_), .ZN(
        ctrl_seq6_SFF_3_n10) );
  DFF_X1 ctrl_seq6_SFF_3_Q_reg_FF_FF ( .D(ctrl_seq6_SFF_3_n5), .CK(clk), .Q(
        ctrl_seq6In_4_), .QN() );
  NAND2_X1 ctrl_seq6_SFF_4_U3 ( .A1(ctrl_seq6_SFF_4_n2), .A2(
        ctrl_seq6_SFF_4_n1), .ZN(ctrl_seq6_SFF_4_n5) );
  OR2_X1 ctrl_seq6_SFF_4_U2 ( .A1(ctrl_n23), .A2(ctrl_seq6_SFF_4_n10), .ZN(
        ctrl_seq6_SFF_4_n1) );
  NAND2_X1 ctrl_seq6_SFF_4_U1 ( .A1(ctrl_seq6_SFF_4_QD), .A2(ctrl_n23), .ZN(
        ctrl_seq6_SFF_4_n2) );
  XOR2_X1 ctrl_seq6_SFF_4_MUXInst_XOR1_U1 ( .A(1'b1), .B(ctrl_seq6In_4_), .Z(
        ctrl_seq6_SFF_4_MUXInst_X) );
  AND2_X1 ctrl_seq6_SFF_4_MUXInst_AND1_U1 ( .A1(ctrl_n6), .A2(
        ctrl_seq6_SFF_4_MUXInst_X), .ZN(ctrl_seq6_SFF_4_MUXInst_Y) );
  XOR2_X1 ctrl_seq6_SFF_4_MUXInst_XOR2_U1 ( .A(ctrl_seq6_SFF_4_MUXInst_Y), .B(
        1'b1), .Z(ctrl_seq6_SFF_4_QD) );
  INV_X1 ctrl_seq6_SFF_4_Q_reg_U1 ( .A(ctrl_seq6Out_4_), .ZN(
        ctrl_seq6_SFF_4_n10) );
  DFF_X1 ctrl_seq6_SFF_4_Q_reg_FF_FF ( .D(ctrl_seq6_SFF_4_n5), .CK(clk), .Q(
        ctrl_seq6Out_4_), .QN() );
  NAND2_X1 ctrl_seq4_SFF_0_U3 ( .A1(ctrl_seq4_SFF_0_n2), .A2(
        ctrl_seq4_SFF_0_n1), .ZN(ctrl_seq4_SFF_0_n5) );
  OR2_X1 ctrl_seq4_SFF_0_U2 ( .A1(ctrl_n23), .A2(ctrl_seq4_SFF_0_n10), .ZN(
        ctrl_seq4_SFF_0_n1) );
  NAND2_X1 ctrl_seq4_SFF_0_U1 ( .A1(ctrl_seq4_SFF_0_QD), .A2(ctrl_n23), .ZN(
        ctrl_seq4_SFF_0_n2) );
  XOR2_X1 ctrl_seq4_SFF_0_MUXInst_XOR1_U1 ( .A(1'b1), .B(ctrl_n2), .Z(
        ctrl_seq4_SFF_0_MUXInst_X) );
  AND2_X1 ctrl_seq4_SFF_0_MUXInst_AND1_U1 ( .A1(ctrl_nRstSeq4), .A2(
        ctrl_seq4_SFF_0_MUXInst_X), .ZN(ctrl_seq4_SFF_0_MUXInst_Y) );
  XOR2_X1 ctrl_seq4_SFF_0_MUXInst_XOR2_U1 ( .A(ctrl_seq4_SFF_0_MUXInst_Y), .B(
        1'b1), .Z(ctrl_seq4_SFF_0_QD) );
  INV_X1 ctrl_seq4_SFF_0_Q_reg_U1 ( .A(ctrl_seq4In_1_), .ZN(
        ctrl_seq4_SFF_0_n10) );
  DFF_X1 ctrl_seq4_SFF_0_Q_reg_FF_FF ( .D(ctrl_seq4_SFF_0_n5), .CK(clk), .Q(
        ctrl_seq4In_1_), .QN() );
  NAND2_X1 ctrl_seq4_SFF_1_U3 ( .A1(ctrl_seq4_SFF_1_n2), .A2(
        ctrl_seq4_SFF_1_n1), .ZN(ctrl_seq4_SFF_1_n5) );
  OR2_X1 ctrl_seq4_SFF_1_U2 ( .A1(ctrl_n23), .A2(ctrl_seq4_SFF_1_n10), .ZN(
        ctrl_seq4_SFF_1_n1) );
  NAND2_X1 ctrl_seq4_SFF_1_U1 ( .A1(ctrl_seq4_SFF_1_QD), .A2(ctrl_n23), .ZN(
        ctrl_seq4_SFF_1_n2) );
  XOR2_X1 ctrl_seq4_SFF_1_MUXInst_XOR1_U1 ( .A(1'b0), .B(ctrl_seq4In_1_), .Z(
        ctrl_seq4_SFF_1_MUXInst_X) );
  AND2_X1 ctrl_seq4_SFF_1_MUXInst_AND1_U1 ( .A1(ctrl_nRstSeq4), .A2(
        ctrl_seq4_SFF_1_MUXInst_X), .ZN(ctrl_seq4_SFF_1_MUXInst_Y) );
  XOR2_X1 ctrl_seq4_SFF_1_MUXInst_XOR2_U1 ( .A(ctrl_seq4_SFF_1_MUXInst_Y), .B(
        1'b0), .Z(ctrl_seq4_SFF_1_QD) );
  INV_X1 ctrl_seq4_SFF_1_Q_reg_U1 ( .A(ctrl_seq4Out_1_), .ZN(
        ctrl_seq4_SFF_1_n10) );
  DFF_X1 ctrl_seq4_SFF_1_Q_reg_FF_FF ( .D(ctrl_seq4_SFF_1_n5), .CK(clk), .Q(
        ctrl_seq4Out_1_), .QN() );
  INV_X1 ctrl_CSselMC_reg_U1 ( .A(ctrl_n5), .ZN(ctrl_n16) );
  DFF_X1 ctrl_CSselMC_reg_FF_FF ( .D(ctrl_n21), .CK(clk), .Q(ctrl_n5), .QN()
         );
  INV_X1 ctrl_CSenRC_reg_U1 ( .A(enRCon), .ZN(ctrl_n15) );
  DFF_X1 ctrl_CSenRC_reg_FF_FF ( .D(ctrl_n20), .CK(clk), .Q(enRCon), .QN() );
  XOR2_X1 MUX_StateIn_mux_inst_0_XOR1_U1 ( .A(SboxOut[0]), .B(
        StateOutXORroundKey[0]), .Z(MUX_StateIn_mux_inst_0_X) );
  AND2_X1 MUX_StateIn_mux_inst_0_AND1_U1 ( .A1(intFinal), .A2(
        MUX_StateIn_mux_inst_0_X), .ZN(MUX_StateIn_mux_inst_0_Y) );
  XOR2_X1 MUX_StateIn_mux_inst_0_XOR2_U1 ( .A(MUX_StateIn_mux_inst_0_Y), .B(
        SboxOut[0]), .Z(StateIn[0]) );
  XOR2_X1 MUX_StateIn_mux_inst_1_XOR1_U1 ( .A(SboxOut[1]), .B(
        StateOutXORroundKey[1]), .Z(MUX_StateIn_mux_inst_1_X) );
  AND2_X1 MUX_StateIn_mux_inst_1_AND1_U1 ( .A1(intFinal), .A2(
        MUX_StateIn_mux_inst_1_X), .ZN(MUX_StateIn_mux_inst_1_Y) );
  XOR2_X1 MUX_StateIn_mux_inst_1_XOR2_U1 ( .A(MUX_StateIn_mux_inst_1_Y), .B(
        SboxOut[1]), .Z(StateIn[1]) );
  XOR2_X1 MUX_StateIn_mux_inst_2_XOR1_U1 ( .A(SboxOut[2]), .B(
        StateOutXORroundKey[2]), .Z(MUX_StateIn_mux_inst_2_X) );
  AND2_X1 MUX_StateIn_mux_inst_2_AND1_U1 ( .A1(intFinal), .A2(
        MUX_StateIn_mux_inst_2_X), .ZN(MUX_StateIn_mux_inst_2_Y) );
  XOR2_X1 MUX_StateIn_mux_inst_2_XOR2_U1 ( .A(MUX_StateIn_mux_inst_2_Y), .B(
        SboxOut[2]), .Z(StateIn[2]) );
  XOR2_X1 MUX_StateIn_mux_inst_3_XOR1_U1 ( .A(SboxOut[3]), .B(
        StateOutXORroundKey[3]), .Z(MUX_StateIn_mux_inst_3_X) );
  AND2_X1 MUX_StateIn_mux_inst_3_AND1_U1 ( .A1(intFinal), .A2(
        MUX_StateIn_mux_inst_3_X), .ZN(MUX_StateIn_mux_inst_3_Y) );
  XOR2_X1 MUX_StateIn_mux_inst_3_XOR2_U1 ( .A(MUX_StateIn_mux_inst_3_Y), .B(
        SboxOut[3]), .Z(StateIn[3]) );
  XOR2_X1 MUX_StateIn_mux_inst_4_XOR1_U1 ( .A(SboxOut[4]), .B(
        StateOutXORroundKey[4]), .Z(MUX_StateIn_mux_inst_4_X) );
  AND2_X1 MUX_StateIn_mux_inst_4_AND1_U1 ( .A1(intFinal), .A2(
        MUX_StateIn_mux_inst_4_X), .ZN(MUX_StateIn_mux_inst_4_Y) );
  XOR2_X1 MUX_StateIn_mux_inst_4_XOR2_U1 ( .A(MUX_StateIn_mux_inst_4_Y), .B(
        SboxOut[4]), .Z(StateIn[4]) );
  XOR2_X1 MUX_StateIn_mux_inst_5_XOR1_U1 ( .A(SboxOut[5]), .B(
        StateOutXORroundKey[5]), .Z(MUX_StateIn_mux_inst_5_X) );
  AND2_X1 MUX_StateIn_mux_inst_5_AND1_U1 ( .A1(intFinal), .A2(
        MUX_StateIn_mux_inst_5_X), .ZN(MUX_StateIn_mux_inst_5_Y) );
  XOR2_X1 MUX_StateIn_mux_inst_5_XOR2_U1 ( .A(MUX_StateIn_mux_inst_5_Y), .B(
        SboxOut[5]), .Z(StateIn[5]) );
  XOR2_X1 MUX_StateIn_mux_inst_6_XOR1_U1 ( .A(SboxOut[6]), .B(
        StateOutXORroundKey[6]), .Z(MUX_StateIn_mux_inst_6_X) );
  AND2_X1 MUX_StateIn_mux_inst_6_AND1_U1 ( .A1(intFinal), .A2(
        MUX_StateIn_mux_inst_6_X), .ZN(MUX_StateIn_mux_inst_6_Y) );
  XOR2_X1 MUX_StateIn_mux_inst_6_XOR2_U1 ( .A(MUX_StateIn_mux_inst_6_Y), .B(
        SboxOut[6]), .Z(StateIn[6]) );
  XOR2_X1 MUX_StateIn_mux_inst_7_XOR1_U1 ( .A(SboxOut[7]), .B(
        StateOutXORroundKey[7]), .Z(MUX_StateIn_mux_inst_7_X) );
  AND2_X1 MUX_StateIn_mux_inst_7_AND1_U1 ( .A1(intFinal), .A2(
        MUX_StateIn_mux_inst_7_X), .ZN(MUX_StateIn_mux_inst_7_Y) );
  XOR2_X1 MUX_StateIn_mux_inst_7_XOR2_U1 ( .A(MUX_StateIn_mux_inst_7_Y), .B(
        SboxOut[7]), .Z(StateIn[7]) );
  INV_X2 stateArray_U4 ( .A(stateArray_n8), .ZN(stateArray_n6) );
  AND2_X1 stateArray_U3 ( .A1(n2), .A2(selMC), .ZN(stateArray_nReset_selMC) );
  INV_X2 stateArray_U2 ( .A(stateArray_n8), .ZN(stateArray_n7) );
  INV_X1 stateArray_U1 ( .A(selSR), .ZN(stateArray_n8) );
  XOR2_X1 stateArray_S00reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A(
        stateArray_outS01ser[0]), .B(port_out[0]), .Z(
        stateArray_S00reg_gff_1_SFF_0_MUXInst_X) );
  AND2_X1 stateArray_S00reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A1(stateArray_n7), 
        .A2(stateArray_S00reg_gff_1_SFF_0_MUXInst_X), .ZN(
        stateArray_S00reg_gff_1_SFF_0_MUXInst_Y) );
  XOR2_X1 stateArray_S00reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A(
        stateArray_S00reg_gff_1_SFF_0_MUXInst_Y), .B(stateArray_outS01ser[0]), 
        .Z(stateArray_S00reg_gff_1_SFF_0_QD) );
  INV_X1 stateArray_S00reg_gff_1_SFF_0_Q_reg_U1 ( .A(port_out[0]), .ZN(
        stateArray_S00reg_gff_1_SFF_0_Q_reg_QN) );
  DFF_X1 stateArray_S00reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        stateArray_S00reg_gff_1_SFF_0_QD), .CK(clk), .Q(port_out[0]), .QN() );
  XOR2_X1 stateArray_S00reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A(
        stateArray_outS01ser[1]), .B(port_out[1]), .Z(
        stateArray_S00reg_gff_1_SFF_1_MUXInst_X) );
  AND2_X1 stateArray_S00reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A1(stateArray_n7), 
        .A2(stateArray_S00reg_gff_1_SFF_1_MUXInst_X), .ZN(
        stateArray_S00reg_gff_1_SFF_1_MUXInst_Y) );
  XOR2_X1 stateArray_S00reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A(
        stateArray_S00reg_gff_1_SFF_1_MUXInst_Y), .B(stateArray_outS01ser[1]), 
        .Z(stateArray_S00reg_gff_1_SFF_1_QD) );
  INV_X1 stateArray_S00reg_gff_1_SFF_1_Q_reg_U1 ( .A(port_out[1]), .ZN(
        stateArray_S00reg_gff_1_SFF_1_Q_reg_QN) );
  DFF_X1 stateArray_S00reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        stateArray_S00reg_gff_1_SFF_1_QD), .CK(clk), .Q(port_out[1]), .QN() );
  XOR2_X1 stateArray_S00reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A(
        stateArray_outS01ser[2]), .B(port_out[2]), .Z(
        stateArray_S00reg_gff_1_SFF_2_MUXInst_X) );
  AND2_X1 stateArray_S00reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A1(stateArray_n7), 
        .A2(stateArray_S00reg_gff_1_SFF_2_MUXInst_X), .ZN(
        stateArray_S00reg_gff_1_SFF_2_MUXInst_Y) );
  XOR2_X1 stateArray_S00reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A(
        stateArray_S00reg_gff_1_SFF_2_MUXInst_Y), .B(stateArray_outS01ser[2]), 
        .Z(stateArray_S00reg_gff_1_SFF_2_QD) );
  INV_X1 stateArray_S00reg_gff_1_SFF_2_Q_reg_U1 ( .A(port_out[2]), .ZN(
        stateArray_S00reg_gff_1_SFF_2_Q_reg_QN) );
  DFF_X1 stateArray_S00reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        stateArray_S00reg_gff_1_SFF_2_QD), .CK(clk), .Q(port_out[2]), .QN() );
  XOR2_X1 stateArray_S00reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A(
        stateArray_outS01ser[3]), .B(port_out[3]), .Z(
        stateArray_S00reg_gff_1_SFF_3_MUXInst_X) );
  AND2_X1 stateArray_S00reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A1(stateArray_n7), 
        .A2(stateArray_S00reg_gff_1_SFF_3_MUXInst_X), .ZN(
        stateArray_S00reg_gff_1_SFF_3_MUXInst_Y) );
  XOR2_X1 stateArray_S00reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A(
        stateArray_S00reg_gff_1_SFF_3_MUXInst_Y), .B(stateArray_outS01ser[3]), 
        .Z(stateArray_S00reg_gff_1_SFF_3_QD) );
  INV_X1 stateArray_S00reg_gff_1_SFF_3_Q_reg_U1 ( .A(port_out[3]), .ZN(
        stateArray_S00reg_gff_1_SFF_3_Q_reg_QN) );
  DFF_X1 stateArray_S00reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        stateArray_S00reg_gff_1_SFF_3_QD), .CK(clk), .Q(port_out[3]), .QN() );
  XOR2_X1 stateArray_S00reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A(
        stateArray_outS01ser[4]), .B(port_out[4]), .Z(
        stateArray_S00reg_gff_1_SFF_4_MUXInst_X) );
  AND2_X1 stateArray_S00reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A1(stateArray_n7), 
        .A2(stateArray_S00reg_gff_1_SFF_4_MUXInst_X), .ZN(
        stateArray_S00reg_gff_1_SFF_4_MUXInst_Y) );
  XOR2_X1 stateArray_S00reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A(
        stateArray_S00reg_gff_1_SFF_4_MUXInst_Y), .B(stateArray_outS01ser[4]), 
        .Z(stateArray_S00reg_gff_1_SFF_4_QD) );
  INV_X1 stateArray_S00reg_gff_1_SFF_4_Q_reg_U1 ( .A(port_out[4]), .ZN(
        stateArray_S00reg_gff_1_SFF_4_Q_reg_QN) );
  DFF_X1 stateArray_S00reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        stateArray_S00reg_gff_1_SFF_4_QD), .CK(clk), .Q(port_out[4]), .QN() );
  XOR2_X1 stateArray_S00reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A(
        stateArray_outS01ser[5]), .B(port_out[5]), .Z(
        stateArray_S00reg_gff_1_SFF_5_MUXInst_X) );
  AND2_X1 stateArray_S00reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A1(stateArray_n7), 
        .A2(stateArray_S00reg_gff_1_SFF_5_MUXInst_X), .ZN(
        stateArray_S00reg_gff_1_SFF_5_MUXInst_Y) );
  XOR2_X1 stateArray_S00reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A(
        stateArray_S00reg_gff_1_SFF_5_MUXInst_Y), .B(stateArray_outS01ser[5]), 
        .Z(stateArray_S00reg_gff_1_SFF_5_QD) );
  INV_X1 stateArray_S00reg_gff_1_SFF_5_Q_reg_U1 ( .A(port_out[5]), .ZN(
        stateArray_S00reg_gff_1_SFF_5_Q_reg_QN) );
  DFF_X1 stateArray_S00reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        stateArray_S00reg_gff_1_SFF_5_QD), .CK(clk), .Q(port_out[5]), .QN() );
  XOR2_X1 stateArray_S00reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A(
        stateArray_outS01ser[6]), .B(port_out[6]), .Z(
        stateArray_S00reg_gff_1_SFF_6_MUXInst_X) );
  AND2_X1 stateArray_S00reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A1(stateArray_n7), 
        .A2(stateArray_S00reg_gff_1_SFF_6_MUXInst_X), .ZN(
        stateArray_S00reg_gff_1_SFF_6_MUXInst_Y) );
  XOR2_X1 stateArray_S00reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A(
        stateArray_S00reg_gff_1_SFF_6_MUXInst_Y), .B(stateArray_outS01ser[6]), 
        .Z(stateArray_S00reg_gff_1_SFF_6_QD) );
  INV_X1 stateArray_S00reg_gff_1_SFF_6_Q_reg_U1 ( .A(port_out[6]), .ZN(
        stateArray_S00reg_gff_1_SFF_6_Q_reg_QN) );
  DFF_X1 stateArray_S00reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        stateArray_S00reg_gff_1_SFF_6_QD), .CK(clk), .Q(port_out[6]), .QN() );
  XOR2_X1 stateArray_S00reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A(
        stateArray_outS01ser[7]), .B(port_out[7]), .Z(
        stateArray_S00reg_gff_1_SFF_7_MUXInst_X) );
  AND2_X1 stateArray_S00reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A1(stateArray_n7), 
        .A2(stateArray_S00reg_gff_1_SFF_7_MUXInst_X), .ZN(
        stateArray_S00reg_gff_1_SFF_7_MUXInst_Y) );
  XOR2_X1 stateArray_S00reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A(
        stateArray_S00reg_gff_1_SFF_7_MUXInst_Y), .B(stateArray_outS01ser[7]), 
        .Z(stateArray_S00reg_gff_1_SFF_7_QD) );
  INV_X1 stateArray_S00reg_gff_1_SFF_7_Q_reg_U1 ( .A(port_out[7]), .ZN(
        stateArray_S00reg_gff_1_SFF_7_Q_reg_QN) );
  DFF_X1 stateArray_S00reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        stateArray_S00reg_gff_1_SFF_7_QD), .CK(clk), .Q(port_out[7]), .QN() );
  XOR2_X1 stateArray_S01reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A(
        stateArray_outS02ser[0]), .B(stateArray_outS01ser[0]), .Z(
        stateArray_S01reg_gff_1_SFF_0_MUXInst_X) );
  AND2_X1 stateArray_S01reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A1(selSR), .A2(
        stateArray_S01reg_gff_1_SFF_0_MUXInst_X), .ZN(
        stateArray_S01reg_gff_1_SFF_0_MUXInst_Y) );
  XOR2_X1 stateArray_S01reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A(
        stateArray_S01reg_gff_1_SFF_0_MUXInst_Y), .B(stateArray_outS02ser[0]), 
        .Z(stateArray_S01reg_gff_1_SFF_0_QD) );
  INV_X1 stateArray_S01reg_gff_1_SFF_0_Q_reg_U1 ( .A(stateArray_outS01ser[0]), 
        .ZN(stateArray_S01reg_gff_1_SFF_0_Q_reg_QN) );
  DFF_X1 stateArray_S01reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        stateArray_S01reg_gff_1_SFF_0_QD), .CK(clk), .Q(
        stateArray_outS01ser[0]), .QN() );
  XOR2_X1 stateArray_S01reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A(
        stateArray_outS02ser[1]), .B(stateArray_outS01ser[1]), .Z(
        stateArray_S01reg_gff_1_SFF_1_MUXInst_X) );
  AND2_X1 stateArray_S01reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A1(selSR), .A2(
        stateArray_S01reg_gff_1_SFF_1_MUXInst_X), .ZN(
        stateArray_S01reg_gff_1_SFF_1_MUXInst_Y) );
  XOR2_X1 stateArray_S01reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A(
        stateArray_S01reg_gff_1_SFF_1_MUXInst_Y), .B(stateArray_outS02ser[1]), 
        .Z(stateArray_S01reg_gff_1_SFF_1_QD) );
  INV_X1 stateArray_S01reg_gff_1_SFF_1_Q_reg_U1 ( .A(stateArray_outS01ser[1]), 
        .ZN(stateArray_S01reg_gff_1_SFF_1_Q_reg_QN) );
  DFF_X1 stateArray_S01reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        stateArray_S01reg_gff_1_SFF_1_QD), .CK(clk), .Q(
        stateArray_outS01ser[1]), .QN() );
  XOR2_X1 stateArray_S01reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A(
        stateArray_outS02ser[2]), .B(stateArray_outS01ser[2]), .Z(
        stateArray_S01reg_gff_1_SFF_2_MUXInst_X) );
  AND2_X1 stateArray_S01reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A1(selSR), .A2(
        stateArray_S01reg_gff_1_SFF_2_MUXInst_X), .ZN(
        stateArray_S01reg_gff_1_SFF_2_MUXInst_Y) );
  XOR2_X1 stateArray_S01reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A(
        stateArray_S01reg_gff_1_SFF_2_MUXInst_Y), .B(stateArray_outS02ser[2]), 
        .Z(stateArray_S01reg_gff_1_SFF_2_QD) );
  INV_X1 stateArray_S01reg_gff_1_SFF_2_Q_reg_U1 ( .A(stateArray_outS01ser[2]), 
        .ZN(stateArray_S01reg_gff_1_SFF_2_Q_reg_QN) );
  DFF_X1 stateArray_S01reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        stateArray_S01reg_gff_1_SFF_2_QD), .CK(clk), .Q(
        stateArray_outS01ser[2]), .QN() );
  XOR2_X1 stateArray_S01reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A(
        stateArray_outS02ser[3]), .B(stateArray_outS01ser[3]), .Z(
        stateArray_S01reg_gff_1_SFF_3_MUXInst_X) );
  AND2_X1 stateArray_S01reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A1(selSR), .A2(
        stateArray_S01reg_gff_1_SFF_3_MUXInst_X), .ZN(
        stateArray_S01reg_gff_1_SFF_3_MUXInst_Y) );
  XOR2_X1 stateArray_S01reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A(
        stateArray_S01reg_gff_1_SFF_3_MUXInst_Y), .B(stateArray_outS02ser[3]), 
        .Z(stateArray_S01reg_gff_1_SFF_3_QD) );
  INV_X1 stateArray_S01reg_gff_1_SFF_3_Q_reg_U1 ( .A(stateArray_outS01ser[3]), 
        .ZN(stateArray_S01reg_gff_1_SFF_3_Q_reg_QN) );
  DFF_X1 stateArray_S01reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        stateArray_S01reg_gff_1_SFF_3_QD), .CK(clk), .Q(
        stateArray_outS01ser[3]), .QN() );
  XOR2_X1 stateArray_S01reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A(
        stateArray_outS02ser[4]), .B(stateArray_outS01ser[4]), .Z(
        stateArray_S01reg_gff_1_SFF_4_MUXInst_X) );
  AND2_X1 stateArray_S01reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A1(selSR), .A2(
        stateArray_S01reg_gff_1_SFF_4_MUXInst_X), .ZN(
        stateArray_S01reg_gff_1_SFF_4_MUXInst_Y) );
  XOR2_X1 stateArray_S01reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A(
        stateArray_S01reg_gff_1_SFF_4_MUXInst_Y), .B(stateArray_outS02ser[4]), 
        .Z(stateArray_S01reg_gff_1_SFF_4_QD) );
  INV_X1 stateArray_S01reg_gff_1_SFF_4_Q_reg_U1 ( .A(stateArray_outS01ser[4]), 
        .ZN(stateArray_S01reg_gff_1_SFF_4_Q_reg_QN) );
  DFF_X1 stateArray_S01reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        stateArray_S01reg_gff_1_SFF_4_QD), .CK(clk), .Q(
        stateArray_outS01ser[4]), .QN() );
  XOR2_X1 stateArray_S01reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A(
        stateArray_outS02ser[5]), .B(stateArray_outS01ser[5]), .Z(
        stateArray_S01reg_gff_1_SFF_5_MUXInst_X) );
  AND2_X1 stateArray_S01reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A1(selSR), .A2(
        stateArray_S01reg_gff_1_SFF_5_MUXInst_X), .ZN(
        stateArray_S01reg_gff_1_SFF_5_MUXInst_Y) );
  XOR2_X1 stateArray_S01reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A(
        stateArray_S01reg_gff_1_SFF_5_MUXInst_Y), .B(stateArray_outS02ser[5]), 
        .Z(stateArray_S01reg_gff_1_SFF_5_QD) );
  INV_X1 stateArray_S01reg_gff_1_SFF_5_Q_reg_U1 ( .A(stateArray_outS01ser[5]), 
        .ZN(stateArray_S01reg_gff_1_SFF_5_Q_reg_QN) );
  DFF_X1 stateArray_S01reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        stateArray_S01reg_gff_1_SFF_5_QD), .CK(clk), .Q(
        stateArray_outS01ser[5]), .QN() );
  XOR2_X1 stateArray_S01reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A(
        stateArray_outS02ser[6]), .B(stateArray_outS01ser[6]), .Z(
        stateArray_S01reg_gff_1_SFF_6_MUXInst_X) );
  AND2_X1 stateArray_S01reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A1(selSR), .A2(
        stateArray_S01reg_gff_1_SFF_6_MUXInst_X), .ZN(
        stateArray_S01reg_gff_1_SFF_6_MUXInst_Y) );
  XOR2_X1 stateArray_S01reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A(
        stateArray_S01reg_gff_1_SFF_6_MUXInst_Y), .B(stateArray_outS02ser[6]), 
        .Z(stateArray_S01reg_gff_1_SFF_6_QD) );
  INV_X1 stateArray_S01reg_gff_1_SFF_6_Q_reg_U1 ( .A(stateArray_outS01ser[6]), 
        .ZN(stateArray_S01reg_gff_1_SFF_6_Q_reg_QN) );
  DFF_X1 stateArray_S01reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        stateArray_S01reg_gff_1_SFF_6_QD), .CK(clk), .Q(
        stateArray_outS01ser[6]), .QN() );
  XOR2_X1 stateArray_S01reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A(
        stateArray_outS02ser[7]), .B(stateArray_outS01ser[7]), .Z(
        stateArray_S01reg_gff_1_SFF_7_MUXInst_X) );
  AND2_X1 stateArray_S01reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A1(selSR), .A2(
        stateArray_S01reg_gff_1_SFF_7_MUXInst_X), .ZN(
        stateArray_S01reg_gff_1_SFF_7_MUXInst_Y) );
  XOR2_X1 stateArray_S01reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A(
        stateArray_S01reg_gff_1_SFF_7_MUXInst_Y), .B(stateArray_outS02ser[7]), 
        .Z(stateArray_S01reg_gff_1_SFF_7_QD) );
  INV_X1 stateArray_S01reg_gff_1_SFF_7_Q_reg_U1 ( .A(stateArray_outS01ser[7]), 
        .ZN(stateArray_S01reg_gff_1_SFF_7_Q_reg_QN) );
  DFF_X1 stateArray_S01reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        stateArray_S01reg_gff_1_SFF_7_QD), .CK(clk), .Q(
        stateArray_outS01ser[7]), .QN() );
  XOR2_X1 stateArray_S02reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A(
        stateArray_outS03ser[0]), .B(stateArray_outS02ser[0]), .Z(
        stateArray_S02reg_gff_1_SFF_0_MUXInst_X) );
  AND2_X1 stateArray_S02reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A1(selSR), .A2(
        stateArray_S02reg_gff_1_SFF_0_MUXInst_X), .ZN(
        stateArray_S02reg_gff_1_SFF_0_MUXInst_Y) );
  XOR2_X1 stateArray_S02reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A(
        stateArray_S02reg_gff_1_SFF_0_MUXInst_Y), .B(stateArray_outS03ser[0]), 
        .Z(stateArray_S02reg_gff_1_SFF_0_QD) );
  INV_X1 stateArray_S02reg_gff_1_SFF_0_Q_reg_U1 ( .A(stateArray_outS02ser[0]), 
        .ZN(stateArray_S02reg_gff_1_SFF_0_Q_reg_QN) );
  DFF_X1 stateArray_S02reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        stateArray_S02reg_gff_1_SFF_0_QD), .CK(clk), .Q(
        stateArray_outS02ser[0]), .QN() );
  XOR2_X1 stateArray_S02reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A(
        stateArray_outS03ser[1]), .B(stateArray_outS02ser[1]), .Z(
        stateArray_S02reg_gff_1_SFF_1_MUXInst_X) );
  AND2_X1 stateArray_S02reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A1(selSR), .A2(
        stateArray_S02reg_gff_1_SFF_1_MUXInst_X), .ZN(
        stateArray_S02reg_gff_1_SFF_1_MUXInst_Y) );
  XOR2_X1 stateArray_S02reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A(
        stateArray_S02reg_gff_1_SFF_1_MUXInst_Y), .B(stateArray_outS03ser[1]), 
        .Z(stateArray_S02reg_gff_1_SFF_1_QD) );
  INV_X1 stateArray_S02reg_gff_1_SFF_1_Q_reg_U1 ( .A(stateArray_outS02ser[1]), 
        .ZN(stateArray_S02reg_gff_1_SFF_1_Q_reg_QN) );
  DFF_X1 stateArray_S02reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        stateArray_S02reg_gff_1_SFF_1_QD), .CK(clk), .Q(
        stateArray_outS02ser[1]), .QN() );
  XOR2_X1 stateArray_S02reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A(
        stateArray_outS03ser[2]), .B(stateArray_outS02ser[2]), .Z(
        stateArray_S02reg_gff_1_SFF_2_MUXInst_X) );
  AND2_X1 stateArray_S02reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A1(selSR), .A2(
        stateArray_S02reg_gff_1_SFF_2_MUXInst_X), .ZN(
        stateArray_S02reg_gff_1_SFF_2_MUXInst_Y) );
  XOR2_X1 stateArray_S02reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A(
        stateArray_S02reg_gff_1_SFF_2_MUXInst_Y), .B(stateArray_outS03ser[2]), 
        .Z(stateArray_S02reg_gff_1_SFF_2_QD) );
  INV_X1 stateArray_S02reg_gff_1_SFF_2_Q_reg_U1 ( .A(stateArray_outS02ser[2]), 
        .ZN(stateArray_S02reg_gff_1_SFF_2_Q_reg_QN) );
  DFF_X1 stateArray_S02reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        stateArray_S02reg_gff_1_SFF_2_QD), .CK(clk), .Q(
        stateArray_outS02ser[2]), .QN() );
  XOR2_X1 stateArray_S02reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A(
        stateArray_outS03ser[3]), .B(stateArray_outS02ser[3]), .Z(
        stateArray_S02reg_gff_1_SFF_3_MUXInst_X) );
  AND2_X1 stateArray_S02reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A1(selSR), .A2(
        stateArray_S02reg_gff_1_SFF_3_MUXInst_X), .ZN(
        stateArray_S02reg_gff_1_SFF_3_MUXInst_Y) );
  XOR2_X1 stateArray_S02reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A(
        stateArray_S02reg_gff_1_SFF_3_MUXInst_Y), .B(stateArray_outS03ser[3]), 
        .Z(stateArray_S02reg_gff_1_SFF_3_QD) );
  INV_X1 stateArray_S02reg_gff_1_SFF_3_Q_reg_U1 ( .A(stateArray_outS02ser[3]), 
        .ZN(stateArray_S02reg_gff_1_SFF_3_Q_reg_QN) );
  DFF_X1 stateArray_S02reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        stateArray_S02reg_gff_1_SFF_3_QD), .CK(clk), .Q(
        stateArray_outS02ser[3]), .QN() );
  XOR2_X1 stateArray_S02reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A(
        stateArray_outS03ser[4]), .B(stateArray_outS02ser[4]), .Z(
        stateArray_S02reg_gff_1_SFF_4_MUXInst_X) );
  AND2_X1 stateArray_S02reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A1(selSR), .A2(
        stateArray_S02reg_gff_1_SFF_4_MUXInst_X), .ZN(
        stateArray_S02reg_gff_1_SFF_4_MUXInst_Y) );
  XOR2_X1 stateArray_S02reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A(
        stateArray_S02reg_gff_1_SFF_4_MUXInst_Y), .B(stateArray_outS03ser[4]), 
        .Z(stateArray_S02reg_gff_1_SFF_4_QD) );
  INV_X1 stateArray_S02reg_gff_1_SFF_4_Q_reg_U1 ( .A(stateArray_outS02ser[4]), 
        .ZN(stateArray_S02reg_gff_1_SFF_4_Q_reg_QN) );
  DFF_X1 stateArray_S02reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        stateArray_S02reg_gff_1_SFF_4_QD), .CK(clk), .Q(
        stateArray_outS02ser[4]), .QN() );
  XOR2_X1 stateArray_S02reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A(
        stateArray_outS03ser[5]), .B(stateArray_outS02ser[5]), .Z(
        stateArray_S02reg_gff_1_SFF_5_MUXInst_X) );
  AND2_X1 stateArray_S02reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A1(selSR), .A2(
        stateArray_S02reg_gff_1_SFF_5_MUXInst_X), .ZN(
        stateArray_S02reg_gff_1_SFF_5_MUXInst_Y) );
  XOR2_X1 stateArray_S02reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A(
        stateArray_S02reg_gff_1_SFF_5_MUXInst_Y), .B(stateArray_outS03ser[5]), 
        .Z(stateArray_S02reg_gff_1_SFF_5_QD) );
  INV_X1 stateArray_S02reg_gff_1_SFF_5_Q_reg_U1 ( .A(stateArray_outS02ser[5]), 
        .ZN(stateArray_S02reg_gff_1_SFF_5_Q_reg_QN) );
  DFF_X1 stateArray_S02reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        stateArray_S02reg_gff_1_SFF_5_QD), .CK(clk), .Q(
        stateArray_outS02ser[5]), .QN() );
  XOR2_X1 stateArray_S02reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A(
        stateArray_outS03ser[6]), .B(stateArray_outS02ser[6]), .Z(
        stateArray_S02reg_gff_1_SFF_6_MUXInst_X) );
  AND2_X1 stateArray_S02reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A1(selSR), .A2(
        stateArray_S02reg_gff_1_SFF_6_MUXInst_X), .ZN(
        stateArray_S02reg_gff_1_SFF_6_MUXInst_Y) );
  XOR2_X1 stateArray_S02reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A(
        stateArray_S02reg_gff_1_SFF_6_MUXInst_Y), .B(stateArray_outS03ser[6]), 
        .Z(stateArray_S02reg_gff_1_SFF_6_QD) );
  INV_X1 stateArray_S02reg_gff_1_SFF_6_Q_reg_U1 ( .A(stateArray_outS02ser[6]), 
        .ZN(stateArray_S02reg_gff_1_SFF_6_Q_reg_QN) );
  DFF_X1 stateArray_S02reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        stateArray_S02reg_gff_1_SFF_6_QD), .CK(clk), .Q(
        stateArray_outS02ser[6]), .QN() );
  XOR2_X1 stateArray_S02reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A(
        stateArray_outS03ser[7]), .B(stateArray_outS02ser[7]), .Z(
        stateArray_S02reg_gff_1_SFF_7_MUXInst_X) );
  AND2_X1 stateArray_S02reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A1(selSR), .A2(
        stateArray_S02reg_gff_1_SFF_7_MUXInst_X), .ZN(
        stateArray_S02reg_gff_1_SFF_7_MUXInst_Y) );
  XOR2_X1 stateArray_S02reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A(
        stateArray_S02reg_gff_1_SFF_7_MUXInst_Y), .B(stateArray_outS03ser[7]), 
        .Z(stateArray_S02reg_gff_1_SFF_7_QD) );
  INV_X1 stateArray_S02reg_gff_1_SFF_7_Q_reg_U1 ( .A(stateArray_outS02ser[7]), 
        .ZN(stateArray_S02reg_gff_1_SFF_7_Q_reg_QN) );
  DFF_X1 stateArray_S02reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        stateArray_S02reg_gff_1_SFF_7_QD), .CK(clk), .Q(
        stateArray_outS02ser[7]), .QN() );
  XOR2_X1 stateArray_S03reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A(
        stateArray_inS03ser[0]), .B(stateArray_outS03ser[0]), .Z(
        stateArray_S03reg_gff_1_SFF_0_MUXInst_X) );
  AND2_X1 stateArray_S03reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A1(stateArray_n6), 
        .A2(stateArray_S03reg_gff_1_SFF_0_MUXInst_X), .ZN(
        stateArray_S03reg_gff_1_SFF_0_MUXInst_Y) );
  XOR2_X1 stateArray_S03reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A(
        stateArray_S03reg_gff_1_SFF_0_MUXInst_Y), .B(stateArray_inS03ser[0]), 
        .Z(stateArray_S03reg_gff_1_SFF_0_QD) );
  INV_X1 stateArray_S03reg_gff_1_SFF_0_Q_reg_U1 ( .A(stateArray_outS03ser[0]), 
        .ZN(stateArray_S03reg_gff_1_SFF_0_Q_reg_QN) );
  DFF_X1 stateArray_S03reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        stateArray_S03reg_gff_1_SFF_0_QD), .CK(clk), .Q(
        stateArray_outS03ser[0]), .QN() );
  XOR2_X1 stateArray_S03reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A(
        stateArray_inS03ser[1]), .B(stateArray_outS03ser[1]), .Z(
        stateArray_S03reg_gff_1_SFF_1_MUXInst_X) );
  AND2_X1 stateArray_S03reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A1(stateArray_n6), 
        .A2(stateArray_S03reg_gff_1_SFF_1_MUXInst_X), .ZN(
        stateArray_S03reg_gff_1_SFF_1_MUXInst_Y) );
  XOR2_X1 stateArray_S03reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A(
        stateArray_S03reg_gff_1_SFF_1_MUXInst_Y), .B(stateArray_inS03ser[1]), 
        .Z(stateArray_S03reg_gff_1_SFF_1_QD) );
  INV_X1 stateArray_S03reg_gff_1_SFF_1_Q_reg_U1 ( .A(stateArray_outS03ser[1]), 
        .ZN(stateArray_S03reg_gff_1_SFF_1_Q_reg_QN) );
  DFF_X1 stateArray_S03reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        stateArray_S03reg_gff_1_SFF_1_QD), .CK(clk), .Q(
        stateArray_outS03ser[1]), .QN() );
  XOR2_X1 stateArray_S03reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A(
        stateArray_inS03ser[2]), .B(stateArray_outS03ser[2]), .Z(
        stateArray_S03reg_gff_1_SFF_2_MUXInst_X) );
  AND2_X1 stateArray_S03reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A1(stateArray_n6), 
        .A2(stateArray_S03reg_gff_1_SFF_2_MUXInst_X), .ZN(
        stateArray_S03reg_gff_1_SFF_2_MUXInst_Y) );
  XOR2_X1 stateArray_S03reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A(
        stateArray_S03reg_gff_1_SFF_2_MUXInst_Y), .B(stateArray_inS03ser[2]), 
        .Z(stateArray_S03reg_gff_1_SFF_2_QD) );
  INV_X1 stateArray_S03reg_gff_1_SFF_2_Q_reg_U1 ( .A(stateArray_outS03ser[2]), 
        .ZN(stateArray_S03reg_gff_1_SFF_2_Q_reg_QN) );
  DFF_X1 stateArray_S03reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        stateArray_S03reg_gff_1_SFF_2_QD), .CK(clk), .Q(
        stateArray_outS03ser[2]), .QN() );
  XOR2_X1 stateArray_S03reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A(
        stateArray_inS03ser[3]), .B(stateArray_outS03ser[3]), .Z(
        stateArray_S03reg_gff_1_SFF_3_MUXInst_X) );
  AND2_X1 stateArray_S03reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A1(stateArray_n6), 
        .A2(stateArray_S03reg_gff_1_SFF_3_MUXInst_X), .ZN(
        stateArray_S03reg_gff_1_SFF_3_MUXInst_Y) );
  XOR2_X1 stateArray_S03reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A(
        stateArray_S03reg_gff_1_SFF_3_MUXInst_Y), .B(stateArray_inS03ser[3]), 
        .Z(stateArray_S03reg_gff_1_SFF_3_QD) );
  INV_X1 stateArray_S03reg_gff_1_SFF_3_Q_reg_U1 ( .A(stateArray_outS03ser[3]), 
        .ZN(stateArray_S03reg_gff_1_SFF_3_Q_reg_QN) );
  DFF_X1 stateArray_S03reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        stateArray_S03reg_gff_1_SFF_3_QD), .CK(clk), .Q(
        stateArray_outS03ser[3]), .QN() );
  XOR2_X1 stateArray_S03reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A(
        stateArray_inS03ser[4]), .B(stateArray_outS03ser[4]), .Z(
        stateArray_S03reg_gff_1_SFF_4_MUXInst_X) );
  AND2_X1 stateArray_S03reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A1(stateArray_n6), 
        .A2(stateArray_S03reg_gff_1_SFF_4_MUXInst_X), .ZN(
        stateArray_S03reg_gff_1_SFF_4_MUXInst_Y) );
  XOR2_X1 stateArray_S03reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A(
        stateArray_S03reg_gff_1_SFF_4_MUXInst_Y), .B(stateArray_inS03ser[4]), 
        .Z(stateArray_S03reg_gff_1_SFF_4_QD) );
  INV_X1 stateArray_S03reg_gff_1_SFF_4_Q_reg_U1 ( .A(stateArray_outS03ser[4]), 
        .ZN(stateArray_S03reg_gff_1_SFF_4_Q_reg_QN) );
  DFF_X1 stateArray_S03reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        stateArray_S03reg_gff_1_SFF_4_QD), .CK(clk), .Q(
        stateArray_outS03ser[4]), .QN() );
  XOR2_X1 stateArray_S03reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A(
        stateArray_inS03ser[5]), .B(stateArray_outS03ser[5]), .Z(
        stateArray_S03reg_gff_1_SFF_5_MUXInst_X) );
  AND2_X1 stateArray_S03reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A1(stateArray_n6), 
        .A2(stateArray_S03reg_gff_1_SFF_5_MUXInst_X), .ZN(
        stateArray_S03reg_gff_1_SFF_5_MUXInst_Y) );
  XOR2_X1 stateArray_S03reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A(
        stateArray_S03reg_gff_1_SFF_5_MUXInst_Y), .B(stateArray_inS03ser[5]), 
        .Z(stateArray_S03reg_gff_1_SFF_5_QD) );
  INV_X1 stateArray_S03reg_gff_1_SFF_5_Q_reg_U1 ( .A(stateArray_outS03ser[5]), 
        .ZN(stateArray_S03reg_gff_1_SFF_5_Q_reg_QN) );
  DFF_X1 stateArray_S03reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        stateArray_S03reg_gff_1_SFF_5_QD), .CK(clk), .Q(
        stateArray_outS03ser[5]), .QN() );
  XOR2_X1 stateArray_S03reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A(
        stateArray_inS03ser[6]), .B(stateArray_outS03ser[6]), .Z(
        stateArray_S03reg_gff_1_SFF_6_MUXInst_X) );
  AND2_X1 stateArray_S03reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A1(stateArray_n6), 
        .A2(stateArray_S03reg_gff_1_SFF_6_MUXInst_X), .ZN(
        stateArray_S03reg_gff_1_SFF_6_MUXInst_Y) );
  XOR2_X1 stateArray_S03reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A(
        stateArray_S03reg_gff_1_SFF_6_MUXInst_Y), .B(stateArray_inS03ser[6]), 
        .Z(stateArray_S03reg_gff_1_SFF_6_QD) );
  INV_X1 stateArray_S03reg_gff_1_SFF_6_Q_reg_U1 ( .A(stateArray_outS03ser[6]), 
        .ZN(stateArray_S03reg_gff_1_SFF_6_Q_reg_QN) );
  DFF_X1 stateArray_S03reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        stateArray_S03reg_gff_1_SFF_6_QD), .CK(clk), .Q(
        stateArray_outS03ser[6]), .QN() );
  XOR2_X1 stateArray_S03reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A(
        stateArray_inS03ser[7]), .B(stateArray_outS03ser[7]), .Z(
        stateArray_S03reg_gff_1_SFF_7_MUXInst_X) );
  AND2_X1 stateArray_S03reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A1(stateArray_n6), 
        .A2(stateArray_S03reg_gff_1_SFF_7_MUXInst_X), .ZN(
        stateArray_S03reg_gff_1_SFF_7_MUXInst_Y) );
  XOR2_X1 stateArray_S03reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A(
        stateArray_S03reg_gff_1_SFF_7_MUXInst_Y), .B(stateArray_inS03ser[7]), 
        .Z(stateArray_S03reg_gff_1_SFF_7_QD) );
  INV_X1 stateArray_S03reg_gff_1_SFF_7_Q_reg_U1 ( .A(stateArray_outS03ser[7]), 
        .ZN(stateArray_S03reg_gff_1_SFF_7_Q_reg_QN) );
  DFF_X1 stateArray_S03reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        stateArray_S03reg_gff_1_SFF_7_QD), .CK(clk), .Q(
        stateArray_outS03ser[7]), .QN() );
  XOR2_X1 stateArray_S10reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A(
        stateArray_outS11ser[0]), .B(stateArray_outS11ser[0]), .Z(
        stateArray_S10reg_gff_1_SFF_0_MUXInst_X) );
  AND2_X1 stateArray_S10reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A1(stateArray_n7), 
        .A2(stateArray_S10reg_gff_1_SFF_0_MUXInst_X), .ZN(
        stateArray_S10reg_gff_1_SFF_0_MUXInst_Y) );
  XOR2_X1 stateArray_S10reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A(
        stateArray_S10reg_gff_1_SFF_0_MUXInst_Y), .B(stateArray_outS11ser[0]), 
        .Z(stateArray_S10reg_gff_1_SFF_0_QD) );
  INV_X1 stateArray_S10reg_gff_1_SFF_0_Q_reg_U1 ( .A(MCin[16]), .ZN(
        stateArray_S10reg_gff_1_SFF_0_Q_reg_QN) );
  DFF_X1 stateArray_S10reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        stateArray_S10reg_gff_1_SFF_0_QD), .CK(clk), .Q(MCin[16]), .QN() );
  XOR2_X1 stateArray_S10reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A(
        stateArray_outS11ser[1]), .B(stateArray_outS11ser[1]), .Z(
        stateArray_S10reg_gff_1_SFF_1_MUXInst_X) );
  AND2_X1 stateArray_S10reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A1(stateArray_n7), 
        .A2(stateArray_S10reg_gff_1_SFF_1_MUXInst_X), .ZN(
        stateArray_S10reg_gff_1_SFF_1_MUXInst_Y) );
  XOR2_X1 stateArray_S10reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A(
        stateArray_S10reg_gff_1_SFF_1_MUXInst_Y), .B(stateArray_outS11ser[1]), 
        .Z(stateArray_S10reg_gff_1_SFF_1_QD) );
  INV_X1 stateArray_S10reg_gff_1_SFF_1_Q_reg_U1 ( .A(MixColumns_line1_S02[2]), 
        .ZN(stateArray_S10reg_gff_1_SFF_1_Q_reg_QN) );
  DFF_X1 stateArray_S10reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        stateArray_S10reg_gff_1_SFF_1_QD), .CK(clk), .Q(
        MixColumns_line1_S02[2]), .QN() );
  XOR2_X1 stateArray_S10reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A(
        stateArray_outS11ser[2]), .B(stateArray_outS11ser[2]), .Z(
        stateArray_S10reg_gff_1_SFF_2_MUXInst_X) );
  AND2_X1 stateArray_S10reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A1(stateArray_n7), 
        .A2(stateArray_S10reg_gff_1_SFF_2_MUXInst_X), .ZN(
        stateArray_S10reg_gff_1_SFF_2_MUXInst_Y) );
  XOR2_X1 stateArray_S10reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A(
        stateArray_S10reg_gff_1_SFF_2_MUXInst_Y), .B(stateArray_outS11ser[2]), 
        .Z(stateArray_S10reg_gff_1_SFF_2_QD) );
  INV_X1 stateArray_S10reg_gff_1_SFF_2_Q_reg_U1 ( .A(MCin[18]), .ZN(
        stateArray_S10reg_gff_1_SFF_2_Q_reg_QN) );
  DFF_X1 stateArray_S10reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        stateArray_S10reg_gff_1_SFF_2_QD), .CK(clk), .Q(MCin[18]), .QN() );
  XOR2_X1 stateArray_S10reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A(
        stateArray_outS11ser[3]), .B(stateArray_outS11ser[3]), .Z(
        stateArray_S10reg_gff_1_SFF_3_MUXInst_X) );
  AND2_X1 stateArray_S10reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A1(stateArray_n7), 
        .A2(stateArray_S10reg_gff_1_SFF_3_MUXInst_X), .ZN(
        stateArray_S10reg_gff_1_SFF_3_MUXInst_Y) );
  XOR2_X1 stateArray_S10reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A(
        stateArray_S10reg_gff_1_SFF_3_MUXInst_Y), .B(stateArray_outS11ser[3]), 
        .Z(stateArray_S10reg_gff_1_SFF_3_QD) );
  INV_X1 stateArray_S10reg_gff_1_SFF_3_Q_reg_U1 ( .A(MCin[19]), .ZN(
        stateArray_S10reg_gff_1_SFF_3_Q_reg_QN) );
  DFF_X1 stateArray_S10reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        stateArray_S10reg_gff_1_SFF_3_QD), .CK(clk), .Q(MCin[19]), .QN() );
  XOR2_X1 stateArray_S10reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A(
        stateArray_outS11ser[4]), .B(stateArray_outS11ser[4]), .Z(
        stateArray_S10reg_gff_1_SFF_4_MUXInst_X) );
  AND2_X1 stateArray_S10reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A1(stateArray_n7), 
        .A2(stateArray_S10reg_gff_1_SFF_4_MUXInst_X), .ZN(
        stateArray_S10reg_gff_1_SFF_4_MUXInst_Y) );
  XOR2_X1 stateArray_S10reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A(
        stateArray_S10reg_gff_1_SFF_4_MUXInst_Y), .B(stateArray_outS11ser[4]), 
        .Z(stateArray_S10reg_gff_1_SFF_4_QD) );
  INV_X1 stateArray_S10reg_gff_1_SFF_4_Q_reg_U1 ( .A(MixColumns_line1_S02[5]), 
        .ZN(stateArray_S10reg_gff_1_SFF_4_Q_reg_QN) );
  DFF_X1 stateArray_S10reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        stateArray_S10reg_gff_1_SFF_4_QD), .CK(clk), .Q(
        MixColumns_line1_S02[5]), .QN() );
  XOR2_X1 stateArray_S10reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A(
        stateArray_outS11ser[5]), .B(stateArray_outS11ser[5]), .Z(
        stateArray_S10reg_gff_1_SFF_5_MUXInst_X) );
  AND2_X1 stateArray_S10reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A1(stateArray_n7), 
        .A2(stateArray_S10reg_gff_1_SFF_5_MUXInst_X), .ZN(
        stateArray_S10reg_gff_1_SFF_5_MUXInst_Y) );
  XOR2_X1 stateArray_S10reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A(
        stateArray_S10reg_gff_1_SFF_5_MUXInst_Y), .B(stateArray_outS11ser[5]), 
        .Z(stateArray_S10reg_gff_1_SFF_5_QD) );
  INV_X1 stateArray_S10reg_gff_1_SFF_5_Q_reg_U1 ( .A(MixColumns_line1_S02[6]), 
        .ZN(stateArray_S10reg_gff_1_SFF_5_Q_reg_QN) );
  DFF_X1 stateArray_S10reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        stateArray_S10reg_gff_1_SFF_5_QD), .CK(clk), .Q(
        MixColumns_line1_S02[6]), .QN() );
  XOR2_X1 stateArray_S10reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A(
        stateArray_outS11ser[6]), .B(stateArray_outS11ser[6]), .Z(
        stateArray_S10reg_gff_1_SFF_6_MUXInst_X) );
  AND2_X1 stateArray_S10reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A1(stateArray_n7), 
        .A2(stateArray_S10reg_gff_1_SFF_6_MUXInst_X), .ZN(
        stateArray_S10reg_gff_1_SFF_6_MUXInst_Y) );
  XOR2_X1 stateArray_S10reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A(
        stateArray_S10reg_gff_1_SFF_6_MUXInst_Y), .B(stateArray_outS11ser[6]), 
        .Z(stateArray_S10reg_gff_1_SFF_6_QD) );
  INV_X1 stateArray_S10reg_gff_1_SFF_6_Q_reg_U1 ( .A(MixColumns_line1_S02[7]), 
        .ZN(stateArray_S10reg_gff_1_SFF_6_Q_reg_QN) );
  DFF_X1 stateArray_S10reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        stateArray_S10reg_gff_1_SFF_6_QD), .CK(clk), .Q(
        MixColumns_line1_S02[7]), .QN() );
  XOR2_X1 stateArray_S10reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A(
        stateArray_outS11ser[7]), .B(stateArray_outS11ser[7]), .Z(
        stateArray_S10reg_gff_1_SFF_7_MUXInst_X) );
  AND2_X1 stateArray_S10reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A1(stateArray_n7), 
        .A2(stateArray_S10reg_gff_1_SFF_7_MUXInst_X), .ZN(
        stateArray_S10reg_gff_1_SFF_7_MUXInst_Y) );
  XOR2_X1 stateArray_S10reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A(
        stateArray_S10reg_gff_1_SFF_7_MUXInst_Y), .B(stateArray_outS11ser[7]), 
        .Z(stateArray_S10reg_gff_1_SFF_7_QD) );
  INV_X1 stateArray_S10reg_gff_1_SFF_7_Q_reg_U1 ( .A(MixColumns_line1_S02[0]), 
        .ZN(stateArray_S10reg_gff_1_SFF_7_Q_reg_QN) );
  DFF_X1 stateArray_S10reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        stateArray_S10reg_gff_1_SFF_7_QD), .CK(clk), .Q(
        MixColumns_line1_S02[0]), .QN() );
  XOR2_X1 stateArray_S11reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A(
        stateArray_outS12ser[0]), .B(stateArray_outS12ser[0]), .Z(
        stateArray_S11reg_gff_1_SFF_0_MUXInst_X) );
  AND2_X1 stateArray_S11reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A1(stateArray_n7), 
        .A2(stateArray_S11reg_gff_1_SFF_0_MUXInst_X), .ZN(
        stateArray_S11reg_gff_1_SFF_0_MUXInst_Y) );
  XOR2_X1 stateArray_S11reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A(
        stateArray_S11reg_gff_1_SFF_0_MUXInst_Y), .B(stateArray_outS12ser[0]), 
        .Z(stateArray_S11reg_gff_1_SFF_0_QD) );
  INV_X1 stateArray_S11reg_gff_1_SFF_0_Q_reg_U1 ( .A(stateArray_outS11ser[0]), 
        .ZN(stateArray_S11reg_gff_1_SFF_0_Q_reg_QN) );
  DFF_X1 stateArray_S11reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        stateArray_S11reg_gff_1_SFF_0_QD), .CK(clk), .Q(
        stateArray_outS11ser[0]), .QN() );
  XOR2_X1 stateArray_S11reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A(
        stateArray_outS12ser[1]), .B(stateArray_outS12ser[1]), .Z(
        stateArray_S11reg_gff_1_SFF_1_MUXInst_X) );
  AND2_X1 stateArray_S11reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A1(stateArray_n7), 
        .A2(stateArray_S11reg_gff_1_SFF_1_MUXInst_X), .ZN(
        stateArray_S11reg_gff_1_SFF_1_MUXInst_Y) );
  XOR2_X1 stateArray_S11reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A(
        stateArray_S11reg_gff_1_SFF_1_MUXInst_Y), .B(stateArray_outS12ser[1]), 
        .Z(stateArray_S11reg_gff_1_SFF_1_QD) );
  INV_X1 stateArray_S11reg_gff_1_SFF_1_Q_reg_U1 ( .A(stateArray_outS11ser[1]), 
        .ZN(stateArray_S11reg_gff_1_SFF_1_Q_reg_QN) );
  DFF_X1 stateArray_S11reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        stateArray_S11reg_gff_1_SFF_1_QD), .CK(clk), .Q(
        stateArray_outS11ser[1]), .QN() );
  XOR2_X1 stateArray_S11reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A(
        stateArray_outS12ser[2]), .B(stateArray_outS12ser[2]), .Z(
        stateArray_S11reg_gff_1_SFF_2_MUXInst_X) );
  AND2_X1 stateArray_S11reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A1(stateArray_n7), 
        .A2(stateArray_S11reg_gff_1_SFF_2_MUXInst_X), .ZN(
        stateArray_S11reg_gff_1_SFF_2_MUXInst_Y) );
  XOR2_X1 stateArray_S11reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A(
        stateArray_S11reg_gff_1_SFF_2_MUXInst_Y), .B(stateArray_outS12ser[2]), 
        .Z(stateArray_S11reg_gff_1_SFF_2_QD) );
  INV_X1 stateArray_S11reg_gff_1_SFF_2_Q_reg_U1 ( .A(stateArray_outS11ser[2]), 
        .ZN(stateArray_S11reg_gff_1_SFF_2_Q_reg_QN) );
  DFF_X1 stateArray_S11reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        stateArray_S11reg_gff_1_SFF_2_QD), .CK(clk), .Q(
        stateArray_outS11ser[2]), .QN() );
  XOR2_X1 stateArray_S11reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A(
        stateArray_outS12ser[3]), .B(stateArray_outS12ser[3]), .Z(
        stateArray_S11reg_gff_1_SFF_3_MUXInst_X) );
  AND2_X1 stateArray_S11reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A1(stateArray_n7), 
        .A2(stateArray_S11reg_gff_1_SFF_3_MUXInst_X), .ZN(
        stateArray_S11reg_gff_1_SFF_3_MUXInst_Y) );
  XOR2_X1 stateArray_S11reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A(
        stateArray_S11reg_gff_1_SFF_3_MUXInst_Y), .B(stateArray_outS12ser[3]), 
        .Z(stateArray_S11reg_gff_1_SFF_3_QD) );
  INV_X1 stateArray_S11reg_gff_1_SFF_3_Q_reg_U1 ( .A(stateArray_outS11ser[3]), 
        .ZN(stateArray_S11reg_gff_1_SFF_3_Q_reg_QN) );
  DFF_X1 stateArray_S11reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        stateArray_S11reg_gff_1_SFF_3_QD), .CK(clk), .Q(
        stateArray_outS11ser[3]), .QN() );
  XOR2_X1 stateArray_S11reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A(
        stateArray_outS12ser[4]), .B(stateArray_outS12ser[4]), .Z(
        stateArray_S11reg_gff_1_SFF_4_MUXInst_X) );
  AND2_X1 stateArray_S11reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A1(stateArray_n7), 
        .A2(stateArray_S11reg_gff_1_SFF_4_MUXInst_X), .ZN(
        stateArray_S11reg_gff_1_SFF_4_MUXInst_Y) );
  XOR2_X1 stateArray_S11reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A(
        stateArray_S11reg_gff_1_SFF_4_MUXInst_Y), .B(stateArray_outS12ser[4]), 
        .Z(stateArray_S11reg_gff_1_SFF_4_QD) );
  INV_X1 stateArray_S11reg_gff_1_SFF_4_Q_reg_U1 ( .A(stateArray_outS11ser[4]), 
        .ZN(stateArray_S11reg_gff_1_SFF_4_Q_reg_QN) );
  DFF_X1 stateArray_S11reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        stateArray_S11reg_gff_1_SFF_4_QD), .CK(clk), .Q(
        stateArray_outS11ser[4]), .QN() );
  XOR2_X1 stateArray_S11reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A(
        stateArray_outS12ser[5]), .B(stateArray_outS12ser[5]), .Z(
        stateArray_S11reg_gff_1_SFF_5_MUXInst_X) );
  AND2_X1 stateArray_S11reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A1(stateArray_n7), 
        .A2(stateArray_S11reg_gff_1_SFF_5_MUXInst_X), .ZN(
        stateArray_S11reg_gff_1_SFF_5_MUXInst_Y) );
  XOR2_X1 stateArray_S11reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A(
        stateArray_S11reg_gff_1_SFF_5_MUXInst_Y), .B(stateArray_outS12ser[5]), 
        .Z(stateArray_S11reg_gff_1_SFF_5_QD) );
  INV_X1 stateArray_S11reg_gff_1_SFF_5_Q_reg_U1 ( .A(stateArray_outS11ser[5]), 
        .ZN(stateArray_S11reg_gff_1_SFF_5_Q_reg_QN) );
  DFF_X1 stateArray_S11reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        stateArray_S11reg_gff_1_SFF_5_QD), .CK(clk), .Q(
        stateArray_outS11ser[5]), .QN() );
  XOR2_X1 stateArray_S11reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A(
        stateArray_outS12ser[6]), .B(stateArray_outS12ser[6]), .Z(
        stateArray_S11reg_gff_1_SFF_6_MUXInst_X) );
  AND2_X1 stateArray_S11reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A1(stateArray_n7), 
        .A2(stateArray_S11reg_gff_1_SFF_6_MUXInst_X), .ZN(
        stateArray_S11reg_gff_1_SFF_6_MUXInst_Y) );
  XOR2_X1 stateArray_S11reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A(
        stateArray_S11reg_gff_1_SFF_6_MUXInst_Y), .B(stateArray_outS12ser[6]), 
        .Z(stateArray_S11reg_gff_1_SFF_6_QD) );
  INV_X1 stateArray_S11reg_gff_1_SFF_6_Q_reg_U1 ( .A(stateArray_outS11ser[6]), 
        .ZN(stateArray_S11reg_gff_1_SFF_6_Q_reg_QN) );
  DFF_X1 stateArray_S11reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        stateArray_S11reg_gff_1_SFF_6_QD), .CK(clk), .Q(
        stateArray_outS11ser[6]), .QN() );
  XOR2_X1 stateArray_S11reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A(
        stateArray_outS12ser[7]), .B(stateArray_outS12ser[7]), .Z(
        stateArray_S11reg_gff_1_SFF_7_MUXInst_X) );
  AND2_X1 stateArray_S11reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A1(stateArray_n7), 
        .A2(stateArray_S11reg_gff_1_SFF_7_MUXInst_X), .ZN(
        stateArray_S11reg_gff_1_SFF_7_MUXInst_Y) );
  XOR2_X1 stateArray_S11reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A(
        stateArray_S11reg_gff_1_SFF_7_MUXInst_Y), .B(stateArray_outS12ser[7]), 
        .Z(stateArray_S11reg_gff_1_SFF_7_QD) );
  INV_X1 stateArray_S11reg_gff_1_SFF_7_Q_reg_U1 ( .A(stateArray_outS11ser[7]), 
        .ZN(stateArray_S11reg_gff_1_SFF_7_Q_reg_QN) );
  DFF_X1 stateArray_S11reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        stateArray_S11reg_gff_1_SFF_7_QD), .CK(clk), .Q(
        stateArray_outS11ser[7]), .QN() );
  XOR2_X1 stateArray_S12reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A(
        stateArray_outS13ser[0]), .B(stateArray_outS13ser[0]), .Z(
        stateArray_S12reg_gff_1_SFF_0_MUXInst_X) );
  AND2_X1 stateArray_S12reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A1(stateArray_n7), 
        .A2(stateArray_S12reg_gff_1_SFF_0_MUXInst_X), .ZN(
        stateArray_S12reg_gff_1_SFF_0_MUXInst_Y) );
  XOR2_X1 stateArray_S12reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A(
        stateArray_S12reg_gff_1_SFF_0_MUXInst_Y), .B(stateArray_outS13ser[0]), 
        .Z(stateArray_S12reg_gff_1_SFF_0_QD) );
  INV_X1 stateArray_S12reg_gff_1_SFF_0_Q_reg_U1 ( .A(stateArray_outS12ser[0]), 
        .ZN(stateArray_S12reg_gff_1_SFF_0_Q_reg_QN) );
  DFF_X1 stateArray_S12reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        stateArray_S12reg_gff_1_SFF_0_QD), .CK(clk), .Q(
        stateArray_outS12ser[0]), .QN() );
  XOR2_X1 stateArray_S12reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A(
        stateArray_outS13ser[1]), .B(stateArray_outS13ser[1]), .Z(
        stateArray_S12reg_gff_1_SFF_1_MUXInst_X) );
  AND2_X1 stateArray_S12reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A1(stateArray_n7), 
        .A2(stateArray_S12reg_gff_1_SFF_1_MUXInst_X), .ZN(
        stateArray_S12reg_gff_1_SFF_1_MUXInst_Y) );
  XOR2_X1 stateArray_S12reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A(
        stateArray_S12reg_gff_1_SFF_1_MUXInst_Y), .B(stateArray_outS13ser[1]), 
        .Z(stateArray_S12reg_gff_1_SFF_1_QD) );
  INV_X1 stateArray_S12reg_gff_1_SFF_1_Q_reg_U1 ( .A(stateArray_outS12ser[1]), 
        .ZN(stateArray_S12reg_gff_1_SFF_1_Q_reg_QN) );
  DFF_X1 stateArray_S12reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        stateArray_S12reg_gff_1_SFF_1_QD), .CK(clk), .Q(
        stateArray_outS12ser[1]), .QN() );
  XOR2_X1 stateArray_S12reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A(
        stateArray_outS13ser[2]), .B(stateArray_outS13ser[2]), .Z(
        stateArray_S12reg_gff_1_SFF_2_MUXInst_X) );
  AND2_X1 stateArray_S12reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A1(stateArray_n7), 
        .A2(stateArray_S12reg_gff_1_SFF_2_MUXInst_X), .ZN(
        stateArray_S12reg_gff_1_SFF_2_MUXInst_Y) );
  XOR2_X1 stateArray_S12reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A(
        stateArray_S12reg_gff_1_SFF_2_MUXInst_Y), .B(stateArray_outS13ser[2]), 
        .Z(stateArray_S12reg_gff_1_SFF_2_QD) );
  INV_X1 stateArray_S12reg_gff_1_SFF_2_Q_reg_U1 ( .A(stateArray_outS12ser[2]), 
        .ZN(stateArray_S12reg_gff_1_SFF_2_Q_reg_QN) );
  DFF_X1 stateArray_S12reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        stateArray_S12reg_gff_1_SFF_2_QD), .CK(clk), .Q(
        stateArray_outS12ser[2]), .QN() );
  XOR2_X1 stateArray_S12reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A(
        stateArray_outS13ser[3]), .B(stateArray_outS13ser[3]), .Z(
        stateArray_S12reg_gff_1_SFF_3_MUXInst_X) );
  AND2_X1 stateArray_S12reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A1(stateArray_n7), 
        .A2(stateArray_S12reg_gff_1_SFF_3_MUXInst_X), .ZN(
        stateArray_S12reg_gff_1_SFF_3_MUXInst_Y) );
  XOR2_X1 stateArray_S12reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A(
        stateArray_S12reg_gff_1_SFF_3_MUXInst_Y), .B(stateArray_outS13ser[3]), 
        .Z(stateArray_S12reg_gff_1_SFF_3_QD) );
  INV_X1 stateArray_S12reg_gff_1_SFF_3_Q_reg_U1 ( .A(stateArray_outS12ser[3]), 
        .ZN(stateArray_S12reg_gff_1_SFF_3_Q_reg_QN) );
  DFF_X1 stateArray_S12reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        stateArray_S12reg_gff_1_SFF_3_QD), .CK(clk), .Q(
        stateArray_outS12ser[3]), .QN() );
  XOR2_X1 stateArray_S12reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A(
        stateArray_outS13ser[4]), .B(stateArray_outS13ser[4]), .Z(
        stateArray_S12reg_gff_1_SFF_4_MUXInst_X) );
  AND2_X1 stateArray_S12reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A1(stateArray_n7), 
        .A2(stateArray_S12reg_gff_1_SFF_4_MUXInst_X), .ZN(
        stateArray_S12reg_gff_1_SFF_4_MUXInst_Y) );
  XOR2_X1 stateArray_S12reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A(
        stateArray_S12reg_gff_1_SFF_4_MUXInst_Y), .B(stateArray_outS13ser[4]), 
        .Z(stateArray_S12reg_gff_1_SFF_4_QD) );
  INV_X1 stateArray_S12reg_gff_1_SFF_4_Q_reg_U1 ( .A(stateArray_outS12ser[4]), 
        .ZN(stateArray_S12reg_gff_1_SFF_4_Q_reg_QN) );
  DFF_X1 stateArray_S12reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        stateArray_S12reg_gff_1_SFF_4_QD), .CK(clk), .Q(
        stateArray_outS12ser[4]), .QN() );
  XOR2_X1 stateArray_S12reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A(
        stateArray_outS13ser[5]), .B(stateArray_outS13ser[5]), .Z(
        stateArray_S12reg_gff_1_SFF_5_MUXInst_X) );
  AND2_X1 stateArray_S12reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A1(stateArray_n7), 
        .A2(stateArray_S12reg_gff_1_SFF_5_MUXInst_X), .ZN(
        stateArray_S12reg_gff_1_SFF_5_MUXInst_Y) );
  XOR2_X1 stateArray_S12reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A(
        stateArray_S12reg_gff_1_SFF_5_MUXInst_Y), .B(stateArray_outS13ser[5]), 
        .Z(stateArray_S12reg_gff_1_SFF_5_QD) );
  INV_X1 stateArray_S12reg_gff_1_SFF_5_Q_reg_U1 ( .A(stateArray_outS12ser[5]), 
        .ZN(stateArray_S12reg_gff_1_SFF_5_Q_reg_QN) );
  DFF_X1 stateArray_S12reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        stateArray_S12reg_gff_1_SFF_5_QD), .CK(clk), .Q(
        stateArray_outS12ser[5]), .QN() );
  XOR2_X1 stateArray_S12reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A(
        stateArray_outS13ser[6]), .B(stateArray_outS13ser[6]), .Z(
        stateArray_S12reg_gff_1_SFF_6_MUXInst_X) );
  AND2_X1 stateArray_S12reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A1(stateArray_n7), 
        .A2(stateArray_S12reg_gff_1_SFF_6_MUXInst_X), .ZN(
        stateArray_S12reg_gff_1_SFF_6_MUXInst_Y) );
  XOR2_X1 stateArray_S12reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A(
        stateArray_S12reg_gff_1_SFF_6_MUXInst_Y), .B(stateArray_outS13ser[6]), 
        .Z(stateArray_S12reg_gff_1_SFF_6_QD) );
  INV_X1 stateArray_S12reg_gff_1_SFF_6_Q_reg_U1 ( .A(stateArray_outS12ser[6]), 
        .ZN(stateArray_S12reg_gff_1_SFF_6_Q_reg_QN) );
  DFF_X1 stateArray_S12reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        stateArray_S12reg_gff_1_SFF_6_QD), .CK(clk), .Q(
        stateArray_outS12ser[6]), .QN() );
  XOR2_X1 stateArray_S12reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A(
        stateArray_outS13ser[7]), .B(stateArray_outS13ser[7]), .Z(
        stateArray_S12reg_gff_1_SFF_7_MUXInst_X) );
  AND2_X1 stateArray_S12reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A1(stateArray_n7), 
        .A2(stateArray_S12reg_gff_1_SFF_7_MUXInst_X), .ZN(
        stateArray_S12reg_gff_1_SFF_7_MUXInst_Y) );
  XOR2_X1 stateArray_S12reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A(
        stateArray_S12reg_gff_1_SFF_7_MUXInst_Y), .B(stateArray_outS13ser[7]), 
        .Z(stateArray_S12reg_gff_1_SFF_7_QD) );
  INV_X1 stateArray_S12reg_gff_1_SFF_7_Q_reg_U1 ( .A(stateArray_outS12ser[7]), 
        .ZN(stateArray_S12reg_gff_1_SFF_7_Q_reg_QN) );
  DFF_X1 stateArray_S12reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        stateArray_S12reg_gff_1_SFF_7_QD), .CK(clk), .Q(
        stateArray_outS12ser[7]), .QN() );
  XOR2_X1 stateArray_S13reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A(
        stateArray_inS13ser[0]), .B(MCin[16]), .Z(
        stateArray_S13reg_gff_1_SFF_0_MUXInst_X) );
  AND2_X1 stateArray_S13reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A1(stateArray_n7), 
        .A2(stateArray_S13reg_gff_1_SFF_0_MUXInst_X), .ZN(
        stateArray_S13reg_gff_1_SFF_0_MUXInst_Y) );
  XOR2_X1 stateArray_S13reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A(
        stateArray_S13reg_gff_1_SFF_0_MUXInst_Y), .B(stateArray_inS13ser[0]), 
        .Z(stateArray_S13reg_gff_1_SFF_0_QD) );
  INV_X1 stateArray_S13reg_gff_1_SFF_0_Q_reg_U1 ( .A(stateArray_outS13ser[0]), 
        .ZN(stateArray_S13reg_gff_1_SFF_0_Q_reg_QN) );
  DFF_X1 stateArray_S13reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        stateArray_S13reg_gff_1_SFF_0_QD), .CK(clk), .Q(
        stateArray_outS13ser[0]), .QN() );
  XOR2_X1 stateArray_S13reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A(
        stateArray_inS13ser[1]), .B(MixColumns_line1_S02[2]), .Z(
        stateArray_S13reg_gff_1_SFF_1_MUXInst_X) );
  AND2_X1 stateArray_S13reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A1(stateArray_n7), 
        .A2(stateArray_S13reg_gff_1_SFF_1_MUXInst_X), .ZN(
        stateArray_S13reg_gff_1_SFF_1_MUXInst_Y) );
  XOR2_X1 stateArray_S13reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A(
        stateArray_S13reg_gff_1_SFF_1_MUXInst_Y), .B(stateArray_inS13ser[1]), 
        .Z(stateArray_S13reg_gff_1_SFF_1_QD) );
  INV_X1 stateArray_S13reg_gff_1_SFF_1_Q_reg_U1 ( .A(stateArray_outS13ser[1]), 
        .ZN(stateArray_S13reg_gff_1_SFF_1_Q_reg_QN) );
  DFF_X1 stateArray_S13reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        stateArray_S13reg_gff_1_SFF_1_QD), .CK(clk), .Q(
        stateArray_outS13ser[1]), .QN() );
  XOR2_X1 stateArray_S13reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A(
        stateArray_inS13ser[2]), .B(MCin[18]), .Z(
        stateArray_S13reg_gff_1_SFF_2_MUXInst_X) );
  AND2_X1 stateArray_S13reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A1(stateArray_n7), 
        .A2(stateArray_S13reg_gff_1_SFF_2_MUXInst_X), .ZN(
        stateArray_S13reg_gff_1_SFF_2_MUXInst_Y) );
  XOR2_X1 stateArray_S13reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A(
        stateArray_S13reg_gff_1_SFF_2_MUXInst_Y), .B(stateArray_inS13ser[2]), 
        .Z(stateArray_S13reg_gff_1_SFF_2_QD) );
  INV_X1 stateArray_S13reg_gff_1_SFF_2_Q_reg_U1 ( .A(stateArray_outS13ser[2]), 
        .ZN(stateArray_S13reg_gff_1_SFF_2_Q_reg_QN) );
  DFF_X1 stateArray_S13reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        stateArray_S13reg_gff_1_SFF_2_QD), .CK(clk), .Q(
        stateArray_outS13ser[2]), .QN() );
  XOR2_X1 stateArray_S13reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A(
        stateArray_inS13ser[3]), .B(MCin[19]), .Z(
        stateArray_S13reg_gff_1_SFF_3_MUXInst_X) );
  AND2_X1 stateArray_S13reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A1(stateArray_n7), 
        .A2(stateArray_S13reg_gff_1_SFF_3_MUXInst_X), .ZN(
        stateArray_S13reg_gff_1_SFF_3_MUXInst_Y) );
  XOR2_X1 stateArray_S13reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A(
        stateArray_S13reg_gff_1_SFF_3_MUXInst_Y), .B(stateArray_inS13ser[3]), 
        .Z(stateArray_S13reg_gff_1_SFF_3_QD) );
  INV_X1 stateArray_S13reg_gff_1_SFF_3_Q_reg_U1 ( .A(stateArray_outS13ser[3]), 
        .ZN(stateArray_S13reg_gff_1_SFF_3_Q_reg_QN) );
  DFF_X1 stateArray_S13reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        stateArray_S13reg_gff_1_SFF_3_QD), .CK(clk), .Q(
        stateArray_outS13ser[3]), .QN() );
  XOR2_X1 stateArray_S13reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A(
        stateArray_inS13ser[4]), .B(MixColumns_line1_S02[5]), .Z(
        stateArray_S13reg_gff_1_SFF_4_MUXInst_X) );
  AND2_X1 stateArray_S13reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A1(stateArray_n7), 
        .A2(stateArray_S13reg_gff_1_SFF_4_MUXInst_X), .ZN(
        stateArray_S13reg_gff_1_SFF_4_MUXInst_Y) );
  XOR2_X1 stateArray_S13reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A(
        stateArray_S13reg_gff_1_SFF_4_MUXInst_Y), .B(stateArray_inS13ser[4]), 
        .Z(stateArray_S13reg_gff_1_SFF_4_QD) );
  INV_X1 stateArray_S13reg_gff_1_SFF_4_Q_reg_U1 ( .A(stateArray_outS13ser[4]), 
        .ZN(stateArray_S13reg_gff_1_SFF_4_Q_reg_QN) );
  DFF_X1 stateArray_S13reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        stateArray_S13reg_gff_1_SFF_4_QD), .CK(clk), .Q(
        stateArray_outS13ser[4]), .QN() );
  XOR2_X1 stateArray_S13reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A(
        stateArray_inS13ser[5]), .B(MixColumns_line1_S02[6]), .Z(
        stateArray_S13reg_gff_1_SFF_5_MUXInst_X) );
  AND2_X1 stateArray_S13reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A1(stateArray_n7), 
        .A2(stateArray_S13reg_gff_1_SFF_5_MUXInst_X), .ZN(
        stateArray_S13reg_gff_1_SFF_5_MUXInst_Y) );
  XOR2_X1 stateArray_S13reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A(
        stateArray_S13reg_gff_1_SFF_5_MUXInst_Y), .B(stateArray_inS13ser[5]), 
        .Z(stateArray_S13reg_gff_1_SFF_5_QD) );
  INV_X1 stateArray_S13reg_gff_1_SFF_5_Q_reg_U1 ( .A(stateArray_outS13ser[5]), 
        .ZN(stateArray_S13reg_gff_1_SFF_5_Q_reg_QN) );
  DFF_X1 stateArray_S13reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        stateArray_S13reg_gff_1_SFF_5_QD), .CK(clk), .Q(
        stateArray_outS13ser[5]), .QN() );
  XOR2_X1 stateArray_S13reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A(
        stateArray_inS13ser[6]), .B(MixColumns_line1_S02[7]), .Z(
        stateArray_S13reg_gff_1_SFF_6_MUXInst_X) );
  AND2_X1 stateArray_S13reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A1(stateArray_n7), 
        .A2(stateArray_S13reg_gff_1_SFF_6_MUXInst_X), .ZN(
        stateArray_S13reg_gff_1_SFF_6_MUXInst_Y) );
  XOR2_X1 stateArray_S13reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A(
        stateArray_S13reg_gff_1_SFF_6_MUXInst_Y), .B(stateArray_inS13ser[6]), 
        .Z(stateArray_S13reg_gff_1_SFF_6_QD) );
  INV_X1 stateArray_S13reg_gff_1_SFF_6_Q_reg_U1 ( .A(stateArray_outS13ser[6]), 
        .ZN(stateArray_S13reg_gff_1_SFF_6_Q_reg_QN) );
  DFF_X1 stateArray_S13reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        stateArray_S13reg_gff_1_SFF_6_QD), .CK(clk), .Q(
        stateArray_outS13ser[6]), .QN() );
  XOR2_X1 stateArray_S13reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A(
        stateArray_inS13ser[7]), .B(MixColumns_line1_S02[0]), .Z(
        stateArray_S13reg_gff_1_SFF_7_MUXInst_X) );
  AND2_X1 stateArray_S13reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A1(stateArray_n7), 
        .A2(stateArray_S13reg_gff_1_SFF_7_MUXInst_X), .ZN(
        stateArray_S13reg_gff_1_SFF_7_MUXInst_Y) );
  XOR2_X1 stateArray_S13reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A(
        stateArray_S13reg_gff_1_SFF_7_MUXInst_Y), .B(stateArray_inS13ser[7]), 
        .Z(stateArray_S13reg_gff_1_SFF_7_QD) );
  INV_X1 stateArray_S13reg_gff_1_SFF_7_Q_reg_U1 ( .A(stateArray_outS13ser[7]), 
        .ZN(stateArray_S13reg_gff_1_SFF_7_Q_reg_QN) );
  DFF_X1 stateArray_S13reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        stateArray_S13reg_gff_1_SFF_7_QD), .CK(clk), .Q(
        stateArray_outS13ser[7]), .QN() );
  XOR2_X1 stateArray_S20reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A(
        stateArray_outS21ser[0]), .B(stateArray_outS22ser[0]), .Z(
        stateArray_S20reg_gff_1_SFF_0_MUXInst_X) );
  AND2_X1 stateArray_S20reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A1(stateArray_n7), 
        .A2(stateArray_S20reg_gff_1_SFF_0_MUXInst_X), .ZN(
        stateArray_S20reg_gff_1_SFF_0_MUXInst_Y) );
  XOR2_X1 stateArray_S20reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A(
        stateArray_S20reg_gff_1_SFF_0_MUXInst_Y), .B(stateArray_outS21ser[0]), 
        .Z(stateArray_S20reg_gff_1_SFF_0_QD) );
  INV_X1 stateArray_S20reg_gff_1_SFF_0_Q_reg_U1 ( .A(MCin[8]), .ZN(
        stateArray_S20reg_gff_1_SFF_0_Q_reg_QN) );
  DFF_X1 stateArray_S20reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        stateArray_S20reg_gff_1_SFF_0_QD), .CK(clk), .Q(MCin[8]), .QN() );
  XOR2_X1 stateArray_S20reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A(
        stateArray_outS21ser[1]), .B(stateArray_outS22ser[1]), .Z(
        stateArray_S20reg_gff_1_SFF_1_MUXInst_X) );
  AND2_X1 stateArray_S20reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A1(stateArray_n7), 
        .A2(stateArray_S20reg_gff_1_SFF_1_MUXInst_X), .ZN(
        stateArray_S20reg_gff_1_SFF_1_MUXInst_Y) );
  XOR2_X1 stateArray_S20reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A(
        stateArray_S20reg_gff_1_SFF_1_MUXInst_Y), .B(stateArray_outS21ser[1]), 
        .Z(stateArray_S20reg_gff_1_SFF_1_QD) );
  INV_X1 stateArray_S20reg_gff_1_SFF_1_Q_reg_U1 ( .A(MixColumns_line2_S02[2]), 
        .ZN(stateArray_S20reg_gff_1_SFF_1_Q_reg_QN) );
  DFF_X1 stateArray_S20reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        stateArray_S20reg_gff_1_SFF_1_QD), .CK(clk), .Q(
        MixColumns_line2_S02[2]), .QN() );
  XOR2_X1 stateArray_S20reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A(
        stateArray_outS21ser[2]), .B(stateArray_outS22ser[2]), .Z(
        stateArray_S20reg_gff_1_SFF_2_MUXInst_X) );
  AND2_X1 stateArray_S20reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A1(stateArray_n7), 
        .A2(stateArray_S20reg_gff_1_SFF_2_MUXInst_X), .ZN(
        stateArray_S20reg_gff_1_SFF_2_MUXInst_Y) );
  XOR2_X1 stateArray_S20reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A(
        stateArray_S20reg_gff_1_SFF_2_MUXInst_Y), .B(stateArray_outS21ser[2]), 
        .Z(stateArray_S20reg_gff_1_SFF_2_QD) );
  INV_X1 stateArray_S20reg_gff_1_SFF_2_Q_reg_U1 ( .A(MCin[10]), .ZN(
        stateArray_S20reg_gff_1_SFF_2_Q_reg_QN) );
  DFF_X1 stateArray_S20reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        stateArray_S20reg_gff_1_SFF_2_QD), .CK(clk), .Q(MCin[10]), .QN() );
  XOR2_X1 stateArray_S20reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A(
        stateArray_outS21ser[3]), .B(stateArray_outS22ser[3]), .Z(
        stateArray_S20reg_gff_1_SFF_3_MUXInst_X) );
  AND2_X1 stateArray_S20reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A1(stateArray_n7), 
        .A2(stateArray_S20reg_gff_1_SFF_3_MUXInst_X), .ZN(
        stateArray_S20reg_gff_1_SFF_3_MUXInst_Y) );
  XOR2_X1 stateArray_S20reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A(
        stateArray_S20reg_gff_1_SFF_3_MUXInst_Y), .B(stateArray_outS21ser[3]), 
        .Z(stateArray_S20reg_gff_1_SFF_3_QD) );
  INV_X1 stateArray_S20reg_gff_1_SFF_3_Q_reg_U1 ( .A(MCin[11]), .ZN(
        stateArray_S20reg_gff_1_SFF_3_Q_reg_QN) );
  DFF_X1 stateArray_S20reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        stateArray_S20reg_gff_1_SFF_3_QD), .CK(clk), .Q(MCin[11]), .QN() );
  XOR2_X1 stateArray_S20reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A(
        stateArray_outS21ser[4]), .B(stateArray_outS22ser[4]), .Z(
        stateArray_S20reg_gff_1_SFF_4_MUXInst_X) );
  AND2_X1 stateArray_S20reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A1(stateArray_n7), 
        .A2(stateArray_S20reg_gff_1_SFF_4_MUXInst_X), .ZN(
        stateArray_S20reg_gff_1_SFF_4_MUXInst_Y) );
  XOR2_X1 stateArray_S20reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A(
        stateArray_S20reg_gff_1_SFF_4_MUXInst_Y), .B(stateArray_outS21ser[4]), 
        .Z(stateArray_S20reg_gff_1_SFF_4_QD) );
  INV_X1 stateArray_S20reg_gff_1_SFF_4_Q_reg_U1 ( .A(MixColumns_line2_S02[5]), 
        .ZN(stateArray_S20reg_gff_1_SFF_4_Q_reg_QN) );
  DFF_X1 stateArray_S20reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        stateArray_S20reg_gff_1_SFF_4_QD), .CK(clk), .Q(
        MixColumns_line2_S02[5]), .QN() );
  XOR2_X1 stateArray_S20reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A(
        stateArray_outS21ser[5]), .B(stateArray_outS22ser[5]), .Z(
        stateArray_S20reg_gff_1_SFF_5_MUXInst_X) );
  AND2_X1 stateArray_S20reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A1(stateArray_n7), 
        .A2(stateArray_S20reg_gff_1_SFF_5_MUXInst_X), .ZN(
        stateArray_S20reg_gff_1_SFF_5_MUXInst_Y) );
  XOR2_X1 stateArray_S20reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A(
        stateArray_S20reg_gff_1_SFF_5_MUXInst_Y), .B(stateArray_outS21ser[5]), 
        .Z(stateArray_S20reg_gff_1_SFF_5_QD) );
  INV_X1 stateArray_S20reg_gff_1_SFF_5_Q_reg_U1 ( .A(MixColumns_line2_S02[6]), 
        .ZN(stateArray_S20reg_gff_1_SFF_5_Q_reg_QN) );
  DFF_X1 stateArray_S20reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        stateArray_S20reg_gff_1_SFF_5_QD), .CK(clk), .Q(
        MixColumns_line2_S02[6]), .QN() );
  XOR2_X1 stateArray_S20reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A(
        stateArray_outS21ser[6]), .B(stateArray_outS22ser[6]), .Z(
        stateArray_S20reg_gff_1_SFF_6_MUXInst_X) );
  AND2_X1 stateArray_S20reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A1(stateArray_n7), 
        .A2(stateArray_S20reg_gff_1_SFF_6_MUXInst_X), .ZN(
        stateArray_S20reg_gff_1_SFF_6_MUXInst_Y) );
  XOR2_X1 stateArray_S20reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A(
        stateArray_S20reg_gff_1_SFF_6_MUXInst_Y), .B(stateArray_outS21ser[6]), 
        .Z(stateArray_S20reg_gff_1_SFF_6_QD) );
  INV_X1 stateArray_S20reg_gff_1_SFF_6_Q_reg_U1 ( .A(MixColumns_line2_S02[7]), 
        .ZN(stateArray_S20reg_gff_1_SFF_6_Q_reg_QN) );
  DFF_X1 stateArray_S20reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        stateArray_S20reg_gff_1_SFF_6_QD), .CK(clk), .Q(
        MixColumns_line2_S02[7]), .QN() );
  XOR2_X1 stateArray_S20reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A(
        stateArray_outS21ser[7]), .B(stateArray_outS22ser[7]), .Z(
        stateArray_S20reg_gff_1_SFF_7_MUXInst_X) );
  AND2_X1 stateArray_S20reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A1(stateArray_n7), 
        .A2(stateArray_S20reg_gff_1_SFF_7_MUXInst_X), .ZN(
        stateArray_S20reg_gff_1_SFF_7_MUXInst_Y) );
  XOR2_X1 stateArray_S20reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A(
        stateArray_S20reg_gff_1_SFF_7_MUXInst_Y), .B(stateArray_outS21ser[7]), 
        .Z(stateArray_S20reg_gff_1_SFF_7_QD) );
  INV_X1 stateArray_S20reg_gff_1_SFF_7_Q_reg_U1 ( .A(MixColumns_line2_S02[0]), 
        .ZN(stateArray_S20reg_gff_1_SFF_7_Q_reg_QN) );
  DFF_X1 stateArray_S20reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        stateArray_S20reg_gff_1_SFF_7_QD), .CK(clk), .Q(
        MixColumns_line2_S02[0]), .QN() );
  XOR2_X1 stateArray_S21reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A(
        stateArray_outS22ser[0]), .B(stateArray_outS23ser[0]), .Z(
        stateArray_S21reg_gff_1_SFF_0_MUXInst_X) );
  AND2_X1 stateArray_S21reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A1(stateArray_n7), 
        .A2(stateArray_S21reg_gff_1_SFF_0_MUXInst_X), .ZN(
        stateArray_S21reg_gff_1_SFF_0_MUXInst_Y) );
  XOR2_X1 stateArray_S21reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A(
        stateArray_S21reg_gff_1_SFF_0_MUXInst_Y), .B(stateArray_outS22ser[0]), 
        .Z(stateArray_S21reg_gff_1_SFF_0_QD) );
  INV_X1 stateArray_S21reg_gff_1_SFF_0_Q_reg_U1 ( .A(stateArray_outS21ser[0]), 
        .ZN(stateArray_S21reg_gff_1_SFF_0_Q_reg_QN) );
  DFF_X1 stateArray_S21reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        stateArray_S21reg_gff_1_SFF_0_QD), .CK(clk), .Q(
        stateArray_outS21ser[0]), .QN() );
  XOR2_X1 stateArray_S21reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A(
        stateArray_outS22ser[1]), .B(stateArray_outS23ser[1]), .Z(
        stateArray_S21reg_gff_1_SFF_1_MUXInst_X) );
  AND2_X1 stateArray_S21reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A1(stateArray_n7), 
        .A2(stateArray_S21reg_gff_1_SFF_1_MUXInst_X), .ZN(
        stateArray_S21reg_gff_1_SFF_1_MUXInst_Y) );
  XOR2_X1 stateArray_S21reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A(
        stateArray_S21reg_gff_1_SFF_1_MUXInst_Y), .B(stateArray_outS22ser[1]), 
        .Z(stateArray_S21reg_gff_1_SFF_1_QD) );
  INV_X1 stateArray_S21reg_gff_1_SFF_1_Q_reg_U1 ( .A(stateArray_outS21ser[1]), 
        .ZN(stateArray_S21reg_gff_1_SFF_1_Q_reg_QN) );
  DFF_X1 stateArray_S21reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        stateArray_S21reg_gff_1_SFF_1_QD), .CK(clk), .Q(
        stateArray_outS21ser[1]), .QN() );
  XOR2_X1 stateArray_S21reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A(
        stateArray_outS22ser[2]), .B(stateArray_outS23ser[2]), .Z(
        stateArray_S21reg_gff_1_SFF_2_MUXInst_X) );
  AND2_X1 stateArray_S21reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A1(stateArray_n7), 
        .A2(stateArray_S21reg_gff_1_SFF_2_MUXInst_X), .ZN(
        stateArray_S21reg_gff_1_SFF_2_MUXInst_Y) );
  XOR2_X1 stateArray_S21reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A(
        stateArray_S21reg_gff_1_SFF_2_MUXInst_Y), .B(stateArray_outS22ser[2]), 
        .Z(stateArray_S21reg_gff_1_SFF_2_QD) );
  INV_X1 stateArray_S21reg_gff_1_SFF_2_Q_reg_U1 ( .A(stateArray_outS21ser[2]), 
        .ZN(stateArray_S21reg_gff_1_SFF_2_Q_reg_QN) );
  DFF_X1 stateArray_S21reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        stateArray_S21reg_gff_1_SFF_2_QD), .CK(clk), .Q(
        stateArray_outS21ser[2]), .QN() );
  XOR2_X1 stateArray_S21reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A(
        stateArray_outS22ser[3]), .B(stateArray_outS23ser[3]), .Z(
        stateArray_S21reg_gff_1_SFF_3_MUXInst_X) );
  AND2_X1 stateArray_S21reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A1(stateArray_n7), 
        .A2(stateArray_S21reg_gff_1_SFF_3_MUXInst_X), .ZN(
        stateArray_S21reg_gff_1_SFF_3_MUXInst_Y) );
  XOR2_X1 stateArray_S21reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A(
        stateArray_S21reg_gff_1_SFF_3_MUXInst_Y), .B(stateArray_outS22ser[3]), 
        .Z(stateArray_S21reg_gff_1_SFF_3_QD) );
  INV_X1 stateArray_S21reg_gff_1_SFF_3_Q_reg_U1 ( .A(stateArray_outS21ser[3]), 
        .ZN(stateArray_S21reg_gff_1_SFF_3_Q_reg_QN) );
  DFF_X1 stateArray_S21reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        stateArray_S21reg_gff_1_SFF_3_QD), .CK(clk), .Q(
        stateArray_outS21ser[3]), .QN() );
  XOR2_X1 stateArray_S21reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A(
        stateArray_outS22ser[4]), .B(stateArray_outS23ser[4]), .Z(
        stateArray_S21reg_gff_1_SFF_4_MUXInst_X) );
  AND2_X1 stateArray_S21reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A1(stateArray_n7), 
        .A2(stateArray_S21reg_gff_1_SFF_4_MUXInst_X), .ZN(
        stateArray_S21reg_gff_1_SFF_4_MUXInst_Y) );
  XOR2_X1 stateArray_S21reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A(
        stateArray_S21reg_gff_1_SFF_4_MUXInst_Y), .B(stateArray_outS22ser[4]), 
        .Z(stateArray_S21reg_gff_1_SFF_4_QD) );
  INV_X1 stateArray_S21reg_gff_1_SFF_4_Q_reg_U1 ( .A(stateArray_outS21ser[4]), 
        .ZN(stateArray_S21reg_gff_1_SFF_4_Q_reg_QN) );
  DFF_X1 stateArray_S21reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        stateArray_S21reg_gff_1_SFF_4_QD), .CK(clk), .Q(
        stateArray_outS21ser[4]), .QN() );
  XOR2_X1 stateArray_S21reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A(
        stateArray_outS22ser[5]), .B(stateArray_outS23ser[5]), .Z(
        stateArray_S21reg_gff_1_SFF_5_MUXInst_X) );
  AND2_X1 stateArray_S21reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A1(stateArray_n7), 
        .A2(stateArray_S21reg_gff_1_SFF_5_MUXInst_X), .ZN(
        stateArray_S21reg_gff_1_SFF_5_MUXInst_Y) );
  XOR2_X1 stateArray_S21reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A(
        stateArray_S21reg_gff_1_SFF_5_MUXInst_Y), .B(stateArray_outS22ser[5]), 
        .Z(stateArray_S21reg_gff_1_SFF_5_QD) );
  INV_X1 stateArray_S21reg_gff_1_SFF_5_Q_reg_U1 ( .A(stateArray_outS21ser[5]), 
        .ZN(stateArray_S21reg_gff_1_SFF_5_Q_reg_QN) );
  DFF_X1 stateArray_S21reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        stateArray_S21reg_gff_1_SFF_5_QD), .CK(clk), .Q(
        stateArray_outS21ser[5]), .QN() );
  XOR2_X1 stateArray_S21reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A(
        stateArray_outS22ser[6]), .B(stateArray_outS23ser[6]), .Z(
        stateArray_S21reg_gff_1_SFF_6_MUXInst_X) );
  AND2_X1 stateArray_S21reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A1(stateArray_n7), 
        .A2(stateArray_S21reg_gff_1_SFF_6_MUXInst_X), .ZN(
        stateArray_S21reg_gff_1_SFF_6_MUXInst_Y) );
  XOR2_X1 stateArray_S21reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A(
        stateArray_S21reg_gff_1_SFF_6_MUXInst_Y), .B(stateArray_outS22ser[6]), 
        .Z(stateArray_S21reg_gff_1_SFF_6_QD) );
  INV_X1 stateArray_S21reg_gff_1_SFF_6_Q_reg_U1 ( .A(stateArray_outS21ser[6]), 
        .ZN(stateArray_S21reg_gff_1_SFF_6_Q_reg_QN) );
  DFF_X1 stateArray_S21reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        stateArray_S21reg_gff_1_SFF_6_QD), .CK(clk), .Q(
        stateArray_outS21ser[6]), .QN() );
  XOR2_X1 stateArray_S21reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A(
        stateArray_outS22ser[7]), .B(stateArray_outS23ser[7]), .Z(
        stateArray_S21reg_gff_1_SFF_7_MUXInst_X) );
  AND2_X1 stateArray_S21reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A1(stateArray_n7), 
        .A2(stateArray_S21reg_gff_1_SFF_7_MUXInst_X), .ZN(
        stateArray_S21reg_gff_1_SFF_7_MUXInst_Y) );
  XOR2_X1 stateArray_S21reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A(
        stateArray_S21reg_gff_1_SFF_7_MUXInst_Y), .B(stateArray_outS22ser[7]), 
        .Z(stateArray_S21reg_gff_1_SFF_7_QD) );
  INV_X1 stateArray_S21reg_gff_1_SFF_7_Q_reg_U1 ( .A(stateArray_outS21ser[7]), 
        .ZN(stateArray_S21reg_gff_1_SFF_7_Q_reg_QN) );
  DFF_X1 stateArray_S21reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        stateArray_S21reg_gff_1_SFF_7_QD), .CK(clk), .Q(
        stateArray_outS21ser[7]), .QN() );
  XOR2_X1 stateArray_S22reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A(
        stateArray_outS23ser[0]), .B(MCin[8]), .Z(
        stateArray_S22reg_gff_1_SFF_0_MUXInst_X) );
  AND2_X1 stateArray_S22reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A1(stateArray_n6), 
        .A2(stateArray_S22reg_gff_1_SFF_0_MUXInst_X), .ZN(
        stateArray_S22reg_gff_1_SFF_0_MUXInst_Y) );
  XOR2_X1 stateArray_S22reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A(
        stateArray_S22reg_gff_1_SFF_0_MUXInst_Y), .B(stateArray_outS23ser[0]), 
        .Z(stateArray_S22reg_gff_1_SFF_0_QD) );
  INV_X1 stateArray_S22reg_gff_1_SFF_0_Q_reg_U1 ( .A(stateArray_outS22ser[0]), 
        .ZN(stateArray_S22reg_gff_1_SFF_0_Q_reg_QN) );
  DFF_X1 stateArray_S22reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        stateArray_S22reg_gff_1_SFF_0_QD), .CK(clk), .Q(
        stateArray_outS22ser[0]), .QN() );
  XOR2_X1 stateArray_S22reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A(
        stateArray_outS23ser[1]), .B(MixColumns_line2_S02[2]), .Z(
        stateArray_S22reg_gff_1_SFF_1_MUXInst_X) );
  AND2_X1 stateArray_S22reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A1(stateArray_n6), 
        .A2(stateArray_S22reg_gff_1_SFF_1_MUXInst_X), .ZN(
        stateArray_S22reg_gff_1_SFF_1_MUXInst_Y) );
  XOR2_X1 stateArray_S22reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A(
        stateArray_S22reg_gff_1_SFF_1_MUXInst_Y), .B(stateArray_outS23ser[1]), 
        .Z(stateArray_S22reg_gff_1_SFF_1_QD) );
  INV_X1 stateArray_S22reg_gff_1_SFF_1_Q_reg_U1 ( .A(stateArray_outS22ser[1]), 
        .ZN(stateArray_S22reg_gff_1_SFF_1_Q_reg_QN) );
  DFF_X1 stateArray_S22reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        stateArray_S22reg_gff_1_SFF_1_QD), .CK(clk), .Q(
        stateArray_outS22ser[1]), .QN() );
  XOR2_X1 stateArray_S22reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A(
        stateArray_outS23ser[2]), .B(MCin[10]), .Z(
        stateArray_S22reg_gff_1_SFF_2_MUXInst_X) );
  AND2_X1 stateArray_S22reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A1(stateArray_n6), 
        .A2(stateArray_S22reg_gff_1_SFF_2_MUXInst_X), .ZN(
        stateArray_S22reg_gff_1_SFF_2_MUXInst_Y) );
  XOR2_X1 stateArray_S22reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A(
        stateArray_S22reg_gff_1_SFF_2_MUXInst_Y), .B(stateArray_outS23ser[2]), 
        .Z(stateArray_S22reg_gff_1_SFF_2_QD) );
  INV_X1 stateArray_S22reg_gff_1_SFF_2_Q_reg_U1 ( .A(stateArray_outS22ser[2]), 
        .ZN(stateArray_S22reg_gff_1_SFF_2_Q_reg_QN) );
  DFF_X1 stateArray_S22reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        stateArray_S22reg_gff_1_SFF_2_QD), .CK(clk), .Q(
        stateArray_outS22ser[2]), .QN() );
  XOR2_X1 stateArray_S22reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A(
        stateArray_outS23ser[3]), .B(MCin[11]), .Z(
        stateArray_S22reg_gff_1_SFF_3_MUXInst_X) );
  AND2_X1 stateArray_S22reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A1(stateArray_n6), 
        .A2(stateArray_S22reg_gff_1_SFF_3_MUXInst_X), .ZN(
        stateArray_S22reg_gff_1_SFF_3_MUXInst_Y) );
  XOR2_X1 stateArray_S22reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A(
        stateArray_S22reg_gff_1_SFF_3_MUXInst_Y), .B(stateArray_outS23ser[3]), 
        .Z(stateArray_S22reg_gff_1_SFF_3_QD) );
  INV_X1 stateArray_S22reg_gff_1_SFF_3_Q_reg_U1 ( .A(stateArray_outS22ser[3]), 
        .ZN(stateArray_S22reg_gff_1_SFF_3_Q_reg_QN) );
  DFF_X1 stateArray_S22reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        stateArray_S22reg_gff_1_SFF_3_QD), .CK(clk), .Q(
        stateArray_outS22ser[3]), .QN() );
  XOR2_X1 stateArray_S22reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A(
        stateArray_outS23ser[4]), .B(MixColumns_line2_S02[5]), .Z(
        stateArray_S22reg_gff_1_SFF_4_MUXInst_X) );
  AND2_X1 stateArray_S22reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A1(stateArray_n6), 
        .A2(stateArray_S22reg_gff_1_SFF_4_MUXInst_X), .ZN(
        stateArray_S22reg_gff_1_SFF_4_MUXInst_Y) );
  XOR2_X1 stateArray_S22reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A(
        stateArray_S22reg_gff_1_SFF_4_MUXInst_Y), .B(stateArray_outS23ser[4]), 
        .Z(stateArray_S22reg_gff_1_SFF_4_QD) );
  INV_X1 stateArray_S22reg_gff_1_SFF_4_Q_reg_U1 ( .A(stateArray_outS22ser[4]), 
        .ZN(stateArray_S22reg_gff_1_SFF_4_Q_reg_QN) );
  DFF_X1 stateArray_S22reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        stateArray_S22reg_gff_1_SFF_4_QD), .CK(clk), .Q(
        stateArray_outS22ser[4]), .QN() );
  XOR2_X1 stateArray_S22reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A(
        stateArray_outS23ser[5]), .B(MixColumns_line2_S02[6]), .Z(
        stateArray_S22reg_gff_1_SFF_5_MUXInst_X) );
  AND2_X1 stateArray_S22reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A1(stateArray_n6), 
        .A2(stateArray_S22reg_gff_1_SFF_5_MUXInst_X), .ZN(
        stateArray_S22reg_gff_1_SFF_5_MUXInst_Y) );
  XOR2_X1 stateArray_S22reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A(
        stateArray_S22reg_gff_1_SFF_5_MUXInst_Y), .B(stateArray_outS23ser[5]), 
        .Z(stateArray_S22reg_gff_1_SFF_5_QD) );
  INV_X1 stateArray_S22reg_gff_1_SFF_5_Q_reg_U1 ( .A(stateArray_outS22ser[5]), 
        .ZN(stateArray_S22reg_gff_1_SFF_5_Q_reg_QN) );
  DFF_X1 stateArray_S22reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        stateArray_S22reg_gff_1_SFF_5_QD), .CK(clk), .Q(
        stateArray_outS22ser[5]), .QN() );
  XOR2_X1 stateArray_S22reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A(
        stateArray_outS23ser[6]), .B(MixColumns_line2_S02[7]), .Z(
        stateArray_S22reg_gff_1_SFF_6_MUXInst_X) );
  AND2_X1 stateArray_S22reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A1(stateArray_n6), 
        .A2(stateArray_S22reg_gff_1_SFF_6_MUXInst_X), .ZN(
        stateArray_S22reg_gff_1_SFF_6_MUXInst_Y) );
  XOR2_X1 stateArray_S22reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A(
        stateArray_S22reg_gff_1_SFF_6_MUXInst_Y), .B(stateArray_outS23ser[6]), 
        .Z(stateArray_S22reg_gff_1_SFF_6_QD) );
  INV_X1 stateArray_S22reg_gff_1_SFF_6_Q_reg_U1 ( .A(stateArray_outS22ser[6]), 
        .ZN(stateArray_S22reg_gff_1_SFF_6_Q_reg_QN) );
  DFF_X1 stateArray_S22reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        stateArray_S22reg_gff_1_SFF_6_QD), .CK(clk), .Q(
        stateArray_outS22ser[6]), .QN() );
  XOR2_X1 stateArray_S22reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A(
        stateArray_outS23ser[7]), .B(MixColumns_line2_S02[0]), .Z(
        stateArray_S22reg_gff_1_SFF_7_MUXInst_X) );
  AND2_X1 stateArray_S22reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A1(stateArray_n6), 
        .A2(stateArray_S22reg_gff_1_SFF_7_MUXInst_X), .ZN(
        stateArray_S22reg_gff_1_SFF_7_MUXInst_Y) );
  XOR2_X1 stateArray_S22reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A(
        stateArray_S22reg_gff_1_SFF_7_MUXInst_Y), .B(stateArray_outS23ser[7]), 
        .Z(stateArray_S22reg_gff_1_SFF_7_QD) );
  INV_X1 stateArray_S22reg_gff_1_SFF_7_Q_reg_U1 ( .A(stateArray_outS22ser[7]), 
        .ZN(stateArray_S22reg_gff_1_SFF_7_Q_reg_QN) );
  DFF_X1 stateArray_S22reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        stateArray_S22reg_gff_1_SFF_7_QD), .CK(clk), .Q(
        stateArray_outS22ser[7]), .QN() );
  XOR2_X1 stateArray_S23reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A(
        stateArray_inS23ser[0]), .B(stateArray_outS21ser[0]), .Z(
        stateArray_S23reg_gff_1_SFF_0_MUXInst_X) );
  AND2_X1 stateArray_S23reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A1(stateArray_n6), 
        .A2(stateArray_S23reg_gff_1_SFF_0_MUXInst_X), .ZN(
        stateArray_S23reg_gff_1_SFF_0_MUXInst_Y) );
  XOR2_X1 stateArray_S23reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A(
        stateArray_S23reg_gff_1_SFF_0_MUXInst_Y), .B(stateArray_inS23ser[0]), 
        .Z(stateArray_S23reg_gff_1_SFF_0_QD) );
  INV_X1 stateArray_S23reg_gff_1_SFF_0_Q_reg_U1 ( .A(stateArray_outS23ser[0]), 
        .ZN(stateArray_S23reg_gff_1_SFF_0_Q_reg_QN) );
  DFF_X1 stateArray_S23reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        stateArray_S23reg_gff_1_SFF_0_QD), .CK(clk), .Q(
        stateArray_outS23ser[0]), .QN() );
  XOR2_X1 stateArray_S23reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A(
        stateArray_inS23ser[1]), .B(stateArray_outS21ser[1]), .Z(
        stateArray_S23reg_gff_1_SFF_1_MUXInst_X) );
  AND2_X1 stateArray_S23reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A1(stateArray_n6), 
        .A2(stateArray_S23reg_gff_1_SFF_1_MUXInst_X), .ZN(
        stateArray_S23reg_gff_1_SFF_1_MUXInst_Y) );
  XOR2_X1 stateArray_S23reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A(
        stateArray_S23reg_gff_1_SFF_1_MUXInst_Y), .B(stateArray_inS23ser[1]), 
        .Z(stateArray_S23reg_gff_1_SFF_1_QD) );
  INV_X1 stateArray_S23reg_gff_1_SFF_1_Q_reg_U1 ( .A(stateArray_outS23ser[1]), 
        .ZN(stateArray_S23reg_gff_1_SFF_1_Q_reg_QN) );
  DFF_X1 stateArray_S23reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        stateArray_S23reg_gff_1_SFF_1_QD), .CK(clk), .Q(
        stateArray_outS23ser[1]), .QN() );
  XOR2_X1 stateArray_S23reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A(
        stateArray_inS23ser[2]), .B(stateArray_outS21ser[2]), .Z(
        stateArray_S23reg_gff_1_SFF_2_MUXInst_X) );
  AND2_X1 stateArray_S23reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A1(stateArray_n6), 
        .A2(stateArray_S23reg_gff_1_SFF_2_MUXInst_X), .ZN(
        stateArray_S23reg_gff_1_SFF_2_MUXInst_Y) );
  XOR2_X1 stateArray_S23reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A(
        stateArray_S23reg_gff_1_SFF_2_MUXInst_Y), .B(stateArray_inS23ser[2]), 
        .Z(stateArray_S23reg_gff_1_SFF_2_QD) );
  INV_X1 stateArray_S23reg_gff_1_SFF_2_Q_reg_U1 ( .A(stateArray_outS23ser[2]), 
        .ZN(stateArray_S23reg_gff_1_SFF_2_Q_reg_QN) );
  DFF_X1 stateArray_S23reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        stateArray_S23reg_gff_1_SFF_2_QD), .CK(clk), .Q(
        stateArray_outS23ser[2]), .QN() );
  XOR2_X1 stateArray_S23reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A(
        stateArray_inS23ser[3]), .B(stateArray_outS21ser[3]), .Z(
        stateArray_S23reg_gff_1_SFF_3_MUXInst_X) );
  AND2_X1 stateArray_S23reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A1(stateArray_n6), 
        .A2(stateArray_S23reg_gff_1_SFF_3_MUXInst_X), .ZN(
        stateArray_S23reg_gff_1_SFF_3_MUXInst_Y) );
  XOR2_X1 stateArray_S23reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A(
        stateArray_S23reg_gff_1_SFF_3_MUXInst_Y), .B(stateArray_inS23ser[3]), 
        .Z(stateArray_S23reg_gff_1_SFF_3_QD) );
  INV_X1 stateArray_S23reg_gff_1_SFF_3_Q_reg_U1 ( .A(stateArray_outS23ser[3]), 
        .ZN(stateArray_S23reg_gff_1_SFF_3_Q_reg_QN) );
  DFF_X1 stateArray_S23reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        stateArray_S23reg_gff_1_SFF_3_QD), .CK(clk), .Q(
        stateArray_outS23ser[3]), .QN() );
  XOR2_X1 stateArray_S23reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A(
        stateArray_inS23ser[4]), .B(stateArray_outS21ser[4]), .Z(
        stateArray_S23reg_gff_1_SFF_4_MUXInst_X) );
  AND2_X1 stateArray_S23reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A1(stateArray_n6), 
        .A2(stateArray_S23reg_gff_1_SFF_4_MUXInst_X), .ZN(
        stateArray_S23reg_gff_1_SFF_4_MUXInst_Y) );
  XOR2_X1 stateArray_S23reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A(
        stateArray_S23reg_gff_1_SFF_4_MUXInst_Y), .B(stateArray_inS23ser[4]), 
        .Z(stateArray_S23reg_gff_1_SFF_4_QD) );
  INV_X1 stateArray_S23reg_gff_1_SFF_4_Q_reg_U1 ( .A(stateArray_outS23ser[4]), 
        .ZN(stateArray_S23reg_gff_1_SFF_4_Q_reg_QN) );
  DFF_X1 stateArray_S23reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        stateArray_S23reg_gff_1_SFF_4_QD), .CK(clk), .Q(
        stateArray_outS23ser[4]), .QN() );
  XOR2_X1 stateArray_S23reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A(
        stateArray_inS23ser[5]), .B(stateArray_outS21ser[5]), .Z(
        stateArray_S23reg_gff_1_SFF_5_MUXInst_X) );
  AND2_X1 stateArray_S23reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A1(stateArray_n6), 
        .A2(stateArray_S23reg_gff_1_SFF_5_MUXInst_X), .ZN(
        stateArray_S23reg_gff_1_SFF_5_MUXInst_Y) );
  XOR2_X1 stateArray_S23reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A(
        stateArray_S23reg_gff_1_SFF_5_MUXInst_Y), .B(stateArray_inS23ser[5]), 
        .Z(stateArray_S23reg_gff_1_SFF_5_QD) );
  INV_X1 stateArray_S23reg_gff_1_SFF_5_Q_reg_U1 ( .A(stateArray_outS23ser[5]), 
        .ZN(stateArray_S23reg_gff_1_SFF_5_Q_reg_QN) );
  DFF_X1 stateArray_S23reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        stateArray_S23reg_gff_1_SFF_5_QD), .CK(clk), .Q(
        stateArray_outS23ser[5]), .QN() );
  XOR2_X1 stateArray_S23reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A(
        stateArray_inS23ser[6]), .B(stateArray_outS21ser[6]), .Z(
        stateArray_S23reg_gff_1_SFF_6_MUXInst_X) );
  AND2_X1 stateArray_S23reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A1(stateArray_n6), 
        .A2(stateArray_S23reg_gff_1_SFF_6_MUXInst_X), .ZN(
        stateArray_S23reg_gff_1_SFF_6_MUXInst_Y) );
  XOR2_X1 stateArray_S23reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A(
        stateArray_S23reg_gff_1_SFF_6_MUXInst_Y), .B(stateArray_inS23ser[6]), 
        .Z(stateArray_S23reg_gff_1_SFF_6_QD) );
  INV_X1 stateArray_S23reg_gff_1_SFF_6_Q_reg_U1 ( .A(stateArray_outS23ser[6]), 
        .ZN(stateArray_S23reg_gff_1_SFF_6_Q_reg_QN) );
  DFF_X1 stateArray_S23reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        stateArray_S23reg_gff_1_SFF_6_QD), .CK(clk), .Q(
        stateArray_outS23ser[6]), .QN() );
  XOR2_X1 stateArray_S23reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A(
        stateArray_inS23ser[7]), .B(stateArray_outS21ser[7]), .Z(
        stateArray_S23reg_gff_1_SFF_7_MUXInst_X) );
  AND2_X1 stateArray_S23reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A1(stateArray_n6), 
        .A2(stateArray_S23reg_gff_1_SFF_7_MUXInst_X), .ZN(
        stateArray_S23reg_gff_1_SFF_7_MUXInst_Y) );
  XOR2_X1 stateArray_S23reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A(
        stateArray_S23reg_gff_1_SFF_7_MUXInst_Y), .B(stateArray_inS23ser[7]), 
        .Z(stateArray_S23reg_gff_1_SFF_7_QD) );
  INV_X1 stateArray_S23reg_gff_1_SFF_7_Q_reg_U1 ( .A(stateArray_outS23ser[7]), 
        .ZN(stateArray_S23reg_gff_1_SFF_7_Q_reg_QN) );
  DFF_X1 stateArray_S23reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        stateArray_S23reg_gff_1_SFF_7_QD), .CK(clk), .Q(
        stateArray_outS23ser[7]), .QN() );
  XOR2_X1 stateArray_S30reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A(
        stateArray_outS31ser[0]), .B(stateArray_outS33ser[0]), .Z(
        stateArray_S30reg_gff_1_SFF_0_MUXInst_X) );
  AND2_X1 stateArray_S30reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A1(stateArray_n6), 
        .A2(stateArray_S30reg_gff_1_SFF_0_MUXInst_X), .ZN(
        stateArray_S30reg_gff_1_SFF_0_MUXInst_Y) );
  XOR2_X1 stateArray_S30reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A(
        stateArray_S30reg_gff_1_SFF_0_MUXInst_Y), .B(stateArray_outS31ser[0]), 
        .Z(stateArray_S30reg_gff_1_SFF_0_QD) );
  INV_X1 stateArray_S30reg_gff_1_SFF_0_Q_reg_U1 ( .A(MCin[0]), .ZN(
        stateArray_S30reg_gff_1_SFF_0_Q_reg_QN) );
  DFF_X1 stateArray_S30reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        stateArray_S30reg_gff_1_SFF_0_QD), .CK(clk), .Q(MCin[0]), .QN() );
  XOR2_X1 stateArray_S30reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A(
        stateArray_outS31ser[1]), .B(stateArray_outS33ser[1]), .Z(
        stateArray_S30reg_gff_1_SFF_1_MUXInst_X) );
  AND2_X1 stateArray_S30reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A1(stateArray_n6), 
        .A2(stateArray_S30reg_gff_1_SFF_1_MUXInst_X), .ZN(
        stateArray_S30reg_gff_1_SFF_1_MUXInst_Y) );
  XOR2_X1 stateArray_S30reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A(
        stateArray_S30reg_gff_1_SFF_1_MUXInst_Y), .B(stateArray_outS31ser[1]), 
        .Z(stateArray_S30reg_gff_1_SFF_1_QD) );
  INV_X1 stateArray_S30reg_gff_1_SFF_1_Q_reg_U1 ( .A(MixColumns_line3_S02[2]), 
        .ZN(stateArray_S30reg_gff_1_SFF_1_Q_reg_QN) );
  DFF_X1 stateArray_S30reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        stateArray_S30reg_gff_1_SFF_1_QD), .CK(clk), .Q(
        MixColumns_line3_S02[2]), .QN() );
  XOR2_X1 stateArray_S30reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A(
        stateArray_outS31ser[2]), .B(stateArray_outS33ser[2]), .Z(
        stateArray_S30reg_gff_1_SFF_2_MUXInst_X) );
  AND2_X1 stateArray_S30reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A1(stateArray_n6), 
        .A2(stateArray_S30reg_gff_1_SFF_2_MUXInst_X), .ZN(
        stateArray_S30reg_gff_1_SFF_2_MUXInst_Y) );
  XOR2_X1 stateArray_S30reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A(
        stateArray_S30reg_gff_1_SFF_2_MUXInst_Y), .B(stateArray_outS31ser[2]), 
        .Z(stateArray_S30reg_gff_1_SFF_2_QD) );
  INV_X1 stateArray_S30reg_gff_1_SFF_2_Q_reg_U1 ( .A(MCin[2]), .ZN(
        stateArray_S30reg_gff_1_SFF_2_Q_reg_QN) );
  DFF_X1 stateArray_S30reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        stateArray_S30reg_gff_1_SFF_2_QD), .CK(clk), .Q(MCin[2]), .QN() );
  XOR2_X1 stateArray_S30reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A(
        stateArray_outS31ser[3]), .B(stateArray_outS33ser[3]), .Z(
        stateArray_S30reg_gff_1_SFF_3_MUXInst_X) );
  AND2_X1 stateArray_S30reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A1(stateArray_n6), 
        .A2(stateArray_S30reg_gff_1_SFF_3_MUXInst_X), .ZN(
        stateArray_S30reg_gff_1_SFF_3_MUXInst_Y) );
  XOR2_X1 stateArray_S30reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A(
        stateArray_S30reg_gff_1_SFF_3_MUXInst_Y), .B(stateArray_outS31ser[3]), 
        .Z(stateArray_S30reg_gff_1_SFF_3_QD) );
  INV_X1 stateArray_S30reg_gff_1_SFF_3_Q_reg_U1 ( .A(MCin[3]), .ZN(
        stateArray_S30reg_gff_1_SFF_3_Q_reg_QN) );
  DFF_X1 stateArray_S30reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        stateArray_S30reg_gff_1_SFF_3_QD), .CK(clk), .Q(MCin[3]), .QN() );
  XOR2_X1 stateArray_S30reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A(
        stateArray_outS31ser[4]), .B(stateArray_outS33ser[4]), .Z(
        stateArray_S30reg_gff_1_SFF_4_MUXInst_X) );
  AND2_X1 stateArray_S30reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A1(stateArray_n6), 
        .A2(stateArray_S30reg_gff_1_SFF_4_MUXInst_X), .ZN(
        stateArray_S30reg_gff_1_SFF_4_MUXInst_Y) );
  XOR2_X1 stateArray_S30reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A(
        stateArray_S30reg_gff_1_SFF_4_MUXInst_Y), .B(stateArray_outS31ser[4]), 
        .Z(stateArray_S30reg_gff_1_SFF_4_QD) );
  INV_X1 stateArray_S30reg_gff_1_SFF_4_Q_reg_U1 ( .A(MixColumns_line3_S02[5]), 
        .ZN(stateArray_S30reg_gff_1_SFF_4_Q_reg_QN) );
  DFF_X1 stateArray_S30reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        stateArray_S30reg_gff_1_SFF_4_QD), .CK(clk), .Q(
        MixColumns_line3_S02[5]), .QN() );
  XOR2_X1 stateArray_S30reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A(
        stateArray_outS31ser[5]), .B(stateArray_outS33ser[5]), .Z(
        stateArray_S30reg_gff_1_SFF_5_MUXInst_X) );
  AND2_X1 stateArray_S30reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A1(stateArray_n6), 
        .A2(stateArray_S30reg_gff_1_SFF_5_MUXInst_X), .ZN(
        stateArray_S30reg_gff_1_SFF_5_MUXInst_Y) );
  XOR2_X1 stateArray_S30reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A(
        stateArray_S30reg_gff_1_SFF_5_MUXInst_Y), .B(stateArray_outS31ser[5]), 
        .Z(stateArray_S30reg_gff_1_SFF_5_QD) );
  INV_X1 stateArray_S30reg_gff_1_SFF_5_Q_reg_U1 ( .A(MixColumns_line3_S02[6]), 
        .ZN(stateArray_S30reg_gff_1_SFF_5_Q_reg_QN) );
  DFF_X1 stateArray_S30reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        stateArray_S30reg_gff_1_SFF_5_QD), .CK(clk), .Q(
        MixColumns_line3_S02[6]), .QN() );
  XOR2_X1 stateArray_S30reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A(
        stateArray_outS31ser[6]), .B(stateArray_outS33ser[6]), .Z(
        stateArray_S30reg_gff_1_SFF_6_MUXInst_X) );
  AND2_X1 stateArray_S30reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A1(stateArray_n6), 
        .A2(stateArray_S30reg_gff_1_SFF_6_MUXInst_X), .ZN(
        stateArray_S30reg_gff_1_SFF_6_MUXInst_Y) );
  XOR2_X1 stateArray_S30reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A(
        stateArray_S30reg_gff_1_SFF_6_MUXInst_Y), .B(stateArray_outS31ser[6]), 
        .Z(stateArray_S30reg_gff_1_SFF_6_QD) );
  INV_X1 stateArray_S30reg_gff_1_SFF_6_Q_reg_U1 ( .A(MixColumns_line3_S02[7]), 
        .ZN(stateArray_S30reg_gff_1_SFF_6_Q_reg_QN) );
  DFF_X1 stateArray_S30reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        stateArray_S30reg_gff_1_SFF_6_QD), .CK(clk), .Q(
        MixColumns_line3_S02[7]), .QN() );
  XOR2_X1 stateArray_S30reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A(
        stateArray_outS31ser[7]), .B(stateArray_outS33ser[7]), .Z(
        stateArray_S30reg_gff_1_SFF_7_MUXInst_X) );
  AND2_X1 stateArray_S30reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A1(stateArray_n6), 
        .A2(stateArray_S30reg_gff_1_SFF_7_MUXInst_X), .ZN(
        stateArray_S30reg_gff_1_SFF_7_MUXInst_Y) );
  XOR2_X1 stateArray_S30reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A(
        stateArray_S30reg_gff_1_SFF_7_MUXInst_Y), .B(stateArray_outS31ser[7]), 
        .Z(stateArray_S30reg_gff_1_SFF_7_QD) );
  INV_X1 stateArray_S30reg_gff_1_SFF_7_Q_reg_U1 ( .A(MixColumns_line3_S02[0]), 
        .ZN(stateArray_S30reg_gff_1_SFF_7_Q_reg_QN) );
  DFF_X1 stateArray_S30reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        stateArray_S30reg_gff_1_SFF_7_QD), .CK(clk), .Q(
        MixColumns_line3_S02[0]), .QN() );
  XOR2_X1 stateArray_S31reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A(
        stateArray_outS32ser[0]), .B(MCin[0]), .Z(
        stateArray_S31reg_gff_1_SFF_0_MUXInst_X) );
  AND2_X1 stateArray_S31reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A1(stateArray_n6), 
        .A2(stateArray_S31reg_gff_1_SFF_0_MUXInst_X), .ZN(
        stateArray_S31reg_gff_1_SFF_0_MUXInst_Y) );
  XOR2_X1 stateArray_S31reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A(
        stateArray_S31reg_gff_1_SFF_0_MUXInst_Y), .B(stateArray_outS32ser[0]), 
        .Z(stateArray_S31reg_gff_1_SFF_0_QD) );
  INV_X1 stateArray_S31reg_gff_1_SFF_0_Q_reg_U1 ( .A(stateArray_outS31ser[0]), 
        .ZN(stateArray_S31reg_gff_1_SFF_0_Q_reg_QN) );
  DFF_X1 stateArray_S31reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        stateArray_S31reg_gff_1_SFF_0_QD), .CK(clk), .Q(
        stateArray_outS31ser[0]), .QN() );
  XOR2_X1 stateArray_S31reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A(
        stateArray_outS32ser[1]), .B(MixColumns_line3_S02[2]), .Z(
        stateArray_S31reg_gff_1_SFF_1_MUXInst_X) );
  AND2_X1 stateArray_S31reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A1(stateArray_n6), 
        .A2(stateArray_S31reg_gff_1_SFF_1_MUXInst_X), .ZN(
        stateArray_S31reg_gff_1_SFF_1_MUXInst_Y) );
  XOR2_X1 stateArray_S31reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A(
        stateArray_S31reg_gff_1_SFF_1_MUXInst_Y), .B(stateArray_outS32ser[1]), 
        .Z(stateArray_S31reg_gff_1_SFF_1_QD) );
  INV_X1 stateArray_S31reg_gff_1_SFF_1_Q_reg_U1 ( .A(stateArray_outS31ser[1]), 
        .ZN(stateArray_S31reg_gff_1_SFF_1_Q_reg_QN) );
  DFF_X1 stateArray_S31reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        stateArray_S31reg_gff_1_SFF_1_QD), .CK(clk), .Q(
        stateArray_outS31ser[1]), .QN() );
  XOR2_X1 stateArray_S31reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A(
        stateArray_outS32ser[2]), .B(MCin[2]), .Z(
        stateArray_S31reg_gff_1_SFF_2_MUXInst_X) );
  AND2_X1 stateArray_S31reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A1(stateArray_n6), 
        .A2(stateArray_S31reg_gff_1_SFF_2_MUXInst_X), .ZN(
        stateArray_S31reg_gff_1_SFF_2_MUXInst_Y) );
  XOR2_X1 stateArray_S31reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A(
        stateArray_S31reg_gff_1_SFF_2_MUXInst_Y), .B(stateArray_outS32ser[2]), 
        .Z(stateArray_S31reg_gff_1_SFF_2_QD) );
  INV_X1 stateArray_S31reg_gff_1_SFF_2_Q_reg_U1 ( .A(stateArray_outS31ser[2]), 
        .ZN(stateArray_S31reg_gff_1_SFF_2_Q_reg_QN) );
  DFF_X1 stateArray_S31reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        stateArray_S31reg_gff_1_SFF_2_QD), .CK(clk), .Q(
        stateArray_outS31ser[2]), .QN() );
  XOR2_X1 stateArray_S31reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A(
        stateArray_outS32ser[3]), .B(MCin[3]), .Z(
        stateArray_S31reg_gff_1_SFF_3_MUXInst_X) );
  AND2_X1 stateArray_S31reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A1(stateArray_n6), 
        .A2(stateArray_S31reg_gff_1_SFF_3_MUXInst_X), .ZN(
        stateArray_S31reg_gff_1_SFF_3_MUXInst_Y) );
  XOR2_X1 stateArray_S31reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A(
        stateArray_S31reg_gff_1_SFF_3_MUXInst_Y), .B(stateArray_outS32ser[3]), 
        .Z(stateArray_S31reg_gff_1_SFF_3_QD) );
  INV_X1 stateArray_S31reg_gff_1_SFF_3_Q_reg_U1 ( .A(stateArray_outS31ser[3]), 
        .ZN(stateArray_S31reg_gff_1_SFF_3_Q_reg_QN) );
  DFF_X1 stateArray_S31reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        stateArray_S31reg_gff_1_SFF_3_QD), .CK(clk), .Q(
        stateArray_outS31ser[3]), .QN() );
  XOR2_X1 stateArray_S31reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A(
        stateArray_outS32ser[4]), .B(MixColumns_line3_S02[5]), .Z(
        stateArray_S31reg_gff_1_SFF_4_MUXInst_X) );
  AND2_X1 stateArray_S31reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A1(stateArray_n6), 
        .A2(stateArray_S31reg_gff_1_SFF_4_MUXInst_X), .ZN(
        stateArray_S31reg_gff_1_SFF_4_MUXInst_Y) );
  XOR2_X1 stateArray_S31reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A(
        stateArray_S31reg_gff_1_SFF_4_MUXInst_Y), .B(stateArray_outS32ser[4]), 
        .Z(stateArray_S31reg_gff_1_SFF_4_QD) );
  INV_X1 stateArray_S31reg_gff_1_SFF_4_Q_reg_U1 ( .A(stateArray_outS31ser[4]), 
        .ZN(stateArray_S31reg_gff_1_SFF_4_Q_reg_QN) );
  DFF_X1 stateArray_S31reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        stateArray_S31reg_gff_1_SFF_4_QD), .CK(clk), .Q(
        stateArray_outS31ser[4]), .QN() );
  XOR2_X1 stateArray_S31reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A(
        stateArray_outS32ser[5]), .B(MixColumns_line3_S02[6]), .Z(
        stateArray_S31reg_gff_1_SFF_5_MUXInst_X) );
  AND2_X1 stateArray_S31reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A1(stateArray_n6), 
        .A2(stateArray_S31reg_gff_1_SFF_5_MUXInst_X), .ZN(
        stateArray_S31reg_gff_1_SFF_5_MUXInst_Y) );
  XOR2_X1 stateArray_S31reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A(
        stateArray_S31reg_gff_1_SFF_5_MUXInst_Y), .B(stateArray_outS32ser[5]), 
        .Z(stateArray_S31reg_gff_1_SFF_5_QD) );
  INV_X1 stateArray_S31reg_gff_1_SFF_5_Q_reg_U1 ( .A(stateArray_outS31ser[5]), 
        .ZN(stateArray_S31reg_gff_1_SFF_5_Q_reg_QN) );
  DFF_X1 stateArray_S31reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        stateArray_S31reg_gff_1_SFF_5_QD), .CK(clk), .Q(
        stateArray_outS31ser[5]), .QN() );
  XOR2_X1 stateArray_S31reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A(
        stateArray_outS32ser[6]), .B(MixColumns_line3_S02[7]), .Z(
        stateArray_S31reg_gff_1_SFF_6_MUXInst_X) );
  AND2_X1 stateArray_S31reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A1(stateArray_n6), 
        .A2(stateArray_S31reg_gff_1_SFF_6_MUXInst_X), .ZN(
        stateArray_S31reg_gff_1_SFF_6_MUXInst_Y) );
  XOR2_X1 stateArray_S31reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A(
        stateArray_S31reg_gff_1_SFF_6_MUXInst_Y), .B(stateArray_outS32ser[6]), 
        .Z(stateArray_S31reg_gff_1_SFF_6_QD) );
  INV_X1 stateArray_S31reg_gff_1_SFF_6_Q_reg_U1 ( .A(stateArray_outS31ser[6]), 
        .ZN(stateArray_S31reg_gff_1_SFF_6_Q_reg_QN) );
  DFF_X1 stateArray_S31reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        stateArray_S31reg_gff_1_SFF_6_QD), .CK(clk), .Q(
        stateArray_outS31ser[6]), .QN() );
  XOR2_X1 stateArray_S31reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A(
        stateArray_outS32ser[7]), .B(MixColumns_line3_S02[0]), .Z(
        stateArray_S31reg_gff_1_SFF_7_MUXInst_X) );
  AND2_X1 stateArray_S31reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A1(stateArray_n6), 
        .A2(stateArray_S31reg_gff_1_SFF_7_MUXInst_X), .ZN(
        stateArray_S31reg_gff_1_SFF_7_MUXInst_Y) );
  XOR2_X1 stateArray_S31reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A(
        stateArray_S31reg_gff_1_SFF_7_MUXInst_Y), .B(stateArray_outS32ser[7]), 
        .Z(stateArray_S31reg_gff_1_SFF_7_QD) );
  INV_X1 stateArray_S31reg_gff_1_SFF_7_Q_reg_U1 ( .A(stateArray_outS31ser[7]), 
        .ZN(stateArray_S31reg_gff_1_SFF_7_Q_reg_QN) );
  DFF_X1 stateArray_S31reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        stateArray_S31reg_gff_1_SFF_7_QD), .CK(clk), .Q(
        stateArray_outS31ser[7]), .QN() );
  XOR2_X1 stateArray_S32reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A(
        stateArray_outS33ser[0]), .B(stateArray_outS31ser[0]), .Z(
        stateArray_S32reg_gff_1_SFF_0_MUXInst_X) );
  AND2_X1 stateArray_S32reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A1(stateArray_n6), 
        .A2(stateArray_S32reg_gff_1_SFF_0_MUXInst_X), .ZN(
        stateArray_S32reg_gff_1_SFF_0_MUXInst_Y) );
  XOR2_X1 stateArray_S32reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A(
        stateArray_S32reg_gff_1_SFF_0_MUXInst_Y), .B(stateArray_outS33ser[0]), 
        .Z(stateArray_S32reg_gff_1_SFF_0_QD) );
  INV_X1 stateArray_S32reg_gff_1_SFF_0_Q_reg_U1 ( .A(stateArray_outS32ser[0]), 
        .ZN(stateArray_S32reg_gff_1_SFF_0_Q_reg_QN) );
  DFF_X1 stateArray_S32reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        stateArray_S32reg_gff_1_SFF_0_QD), .CK(clk), .Q(
        stateArray_outS32ser[0]), .QN() );
  XOR2_X1 stateArray_S32reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A(
        stateArray_outS33ser[1]), .B(stateArray_outS31ser[1]), .Z(
        stateArray_S32reg_gff_1_SFF_1_MUXInst_X) );
  AND2_X1 stateArray_S32reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A1(stateArray_n6), 
        .A2(stateArray_S32reg_gff_1_SFF_1_MUXInst_X), .ZN(
        stateArray_S32reg_gff_1_SFF_1_MUXInst_Y) );
  XOR2_X1 stateArray_S32reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A(
        stateArray_S32reg_gff_1_SFF_1_MUXInst_Y), .B(stateArray_outS33ser[1]), 
        .Z(stateArray_S32reg_gff_1_SFF_1_QD) );
  INV_X1 stateArray_S32reg_gff_1_SFF_1_Q_reg_U1 ( .A(stateArray_outS32ser[1]), 
        .ZN(stateArray_S32reg_gff_1_SFF_1_Q_reg_QN) );
  DFF_X1 stateArray_S32reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        stateArray_S32reg_gff_1_SFF_1_QD), .CK(clk), .Q(
        stateArray_outS32ser[1]), .QN() );
  XOR2_X1 stateArray_S32reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A(
        stateArray_outS33ser[2]), .B(stateArray_outS31ser[2]), .Z(
        stateArray_S32reg_gff_1_SFF_2_MUXInst_X) );
  AND2_X1 stateArray_S32reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A1(stateArray_n6), 
        .A2(stateArray_S32reg_gff_1_SFF_2_MUXInst_X), .ZN(
        stateArray_S32reg_gff_1_SFF_2_MUXInst_Y) );
  XOR2_X1 stateArray_S32reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A(
        stateArray_S32reg_gff_1_SFF_2_MUXInst_Y), .B(stateArray_outS33ser[2]), 
        .Z(stateArray_S32reg_gff_1_SFF_2_QD) );
  INV_X1 stateArray_S32reg_gff_1_SFF_2_Q_reg_U1 ( .A(stateArray_outS32ser[2]), 
        .ZN(stateArray_S32reg_gff_1_SFF_2_Q_reg_QN) );
  DFF_X1 stateArray_S32reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        stateArray_S32reg_gff_1_SFF_2_QD), .CK(clk), .Q(
        stateArray_outS32ser[2]), .QN() );
  XOR2_X1 stateArray_S32reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A(
        stateArray_outS33ser[3]), .B(stateArray_outS31ser[3]), .Z(
        stateArray_S32reg_gff_1_SFF_3_MUXInst_X) );
  AND2_X1 stateArray_S32reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A1(stateArray_n6), 
        .A2(stateArray_S32reg_gff_1_SFF_3_MUXInst_X), .ZN(
        stateArray_S32reg_gff_1_SFF_3_MUXInst_Y) );
  XOR2_X1 stateArray_S32reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A(
        stateArray_S32reg_gff_1_SFF_3_MUXInst_Y), .B(stateArray_outS33ser[3]), 
        .Z(stateArray_S32reg_gff_1_SFF_3_QD) );
  INV_X1 stateArray_S32reg_gff_1_SFF_3_Q_reg_U1 ( .A(stateArray_outS32ser[3]), 
        .ZN(stateArray_S32reg_gff_1_SFF_3_Q_reg_QN) );
  DFF_X1 stateArray_S32reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        stateArray_S32reg_gff_1_SFF_3_QD), .CK(clk), .Q(
        stateArray_outS32ser[3]), .QN() );
  XOR2_X1 stateArray_S32reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A(
        stateArray_outS33ser[4]), .B(stateArray_outS31ser[4]), .Z(
        stateArray_S32reg_gff_1_SFF_4_MUXInst_X) );
  AND2_X1 stateArray_S32reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A1(stateArray_n6), 
        .A2(stateArray_S32reg_gff_1_SFF_4_MUXInst_X), .ZN(
        stateArray_S32reg_gff_1_SFF_4_MUXInst_Y) );
  XOR2_X1 stateArray_S32reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A(
        stateArray_S32reg_gff_1_SFF_4_MUXInst_Y), .B(stateArray_outS33ser[4]), 
        .Z(stateArray_S32reg_gff_1_SFF_4_QD) );
  INV_X1 stateArray_S32reg_gff_1_SFF_4_Q_reg_U1 ( .A(stateArray_outS32ser[4]), 
        .ZN(stateArray_S32reg_gff_1_SFF_4_Q_reg_QN) );
  DFF_X1 stateArray_S32reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        stateArray_S32reg_gff_1_SFF_4_QD), .CK(clk), .Q(
        stateArray_outS32ser[4]), .QN() );
  XOR2_X1 stateArray_S32reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A(
        stateArray_outS33ser[5]), .B(stateArray_outS31ser[5]), .Z(
        stateArray_S32reg_gff_1_SFF_5_MUXInst_X) );
  AND2_X1 stateArray_S32reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A1(stateArray_n6), 
        .A2(stateArray_S32reg_gff_1_SFF_5_MUXInst_X), .ZN(
        stateArray_S32reg_gff_1_SFF_5_MUXInst_Y) );
  XOR2_X1 stateArray_S32reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A(
        stateArray_S32reg_gff_1_SFF_5_MUXInst_Y), .B(stateArray_outS33ser[5]), 
        .Z(stateArray_S32reg_gff_1_SFF_5_QD) );
  INV_X1 stateArray_S32reg_gff_1_SFF_5_Q_reg_U1 ( .A(stateArray_outS32ser[5]), 
        .ZN(stateArray_S32reg_gff_1_SFF_5_Q_reg_QN) );
  DFF_X1 stateArray_S32reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        stateArray_S32reg_gff_1_SFF_5_QD), .CK(clk), .Q(
        stateArray_outS32ser[5]), .QN() );
  XOR2_X1 stateArray_S32reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A(
        stateArray_outS33ser[6]), .B(stateArray_outS31ser[6]), .Z(
        stateArray_S32reg_gff_1_SFF_6_MUXInst_X) );
  AND2_X1 stateArray_S32reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A1(stateArray_n6), 
        .A2(stateArray_S32reg_gff_1_SFF_6_MUXInst_X), .ZN(
        stateArray_S32reg_gff_1_SFF_6_MUXInst_Y) );
  XOR2_X1 stateArray_S32reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A(
        stateArray_S32reg_gff_1_SFF_6_MUXInst_Y), .B(stateArray_outS33ser[6]), 
        .Z(stateArray_S32reg_gff_1_SFF_6_QD) );
  INV_X1 stateArray_S32reg_gff_1_SFF_6_Q_reg_U1 ( .A(stateArray_outS32ser[6]), 
        .ZN(stateArray_S32reg_gff_1_SFF_6_Q_reg_QN) );
  DFF_X1 stateArray_S32reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        stateArray_S32reg_gff_1_SFF_6_QD), .CK(clk), .Q(
        stateArray_outS32ser[6]), .QN() );
  XOR2_X1 stateArray_S32reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A(
        stateArray_outS33ser[7]), .B(stateArray_outS31ser[7]), .Z(
        stateArray_S32reg_gff_1_SFF_7_MUXInst_X) );
  AND2_X1 stateArray_S32reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A1(stateArray_n6), 
        .A2(stateArray_S32reg_gff_1_SFF_7_MUXInst_X), .ZN(
        stateArray_S32reg_gff_1_SFF_7_MUXInst_Y) );
  XOR2_X1 stateArray_S32reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A(
        stateArray_S32reg_gff_1_SFF_7_MUXInst_Y), .B(stateArray_outS33ser[7]), 
        .Z(stateArray_S32reg_gff_1_SFF_7_QD) );
  INV_X1 stateArray_S32reg_gff_1_SFF_7_Q_reg_U1 ( .A(stateArray_outS32ser[7]), 
        .ZN(stateArray_S32reg_gff_1_SFF_7_Q_reg_QN) );
  DFF_X1 stateArray_S32reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        stateArray_S32reg_gff_1_SFF_7_QD), .CK(clk), .Q(
        stateArray_outS32ser[7]), .QN() );
  XOR2_X1 stateArray_S33reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A(
        stateArray_inS33ser[0]), .B(stateArray_outS32ser[0]), .Z(
        stateArray_S33reg_gff_1_SFF_0_MUXInst_X) );
  AND2_X1 stateArray_S33reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A1(stateArray_n6), 
        .A2(stateArray_S33reg_gff_1_SFF_0_MUXInst_X), .ZN(
        stateArray_S33reg_gff_1_SFF_0_MUXInst_Y) );
  XOR2_X1 stateArray_S33reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A(
        stateArray_S33reg_gff_1_SFF_0_MUXInst_Y), .B(stateArray_inS33ser[0]), 
        .Z(stateArray_S33reg_gff_1_SFF_0_QD) );
  INV_X1 stateArray_S33reg_gff_1_SFF_0_Q_reg_U1 ( .A(stateArray_outS33ser[0]), 
        .ZN(stateArray_S33reg_gff_1_SFF_0_Q_reg_QN) );
  DFF_X1 stateArray_S33reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        stateArray_S33reg_gff_1_SFF_0_QD), .CK(clk), .Q(
        stateArray_outS33ser[0]), .QN() );
  XOR2_X1 stateArray_S33reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A(
        stateArray_inS33ser[1]), .B(stateArray_outS32ser[1]), .Z(
        stateArray_S33reg_gff_1_SFF_1_MUXInst_X) );
  AND2_X1 stateArray_S33reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A1(stateArray_n6), 
        .A2(stateArray_S33reg_gff_1_SFF_1_MUXInst_X), .ZN(
        stateArray_S33reg_gff_1_SFF_1_MUXInst_Y) );
  XOR2_X1 stateArray_S33reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A(
        stateArray_S33reg_gff_1_SFF_1_MUXInst_Y), .B(stateArray_inS33ser[1]), 
        .Z(stateArray_S33reg_gff_1_SFF_1_QD) );
  INV_X1 stateArray_S33reg_gff_1_SFF_1_Q_reg_U1 ( .A(stateArray_outS33ser[1]), 
        .ZN(stateArray_S33reg_gff_1_SFF_1_Q_reg_QN) );
  DFF_X1 stateArray_S33reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        stateArray_S33reg_gff_1_SFF_1_QD), .CK(clk), .Q(
        stateArray_outS33ser[1]), .QN() );
  XOR2_X1 stateArray_S33reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A(
        stateArray_inS33ser[2]), .B(stateArray_outS32ser[2]), .Z(
        stateArray_S33reg_gff_1_SFF_2_MUXInst_X) );
  AND2_X1 stateArray_S33reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A1(stateArray_n6), 
        .A2(stateArray_S33reg_gff_1_SFF_2_MUXInst_X), .ZN(
        stateArray_S33reg_gff_1_SFF_2_MUXInst_Y) );
  XOR2_X1 stateArray_S33reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A(
        stateArray_S33reg_gff_1_SFF_2_MUXInst_Y), .B(stateArray_inS33ser[2]), 
        .Z(stateArray_S33reg_gff_1_SFF_2_QD) );
  INV_X1 stateArray_S33reg_gff_1_SFF_2_Q_reg_U1 ( .A(stateArray_outS33ser[2]), 
        .ZN(stateArray_S33reg_gff_1_SFF_2_Q_reg_QN) );
  DFF_X1 stateArray_S33reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        stateArray_S33reg_gff_1_SFF_2_QD), .CK(clk), .Q(
        stateArray_outS33ser[2]), .QN() );
  XOR2_X1 stateArray_S33reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A(
        stateArray_inS33ser[3]), .B(stateArray_outS32ser[3]), .Z(
        stateArray_S33reg_gff_1_SFF_3_MUXInst_X) );
  AND2_X1 stateArray_S33reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A1(stateArray_n6), 
        .A2(stateArray_S33reg_gff_1_SFF_3_MUXInst_X), .ZN(
        stateArray_S33reg_gff_1_SFF_3_MUXInst_Y) );
  XOR2_X1 stateArray_S33reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A(
        stateArray_S33reg_gff_1_SFF_3_MUXInst_Y), .B(stateArray_inS33ser[3]), 
        .Z(stateArray_S33reg_gff_1_SFF_3_QD) );
  INV_X1 stateArray_S33reg_gff_1_SFF_3_Q_reg_U1 ( .A(stateArray_outS33ser[3]), 
        .ZN(stateArray_S33reg_gff_1_SFF_3_Q_reg_QN) );
  DFF_X1 stateArray_S33reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        stateArray_S33reg_gff_1_SFF_3_QD), .CK(clk), .Q(
        stateArray_outS33ser[3]), .QN() );
  XOR2_X1 stateArray_S33reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A(
        stateArray_inS33ser[4]), .B(stateArray_outS32ser[4]), .Z(
        stateArray_S33reg_gff_1_SFF_4_MUXInst_X) );
  AND2_X1 stateArray_S33reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A1(stateArray_n6), 
        .A2(stateArray_S33reg_gff_1_SFF_4_MUXInst_X), .ZN(
        stateArray_S33reg_gff_1_SFF_4_MUXInst_Y) );
  XOR2_X1 stateArray_S33reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A(
        stateArray_S33reg_gff_1_SFF_4_MUXInst_Y), .B(stateArray_inS33ser[4]), 
        .Z(stateArray_S33reg_gff_1_SFF_4_QD) );
  INV_X1 stateArray_S33reg_gff_1_SFF_4_Q_reg_U1 ( .A(stateArray_outS33ser[4]), 
        .ZN(stateArray_S33reg_gff_1_SFF_4_Q_reg_QN) );
  DFF_X1 stateArray_S33reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        stateArray_S33reg_gff_1_SFF_4_QD), .CK(clk), .Q(
        stateArray_outS33ser[4]), .QN() );
  XOR2_X1 stateArray_S33reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A(
        stateArray_inS33ser[5]), .B(stateArray_outS32ser[5]), .Z(
        stateArray_S33reg_gff_1_SFF_5_MUXInst_X) );
  AND2_X1 stateArray_S33reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A1(stateArray_n6), 
        .A2(stateArray_S33reg_gff_1_SFF_5_MUXInst_X), .ZN(
        stateArray_S33reg_gff_1_SFF_5_MUXInst_Y) );
  XOR2_X1 stateArray_S33reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A(
        stateArray_S33reg_gff_1_SFF_5_MUXInst_Y), .B(stateArray_inS33ser[5]), 
        .Z(stateArray_S33reg_gff_1_SFF_5_QD) );
  INV_X1 stateArray_S33reg_gff_1_SFF_5_Q_reg_U1 ( .A(stateArray_outS33ser[5]), 
        .ZN(stateArray_S33reg_gff_1_SFF_5_Q_reg_QN) );
  DFF_X1 stateArray_S33reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        stateArray_S33reg_gff_1_SFF_5_QD), .CK(clk), .Q(
        stateArray_outS33ser[5]), .QN() );
  XOR2_X1 stateArray_S33reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A(
        stateArray_inS33ser[6]), .B(stateArray_outS32ser[6]), .Z(
        stateArray_S33reg_gff_1_SFF_6_MUXInst_X) );
  AND2_X1 stateArray_S33reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A1(stateArray_n6), 
        .A2(stateArray_S33reg_gff_1_SFF_6_MUXInst_X), .ZN(
        stateArray_S33reg_gff_1_SFF_6_MUXInst_Y) );
  XOR2_X1 stateArray_S33reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A(
        stateArray_S33reg_gff_1_SFF_6_MUXInst_Y), .B(stateArray_inS33ser[6]), 
        .Z(stateArray_S33reg_gff_1_SFF_6_QD) );
  INV_X1 stateArray_S33reg_gff_1_SFF_6_Q_reg_U1 ( .A(stateArray_outS33ser[6]), 
        .ZN(stateArray_S33reg_gff_1_SFF_6_Q_reg_QN) );
  DFF_X1 stateArray_S33reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        stateArray_S33reg_gff_1_SFF_6_QD), .CK(clk), .Q(
        stateArray_outS33ser[6]), .QN() );
  XOR2_X1 stateArray_S33reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A(
        stateArray_inS33ser[7]), .B(stateArray_outS32ser[7]), .Z(
        stateArray_S33reg_gff_1_SFF_7_MUXInst_X) );
  AND2_X1 stateArray_S33reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A1(stateArray_n6), 
        .A2(stateArray_S33reg_gff_1_SFF_7_MUXInst_X), .ZN(
        stateArray_S33reg_gff_1_SFF_7_MUXInst_Y) );
  XOR2_X1 stateArray_S33reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A(
        stateArray_S33reg_gff_1_SFF_7_MUXInst_Y), .B(stateArray_inS33ser[7]), 
        .Z(stateArray_S33reg_gff_1_SFF_7_QD) );
  INV_X1 stateArray_S33reg_gff_1_SFF_7_Q_reg_U1 ( .A(stateArray_outS33ser[7]), 
        .ZN(stateArray_S33reg_gff_1_SFF_7_Q_reg_QN) );
  DFF_X1 stateArray_S33reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        stateArray_S33reg_gff_1_SFF_7_QD), .CK(clk), .Q(
        stateArray_outS33ser[7]), .QN() );
  XOR2_X1 stateArray_MUX_inS03ser_mux_inst_0_XOR1_U1 ( .A(MCin[16]), .B(
        StateInMC[24]), .Z(stateArray_MUX_inS03ser_mux_inst_0_X) );
  AND2_X1 stateArray_MUX_inS03ser_mux_inst_0_AND1_U1 ( .A1(
        stateArray_nReset_selMC), .A2(stateArray_MUX_inS03ser_mux_inst_0_X), 
        .ZN(stateArray_MUX_inS03ser_mux_inst_0_Y) );
  XOR2_X1 stateArray_MUX_inS03ser_mux_inst_0_XOR2_U1 ( .A(
        stateArray_MUX_inS03ser_mux_inst_0_Y), .B(MCin[16]), .Z(
        stateArray_inS03ser[0]) );
  XOR2_X1 stateArray_MUX_inS03ser_mux_inst_1_XOR1_U1 ( .A(
        MixColumns_line1_S02[2]), .B(StateInMC[25]), .Z(
        stateArray_MUX_inS03ser_mux_inst_1_X) );
  AND2_X1 stateArray_MUX_inS03ser_mux_inst_1_AND1_U1 ( .A1(
        stateArray_nReset_selMC), .A2(stateArray_MUX_inS03ser_mux_inst_1_X), 
        .ZN(stateArray_MUX_inS03ser_mux_inst_1_Y) );
  XOR2_X1 stateArray_MUX_inS03ser_mux_inst_1_XOR2_U1 ( .A(
        stateArray_MUX_inS03ser_mux_inst_1_Y), .B(MixColumns_line1_S02[2]), 
        .Z(stateArray_inS03ser[1]) );
  XOR2_X1 stateArray_MUX_inS03ser_mux_inst_2_XOR1_U1 ( .A(MCin[18]), .B(
        StateInMC[26]), .Z(stateArray_MUX_inS03ser_mux_inst_2_X) );
  AND2_X1 stateArray_MUX_inS03ser_mux_inst_2_AND1_U1 ( .A1(
        stateArray_nReset_selMC), .A2(stateArray_MUX_inS03ser_mux_inst_2_X), 
        .ZN(stateArray_MUX_inS03ser_mux_inst_2_Y) );
  XOR2_X1 stateArray_MUX_inS03ser_mux_inst_2_XOR2_U1 ( .A(
        stateArray_MUX_inS03ser_mux_inst_2_Y), .B(MCin[18]), .Z(
        stateArray_inS03ser[2]) );
  XOR2_X1 stateArray_MUX_inS03ser_mux_inst_3_XOR1_U1 ( .A(MCin[19]), .B(
        StateInMC[27]), .Z(stateArray_MUX_inS03ser_mux_inst_3_X) );
  AND2_X1 stateArray_MUX_inS03ser_mux_inst_3_AND1_U1 ( .A1(
        stateArray_nReset_selMC), .A2(stateArray_MUX_inS03ser_mux_inst_3_X), 
        .ZN(stateArray_MUX_inS03ser_mux_inst_3_Y) );
  XOR2_X1 stateArray_MUX_inS03ser_mux_inst_3_XOR2_U1 ( .A(
        stateArray_MUX_inS03ser_mux_inst_3_Y), .B(MCin[19]), .Z(
        stateArray_inS03ser[3]) );
  XOR2_X1 stateArray_MUX_inS03ser_mux_inst_4_XOR1_U1 ( .A(
        MixColumns_line1_S02[5]), .B(StateInMC[28]), .Z(
        stateArray_MUX_inS03ser_mux_inst_4_X) );
  AND2_X1 stateArray_MUX_inS03ser_mux_inst_4_AND1_U1 ( .A1(
        stateArray_nReset_selMC), .A2(stateArray_MUX_inS03ser_mux_inst_4_X), 
        .ZN(stateArray_MUX_inS03ser_mux_inst_4_Y) );
  XOR2_X1 stateArray_MUX_inS03ser_mux_inst_4_XOR2_U1 ( .A(
        stateArray_MUX_inS03ser_mux_inst_4_Y), .B(MixColumns_line1_S02[5]), 
        .Z(stateArray_inS03ser[4]) );
  XOR2_X1 stateArray_MUX_inS03ser_mux_inst_5_XOR1_U1 ( .A(
        MixColumns_line1_S02[6]), .B(StateInMC[29]), .Z(
        stateArray_MUX_inS03ser_mux_inst_5_X) );
  AND2_X1 stateArray_MUX_inS03ser_mux_inst_5_AND1_U1 ( .A1(
        stateArray_nReset_selMC), .A2(stateArray_MUX_inS03ser_mux_inst_5_X), 
        .ZN(stateArray_MUX_inS03ser_mux_inst_5_Y) );
  XOR2_X1 stateArray_MUX_inS03ser_mux_inst_5_XOR2_U1 ( .A(
        stateArray_MUX_inS03ser_mux_inst_5_Y), .B(MixColumns_line1_S02[6]), 
        .Z(stateArray_inS03ser[5]) );
  XOR2_X1 stateArray_MUX_inS03ser_mux_inst_6_XOR1_U1 ( .A(
        MixColumns_line1_S02[7]), .B(StateInMC[30]), .Z(
        stateArray_MUX_inS03ser_mux_inst_6_X) );
  AND2_X1 stateArray_MUX_inS03ser_mux_inst_6_AND1_U1 ( .A1(
        stateArray_nReset_selMC), .A2(stateArray_MUX_inS03ser_mux_inst_6_X), 
        .ZN(stateArray_MUX_inS03ser_mux_inst_6_Y) );
  XOR2_X1 stateArray_MUX_inS03ser_mux_inst_6_XOR2_U1 ( .A(
        stateArray_MUX_inS03ser_mux_inst_6_Y), .B(MixColumns_line1_S02[7]), 
        .Z(stateArray_inS03ser[6]) );
  XOR2_X1 stateArray_MUX_inS03ser_mux_inst_7_XOR1_U1 ( .A(
        MixColumns_line1_S02[0]), .B(StateInMC[31]), .Z(
        stateArray_MUX_inS03ser_mux_inst_7_X) );
  AND2_X1 stateArray_MUX_inS03ser_mux_inst_7_AND1_U1 ( .A1(
        stateArray_nReset_selMC), .A2(stateArray_MUX_inS03ser_mux_inst_7_X), 
        .ZN(stateArray_MUX_inS03ser_mux_inst_7_Y) );
  XOR2_X1 stateArray_MUX_inS03ser_mux_inst_7_XOR2_U1 ( .A(
        stateArray_MUX_inS03ser_mux_inst_7_Y), .B(MixColumns_line1_S02[0]), 
        .Z(stateArray_inS03ser[7]) );
  XOR2_X1 stateArray_MUX_inS13ser_mux_inst_0_XOR1_U1 ( .A(MCin[8]), .B(
        StateInMC[16]), .Z(stateArray_MUX_inS13ser_mux_inst_0_X) );
  AND2_X1 stateArray_MUX_inS13ser_mux_inst_0_AND1_U1 ( .A1(
        stateArray_nReset_selMC), .A2(stateArray_MUX_inS13ser_mux_inst_0_X), 
        .ZN(stateArray_MUX_inS13ser_mux_inst_0_Y) );
  XOR2_X1 stateArray_MUX_inS13ser_mux_inst_0_XOR2_U1 ( .A(
        stateArray_MUX_inS13ser_mux_inst_0_Y), .B(MCin[8]), .Z(
        stateArray_inS13ser[0]) );
  XOR2_X1 stateArray_MUX_inS13ser_mux_inst_1_XOR1_U1 ( .A(
        MixColumns_line2_S02[2]), .B(StateInMC[17]), .Z(
        stateArray_MUX_inS13ser_mux_inst_1_X) );
  AND2_X1 stateArray_MUX_inS13ser_mux_inst_1_AND1_U1 ( .A1(
        stateArray_nReset_selMC), .A2(stateArray_MUX_inS13ser_mux_inst_1_X), 
        .ZN(stateArray_MUX_inS13ser_mux_inst_1_Y) );
  XOR2_X1 stateArray_MUX_inS13ser_mux_inst_1_XOR2_U1 ( .A(
        stateArray_MUX_inS13ser_mux_inst_1_Y), .B(MixColumns_line2_S02[2]), 
        .Z(stateArray_inS13ser[1]) );
  XOR2_X1 stateArray_MUX_inS13ser_mux_inst_2_XOR1_U1 ( .A(MCin[10]), .B(
        StateInMC[18]), .Z(stateArray_MUX_inS13ser_mux_inst_2_X) );
  AND2_X1 stateArray_MUX_inS13ser_mux_inst_2_AND1_U1 ( .A1(
        stateArray_nReset_selMC), .A2(stateArray_MUX_inS13ser_mux_inst_2_X), 
        .ZN(stateArray_MUX_inS13ser_mux_inst_2_Y) );
  XOR2_X1 stateArray_MUX_inS13ser_mux_inst_2_XOR2_U1 ( .A(
        stateArray_MUX_inS13ser_mux_inst_2_Y), .B(MCin[10]), .Z(
        stateArray_inS13ser[2]) );
  XOR2_X1 stateArray_MUX_inS13ser_mux_inst_3_XOR1_U1 ( .A(MCin[11]), .B(
        StateInMC[19]), .Z(stateArray_MUX_inS13ser_mux_inst_3_X) );
  AND2_X1 stateArray_MUX_inS13ser_mux_inst_3_AND1_U1 ( .A1(
        stateArray_nReset_selMC), .A2(stateArray_MUX_inS13ser_mux_inst_3_X), 
        .ZN(stateArray_MUX_inS13ser_mux_inst_3_Y) );
  XOR2_X1 stateArray_MUX_inS13ser_mux_inst_3_XOR2_U1 ( .A(
        stateArray_MUX_inS13ser_mux_inst_3_Y), .B(MCin[11]), .Z(
        stateArray_inS13ser[3]) );
  XOR2_X1 stateArray_MUX_inS13ser_mux_inst_4_XOR1_U1 ( .A(
        MixColumns_line2_S02[5]), .B(StateInMC[20]), .Z(
        stateArray_MUX_inS13ser_mux_inst_4_X) );
  AND2_X1 stateArray_MUX_inS13ser_mux_inst_4_AND1_U1 ( .A1(
        stateArray_nReset_selMC), .A2(stateArray_MUX_inS13ser_mux_inst_4_X), 
        .ZN(stateArray_MUX_inS13ser_mux_inst_4_Y) );
  XOR2_X1 stateArray_MUX_inS13ser_mux_inst_4_XOR2_U1 ( .A(
        stateArray_MUX_inS13ser_mux_inst_4_Y), .B(MixColumns_line2_S02[5]), 
        .Z(stateArray_inS13ser[4]) );
  XOR2_X1 stateArray_MUX_inS13ser_mux_inst_5_XOR1_U1 ( .A(
        MixColumns_line2_S02[6]), .B(StateInMC[21]), .Z(
        stateArray_MUX_inS13ser_mux_inst_5_X) );
  AND2_X1 stateArray_MUX_inS13ser_mux_inst_5_AND1_U1 ( .A1(
        stateArray_nReset_selMC), .A2(stateArray_MUX_inS13ser_mux_inst_5_X), 
        .ZN(stateArray_MUX_inS13ser_mux_inst_5_Y) );
  XOR2_X1 stateArray_MUX_inS13ser_mux_inst_5_XOR2_U1 ( .A(
        stateArray_MUX_inS13ser_mux_inst_5_Y), .B(MixColumns_line2_S02[6]), 
        .Z(stateArray_inS13ser[5]) );
  XOR2_X1 stateArray_MUX_inS13ser_mux_inst_6_XOR1_U1 ( .A(
        MixColumns_line2_S02[7]), .B(StateInMC[22]), .Z(
        stateArray_MUX_inS13ser_mux_inst_6_X) );
  AND2_X1 stateArray_MUX_inS13ser_mux_inst_6_AND1_U1 ( .A1(
        stateArray_nReset_selMC), .A2(stateArray_MUX_inS13ser_mux_inst_6_X), 
        .ZN(stateArray_MUX_inS13ser_mux_inst_6_Y) );
  XOR2_X1 stateArray_MUX_inS13ser_mux_inst_6_XOR2_U1 ( .A(
        stateArray_MUX_inS13ser_mux_inst_6_Y), .B(MixColumns_line2_S02[7]), 
        .Z(stateArray_inS13ser[6]) );
  XOR2_X1 stateArray_MUX_inS13ser_mux_inst_7_XOR1_U1 ( .A(
        MixColumns_line2_S02[0]), .B(StateInMC[23]), .Z(
        stateArray_MUX_inS13ser_mux_inst_7_X) );
  AND2_X1 stateArray_MUX_inS13ser_mux_inst_7_AND1_U1 ( .A1(
        stateArray_nReset_selMC), .A2(stateArray_MUX_inS13ser_mux_inst_7_X), 
        .ZN(stateArray_MUX_inS13ser_mux_inst_7_Y) );
  XOR2_X1 stateArray_MUX_inS13ser_mux_inst_7_XOR2_U1 ( .A(
        stateArray_MUX_inS13ser_mux_inst_7_Y), .B(MixColumns_line2_S02[0]), 
        .Z(stateArray_inS13ser[7]) );
  XOR2_X1 stateArray_MUX_inS23ser_mux_inst_0_XOR1_U1 ( .A(MCin[0]), .B(
        StateInMC[8]), .Z(stateArray_MUX_inS23ser_mux_inst_0_X) );
  AND2_X1 stateArray_MUX_inS23ser_mux_inst_0_AND1_U1 ( .A1(
        stateArray_nReset_selMC), .A2(stateArray_MUX_inS23ser_mux_inst_0_X), 
        .ZN(stateArray_MUX_inS23ser_mux_inst_0_Y) );
  XOR2_X1 stateArray_MUX_inS23ser_mux_inst_0_XOR2_U1 ( .A(
        stateArray_MUX_inS23ser_mux_inst_0_Y), .B(MCin[0]), .Z(
        stateArray_inS23ser[0]) );
  XOR2_X1 stateArray_MUX_inS23ser_mux_inst_1_XOR1_U1 ( .A(
        MixColumns_line3_S02[2]), .B(StateInMC[9]), .Z(
        stateArray_MUX_inS23ser_mux_inst_1_X) );
  AND2_X1 stateArray_MUX_inS23ser_mux_inst_1_AND1_U1 ( .A1(
        stateArray_nReset_selMC), .A2(stateArray_MUX_inS23ser_mux_inst_1_X), 
        .ZN(stateArray_MUX_inS23ser_mux_inst_1_Y) );
  XOR2_X1 stateArray_MUX_inS23ser_mux_inst_1_XOR2_U1 ( .A(
        stateArray_MUX_inS23ser_mux_inst_1_Y), .B(MixColumns_line3_S02[2]), 
        .Z(stateArray_inS23ser[1]) );
  XOR2_X1 stateArray_MUX_inS23ser_mux_inst_2_XOR1_U1 ( .A(MCin[2]), .B(
        StateInMC[10]), .Z(stateArray_MUX_inS23ser_mux_inst_2_X) );
  AND2_X1 stateArray_MUX_inS23ser_mux_inst_2_AND1_U1 ( .A1(
        stateArray_nReset_selMC), .A2(stateArray_MUX_inS23ser_mux_inst_2_X), 
        .ZN(stateArray_MUX_inS23ser_mux_inst_2_Y) );
  XOR2_X1 stateArray_MUX_inS23ser_mux_inst_2_XOR2_U1 ( .A(
        stateArray_MUX_inS23ser_mux_inst_2_Y), .B(MCin[2]), .Z(
        stateArray_inS23ser[2]) );
  XOR2_X1 stateArray_MUX_inS23ser_mux_inst_3_XOR1_U1 ( .A(MCin[3]), .B(
        StateInMC[11]), .Z(stateArray_MUX_inS23ser_mux_inst_3_X) );
  AND2_X1 stateArray_MUX_inS23ser_mux_inst_3_AND1_U1 ( .A1(
        stateArray_nReset_selMC), .A2(stateArray_MUX_inS23ser_mux_inst_3_X), 
        .ZN(stateArray_MUX_inS23ser_mux_inst_3_Y) );
  XOR2_X1 stateArray_MUX_inS23ser_mux_inst_3_XOR2_U1 ( .A(
        stateArray_MUX_inS23ser_mux_inst_3_Y), .B(MCin[3]), .Z(
        stateArray_inS23ser[3]) );
  XOR2_X1 stateArray_MUX_inS23ser_mux_inst_4_XOR1_U1 ( .A(
        MixColumns_line3_S02[5]), .B(StateInMC[12]), .Z(
        stateArray_MUX_inS23ser_mux_inst_4_X) );
  AND2_X1 stateArray_MUX_inS23ser_mux_inst_4_AND1_U1 ( .A1(
        stateArray_nReset_selMC), .A2(stateArray_MUX_inS23ser_mux_inst_4_X), 
        .ZN(stateArray_MUX_inS23ser_mux_inst_4_Y) );
  XOR2_X1 stateArray_MUX_inS23ser_mux_inst_4_XOR2_U1 ( .A(
        stateArray_MUX_inS23ser_mux_inst_4_Y), .B(MixColumns_line3_S02[5]), 
        .Z(stateArray_inS23ser[4]) );
  XOR2_X1 stateArray_MUX_inS23ser_mux_inst_5_XOR1_U1 ( .A(
        MixColumns_line3_S02[6]), .B(StateInMC[13]), .Z(
        stateArray_MUX_inS23ser_mux_inst_5_X) );
  AND2_X1 stateArray_MUX_inS23ser_mux_inst_5_AND1_U1 ( .A1(
        stateArray_nReset_selMC), .A2(stateArray_MUX_inS23ser_mux_inst_5_X), 
        .ZN(stateArray_MUX_inS23ser_mux_inst_5_Y) );
  XOR2_X1 stateArray_MUX_inS23ser_mux_inst_5_XOR2_U1 ( .A(
        stateArray_MUX_inS23ser_mux_inst_5_Y), .B(MixColumns_line3_S02[6]), 
        .Z(stateArray_inS23ser[5]) );
  XOR2_X1 stateArray_MUX_inS23ser_mux_inst_6_XOR1_U1 ( .A(
        MixColumns_line3_S02[7]), .B(StateInMC[14]), .Z(
        stateArray_MUX_inS23ser_mux_inst_6_X) );
  AND2_X1 stateArray_MUX_inS23ser_mux_inst_6_AND1_U1 ( .A1(
        stateArray_nReset_selMC), .A2(stateArray_MUX_inS23ser_mux_inst_6_X), 
        .ZN(stateArray_MUX_inS23ser_mux_inst_6_Y) );
  XOR2_X1 stateArray_MUX_inS23ser_mux_inst_6_XOR2_U1 ( .A(
        stateArray_MUX_inS23ser_mux_inst_6_Y), .B(MixColumns_line3_S02[7]), 
        .Z(stateArray_inS23ser[6]) );
  XOR2_X1 stateArray_MUX_inS23ser_mux_inst_7_XOR1_U1 ( .A(
        MixColumns_line3_S02[0]), .B(StateInMC[15]), .Z(
        stateArray_MUX_inS23ser_mux_inst_7_X) );
  AND2_X1 stateArray_MUX_inS23ser_mux_inst_7_AND1_U1 ( .A1(
        stateArray_nReset_selMC), .A2(stateArray_MUX_inS23ser_mux_inst_7_X), 
        .ZN(stateArray_MUX_inS23ser_mux_inst_7_Y) );
  XOR2_X1 stateArray_MUX_inS23ser_mux_inst_7_XOR2_U1 ( .A(
        stateArray_MUX_inS23ser_mux_inst_7_Y), .B(MixColumns_line3_S02[0]), 
        .Z(stateArray_inS23ser[7]) );
  XOR2_X1 stateArray_MUX_input_MC_mux_inst_0_XOR1_U1 ( .A(StateIn[0]), .B(
        StateInMC[0]), .Z(stateArray_MUX_input_MC_mux_inst_0_X) );
  AND2_X1 stateArray_MUX_input_MC_mux_inst_0_AND1_U1 ( .A1(selMC), .A2(
        stateArray_MUX_input_MC_mux_inst_0_X), .ZN(
        stateArray_MUX_input_MC_mux_inst_0_Y) );
  XOR2_X1 stateArray_MUX_input_MC_mux_inst_0_XOR2_U1 ( .A(
        stateArray_MUX_input_MC_mux_inst_0_Y), .B(StateIn[0]), .Z(
        stateArray_input_MC[0]) );
  XOR2_X1 stateArray_MUX_input_MC_mux_inst_1_XOR1_U1 ( .A(StateIn[1]), .B(
        StateInMC[1]), .Z(stateArray_MUX_input_MC_mux_inst_1_X) );
  AND2_X1 stateArray_MUX_input_MC_mux_inst_1_AND1_U1 ( .A1(selMC), .A2(
        stateArray_MUX_input_MC_mux_inst_1_X), .ZN(
        stateArray_MUX_input_MC_mux_inst_1_Y) );
  XOR2_X1 stateArray_MUX_input_MC_mux_inst_1_XOR2_U1 ( .A(
        stateArray_MUX_input_MC_mux_inst_1_Y), .B(StateIn[1]), .Z(
        stateArray_input_MC[1]) );
  XOR2_X1 stateArray_MUX_input_MC_mux_inst_2_XOR1_U1 ( .A(StateIn[2]), .B(
        StateInMC[2]), .Z(stateArray_MUX_input_MC_mux_inst_2_X) );
  AND2_X1 stateArray_MUX_input_MC_mux_inst_2_AND1_U1 ( .A1(selMC), .A2(
        stateArray_MUX_input_MC_mux_inst_2_X), .ZN(
        stateArray_MUX_input_MC_mux_inst_2_Y) );
  XOR2_X1 stateArray_MUX_input_MC_mux_inst_2_XOR2_U1 ( .A(
        stateArray_MUX_input_MC_mux_inst_2_Y), .B(StateIn[2]), .Z(
        stateArray_input_MC[2]) );
  XOR2_X1 stateArray_MUX_input_MC_mux_inst_3_XOR1_U1 ( .A(StateIn[3]), .B(
        StateInMC[3]), .Z(stateArray_MUX_input_MC_mux_inst_3_X) );
  AND2_X1 stateArray_MUX_input_MC_mux_inst_3_AND1_U1 ( .A1(selMC), .A2(
        stateArray_MUX_input_MC_mux_inst_3_X), .ZN(
        stateArray_MUX_input_MC_mux_inst_3_Y) );
  XOR2_X1 stateArray_MUX_input_MC_mux_inst_3_XOR2_U1 ( .A(
        stateArray_MUX_input_MC_mux_inst_3_Y), .B(StateIn[3]), .Z(
        stateArray_input_MC[3]) );
  XOR2_X1 stateArray_MUX_input_MC_mux_inst_4_XOR1_U1 ( .A(StateIn[4]), .B(
        StateInMC[4]), .Z(stateArray_MUX_input_MC_mux_inst_4_X) );
  AND2_X1 stateArray_MUX_input_MC_mux_inst_4_AND1_U1 ( .A1(selMC), .A2(
        stateArray_MUX_input_MC_mux_inst_4_X), .ZN(
        stateArray_MUX_input_MC_mux_inst_4_Y) );
  XOR2_X1 stateArray_MUX_input_MC_mux_inst_4_XOR2_U1 ( .A(
        stateArray_MUX_input_MC_mux_inst_4_Y), .B(StateIn[4]), .Z(
        stateArray_input_MC[4]) );
  XOR2_X1 stateArray_MUX_input_MC_mux_inst_5_XOR1_U1 ( .A(StateIn[5]), .B(
        StateInMC[5]), .Z(stateArray_MUX_input_MC_mux_inst_5_X) );
  AND2_X1 stateArray_MUX_input_MC_mux_inst_5_AND1_U1 ( .A1(selMC), .A2(
        stateArray_MUX_input_MC_mux_inst_5_X), .ZN(
        stateArray_MUX_input_MC_mux_inst_5_Y) );
  XOR2_X1 stateArray_MUX_input_MC_mux_inst_5_XOR2_U1 ( .A(
        stateArray_MUX_input_MC_mux_inst_5_Y), .B(StateIn[5]), .Z(
        stateArray_input_MC[5]) );
  XOR2_X1 stateArray_MUX_input_MC_mux_inst_6_XOR1_U1 ( .A(StateIn[6]), .B(
        StateInMC[6]), .Z(stateArray_MUX_input_MC_mux_inst_6_X) );
  AND2_X1 stateArray_MUX_input_MC_mux_inst_6_AND1_U1 ( .A1(selMC), .A2(
        stateArray_MUX_input_MC_mux_inst_6_X), .ZN(
        stateArray_MUX_input_MC_mux_inst_6_Y) );
  XOR2_X1 stateArray_MUX_input_MC_mux_inst_6_XOR2_U1 ( .A(
        stateArray_MUX_input_MC_mux_inst_6_Y), .B(StateIn[6]), .Z(
        stateArray_input_MC[6]) );
  XOR2_X1 stateArray_MUX_input_MC_mux_inst_7_XOR1_U1 ( .A(StateIn[7]), .B(
        StateInMC[7]), .Z(stateArray_MUX_input_MC_mux_inst_7_X) );
  AND2_X1 stateArray_MUX_input_MC_mux_inst_7_AND1_U1 ( .A1(selMC), .A2(
        stateArray_MUX_input_MC_mux_inst_7_X), .ZN(
        stateArray_MUX_input_MC_mux_inst_7_Y) );
  XOR2_X1 stateArray_MUX_input_MC_mux_inst_7_XOR2_U1 ( .A(
        stateArray_MUX_input_MC_mux_inst_7_Y), .B(StateIn[7]), .Z(
        stateArray_input_MC[7]) );
  XOR2_X1 stateArray_MUX_inS33ser_mux_inst_0_XOR1_U1 ( .A(port_in[0]), .B(
        stateArray_input_MC[0]), .Z(stateArray_MUX_inS33ser_mux_inst_0_X) );
  AND2_X1 stateArray_MUX_inS33ser_mux_inst_0_AND1_U1 ( .A1(n2), .A2(
        stateArray_MUX_inS33ser_mux_inst_0_X), .ZN(
        stateArray_MUX_inS33ser_mux_inst_0_Y) );
  XOR2_X1 stateArray_MUX_inS33ser_mux_inst_0_XOR2_U1 ( .A(
        stateArray_MUX_inS33ser_mux_inst_0_Y), .B(port_in[0]), .Z(
        stateArray_inS33ser[0]) );
  XOR2_X1 stateArray_MUX_inS33ser_mux_inst_1_XOR1_U1 ( .A(port_in[1]), .B(
        stateArray_input_MC[1]), .Z(stateArray_MUX_inS33ser_mux_inst_1_X) );
  AND2_X1 stateArray_MUX_inS33ser_mux_inst_1_AND1_U1 ( .A1(n2), .A2(
        stateArray_MUX_inS33ser_mux_inst_1_X), .ZN(
        stateArray_MUX_inS33ser_mux_inst_1_Y) );
  XOR2_X1 stateArray_MUX_inS33ser_mux_inst_1_XOR2_U1 ( .A(
        stateArray_MUX_inS33ser_mux_inst_1_Y), .B(port_in[1]), .Z(
        stateArray_inS33ser[1]) );
  XOR2_X1 stateArray_MUX_inS33ser_mux_inst_2_XOR1_U1 ( .A(port_in[2]), .B(
        stateArray_input_MC[2]), .Z(stateArray_MUX_inS33ser_mux_inst_2_X) );
  AND2_X1 stateArray_MUX_inS33ser_mux_inst_2_AND1_U1 ( .A1(n2), .A2(
        stateArray_MUX_inS33ser_mux_inst_2_X), .ZN(
        stateArray_MUX_inS33ser_mux_inst_2_Y) );
  XOR2_X1 stateArray_MUX_inS33ser_mux_inst_2_XOR2_U1 ( .A(
        stateArray_MUX_inS33ser_mux_inst_2_Y), .B(port_in[2]), .Z(
        stateArray_inS33ser[2]) );
  XOR2_X1 stateArray_MUX_inS33ser_mux_inst_3_XOR1_U1 ( .A(port_in[3]), .B(
        stateArray_input_MC[3]), .Z(stateArray_MUX_inS33ser_mux_inst_3_X) );
  AND2_X1 stateArray_MUX_inS33ser_mux_inst_3_AND1_U1 ( .A1(n2), .A2(
        stateArray_MUX_inS33ser_mux_inst_3_X), .ZN(
        stateArray_MUX_inS33ser_mux_inst_3_Y) );
  XOR2_X1 stateArray_MUX_inS33ser_mux_inst_3_XOR2_U1 ( .A(
        stateArray_MUX_inS33ser_mux_inst_3_Y), .B(port_in[3]), .Z(
        stateArray_inS33ser[3]) );
  XOR2_X1 stateArray_MUX_inS33ser_mux_inst_4_XOR1_U1 ( .A(port_in[4]), .B(
        stateArray_input_MC[4]), .Z(stateArray_MUX_inS33ser_mux_inst_4_X) );
  AND2_X1 stateArray_MUX_inS33ser_mux_inst_4_AND1_U1 ( .A1(n2), .A2(
        stateArray_MUX_inS33ser_mux_inst_4_X), .ZN(
        stateArray_MUX_inS33ser_mux_inst_4_Y) );
  XOR2_X1 stateArray_MUX_inS33ser_mux_inst_4_XOR2_U1 ( .A(
        stateArray_MUX_inS33ser_mux_inst_4_Y), .B(port_in[4]), .Z(
        stateArray_inS33ser[4]) );
  XOR2_X1 stateArray_MUX_inS33ser_mux_inst_5_XOR1_U1 ( .A(port_in[5]), .B(
        stateArray_input_MC[5]), .Z(stateArray_MUX_inS33ser_mux_inst_5_X) );
  AND2_X1 stateArray_MUX_inS33ser_mux_inst_5_AND1_U1 ( .A1(n2), .A2(
        stateArray_MUX_inS33ser_mux_inst_5_X), .ZN(
        stateArray_MUX_inS33ser_mux_inst_5_Y) );
  XOR2_X1 stateArray_MUX_inS33ser_mux_inst_5_XOR2_U1 ( .A(
        stateArray_MUX_inS33ser_mux_inst_5_Y), .B(port_in[5]), .Z(
        stateArray_inS33ser[5]) );
  XOR2_X1 stateArray_MUX_inS33ser_mux_inst_6_XOR1_U1 ( .A(port_in[6]), .B(
        stateArray_input_MC[6]), .Z(stateArray_MUX_inS33ser_mux_inst_6_X) );
  AND2_X1 stateArray_MUX_inS33ser_mux_inst_6_AND1_U1 ( .A1(n2), .A2(
        stateArray_MUX_inS33ser_mux_inst_6_X), .ZN(
        stateArray_MUX_inS33ser_mux_inst_6_Y) );
  XOR2_X1 stateArray_MUX_inS33ser_mux_inst_6_XOR2_U1 ( .A(
        stateArray_MUX_inS33ser_mux_inst_6_Y), .B(port_in[6]), .Z(
        stateArray_inS33ser[6]) );
  XOR2_X1 stateArray_MUX_inS33ser_mux_inst_7_XOR1_U1 ( .A(port_in[7]), .B(
        stateArray_input_MC[7]), .Z(stateArray_MUX_inS33ser_mux_inst_7_X) );
  AND2_X1 stateArray_MUX_inS33ser_mux_inst_7_AND1_U1 ( .A1(n2), .A2(
        stateArray_MUX_inS33ser_mux_inst_7_X), .ZN(
        stateArray_MUX_inS33ser_mux_inst_7_Y) );
  XOR2_X1 stateArray_MUX_inS33ser_mux_inst_7_XOR2_U1 ( .A(
        stateArray_MUX_inS33ser_mux_inst_7_Y), .B(port_in[7]), .Z(
        stateArray_inS33ser[7]) );
  INV_X1 MUX_StateInMC_U2 ( .A(intFinal), .ZN(MUX_StateInMC_n4) );
  INV_X1 MUX_StateInMC_U1 ( .A(MUX_StateInMC_n4), .ZN(MUX_StateInMC_n3) );
  XOR2_X1 MUX_StateInMC_mux_inst_0_XOR1_U1 ( .A(MCout[0]), .B(MCin[0]), .Z(
        MUX_StateInMC_mux_inst_0_X) );
  AND2_X1 MUX_StateInMC_mux_inst_0_AND1_U1 ( .A1(MUX_StateInMC_n3), .A2(
        MUX_StateInMC_mux_inst_0_X), .ZN(MUX_StateInMC_mux_inst_0_Y) );
  XOR2_X1 MUX_StateInMC_mux_inst_0_XOR2_U1 ( .A(MUX_StateInMC_mux_inst_0_Y), 
        .B(MCout[0]), .Z(StateInMC[0]) );
  XOR2_X1 MUX_StateInMC_mux_inst_1_XOR1_U1 ( .A(MCout[1]), .B(
        MixColumns_line3_S02[2]), .Z(MUX_StateInMC_mux_inst_1_X) );
  AND2_X1 MUX_StateInMC_mux_inst_1_AND1_U1 ( .A1(MUX_StateInMC_n3), .A2(
        MUX_StateInMC_mux_inst_1_X), .ZN(MUX_StateInMC_mux_inst_1_Y) );
  XOR2_X1 MUX_StateInMC_mux_inst_1_XOR2_U1 ( .A(MUX_StateInMC_mux_inst_1_Y), 
        .B(MCout[1]), .Z(StateInMC[1]) );
  XOR2_X1 MUX_StateInMC_mux_inst_2_XOR1_U1 ( .A(MCout[2]), .B(MCin[2]), .Z(
        MUX_StateInMC_mux_inst_2_X) );
  AND2_X1 MUX_StateInMC_mux_inst_2_AND1_U1 ( .A1(MUX_StateInMC_n3), .A2(
        MUX_StateInMC_mux_inst_2_X), .ZN(MUX_StateInMC_mux_inst_2_Y) );
  XOR2_X1 MUX_StateInMC_mux_inst_2_XOR2_U1 ( .A(MUX_StateInMC_mux_inst_2_Y), 
        .B(MCout[2]), .Z(StateInMC[2]) );
  XOR2_X1 MUX_StateInMC_mux_inst_3_XOR1_U1 ( .A(MCout[3]), .B(MCin[3]), .Z(
        MUX_StateInMC_mux_inst_3_X) );
  AND2_X1 MUX_StateInMC_mux_inst_3_AND1_U1 ( .A1(MUX_StateInMC_n3), .A2(
        MUX_StateInMC_mux_inst_3_X), .ZN(MUX_StateInMC_mux_inst_3_Y) );
  XOR2_X1 MUX_StateInMC_mux_inst_3_XOR2_U1 ( .A(MUX_StateInMC_mux_inst_3_Y), 
        .B(MCout[3]), .Z(StateInMC[3]) );
  XOR2_X1 MUX_StateInMC_mux_inst_4_XOR1_U1 ( .A(MCout[4]), .B(
        MixColumns_line3_S02[5]), .Z(MUX_StateInMC_mux_inst_4_X) );
  AND2_X1 MUX_StateInMC_mux_inst_4_AND1_U1 ( .A1(MUX_StateInMC_n3), .A2(
        MUX_StateInMC_mux_inst_4_X), .ZN(MUX_StateInMC_mux_inst_4_Y) );
  XOR2_X1 MUX_StateInMC_mux_inst_4_XOR2_U1 ( .A(MUX_StateInMC_mux_inst_4_Y), 
        .B(MCout[4]), .Z(StateInMC[4]) );
  XOR2_X1 MUX_StateInMC_mux_inst_5_XOR1_U1 ( .A(MCout[5]), .B(
        MixColumns_line3_S02[6]), .Z(MUX_StateInMC_mux_inst_5_X) );
  AND2_X1 MUX_StateInMC_mux_inst_5_AND1_U1 ( .A1(MUX_StateInMC_n3), .A2(
        MUX_StateInMC_mux_inst_5_X), .ZN(MUX_StateInMC_mux_inst_5_Y) );
  XOR2_X1 MUX_StateInMC_mux_inst_5_XOR2_U1 ( .A(MUX_StateInMC_mux_inst_5_Y), 
        .B(MCout[5]), .Z(StateInMC[5]) );
  XOR2_X1 MUX_StateInMC_mux_inst_6_XOR1_U1 ( .A(MCout[6]), .B(
        MixColumns_line3_S02[7]), .Z(MUX_StateInMC_mux_inst_6_X) );
  AND2_X1 MUX_StateInMC_mux_inst_6_AND1_U1 ( .A1(MUX_StateInMC_n3), .A2(
        MUX_StateInMC_mux_inst_6_X), .ZN(MUX_StateInMC_mux_inst_6_Y) );
  XOR2_X1 MUX_StateInMC_mux_inst_6_XOR2_U1 ( .A(MUX_StateInMC_mux_inst_6_Y), 
        .B(MCout[6]), .Z(StateInMC[6]) );
  XOR2_X1 MUX_StateInMC_mux_inst_7_XOR1_U1 ( .A(MCout[7]), .B(
        MixColumns_line3_S02[0]), .Z(MUX_StateInMC_mux_inst_7_X) );
  AND2_X1 MUX_StateInMC_mux_inst_7_AND1_U1 ( .A1(MUX_StateInMC_n3), .A2(
        MUX_StateInMC_mux_inst_7_X), .ZN(MUX_StateInMC_mux_inst_7_Y) );
  XOR2_X1 MUX_StateInMC_mux_inst_7_XOR2_U1 ( .A(MUX_StateInMC_mux_inst_7_Y), 
        .B(MCout[7]), .Z(StateInMC[7]) );
  XOR2_X1 MUX_StateInMC_mux_inst_8_XOR1_U1 ( .A(MCout[8]), .B(MCin[8]), .Z(
        MUX_StateInMC_mux_inst_8_X) );
  AND2_X1 MUX_StateInMC_mux_inst_8_AND1_U1 ( .A1(MUX_StateInMC_n3), .A2(
        MUX_StateInMC_mux_inst_8_X), .ZN(MUX_StateInMC_mux_inst_8_Y) );
  XOR2_X1 MUX_StateInMC_mux_inst_8_XOR2_U1 ( .A(MUX_StateInMC_mux_inst_8_Y), 
        .B(MCout[8]), .Z(StateInMC[8]) );
  XOR2_X1 MUX_StateInMC_mux_inst_9_XOR1_U1 ( .A(MCout[9]), .B(
        MixColumns_line2_S02[2]), .Z(MUX_StateInMC_mux_inst_9_X) );
  AND2_X1 MUX_StateInMC_mux_inst_9_AND1_U1 ( .A1(MUX_StateInMC_n3), .A2(
        MUX_StateInMC_mux_inst_9_X), .ZN(MUX_StateInMC_mux_inst_9_Y) );
  XOR2_X1 MUX_StateInMC_mux_inst_9_XOR2_U1 ( .A(MUX_StateInMC_mux_inst_9_Y), 
        .B(MCout[9]), .Z(StateInMC[9]) );
  XOR2_X1 MUX_StateInMC_mux_inst_10_XOR1_U1 ( .A(MCout[10]), .B(MCin[10]), .Z(
        MUX_StateInMC_mux_inst_10_X) );
  AND2_X1 MUX_StateInMC_mux_inst_10_AND1_U1 ( .A1(MUX_StateInMC_n3), .A2(
        MUX_StateInMC_mux_inst_10_X), .ZN(MUX_StateInMC_mux_inst_10_Y) );
  XOR2_X1 MUX_StateInMC_mux_inst_10_XOR2_U1 ( .A(MUX_StateInMC_mux_inst_10_Y), 
        .B(MCout[10]), .Z(StateInMC[10]) );
  XOR2_X1 MUX_StateInMC_mux_inst_11_XOR1_U1 ( .A(MCout[11]), .B(MCin[11]), .Z(
        MUX_StateInMC_mux_inst_11_X) );
  AND2_X1 MUX_StateInMC_mux_inst_11_AND1_U1 ( .A1(MUX_StateInMC_n3), .A2(
        MUX_StateInMC_mux_inst_11_X), .ZN(MUX_StateInMC_mux_inst_11_Y) );
  XOR2_X1 MUX_StateInMC_mux_inst_11_XOR2_U1 ( .A(MUX_StateInMC_mux_inst_11_Y), 
        .B(MCout[11]), .Z(StateInMC[11]) );
  XOR2_X1 MUX_StateInMC_mux_inst_12_XOR1_U1 ( .A(MCout[12]), .B(
        MixColumns_line2_S02[5]), .Z(MUX_StateInMC_mux_inst_12_X) );
  AND2_X1 MUX_StateInMC_mux_inst_12_AND1_U1 ( .A1(MUX_StateInMC_n3), .A2(
        MUX_StateInMC_mux_inst_12_X), .ZN(MUX_StateInMC_mux_inst_12_Y) );
  XOR2_X1 MUX_StateInMC_mux_inst_12_XOR2_U1 ( .A(MUX_StateInMC_mux_inst_12_Y), 
        .B(MCout[12]), .Z(StateInMC[12]) );
  XOR2_X1 MUX_StateInMC_mux_inst_13_XOR1_U1 ( .A(MCout[13]), .B(
        MixColumns_line2_S02[6]), .Z(MUX_StateInMC_mux_inst_13_X) );
  AND2_X1 MUX_StateInMC_mux_inst_13_AND1_U1 ( .A1(MUX_StateInMC_n3), .A2(
        MUX_StateInMC_mux_inst_13_X), .ZN(MUX_StateInMC_mux_inst_13_Y) );
  XOR2_X1 MUX_StateInMC_mux_inst_13_XOR2_U1 ( .A(MUX_StateInMC_mux_inst_13_Y), 
        .B(MCout[13]), .Z(StateInMC[13]) );
  XOR2_X1 MUX_StateInMC_mux_inst_14_XOR1_U1 ( .A(MCout[14]), .B(
        MixColumns_line2_S02[7]), .Z(MUX_StateInMC_mux_inst_14_X) );
  AND2_X1 MUX_StateInMC_mux_inst_14_AND1_U1 ( .A1(MUX_StateInMC_n3), .A2(
        MUX_StateInMC_mux_inst_14_X), .ZN(MUX_StateInMC_mux_inst_14_Y) );
  XOR2_X1 MUX_StateInMC_mux_inst_14_XOR2_U1 ( .A(MUX_StateInMC_mux_inst_14_Y), 
        .B(MCout[14]), .Z(StateInMC[14]) );
  XOR2_X1 MUX_StateInMC_mux_inst_15_XOR1_U1 ( .A(MCout[15]), .B(
        MixColumns_line2_S02[0]), .Z(MUX_StateInMC_mux_inst_15_X) );
  AND2_X1 MUX_StateInMC_mux_inst_15_AND1_U1 ( .A1(MUX_StateInMC_n3), .A2(
        MUX_StateInMC_mux_inst_15_X), .ZN(MUX_StateInMC_mux_inst_15_Y) );
  XOR2_X1 MUX_StateInMC_mux_inst_15_XOR2_U1 ( .A(MUX_StateInMC_mux_inst_15_Y), 
        .B(MCout[15]), .Z(StateInMC[15]) );
  XOR2_X1 MUX_StateInMC_mux_inst_16_XOR1_U1 ( .A(MCout[16]), .B(MCin[16]), .Z(
        MUX_StateInMC_mux_inst_16_X) );
  AND2_X1 MUX_StateInMC_mux_inst_16_AND1_U1 ( .A1(MUX_StateInMC_n3), .A2(
        MUX_StateInMC_mux_inst_16_X), .ZN(MUX_StateInMC_mux_inst_16_Y) );
  XOR2_X1 MUX_StateInMC_mux_inst_16_XOR2_U1 ( .A(MUX_StateInMC_mux_inst_16_Y), 
        .B(MCout[16]), .Z(StateInMC[16]) );
  XOR2_X1 MUX_StateInMC_mux_inst_17_XOR1_U1 ( .A(MCout[17]), .B(
        MixColumns_line1_S02[2]), .Z(MUX_StateInMC_mux_inst_17_X) );
  AND2_X1 MUX_StateInMC_mux_inst_17_AND1_U1 ( .A1(MUX_StateInMC_n3), .A2(
        MUX_StateInMC_mux_inst_17_X), .ZN(MUX_StateInMC_mux_inst_17_Y) );
  XOR2_X1 MUX_StateInMC_mux_inst_17_XOR2_U1 ( .A(MUX_StateInMC_mux_inst_17_Y), 
        .B(MCout[17]), .Z(StateInMC[17]) );
  XOR2_X1 MUX_StateInMC_mux_inst_18_XOR1_U1 ( .A(MCout[18]), .B(MCin[18]), .Z(
        MUX_StateInMC_mux_inst_18_X) );
  AND2_X1 MUX_StateInMC_mux_inst_18_AND1_U1 ( .A1(MUX_StateInMC_n3), .A2(
        MUX_StateInMC_mux_inst_18_X), .ZN(MUX_StateInMC_mux_inst_18_Y) );
  XOR2_X1 MUX_StateInMC_mux_inst_18_XOR2_U1 ( .A(MUX_StateInMC_mux_inst_18_Y), 
        .B(MCout[18]), .Z(StateInMC[18]) );
  XOR2_X1 MUX_StateInMC_mux_inst_19_XOR1_U1 ( .A(MCout[19]), .B(MCin[19]), .Z(
        MUX_StateInMC_mux_inst_19_X) );
  AND2_X1 MUX_StateInMC_mux_inst_19_AND1_U1 ( .A1(MUX_StateInMC_n3), .A2(
        MUX_StateInMC_mux_inst_19_X), .ZN(MUX_StateInMC_mux_inst_19_Y) );
  XOR2_X1 MUX_StateInMC_mux_inst_19_XOR2_U1 ( .A(MUX_StateInMC_mux_inst_19_Y), 
        .B(MCout[19]), .Z(StateInMC[19]) );
  XOR2_X1 MUX_StateInMC_mux_inst_20_XOR1_U1 ( .A(MCout[20]), .B(
        MixColumns_line1_S02[5]), .Z(MUX_StateInMC_mux_inst_20_X) );
  AND2_X1 MUX_StateInMC_mux_inst_20_AND1_U1 ( .A1(intFinal), .A2(
        MUX_StateInMC_mux_inst_20_X), .ZN(MUX_StateInMC_mux_inst_20_Y) );
  XOR2_X1 MUX_StateInMC_mux_inst_20_XOR2_U1 ( .A(MUX_StateInMC_mux_inst_20_Y), 
        .B(MCout[20]), .Z(StateInMC[20]) );
  XOR2_X1 MUX_StateInMC_mux_inst_21_XOR1_U1 ( .A(MCout[21]), .B(
        MixColumns_line1_S02[6]), .Z(MUX_StateInMC_mux_inst_21_X) );
  AND2_X1 MUX_StateInMC_mux_inst_21_AND1_U1 ( .A1(MUX_StateInMC_n3), .A2(
        MUX_StateInMC_mux_inst_21_X), .ZN(MUX_StateInMC_mux_inst_21_Y) );
  XOR2_X1 MUX_StateInMC_mux_inst_21_XOR2_U1 ( .A(MUX_StateInMC_mux_inst_21_Y), 
        .B(MCout[21]), .Z(StateInMC[21]) );
  XOR2_X1 MUX_StateInMC_mux_inst_22_XOR1_U1 ( .A(MCout[22]), .B(
        MixColumns_line1_S02[7]), .Z(MUX_StateInMC_mux_inst_22_X) );
  AND2_X1 MUX_StateInMC_mux_inst_22_AND1_U1 ( .A1(MUX_StateInMC_n3), .A2(
        MUX_StateInMC_mux_inst_22_X), .ZN(MUX_StateInMC_mux_inst_22_Y) );
  XOR2_X1 MUX_StateInMC_mux_inst_22_XOR2_U1 ( .A(MUX_StateInMC_mux_inst_22_Y), 
        .B(MCout[22]), .Z(StateInMC[22]) );
  XOR2_X1 MUX_StateInMC_mux_inst_23_XOR1_U1 ( .A(MCout[23]), .B(
        MixColumns_line1_S02[0]), .Z(MUX_StateInMC_mux_inst_23_X) );
  AND2_X1 MUX_StateInMC_mux_inst_23_AND1_U1 ( .A1(MUX_StateInMC_n3), .A2(
        MUX_StateInMC_mux_inst_23_X), .ZN(MUX_StateInMC_mux_inst_23_Y) );
  XOR2_X1 MUX_StateInMC_mux_inst_23_XOR2_U1 ( .A(MUX_StateInMC_mux_inst_23_Y), 
        .B(MCout[23]), .Z(StateInMC[23]) );
  XOR2_X1 MUX_StateInMC_mux_inst_24_XOR1_U1 ( .A(MCout[24]), .B(port_out[0]), 
        .Z(MUX_StateInMC_mux_inst_24_X) );
  AND2_X1 MUX_StateInMC_mux_inst_24_AND1_U1 ( .A1(intFinal), .A2(
        MUX_StateInMC_mux_inst_24_X), .ZN(MUX_StateInMC_mux_inst_24_Y) );
  XOR2_X1 MUX_StateInMC_mux_inst_24_XOR2_U1 ( .A(MUX_StateInMC_mux_inst_24_Y), 
        .B(MCout[24]), .Z(StateInMC[24]) );
  XOR2_X1 MUX_StateInMC_mux_inst_25_XOR1_U1 ( .A(MCout[25]), .B(port_out[1]), 
        .Z(MUX_StateInMC_mux_inst_25_X) );
  AND2_X1 MUX_StateInMC_mux_inst_25_AND1_U1 ( .A1(intFinal), .A2(
        MUX_StateInMC_mux_inst_25_X), .ZN(MUX_StateInMC_mux_inst_25_Y) );
  XOR2_X1 MUX_StateInMC_mux_inst_25_XOR2_U1 ( .A(MUX_StateInMC_mux_inst_25_Y), 
        .B(MCout[25]), .Z(StateInMC[25]) );
  XOR2_X1 MUX_StateInMC_mux_inst_26_XOR1_U1 ( .A(MCout[26]), .B(port_out[2]), 
        .Z(MUX_StateInMC_mux_inst_26_X) );
  AND2_X1 MUX_StateInMC_mux_inst_26_AND1_U1 ( .A1(intFinal), .A2(
        MUX_StateInMC_mux_inst_26_X), .ZN(MUX_StateInMC_mux_inst_26_Y) );
  XOR2_X1 MUX_StateInMC_mux_inst_26_XOR2_U1 ( .A(MUX_StateInMC_mux_inst_26_Y), 
        .B(MCout[26]), .Z(StateInMC[26]) );
  XOR2_X1 MUX_StateInMC_mux_inst_27_XOR1_U1 ( .A(MCout[27]), .B(port_out[3]), 
        .Z(MUX_StateInMC_mux_inst_27_X) );
  AND2_X1 MUX_StateInMC_mux_inst_27_AND1_U1 ( .A1(intFinal), .A2(
        MUX_StateInMC_mux_inst_27_X), .ZN(MUX_StateInMC_mux_inst_27_Y) );
  XOR2_X1 MUX_StateInMC_mux_inst_27_XOR2_U1 ( .A(MUX_StateInMC_mux_inst_27_Y), 
        .B(MCout[27]), .Z(StateInMC[27]) );
  XOR2_X1 MUX_StateInMC_mux_inst_28_XOR1_U1 ( .A(MCout[28]), .B(port_out[4]), 
        .Z(MUX_StateInMC_mux_inst_28_X) );
  AND2_X1 MUX_StateInMC_mux_inst_28_AND1_U1 ( .A1(MUX_StateInMC_n3), .A2(
        MUX_StateInMC_mux_inst_28_X), .ZN(MUX_StateInMC_mux_inst_28_Y) );
  XOR2_X1 MUX_StateInMC_mux_inst_28_XOR2_U1 ( .A(MUX_StateInMC_mux_inst_28_Y), 
        .B(MCout[28]), .Z(StateInMC[28]) );
  XOR2_X1 MUX_StateInMC_mux_inst_29_XOR1_U1 ( .A(MCout[29]), .B(port_out[5]), 
        .Z(MUX_StateInMC_mux_inst_29_X) );
  AND2_X1 MUX_StateInMC_mux_inst_29_AND1_U1 ( .A1(MUX_StateInMC_n3), .A2(
        MUX_StateInMC_mux_inst_29_X), .ZN(MUX_StateInMC_mux_inst_29_Y) );
  XOR2_X1 MUX_StateInMC_mux_inst_29_XOR2_U1 ( .A(MUX_StateInMC_mux_inst_29_Y), 
        .B(MCout[29]), .Z(StateInMC[29]) );
  XOR2_X1 MUX_StateInMC_mux_inst_30_XOR1_U1 ( .A(MCout[30]), .B(port_out[6]), 
        .Z(MUX_StateInMC_mux_inst_30_X) );
  AND2_X1 MUX_StateInMC_mux_inst_30_AND1_U1 ( .A1(MUX_StateInMC_n3), .A2(
        MUX_StateInMC_mux_inst_30_X), .ZN(MUX_StateInMC_mux_inst_30_Y) );
  XOR2_X1 MUX_StateInMC_mux_inst_30_XOR2_U1 ( .A(MUX_StateInMC_mux_inst_30_Y), 
        .B(MCout[30]), .Z(StateInMC[30]) );
  XOR2_X1 MUX_StateInMC_mux_inst_31_XOR1_U1 ( .A(MCout[31]), .B(port_out[7]), 
        .Z(MUX_StateInMC_mux_inst_31_X) );
  AND2_X1 MUX_StateInMC_mux_inst_31_AND1_U1 ( .A1(MUX_StateInMC_n3), .A2(
        MUX_StateInMC_mux_inst_31_X), .ZN(MUX_StateInMC_mux_inst_31_Y) );
  XOR2_X1 MUX_StateInMC_mux_inst_31_XOR2_U1 ( .A(MUX_StateInMC_mux_inst_31_Y), 
        .B(MCout[31]), .Z(StateInMC[31]) );
  XOR2_X1 KeyArray_U32 ( .A(KeyArray_outS01ser_7_), .B(keyStateIn[7]), .Z(
        KeyArray_outS01ser_XOR_00[7]) );
  XOR2_X1 KeyArray_U31 ( .A(KeyArray_outS01ser_6_), .B(keyStateIn[6]), .Z(
        KeyArray_outS01ser_XOR_00[6]) );
  XOR2_X1 KeyArray_U30 ( .A(KeyArray_outS01ser_5_), .B(keyStateIn[5]), .Z(
        KeyArray_outS01ser_XOR_00[5]) );
  XOR2_X1 KeyArray_U29 ( .A(KeyArray_outS01ser_4_), .B(keyStateIn[4]), .Z(
        KeyArray_outS01ser_XOR_00[4]) );
  XOR2_X1 KeyArray_U28 ( .A(KeyArray_outS01ser_3_), .B(keyStateIn[3]), .Z(
        KeyArray_outS01ser_XOR_00[3]) );
  XOR2_X1 KeyArray_U27 ( .A(KeyArray_outS01ser_2_), .B(keyStateIn[2]), .Z(
        KeyArray_outS01ser_XOR_00[2]) );
  XOR2_X1 KeyArray_U26 ( .A(KeyArray_outS01ser_1_), .B(keyStateIn[1]), .Z(
        KeyArray_outS01ser_XOR_00[1]) );
  XOR2_X1 KeyArray_U25 ( .A(KeyArray_outS01ser_0_), .B(keyStateIn[0]), .Z(
        KeyArray_outS01ser_XOR_00[0]) );
  AND2_X1 KeyArray_U24 ( .A1(n2), .A2(intselXOR), .ZN(KeyArray_nReset_selXOR)
         );
  XNOR2_X1 KeyArray_U23 ( .A(KeyArray_n32), .B(keyStateIn[7]), .ZN(
        KeyArray_inS30par[7]) );
  XNOR2_X1 KeyArray_U22 ( .A(roundConstant[7]), .B(SboxOut[7]), .ZN(
        KeyArray_n32) );
  XNOR2_X1 KeyArray_U21 ( .A(KeyArray_n31), .B(keyStateIn[6]), .ZN(
        KeyArray_inS30par[6]) );
  XNOR2_X1 KeyArray_U20 ( .A(roundConstant[6]), .B(SboxOut[6]), .ZN(
        KeyArray_n31) );
  XNOR2_X1 KeyArray_U19 ( .A(KeyArray_n30), .B(keyStateIn[5]), .ZN(
        KeyArray_inS30par[5]) );
  XNOR2_X1 KeyArray_U18 ( .A(roundConstant[5]), .B(SboxOut[5]), .ZN(
        KeyArray_n30) );
  XNOR2_X1 KeyArray_U17 ( .A(KeyArray_n29), .B(keyStateIn[4]), .ZN(
        KeyArray_inS30par[4]) );
  XNOR2_X1 KeyArray_U16 ( .A(roundConstant[4]), .B(SboxOut[4]), .ZN(
        KeyArray_n29) );
  XNOR2_X1 KeyArray_U15 ( .A(KeyArray_n28), .B(keyStateIn[3]), .ZN(
        KeyArray_inS30par[3]) );
  XNOR2_X1 KeyArray_U14 ( .A(roundConstant[3]), .B(SboxOut[3]), .ZN(
        KeyArray_n28) );
  XNOR2_X1 KeyArray_U13 ( .A(KeyArray_n27), .B(keyStateIn[2]), .ZN(
        KeyArray_inS30par[2]) );
  XNOR2_X1 KeyArray_U12 ( .A(roundConstant[2]), .B(SboxOut[2]), .ZN(
        KeyArray_n27) );
  XNOR2_X1 KeyArray_U11 ( .A(KeyArray_n26), .B(keyStateIn[1]), .ZN(
        KeyArray_inS30par[1]) );
  XNOR2_X1 KeyArray_U10 ( .A(roundConstant[1]), .B(SboxOut[1]), .ZN(
        KeyArray_n26) );
  XNOR2_X1 KeyArray_U9 ( .A(KeyArray_n25), .B(keyStateIn[0]), .ZN(
        KeyArray_inS30par[0]) );
  XNOR2_X1 KeyArray_U8 ( .A(roundConstant[0]), .B(SboxOut[0]), .ZN(
        KeyArray_n25) );
  INV_X2 KeyArray_U7 ( .A(KeyArray_n24), .ZN(KeyArray_n21) );
  INV_X2 KeyArray_U6 ( .A(KeyArray_n24), .ZN(KeyArray_n22) );
  INV_X1 KeyArray_U5 ( .A(selMC), .ZN(KeyArray_n24) );
  INV_X1 KeyArray_U4 ( .A(KeyArray_n24), .ZN(KeyArray_n23) );
  INV_X4 KeyArray_U3 ( .A(KeyArray_n20), .ZN(KeyArray_n19) );
  INV_X1 KeyArray_U2 ( .A(enKS), .ZN(KeyArray_n20) );
  INV_X8 KeyArray_U1 ( .A(KeyArray_n20), .ZN(KeyArray_n18) );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_0_U3 ( .A1(KeyArray_S00reg_gff_1_SFF_0_n2), .A2(KeyArray_S00reg_gff_1_SFF_0_n1), .ZN(KeyArray_S00reg_gff_1_SFF_0_n6) );
  OR2_X1 KeyArray_S00reg_gff_1_SFF_0_U2 ( .A1(KeyArray_n19), .A2(
        KeyArray_S00reg_gff_1_SFF_0_n3), .ZN(KeyArray_S00reg_gff_1_SFF_0_n1)
         );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_0_U1 ( .A1(KeyArray_S00reg_gff_1_SFF_0_QD), .A2(KeyArray_n19), .ZN(KeyArray_S00reg_gff_1_SFF_0_n2) );
  XOR2_X1 KeyArray_S00reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A(
        KeyArray_inS00ser[0]), .B(KeyArray_outS10ser[0]), .Z(
        KeyArray_S00reg_gff_1_SFF_0_MUXInst_X) );
  AND2_X1 KeyArray_S00reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A1(KeyArray_n23), 
        .A2(KeyArray_S00reg_gff_1_SFF_0_MUXInst_X), .ZN(
        KeyArray_S00reg_gff_1_SFF_0_MUXInst_Y) );
  XOR2_X1 KeyArray_S00reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A(
        KeyArray_S00reg_gff_1_SFF_0_MUXInst_Y), .B(KeyArray_inS00ser[0]), .Z(
        KeyArray_S00reg_gff_1_SFF_0_QD) );
  INV_X1 KeyArray_S00reg_gff_1_SFF_0_Q_reg_U1 ( .A(keyStateIn[0]), .ZN(
        KeyArray_S00reg_gff_1_SFF_0_n3) );
  DFF_X1 KeyArray_S00reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        KeyArray_S00reg_gff_1_SFF_0_n6), .CK(clk), .Q(keyStateIn[0]), .QN() );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_1_U3 ( .A1(KeyArray_S00reg_gff_1_SFF_1_n2), .A2(KeyArray_S00reg_gff_1_SFF_1_n1), .ZN(KeyArray_S00reg_gff_1_SFF_1_n6) );
  OR2_X1 KeyArray_S00reg_gff_1_SFF_1_U2 ( .A1(KeyArray_n19), .A2(
        KeyArray_S00reg_gff_1_SFF_1_n11), .ZN(KeyArray_S00reg_gff_1_SFF_1_n1)
         );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_1_U1 ( .A1(KeyArray_S00reg_gff_1_SFF_1_QD), .A2(KeyArray_n19), .ZN(KeyArray_S00reg_gff_1_SFF_1_n2) );
  XOR2_X1 KeyArray_S00reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A(
        KeyArray_inS00ser[1]), .B(KeyArray_outS10ser[1]), .Z(
        KeyArray_S00reg_gff_1_SFF_1_MUXInst_X) );
  AND2_X1 KeyArray_S00reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A1(KeyArray_n23), 
        .A2(KeyArray_S00reg_gff_1_SFF_1_MUXInst_X), .ZN(
        KeyArray_S00reg_gff_1_SFF_1_MUXInst_Y) );
  XOR2_X1 KeyArray_S00reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A(
        KeyArray_S00reg_gff_1_SFF_1_MUXInst_Y), .B(KeyArray_inS00ser[1]), .Z(
        KeyArray_S00reg_gff_1_SFF_1_QD) );
  INV_X1 KeyArray_S00reg_gff_1_SFF_1_Q_reg_U1 ( .A(keyStateIn[1]), .ZN(
        KeyArray_S00reg_gff_1_SFF_1_n11) );
  DFF_X1 KeyArray_S00reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        KeyArray_S00reg_gff_1_SFF_1_n6), .CK(clk), .Q(keyStateIn[1]), .QN() );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_2_U3 ( .A1(KeyArray_S00reg_gff_1_SFF_2_n2), .A2(KeyArray_S00reg_gff_1_SFF_2_n1), .ZN(KeyArray_S00reg_gff_1_SFF_2_n6) );
  OR2_X1 KeyArray_S00reg_gff_1_SFF_2_U2 ( .A1(KeyArray_n19), .A2(
        KeyArray_S00reg_gff_1_SFF_2_n11), .ZN(KeyArray_S00reg_gff_1_SFF_2_n1)
         );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_2_U1 ( .A1(KeyArray_S00reg_gff_1_SFF_2_QD), .A2(KeyArray_n19), .ZN(KeyArray_S00reg_gff_1_SFF_2_n2) );
  XOR2_X1 KeyArray_S00reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A(
        KeyArray_inS00ser[2]), .B(KeyArray_outS10ser[2]), .Z(
        KeyArray_S00reg_gff_1_SFF_2_MUXInst_X) );
  AND2_X1 KeyArray_S00reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A1(KeyArray_n23), 
        .A2(KeyArray_S00reg_gff_1_SFF_2_MUXInst_X), .ZN(
        KeyArray_S00reg_gff_1_SFF_2_MUXInst_Y) );
  XOR2_X1 KeyArray_S00reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A(
        KeyArray_S00reg_gff_1_SFF_2_MUXInst_Y), .B(KeyArray_inS00ser[2]), .Z(
        KeyArray_S00reg_gff_1_SFF_2_QD) );
  INV_X1 KeyArray_S00reg_gff_1_SFF_2_Q_reg_U1 ( .A(keyStateIn[2]), .ZN(
        KeyArray_S00reg_gff_1_SFF_2_n11) );
  DFF_X1 KeyArray_S00reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        KeyArray_S00reg_gff_1_SFF_2_n6), .CK(clk), .Q(keyStateIn[2]), .QN() );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_3_U3 ( .A1(KeyArray_S00reg_gff_1_SFF_3_n2), .A2(KeyArray_S00reg_gff_1_SFF_3_n1), .ZN(KeyArray_S00reg_gff_1_SFF_3_n6) );
  OR2_X1 KeyArray_S00reg_gff_1_SFF_3_U2 ( .A1(KeyArray_n19), .A2(
        KeyArray_S00reg_gff_1_SFF_3_n11), .ZN(KeyArray_S00reg_gff_1_SFF_3_n1)
         );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_3_U1 ( .A1(KeyArray_S00reg_gff_1_SFF_3_QD), .A2(KeyArray_n19), .ZN(KeyArray_S00reg_gff_1_SFF_3_n2) );
  XOR2_X1 KeyArray_S00reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A(
        KeyArray_inS00ser[3]), .B(KeyArray_outS10ser[3]), .Z(
        KeyArray_S00reg_gff_1_SFF_3_MUXInst_X) );
  AND2_X1 KeyArray_S00reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A1(KeyArray_n23), 
        .A2(KeyArray_S00reg_gff_1_SFF_3_MUXInst_X), .ZN(
        KeyArray_S00reg_gff_1_SFF_3_MUXInst_Y) );
  XOR2_X1 KeyArray_S00reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A(
        KeyArray_S00reg_gff_1_SFF_3_MUXInst_Y), .B(KeyArray_inS00ser[3]), .Z(
        KeyArray_S00reg_gff_1_SFF_3_QD) );
  INV_X1 KeyArray_S00reg_gff_1_SFF_3_Q_reg_U1 ( .A(keyStateIn[3]), .ZN(
        KeyArray_S00reg_gff_1_SFF_3_n11) );
  DFF_X1 KeyArray_S00reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        KeyArray_S00reg_gff_1_SFF_3_n6), .CK(clk), .Q(keyStateIn[3]), .QN() );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_4_U3 ( .A1(KeyArray_S00reg_gff_1_SFF_4_n2), .A2(KeyArray_S00reg_gff_1_SFF_4_n1), .ZN(KeyArray_S00reg_gff_1_SFF_4_n6) );
  OR2_X1 KeyArray_S00reg_gff_1_SFF_4_U2 ( .A1(KeyArray_n19), .A2(
        KeyArray_S00reg_gff_1_SFF_4_n11), .ZN(KeyArray_S00reg_gff_1_SFF_4_n1)
         );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_4_U1 ( .A1(KeyArray_S00reg_gff_1_SFF_4_QD), .A2(KeyArray_n19), .ZN(KeyArray_S00reg_gff_1_SFF_4_n2) );
  XOR2_X1 KeyArray_S00reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A(
        KeyArray_inS00ser[4]), .B(KeyArray_outS10ser[4]), .Z(
        KeyArray_S00reg_gff_1_SFF_4_MUXInst_X) );
  AND2_X1 KeyArray_S00reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A1(KeyArray_n23), 
        .A2(KeyArray_S00reg_gff_1_SFF_4_MUXInst_X), .ZN(
        KeyArray_S00reg_gff_1_SFF_4_MUXInst_Y) );
  XOR2_X1 KeyArray_S00reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A(
        KeyArray_S00reg_gff_1_SFF_4_MUXInst_Y), .B(KeyArray_inS00ser[4]), .Z(
        KeyArray_S00reg_gff_1_SFF_4_QD) );
  INV_X1 KeyArray_S00reg_gff_1_SFF_4_Q_reg_U1 ( .A(keyStateIn[4]), .ZN(
        KeyArray_S00reg_gff_1_SFF_4_n11) );
  DFF_X1 KeyArray_S00reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        KeyArray_S00reg_gff_1_SFF_4_n6), .CK(clk), .Q(keyStateIn[4]), .QN() );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_5_U3 ( .A1(KeyArray_S00reg_gff_1_SFF_5_n2), .A2(KeyArray_S00reg_gff_1_SFF_5_n1), .ZN(KeyArray_S00reg_gff_1_SFF_5_n6) );
  OR2_X1 KeyArray_S00reg_gff_1_SFF_5_U2 ( .A1(KeyArray_n19), .A2(
        KeyArray_S00reg_gff_1_SFF_5_n11), .ZN(KeyArray_S00reg_gff_1_SFF_5_n1)
         );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_5_U1 ( .A1(KeyArray_S00reg_gff_1_SFF_5_QD), .A2(KeyArray_n19), .ZN(KeyArray_S00reg_gff_1_SFF_5_n2) );
  XOR2_X1 KeyArray_S00reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A(
        KeyArray_inS00ser[5]), .B(KeyArray_outS10ser[5]), .Z(
        KeyArray_S00reg_gff_1_SFF_5_MUXInst_X) );
  AND2_X1 KeyArray_S00reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A1(KeyArray_n23), 
        .A2(KeyArray_S00reg_gff_1_SFF_5_MUXInst_X), .ZN(
        KeyArray_S00reg_gff_1_SFF_5_MUXInst_Y) );
  XOR2_X1 KeyArray_S00reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A(
        KeyArray_S00reg_gff_1_SFF_5_MUXInst_Y), .B(KeyArray_inS00ser[5]), .Z(
        KeyArray_S00reg_gff_1_SFF_5_QD) );
  INV_X1 KeyArray_S00reg_gff_1_SFF_5_Q_reg_U1 ( .A(keyStateIn[5]), .ZN(
        KeyArray_S00reg_gff_1_SFF_5_n11) );
  DFF_X1 KeyArray_S00reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        KeyArray_S00reg_gff_1_SFF_5_n6), .CK(clk), .Q(keyStateIn[5]), .QN() );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_6_U3 ( .A1(KeyArray_S00reg_gff_1_SFF_6_n2), .A2(KeyArray_S00reg_gff_1_SFF_6_n1), .ZN(KeyArray_S00reg_gff_1_SFF_6_n6) );
  OR2_X1 KeyArray_S00reg_gff_1_SFF_6_U2 ( .A1(KeyArray_n19), .A2(
        KeyArray_S00reg_gff_1_SFF_6_n11), .ZN(KeyArray_S00reg_gff_1_SFF_6_n1)
         );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_6_U1 ( .A1(KeyArray_S00reg_gff_1_SFF_6_QD), .A2(KeyArray_n19), .ZN(KeyArray_S00reg_gff_1_SFF_6_n2) );
  XOR2_X1 KeyArray_S00reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A(
        KeyArray_inS00ser[6]), .B(KeyArray_outS10ser[6]), .Z(
        KeyArray_S00reg_gff_1_SFF_6_MUXInst_X) );
  AND2_X1 KeyArray_S00reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A1(KeyArray_n23), 
        .A2(KeyArray_S00reg_gff_1_SFF_6_MUXInst_X), .ZN(
        KeyArray_S00reg_gff_1_SFF_6_MUXInst_Y) );
  XOR2_X1 KeyArray_S00reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A(
        KeyArray_S00reg_gff_1_SFF_6_MUXInst_Y), .B(KeyArray_inS00ser[6]), .Z(
        KeyArray_S00reg_gff_1_SFF_6_QD) );
  INV_X1 KeyArray_S00reg_gff_1_SFF_6_Q_reg_U1 ( .A(keyStateIn[6]), .ZN(
        KeyArray_S00reg_gff_1_SFF_6_n11) );
  DFF_X1 KeyArray_S00reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        KeyArray_S00reg_gff_1_SFF_6_n6), .CK(clk), .Q(keyStateIn[6]), .QN() );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_7_U3 ( .A1(KeyArray_S00reg_gff_1_SFF_7_n2), .A2(KeyArray_S00reg_gff_1_SFF_7_n1), .ZN(KeyArray_S00reg_gff_1_SFF_7_n6) );
  OR2_X1 KeyArray_S00reg_gff_1_SFF_7_U2 ( .A1(KeyArray_n19), .A2(
        KeyArray_S00reg_gff_1_SFF_7_n11), .ZN(KeyArray_S00reg_gff_1_SFF_7_n1)
         );
  NAND2_X1 KeyArray_S00reg_gff_1_SFF_7_U1 ( .A1(KeyArray_S00reg_gff_1_SFF_7_QD), .A2(KeyArray_n19), .ZN(KeyArray_S00reg_gff_1_SFF_7_n2) );
  XOR2_X1 KeyArray_S00reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A(
        KeyArray_inS00ser[7]), .B(KeyArray_outS10ser[7]), .Z(
        KeyArray_S00reg_gff_1_SFF_7_MUXInst_X) );
  AND2_X1 KeyArray_S00reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A1(KeyArray_n23), 
        .A2(KeyArray_S00reg_gff_1_SFF_7_MUXInst_X), .ZN(
        KeyArray_S00reg_gff_1_SFF_7_MUXInst_Y) );
  XOR2_X1 KeyArray_S00reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A(
        KeyArray_S00reg_gff_1_SFF_7_MUXInst_Y), .B(KeyArray_inS00ser[7]), .Z(
        KeyArray_S00reg_gff_1_SFF_7_QD) );
  INV_X1 KeyArray_S00reg_gff_1_SFF_7_Q_reg_U1 ( .A(keyStateIn[7]), .ZN(
        KeyArray_S00reg_gff_1_SFF_7_n11) );
  DFF_X1 KeyArray_S00reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        KeyArray_S00reg_gff_1_SFF_7_n6), .CK(clk), .Q(keyStateIn[7]), .QN() );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_0_U3 ( .A1(KeyArray_S01reg_gff_1_SFF_0_n2), .A2(KeyArray_S01reg_gff_1_SFF_0_n1), .ZN(KeyArray_S01reg_gff_1_SFF_0_n6) );
  OR2_X1 KeyArray_S01reg_gff_1_SFF_0_U2 ( .A1(KeyArray_n19), .A2(
        KeyArray_S01reg_gff_1_SFF_0_n11), .ZN(KeyArray_S01reg_gff_1_SFF_0_n1)
         );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_0_U1 ( .A1(KeyArray_S01reg_gff_1_SFF_0_QD), .A2(KeyArray_n19), .ZN(KeyArray_S01reg_gff_1_SFF_0_n2) );
  XOR2_X1 KeyArray_S01reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS02ser[0]), .B(KeyArray_outS11ser[0]), .Z(
        KeyArray_S01reg_gff_1_SFF_0_MUXInst_X) );
  AND2_X1 KeyArray_S01reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A1(KeyArray_n23), 
        .A2(KeyArray_S01reg_gff_1_SFF_0_MUXInst_X), .ZN(
        KeyArray_S01reg_gff_1_SFF_0_MUXInst_Y) );
  XOR2_X1 KeyArray_S01reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A(
        KeyArray_S01reg_gff_1_SFF_0_MUXInst_Y), .B(KeyArray_outS02ser[0]), .Z(
        KeyArray_S01reg_gff_1_SFF_0_QD) );
  INV_X1 KeyArray_S01reg_gff_1_SFF_0_Q_reg_U1 ( .A(KeyArray_outS01ser_0_), 
        .ZN(KeyArray_S01reg_gff_1_SFF_0_n11) );
  DFF_X1 KeyArray_S01reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        KeyArray_S01reg_gff_1_SFF_0_n6), .CK(clk), .Q(KeyArray_outS01ser_0_), 
        .QN() );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_1_U3 ( .A1(KeyArray_S01reg_gff_1_SFF_1_n2), .A2(KeyArray_S01reg_gff_1_SFF_1_n1), .ZN(KeyArray_S01reg_gff_1_SFF_1_n6) );
  OR2_X1 KeyArray_S01reg_gff_1_SFF_1_U2 ( .A1(KeyArray_n19), .A2(
        KeyArray_S01reg_gff_1_SFF_1_n11), .ZN(KeyArray_S01reg_gff_1_SFF_1_n1)
         );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_1_U1 ( .A1(KeyArray_S01reg_gff_1_SFF_1_QD), .A2(KeyArray_n19), .ZN(KeyArray_S01reg_gff_1_SFF_1_n2) );
  XOR2_X1 KeyArray_S01reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS02ser[1]), .B(KeyArray_outS11ser[1]), .Z(
        KeyArray_S01reg_gff_1_SFF_1_MUXInst_X) );
  AND2_X1 KeyArray_S01reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A1(KeyArray_n23), 
        .A2(KeyArray_S01reg_gff_1_SFF_1_MUXInst_X), .ZN(
        KeyArray_S01reg_gff_1_SFF_1_MUXInst_Y) );
  XOR2_X1 KeyArray_S01reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A(
        KeyArray_S01reg_gff_1_SFF_1_MUXInst_Y), .B(KeyArray_outS02ser[1]), .Z(
        KeyArray_S01reg_gff_1_SFF_1_QD) );
  INV_X1 KeyArray_S01reg_gff_1_SFF_1_Q_reg_U1 ( .A(KeyArray_outS01ser_1_), 
        .ZN(KeyArray_S01reg_gff_1_SFF_1_n11) );
  DFF_X1 KeyArray_S01reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        KeyArray_S01reg_gff_1_SFF_1_n6), .CK(clk), .Q(KeyArray_outS01ser_1_), 
        .QN() );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_2_U3 ( .A1(KeyArray_S01reg_gff_1_SFF_2_n2), .A2(KeyArray_S01reg_gff_1_SFF_2_n1), .ZN(KeyArray_S01reg_gff_1_SFF_2_n6) );
  OR2_X1 KeyArray_S01reg_gff_1_SFF_2_U2 ( .A1(KeyArray_n19), .A2(
        KeyArray_S01reg_gff_1_SFF_2_n11), .ZN(KeyArray_S01reg_gff_1_SFF_2_n1)
         );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_2_U1 ( .A1(KeyArray_S01reg_gff_1_SFF_2_QD), .A2(KeyArray_n19), .ZN(KeyArray_S01reg_gff_1_SFF_2_n2) );
  XOR2_X1 KeyArray_S01reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS02ser[2]), .B(KeyArray_outS11ser[2]), .Z(
        KeyArray_S01reg_gff_1_SFF_2_MUXInst_X) );
  AND2_X1 KeyArray_S01reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A1(KeyArray_n23), 
        .A2(KeyArray_S01reg_gff_1_SFF_2_MUXInst_X), .ZN(
        KeyArray_S01reg_gff_1_SFF_2_MUXInst_Y) );
  XOR2_X1 KeyArray_S01reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A(
        KeyArray_S01reg_gff_1_SFF_2_MUXInst_Y), .B(KeyArray_outS02ser[2]), .Z(
        KeyArray_S01reg_gff_1_SFF_2_QD) );
  INV_X1 KeyArray_S01reg_gff_1_SFF_2_Q_reg_U1 ( .A(KeyArray_outS01ser_2_), 
        .ZN(KeyArray_S01reg_gff_1_SFF_2_n11) );
  DFF_X1 KeyArray_S01reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        KeyArray_S01reg_gff_1_SFF_2_n6), .CK(clk), .Q(KeyArray_outS01ser_2_), 
        .QN() );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_3_U3 ( .A1(KeyArray_S01reg_gff_1_SFF_3_n2), .A2(KeyArray_S01reg_gff_1_SFF_3_n1), .ZN(KeyArray_S01reg_gff_1_SFF_3_n6) );
  OR2_X1 KeyArray_S01reg_gff_1_SFF_3_U2 ( .A1(KeyArray_n19), .A2(
        KeyArray_S01reg_gff_1_SFF_3_n11), .ZN(KeyArray_S01reg_gff_1_SFF_3_n1)
         );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_3_U1 ( .A1(KeyArray_S01reg_gff_1_SFF_3_QD), .A2(KeyArray_n19), .ZN(KeyArray_S01reg_gff_1_SFF_3_n2) );
  XOR2_X1 KeyArray_S01reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS02ser[3]), .B(KeyArray_outS11ser[3]), .Z(
        KeyArray_S01reg_gff_1_SFF_3_MUXInst_X) );
  AND2_X1 KeyArray_S01reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A1(KeyArray_n23), 
        .A2(KeyArray_S01reg_gff_1_SFF_3_MUXInst_X), .ZN(
        KeyArray_S01reg_gff_1_SFF_3_MUXInst_Y) );
  XOR2_X1 KeyArray_S01reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A(
        KeyArray_S01reg_gff_1_SFF_3_MUXInst_Y), .B(KeyArray_outS02ser[3]), .Z(
        KeyArray_S01reg_gff_1_SFF_3_QD) );
  INV_X1 KeyArray_S01reg_gff_1_SFF_3_Q_reg_U1 ( .A(KeyArray_outS01ser_3_), 
        .ZN(KeyArray_S01reg_gff_1_SFF_3_n11) );
  DFF_X1 KeyArray_S01reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        KeyArray_S01reg_gff_1_SFF_3_n6), .CK(clk), .Q(KeyArray_outS01ser_3_), 
        .QN() );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_4_U3 ( .A1(KeyArray_S01reg_gff_1_SFF_4_n2), .A2(KeyArray_S01reg_gff_1_SFF_4_n1), .ZN(KeyArray_S01reg_gff_1_SFF_4_n6) );
  OR2_X1 KeyArray_S01reg_gff_1_SFF_4_U2 ( .A1(KeyArray_n19), .A2(
        KeyArray_S01reg_gff_1_SFF_4_n11), .ZN(KeyArray_S01reg_gff_1_SFF_4_n1)
         );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_4_U1 ( .A1(KeyArray_S01reg_gff_1_SFF_4_QD), .A2(KeyArray_n19), .ZN(KeyArray_S01reg_gff_1_SFF_4_n2) );
  XOR2_X1 KeyArray_S01reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS02ser[4]), .B(KeyArray_outS11ser[4]), .Z(
        KeyArray_S01reg_gff_1_SFF_4_MUXInst_X) );
  AND2_X1 KeyArray_S01reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A1(KeyArray_n23), 
        .A2(KeyArray_S01reg_gff_1_SFF_4_MUXInst_X), .ZN(
        KeyArray_S01reg_gff_1_SFF_4_MUXInst_Y) );
  XOR2_X1 KeyArray_S01reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A(
        KeyArray_S01reg_gff_1_SFF_4_MUXInst_Y), .B(KeyArray_outS02ser[4]), .Z(
        KeyArray_S01reg_gff_1_SFF_4_QD) );
  INV_X1 KeyArray_S01reg_gff_1_SFF_4_Q_reg_U1 ( .A(KeyArray_outS01ser_4_), 
        .ZN(KeyArray_S01reg_gff_1_SFF_4_n11) );
  DFF_X1 KeyArray_S01reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        KeyArray_S01reg_gff_1_SFF_4_n6), .CK(clk), .Q(KeyArray_outS01ser_4_), 
        .QN() );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_5_U3 ( .A1(KeyArray_S01reg_gff_1_SFF_5_n2), .A2(KeyArray_S01reg_gff_1_SFF_5_n1), .ZN(KeyArray_S01reg_gff_1_SFF_5_n6) );
  OR2_X1 KeyArray_S01reg_gff_1_SFF_5_U2 ( .A1(KeyArray_n19), .A2(
        KeyArray_S01reg_gff_1_SFF_5_n11), .ZN(KeyArray_S01reg_gff_1_SFF_5_n1)
         );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_5_U1 ( .A1(KeyArray_S01reg_gff_1_SFF_5_QD), .A2(KeyArray_n19), .ZN(KeyArray_S01reg_gff_1_SFF_5_n2) );
  XOR2_X1 KeyArray_S01reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS02ser[5]), .B(KeyArray_outS11ser[5]), .Z(
        KeyArray_S01reg_gff_1_SFF_5_MUXInst_X) );
  AND2_X1 KeyArray_S01reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A1(KeyArray_n23), 
        .A2(KeyArray_S01reg_gff_1_SFF_5_MUXInst_X), .ZN(
        KeyArray_S01reg_gff_1_SFF_5_MUXInst_Y) );
  XOR2_X1 KeyArray_S01reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A(
        KeyArray_S01reg_gff_1_SFF_5_MUXInst_Y), .B(KeyArray_outS02ser[5]), .Z(
        KeyArray_S01reg_gff_1_SFF_5_QD) );
  INV_X1 KeyArray_S01reg_gff_1_SFF_5_Q_reg_U1 ( .A(KeyArray_outS01ser_5_), 
        .ZN(KeyArray_S01reg_gff_1_SFF_5_n11) );
  DFF_X1 KeyArray_S01reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        KeyArray_S01reg_gff_1_SFF_5_n6), .CK(clk), .Q(KeyArray_outS01ser_5_), 
        .QN() );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_6_U3 ( .A1(KeyArray_S01reg_gff_1_SFF_6_n2), .A2(KeyArray_S01reg_gff_1_SFF_6_n1), .ZN(KeyArray_S01reg_gff_1_SFF_6_n6) );
  OR2_X1 KeyArray_S01reg_gff_1_SFF_6_U2 ( .A1(KeyArray_n19), .A2(
        KeyArray_S01reg_gff_1_SFF_6_n11), .ZN(KeyArray_S01reg_gff_1_SFF_6_n1)
         );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_6_U1 ( .A1(KeyArray_S01reg_gff_1_SFF_6_QD), .A2(KeyArray_n19), .ZN(KeyArray_S01reg_gff_1_SFF_6_n2) );
  XOR2_X1 KeyArray_S01reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS02ser[6]), .B(KeyArray_outS11ser[6]), .Z(
        KeyArray_S01reg_gff_1_SFF_6_MUXInst_X) );
  AND2_X1 KeyArray_S01reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A1(KeyArray_n23), 
        .A2(KeyArray_S01reg_gff_1_SFF_6_MUXInst_X), .ZN(
        KeyArray_S01reg_gff_1_SFF_6_MUXInst_Y) );
  XOR2_X1 KeyArray_S01reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A(
        KeyArray_S01reg_gff_1_SFF_6_MUXInst_Y), .B(KeyArray_outS02ser[6]), .Z(
        KeyArray_S01reg_gff_1_SFF_6_QD) );
  INV_X1 KeyArray_S01reg_gff_1_SFF_6_Q_reg_U1 ( .A(KeyArray_outS01ser_6_), 
        .ZN(KeyArray_S01reg_gff_1_SFF_6_n11) );
  DFF_X1 KeyArray_S01reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        KeyArray_S01reg_gff_1_SFF_6_n6), .CK(clk), .Q(KeyArray_outS01ser_6_), 
        .QN() );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_7_U3 ( .A1(KeyArray_S01reg_gff_1_SFF_7_n2), .A2(KeyArray_S01reg_gff_1_SFF_7_n1), .ZN(KeyArray_S01reg_gff_1_SFF_7_n6) );
  OR2_X1 KeyArray_S01reg_gff_1_SFF_7_U2 ( .A1(KeyArray_n19), .A2(
        KeyArray_S01reg_gff_1_SFF_7_n11), .ZN(KeyArray_S01reg_gff_1_SFF_7_n1)
         );
  NAND2_X1 KeyArray_S01reg_gff_1_SFF_7_U1 ( .A1(KeyArray_S01reg_gff_1_SFF_7_QD), .A2(KeyArray_n19), .ZN(KeyArray_S01reg_gff_1_SFF_7_n2) );
  XOR2_X1 KeyArray_S01reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS02ser[7]), .B(KeyArray_outS11ser[7]), .Z(
        KeyArray_S01reg_gff_1_SFF_7_MUXInst_X) );
  AND2_X1 KeyArray_S01reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A1(KeyArray_n23), 
        .A2(KeyArray_S01reg_gff_1_SFF_7_MUXInst_X), .ZN(
        KeyArray_S01reg_gff_1_SFF_7_MUXInst_Y) );
  XOR2_X1 KeyArray_S01reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A(
        KeyArray_S01reg_gff_1_SFF_7_MUXInst_Y), .B(KeyArray_outS02ser[7]), .Z(
        KeyArray_S01reg_gff_1_SFF_7_QD) );
  INV_X1 KeyArray_S01reg_gff_1_SFF_7_Q_reg_U1 ( .A(KeyArray_outS01ser_7_), 
        .ZN(KeyArray_S01reg_gff_1_SFF_7_n11) );
  DFF_X1 KeyArray_S01reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        KeyArray_S01reg_gff_1_SFF_7_n6), .CK(clk), .Q(KeyArray_outS01ser_7_), 
        .QN() );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_0_U3 ( .A1(KeyArray_S02reg_gff_1_SFF_0_n2), .A2(KeyArray_S02reg_gff_1_SFF_0_n1), .ZN(KeyArray_S02reg_gff_1_SFF_0_n6) );
  OR2_X1 KeyArray_S02reg_gff_1_SFF_0_U2 ( .A1(KeyArray_n19), .A2(
        KeyArray_S02reg_gff_1_SFF_0_n11), .ZN(KeyArray_S02reg_gff_1_SFF_0_n1)
         );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_0_U1 ( .A1(KeyArray_S02reg_gff_1_SFF_0_QD), .A2(KeyArray_n19), .ZN(KeyArray_S02reg_gff_1_SFF_0_n2) );
  XOR2_X1 KeyArray_S02reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS03ser[0]), .B(KeyArray_outS12ser[0]), .Z(
        KeyArray_S02reg_gff_1_SFF_0_MUXInst_X) );
  AND2_X1 KeyArray_S02reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A1(KeyArray_n23), 
        .A2(KeyArray_S02reg_gff_1_SFF_0_MUXInst_X), .ZN(
        KeyArray_S02reg_gff_1_SFF_0_MUXInst_Y) );
  XOR2_X1 KeyArray_S02reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A(
        KeyArray_S02reg_gff_1_SFF_0_MUXInst_Y), .B(KeyArray_outS03ser[0]), .Z(
        KeyArray_S02reg_gff_1_SFF_0_QD) );
  INV_X1 KeyArray_S02reg_gff_1_SFF_0_Q_reg_U1 ( .A(KeyArray_outS02ser[0]), 
        .ZN(KeyArray_S02reg_gff_1_SFF_0_n11) );
  DFF_X1 KeyArray_S02reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        KeyArray_S02reg_gff_1_SFF_0_n6), .CK(clk), .Q(KeyArray_outS02ser[0]), 
        .QN() );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_1_U3 ( .A1(KeyArray_S02reg_gff_1_SFF_1_n2), .A2(KeyArray_S02reg_gff_1_SFF_1_n1), .ZN(KeyArray_S02reg_gff_1_SFF_1_n6) );
  OR2_X1 KeyArray_S02reg_gff_1_SFF_1_U2 ( .A1(KeyArray_n19), .A2(
        KeyArray_S02reg_gff_1_SFF_1_n11), .ZN(KeyArray_S02reg_gff_1_SFF_1_n1)
         );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_1_U1 ( .A1(KeyArray_S02reg_gff_1_SFF_1_QD), .A2(KeyArray_n19), .ZN(KeyArray_S02reg_gff_1_SFF_1_n2) );
  XOR2_X1 KeyArray_S02reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS03ser[1]), .B(KeyArray_outS12ser[1]), .Z(
        KeyArray_S02reg_gff_1_SFF_1_MUXInst_X) );
  AND2_X1 KeyArray_S02reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A1(KeyArray_n23), 
        .A2(KeyArray_S02reg_gff_1_SFF_1_MUXInst_X), .ZN(
        KeyArray_S02reg_gff_1_SFF_1_MUXInst_Y) );
  XOR2_X1 KeyArray_S02reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A(
        KeyArray_S02reg_gff_1_SFF_1_MUXInst_Y), .B(KeyArray_outS03ser[1]), .Z(
        KeyArray_S02reg_gff_1_SFF_1_QD) );
  INV_X1 KeyArray_S02reg_gff_1_SFF_1_Q_reg_U1 ( .A(KeyArray_outS02ser[1]), 
        .ZN(KeyArray_S02reg_gff_1_SFF_1_n11) );
  DFF_X1 KeyArray_S02reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        KeyArray_S02reg_gff_1_SFF_1_n6), .CK(clk), .Q(KeyArray_outS02ser[1]), 
        .QN() );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_2_U3 ( .A1(KeyArray_S02reg_gff_1_SFF_2_n2), .A2(KeyArray_S02reg_gff_1_SFF_2_n1), .ZN(KeyArray_S02reg_gff_1_SFF_2_n6) );
  OR2_X1 KeyArray_S02reg_gff_1_SFF_2_U2 ( .A1(KeyArray_n19), .A2(
        KeyArray_S02reg_gff_1_SFF_2_n11), .ZN(KeyArray_S02reg_gff_1_SFF_2_n1)
         );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_2_U1 ( .A1(KeyArray_S02reg_gff_1_SFF_2_QD), .A2(KeyArray_n19), .ZN(KeyArray_S02reg_gff_1_SFF_2_n2) );
  XOR2_X1 KeyArray_S02reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS03ser[2]), .B(KeyArray_outS12ser[2]), .Z(
        KeyArray_S02reg_gff_1_SFF_2_MUXInst_X) );
  AND2_X1 KeyArray_S02reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A1(KeyArray_n23), 
        .A2(KeyArray_S02reg_gff_1_SFF_2_MUXInst_X), .ZN(
        KeyArray_S02reg_gff_1_SFF_2_MUXInst_Y) );
  XOR2_X1 KeyArray_S02reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A(
        KeyArray_S02reg_gff_1_SFF_2_MUXInst_Y), .B(KeyArray_outS03ser[2]), .Z(
        KeyArray_S02reg_gff_1_SFF_2_QD) );
  INV_X1 KeyArray_S02reg_gff_1_SFF_2_Q_reg_U1 ( .A(KeyArray_outS02ser[2]), 
        .ZN(KeyArray_S02reg_gff_1_SFF_2_n11) );
  DFF_X1 KeyArray_S02reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        KeyArray_S02reg_gff_1_SFF_2_n6), .CK(clk), .Q(KeyArray_outS02ser[2]), 
        .QN() );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_3_U3 ( .A1(KeyArray_S02reg_gff_1_SFF_3_n2), .A2(KeyArray_S02reg_gff_1_SFF_3_n1), .ZN(KeyArray_S02reg_gff_1_SFF_3_n6) );
  OR2_X1 KeyArray_S02reg_gff_1_SFF_3_U2 ( .A1(KeyArray_n19), .A2(
        KeyArray_S02reg_gff_1_SFF_3_n11), .ZN(KeyArray_S02reg_gff_1_SFF_3_n1)
         );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_3_U1 ( .A1(KeyArray_S02reg_gff_1_SFF_3_QD), .A2(KeyArray_n19), .ZN(KeyArray_S02reg_gff_1_SFF_3_n2) );
  XOR2_X1 KeyArray_S02reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS03ser[3]), .B(KeyArray_outS12ser[3]), .Z(
        KeyArray_S02reg_gff_1_SFF_3_MUXInst_X) );
  AND2_X1 KeyArray_S02reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A1(KeyArray_n23), 
        .A2(KeyArray_S02reg_gff_1_SFF_3_MUXInst_X), .ZN(
        KeyArray_S02reg_gff_1_SFF_3_MUXInst_Y) );
  XOR2_X1 KeyArray_S02reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A(
        KeyArray_S02reg_gff_1_SFF_3_MUXInst_Y), .B(KeyArray_outS03ser[3]), .Z(
        KeyArray_S02reg_gff_1_SFF_3_QD) );
  INV_X1 KeyArray_S02reg_gff_1_SFF_3_Q_reg_U1 ( .A(KeyArray_outS02ser[3]), 
        .ZN(KeyArray_S02reg_gff_1_SFF_3_n11) );
  DFF_X1 KeyArray_S02reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        KeyArray_S02reg_gff_1_SFF_3_n6), .CK(clk), .Q(KeyArray_outS02ser[3]), 
        .QN() );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_4_U3 ( .A1(KeyArray_S02reg_gff_1_SFF_4_n2), .A2(KeyArray_S02reg_gff_1_SFF_4_n1), .ZN(KeyArray_S02reg_gff_1_SFF_4_n6) );
  OR2_X1 KeyArray_S02reg_gff_1_SFF_4_U2 ( .A1(KeyArray_n19), .A2(
        KeyArray_S02reg_gff_1_SFF_4_n11), .ZN(KeyArray_S02reg_gff_1_SFF_4_n1)
         );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_4_U1 ( .A1(KeyArray_S02reg_gff_1_SFF_4_QD), .A2(KeyArray_n19), .ZN(KeyArray_S02reg_gff_1_SFF_4_n2) );
  XOR2_X1 KeyArray_S02reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS03ser[4]), .B(KeyArray_outS12ser[4]), .Z(
        KeyArray_S02reg_gff_1_SFF_4_MUXInst_X) );
  AND2_X1 KeyArray_S02reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A1(KeyArray_n23), 
        .A2(KeyArray_S02reg_gff_1_SFF_4_MUXInst_X), .ZN(
        KeyArray_S02reg_gff_1_SFF_4_MUXInst_Y) );
  XOR2_X1 KeyArray_S02reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A(
        KeyArray_S02reg_gff_1_SFF_4_MUXInst_Y), .B(KeyArray_outS03ser[4]), .Z(
        KeyArray_S02reg_gff_1_SFF_4_QD) );
  INV_X1 KeyArray_S02reg_gff_1_SFF_4_Q_reg_U1 ( .A(KeyArray_outS02ser[4]), 
        .ZN(KeyArray_S02reg_gff_1_SFF_4_n11) );
  DFF_X1 KeyArray_S02reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        KeyArray_S02reg_gff_1_SFF_4_n6), .CK(clk), .Q(KeyArray_outS02ser[4]), 
        .QN() );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_5_U3 ( .A1(KeyArray_S02reg_gff_1_SFF_5_n2), .A2(KeyArray_S02reg_gff_1_SFF_5_n1), .ZN(KeyArray_S02reg_gff_1_SFF_5_n6) );
  OR2_X1 KeyArray_S02reg_gff_1_SFF_5_U2 ( .A1(KeyArray_n19), .A2(
        KeyArray_S02reg_gff_1_SFF_5_n11), .ZN(KeyArray_S02reg_gff_1_SFF_5_n1)
         );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_5_U1 ( .A1(KeyArray_S02reg_gff_1_SFF_5_QD), .A2(KeyArray_n19), .ZN(KeyArray_S02reg_gff_1_SFF_5_n2) );
  XOR2_X1 KeyArray_S02reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS03ser[5]), .B(KeyArray_outS12ser[5]), .Z(
        KeyArray_S02reg_gff_1_SFF_5_MUXInst_X) );
  AND2_X1 KeyArray_S02reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A1(KeyArray_n23), 
        .A2(KeyArray_S02reg_gff_1_SFF_5_MUXInst_X), .ZN(
        KeyArray_S02reg_gff_1_SFF_5_MUXInst_Y) );
  XOR2_X1 KeyArray_S02reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A(
        KeyArray_S02reg_gff_1_SFF_5_MUXInst_Y), .B(KeyArray_outS03ser[5]), .Z(
        KeyArray_S02reg_gff_1_SFF_5_QD) );
  INV_X1 KeyArray_S02reg_gff_1_SFF_5_Q_reg_U1 ( .A(KeyArray_outS02ser[5]), 
        .ZN(KeyArray_S02reg_gff_1_SFF_5_n11) );
  DFF_X1 KeyArray_S02reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        KeyArray_S02reg_gff_1_SFF_5_n6), .CK(clk), .Q(KeyArray_outS02ser[5]), 
        .QN() );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_6_U3 ( .A1(KeyArray_S02reg_gff_1_SFF_6_n2), .A2(KeyArray_S02reg_gff_1_SFF_6_n1), .ZN(KeyArray_S02reg_gff_1_SFF_6_n6) );
  OR2_X1 KeyArray_S02reg_gff_1_SFF_6_U2 ( .A1(KeyArray_n19), .A2(
        KeyArray_S02reg_gff_1_SFF_6_n11), .ZN(KeyArray_S02reg_gff_1_SFF_6_n1)
         );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_6_U1 ( .A1(KeyArray_S02reg_gff_1_SFF_6_QD), .A2(KeyArray_n19), .ZN(KeyArray_S02reg_gff_1_SFF_6_n2) );
  XOR2_X1 KeyArray_S02reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS03ser[6]), .B(KeyArray_outS12ser[6]), .Z(
        KeyArray_S02reg_gff_1_SFF_6_MUXInst_X) );
  AND2_X1 KeyArray_S02reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A1(KeyArray_n23), 
        .A2(KeyArray_S02reg_gff_1_SFF_6_MUXInst_X), .ZN(
        KeyArray_S02reg_gff_1_SFF_6_MUXInst_Y) );
  XOR2_X1 KeyArray_S02reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A(
        KeyArray_S02reg_gff_1_SFF_6_MUXInst_Y), .B(KeyArray_outS03ser[6]), .Z(
        KeyArray_S02reg_gff_1_SFF_6_QD) );
  INV_X1 KeyArray_S02reg_gff_1_SFF_6_Q_reg_U1 ( .A(KeyArray_outS02ser[6]), 
        .ZN(KeyArray_S02reg_gff_1_SFF_6_n11) );
  DFF_X1 KeyArray_S02reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        KeyArray_S02reg_gff_1_SFF_6_n6), .CK(clk), .Q(KeyArray_outS02ser[6]), 
        .QN() );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_7_U3 ( .A1(KeyArray_S02reg_gff_1_SFF_7_n2), .A2(KeyArray_S02reg_gff_1_SFF_7_n1), .ZN(KeyArray_S02reg_gff_1_SFF_7_n6) );
  OR2_X1 KeyArray_S02reg_gff_1_SFF_7_U2 ( .A1(KeyArray_n19), .A2(
        KeyArray_S02reg_gff_1_SFF_7_n11), .ZN(KeyArray_S02reg_gff_1_SFF_7_n1)
         );
  NAND2_X1 KeyArray_S02reg_gff_1_SFF_7_U1 ( .A1(KeyArray_S02reg_gff_1_SFF_7_QD), .A2(KeyArray_n19), .ZN(KeyArray_S02reg_gff_1_SFF_7_n2) );
  XOR2_X1 KeyArray_S02reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS03ser[7]), .B(KeyArray_outS12ser[7]), .Z(
        KeyArray_S02reg_gff_1_SFF_7_MUXInst_X) );
  AND2_X1 KeyArray_S02reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A1(KeyArray_n23), 
        .A2(KeyArray_S02reg_gff_1_SFF_7_MUXInst_X), .ZN(
        KeyArray_S02reg_gff_1_SFF_7_MUXInst_Y) );
  XOR2_X1 KeyArray_S02reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A(
        KeyArray_S02reg_gff_1_SFF_7_MUXInst_Y), .B(KeyArray_outS03ser[7]), .Z(
        KeyArray_S02reg_gff_1_SFF_7_QD) );
  INV_X1 KeyArray_S02reg_gff_1_SFF_7_Q_reg_U1 ( .A(KeyArray_outS02ser[7]), 
        .ZN(KeyArray_S02reg_gff_1_SFF_7_n11) );
  DFF_X1 KeyArray_S02reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        KeyArray_S02reg_gff_1_SFF_7_n6), .CK(clk), .Q(KeyArray_outS02ser[7]), 
        .QN() );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_0_U3 ( .A1(KeyArray_S03reg_gff_1_SFF_0_n2), .A2(KeyArray_S03reg_gff_1_SFF_0_n1), .ZN(KeyArray_S03reg_gff_1_SFF_0_n6) );
  OR2_X1 KeyArray_S03reg_gff_1_SFF_0_U2 ( .A1(KeyArray_n19), .A2(
        KeyArray_S03reg_gff_1_SFF_0_n11), .ZN(KeyArray_S03reg_gff_1_SFF_0_n1)
         );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_0_U1 ( .A1(KeyArray_S03reg_gff_1_SFF_0_QD), .A2(KeyArray_n19), .ZN(KeyArray_S03reg_gff_1_SFF_0_n2) );
  XOR2_X1 KeyArray_S03reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS10ser[0]), .B(keySBIn[0]), .Z(
        KeyArray_S03reg_gff_1_SFF_0_MUXInst_X) );
  AND2_X1 KeyArray_S03reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A1(KeyArray_n23), 
        .A2(KeyArray_S03reg_gff_1_SFF_0_MUXInst_X), .ZN(
        KeyArray_S03reg_gff_1_SFF_0_MUXInst_Y) );
  XOR2_X1 KeyArray_S03reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A(
        KeyArray_S03reg_gff_1_SFF_0_MUXInst_Y), .B(KeyArray_outS10ser[0]), .Z(
        KeyArray_S03reg_gff_1_SFF_0_QD) );
  INV_X1 KeyArray_S03reg_gff_1_SFF_0_Q_reg_U1 ( .A(KeyArray_outS03ser[0]), 
        .ZN(KeyArray_S03reg_gff_1_SFF_0_n11) );
  DFF_X1 KeyArray_S03reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        KeyArray_S03reg_gff_1_SFF_0_n6), .CK(clk), .Q(KeyArray_outS03ser[0]), 
        .QN() );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_1_U3 ( .A1(KeyArray_S03reg_gff_1_SFF_1_n2), .A2(KeyArray_S03reg_gff_1_SFF_1_n1), .ZN(KeyArray_S03reg_gff_1_SFF_1_n6) );
  OR2_X1 KeyArray_S03reg_gff_1_SFF_1_U2 ( .A1(KeyArray_n19), .A2(
        KeyArray_S03reg_gff_1_SFF_1_n11), .ZN(KeyArray_S03reg_gff_1_SFF_1_n1)
         );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_1_U1 ( .A1(KeyArray_S03reg_gff_1_SFF_1_QD), .A2(KeyArray_n19), .ZN(KeyArray_S03reg_gff_1_SFF_1_n2) );
  XOR2_X1 KeyArray_S03reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS10ser[1]), .B(keySBIn[1]), .Z(
        KeyArray_S03reg_gff_1_SFF_1_MUXInst_X) );
  AND2_X1 KeyArray_S03reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A1(KeyArray_n23), 
        .A2(KeyArray_S03reg_gff_1_SFF_1_MUXInst_X), .ZN(
        KeyArray_S03reg_gff_1_SFF_1_MUXInst_Y) );
  XOR2_X1 KeyArray_S03reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A(
        KeyArray_S03reg_gff_1_SFF_1_MUXInst_Y), .B(KeyArray_outS10ser[1]), .Z(
        KeyArray_S03reg_gff_1_SFF_1_QD) );
  INV_X1 KeyArray_S03reg_gff_1_SFF_1_Q_reg_U1 ( .A(KeyArray_outS03ser[1]), 
        .ZN(KeyArray_S03reg_gff_1_SFF_1_n11) );
  DFF_X1 KeyArray_S03reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        KeyArray_S03reg_gff_1_SFF_1_n6), .CK(clk), .Q(KeyArray_outS03ser[1]), 
        .QN() );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_2_U3 ( .A1(KeyArray_S03reg_gff_1_SFF_2_n2), .A2(KeyArray_S03reg_gff_1_SFF_2_n1), .ZN(KeyArray_S03reg_gff_1_SFF_2_n6) );
  OR2_X1 KeyArray_S03reg_gff_1_SFF_2_U2 ( .A1(KeyArray_n19), .A2(
        KeyArray_S03reg_gff_1_SFF_2_n11), .ZN(KeyArray_S03reg_gff_1_SFF_2_n1)
         );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_2_U1 ( .A1(KeyArray_S03reg_gff_1_SFF_2_QD), .A2(KeyArray_n19), .ZN(KeyArray_S03reg_gff_1_SFF_2_n2) );
  XOR2_X1 KeyArray_S03reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS10ser[2]), .B(keySBIn[2]), .Z(
        KeyArray_S03reg_gff_1_SFF_2_MUXInst_X) );
  AND2_X1 KeyArray_S03reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A1(KeyArray_n23), 
        .A2(KeyArray_S03reg_gff_1_SFF_2_MUXInst_X), .ZN(
        KeyArray_S03reg_gff_1_SFF_2_MUXInst_Y) );
  XOR2_X1 KeyArray_S03reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A(
        KeyArray_S03reg_gff_1_SFF_2_MUXInst_Y), .B(KeyArray_outS10ser[2]), .Z(
        KeyArray_S03reg_gff_1_SFF_2_QD) );
  INV_X1 KeyArray_S03reg_gff_1_SFF_2_Q_reg_U1 ( .A(KeyArray_outS03ser[2]), 
        .ZN(KeyArray_S03reg_gff_1_SFF_2_n11) );
  DFF_X1 KeyArray_S03reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        KeyArray_S03reg_gff_1_SFF_2_n6), .CK(clk), .Q(KeyArray_outS03ser[2]), 
        .QN() );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_3_U3 ( .A1(KeyArray_S03reg_gff_1_SFF_3_n2), .A2(KeyArray_S03reg_gff_1_SFF_3_n1), .ZN(KeyArray_S03reg_gff_1_SFF_3_n6) );
  OR2_X1 KeyArray_S03reg_gff_1_SFF_3_U2 ( .A1(KeyArray_n19), .A2(
        KeyArray_S03reg_gff_1_SFF_3_n11), .ZN(KeyArray_S03reg_gff_1_SFF_3_n1)
         );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_3_U1 ( .A1(KeyArray_S03reg_gff_1_SFF_3_QD), .A2(KeyArray_n19), .ZN(KeyArray_S03reg_gff_1_SFF_3_n2) );
  XOR2_X1 KeyArray_S03reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS10ser[3]), .B(keySBIn[3]), .Z(
        KeyArray_S03reg_gff_1_SFF_3_MUXInst_X) );
  AND2_X1 KeyArray_S03reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A1(KeyArray_n23), 
        .A2(KeyArray_S03reg_gff_1_SFF_3_MUXInst_X), .ZN(
        KeyArray_S03reg_gff_1_SFF_3_MUXInst_Y) );
  XOR2_X1 KeyArray_S03reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A(
        KeyArray_S03reg_gff_1_SFF_3_MUXInst_Y), .B(KeyArray_outS10ser[3]), .Z(
        KeyArray_S03reg_gff_1_SFF_3_QD) );
  INV_X1 KeyArray_S03reg_gff_1_SFF_3_Q_reg_U1 ( .A(KeyArray_outS03ser[3]), 
        .ZN(KeyArray_S03reg_gff_1_SFF_3_n11) );
  DFF_X1 KeyArray_S03reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        KeyArray_S03reg_gff_1_SFF_3_n6), .CK(clk), .Q(KeyArray_outS03ser[3]), 
        .QN() );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_4_U3 ( .A1(KeyArray_S03reg_gff_1_SFF_4_n2), .A2(KeyArray_S03reg_gff_1_SFF_4_n1), .ZN(KeyArray_S03reg_gff_1_SFF_4_n6) );
  OR2_X1 KeyArray_S03reg_gff_1_SFF_4_U2 ( .A1(KeyArray_n19), .A2(
        KeyArray_S03reg_gff_1_SFF_4_n11), .ZN(KeyArray_S03reg_gff_1_SFF_4_n1)
         );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_4_U1 ( .A1(KeyArray_S03reg_gff_1_SFF_4_QD), .A2(KeyArray_n19), .ZN(KeyArray_S03reg_gff_1_SFF_4_n2) );
  XOR2_X1 KeyArray_S03reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS10ser[4]), .B(keySBIn[4]), .Z(
        KeyArray_S03reg_gff_1_SFF_4_MUXInst_X) );
  AND2_X1 KeyArray_S03reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A1(KeyArray_n23), 
        .A2(KeyArray_S03reg_gff_1_SFF_4_MUXInst_X), .ZN(
        KeyArray_S03reg_gff_1_SFF_4_MUXInst_Y) );
  XOR2_X1 KeyArray_S03reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A(
        KeyArray_S03reg_gff_1_SFF_4_MUXInst_Y), .B(KeyArray_outS10ser[4]), .Z(
        KeyArray_S03reg_gff_1_SFF_4_QD) );
  INV_X1 KeyArray_S03reg_gff_1_SFF_4_Q_reg_U1 ( .A(KeyArray_outS03ser[4]), 
        .ZN(KeyArray_S03reg_gff_1_SFF_4_n11) );
  DFF_X1 KeyArray_S03reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        KeyArray_S03reg_gff_1_SFF_4_n6), .CK(clk), .Q(KeyArray_outS03ser[4]), 
        .QN() );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_5_U3 ( .A1(KeyArray_S03reg_gff_1_SFF_5_n2), .A2(KeyArray_S03reg_gff_1_SFF_5_n1), .ZN(KeyArray_S03reg_gff_1_SFF_5_n5) );
  OR2_X1 KeyArray_S03reg_gff_1_SFF_5_U2 ( .A1(KeyArray_n19), .A2(
        KeyArray_S03reg_gff_1_SFF_5_n3), .ZN(KeyArray_S03reg_gff_1_SFF_5_n1)
         );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_5_U1 ( .A1(KeyArray_S03reg_gff_1_SFF_5_QD), .A2(KeyArray_n19), .ZN(KeyArray_S03reg_gff_1_SFF_5_n2) );
  XOR2_X1 KeyArray_S03reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS10ser[5]), .B(keySBIn[5]), .Z(
        KeyArray_S03reg_gff_1_SFF_5_MUXInst_X) );
  AND2_X1 KeyArray_S03reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A1(KeyArray_n23), 
        .A2(KeyArray_S03reg_gff_1_SFF_5_MUXInst_X), .ZN(
        KeyArray_S03reg_gff_1_SFF_5_MUXInst_Y) );
  XOR2_X1 KeyArray_S03reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A(
        KeyArray_S03reg_gff_1_SFF_5_MUXInst_Y), .B(KeyArray_outS10ser[5]), .Z(
        KeyArray_S03reg_gff_1_SFF_5_QD) );
  INV_X1 KeyArray_S03reg_gff_1_SFF_5_Q_reg_U1 ( .A(KeyArray_outS03ser[5]), 
        .ZN(KeyArray_S03reg_gff_1_SFF_5_n3) );
  DFF_X1 KeyArray_S03reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        KeyArray_S03reg_gff_1_SFF_5_n5), .CK(clk), .Q(KeyArray_outS03ser[5]), 
        .QN() );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_6_U3 ( .A1(KeyArray_S03reg_gff_1_SFF_6_n2), .A2(KeyArray_S03reg_gff_1_SFF_6_n1), .ZN(KeyArray_S03reg_gff_1_SFF_6_n5) );
  OR2_X1 KeyArray_S03reg_gff_1_SFF_6_U2 ( .A1(KeyArray_n19), .A2(
        KeyArray_S03reg_gff_1_SFF_6_n10), .ZN(KeyArray_S03reg_gff_1_SFF_6_n1)
         );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_6_U1 ( .A1(KeyArray_S03reg_gff_1_SFF_6_QD), .A2(KeyArray_n19), .ZN(KeyArray_S03reg_gff_1_SFF_6_n2) );
  XOR2_X1 KeyArray_S03reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS10ser[6]), .B(keySBIn[6]), .Z(
        KeyArray_S03reg_gff_1_SFF_6_MUXInst_X) );
  AND2_X1 KeyArray_S03reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A1(KeyArray_n23), 
        .A2(KeyArray_S03reg_gff_1_SFF_6_MUXInst_X), .ZN(
        KeyArray_S03reg_gff_1_SFF_6_MUXInst_Y) );
  XOR2_X1 KeyArray_S03reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A(
        KeyArray_S03reg_gff_1_SFF_6_MUXInst_Y), .B(KeyArray_outS10ser[6]), .Z(
        KeyArray_S03reg_gff_1_SFF_6_QD) );
  INV_X1 KeyArray_S03reg_gff_1_SFF_6_Q_reg_U1 ( .A(KeyArray_outS03ser[6]), 
        .ZN(KeyArray_S03reg_gff_1_SFF_6_n10) );
  DFF_X1 KeyArray_S03reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        KeyArray_S03reg_gff_1_SFF_6_n5), .CK(clk), .Q(KeyArray_outS03ser[6]), 
        .QN() );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_7_U3 ( .A1(KeyArray_S03reg_gff_1_SFF_7_n2), .A2(KeyArray_S03reg_gff_1_SFF_7_n1), .ZN(KeyArray_S03reg_gff_1_SFF_7_n5) );
  OR2_X1 KeyArray_S03reg_gff_1_SFF_7_U2 ( .A1(KeyArray_n19), .A2(
        KeyArray_S03reg_gff_1_SFF_7_n10), .ZN(KeyArray_S03reg_gff_1_SFF_7_n1)
         );
  NAND2_X1 KeyArray_S03reg_gff_1_SFF_7_U1 ( .A1(KeyArray_S03reg_gff_1_SFF_7_QD), .A2(KeyArray_n19), .ZN(KeyArray_S03reg_gff_1_SFF_7_n2) );
  XOR2_X1 KeyArray_S03reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS10ser[7]), .B(keySBIn[7]), .Z(
        KeyArray_S03reg_gff_1_SFF_7_MUXInst_X) );
  AND2_X1 KeyArray_S03reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A1(KeyArray_n23), 
        .A2(KeyArray_S03reg_gff_1_SFF_7_MUXInst_X), .ZN(
        KeyArray_S03reg_gff_1_SFF_7_MUXInst_Y) );
  XOR2_X1 KeyArray_S03reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A(
        KeyArray_S03reg_gff_1_SFF_7_MUXInst_Y), .B(KeyArray_outS10ser[7]), .Z(
        KeyArray_S03reg_gff_1_SFF_7_QD) );
  INV_X1 KeyArray_S03reg_gff_1_SFF_7_Q_reg_U1 ( .A(KeyArray_outS03ser[7]), 
        .ZN(KeyArray_S03reg_gff_1_SFF_7_n10) );
  DFF_X1 KeyArray_S03reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        KeyArray_S03reg_gff_1_SFF_7_n5), .CK(clk), .Q(KeyArray_outS03ser[7]), 
        .QN() );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_0_U3 ( .A1(KeyArray_S10reg_gff_1_SFF_0_n2), .A2(KeyArray_S10reg_gff_1_SFF_0_n1), .ZN(KeyArray_S10reg_gff_1_SFF_0_n5) );
  OR2_X1 KeyArray_S10reg_gff_1_SFF_0_U2 ( .A1(KeyArray_n19), .A2(
        KeyArray_S10reg_gff_1_SFF_0_n10), .ZN(KeyArray_S10reg_gff_1_SFF_0_n1)
         );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_0_U1 ( .A1(KeyArray_S10reg_gff_1_SFF_0_QD), .A2(KeyArray_n19), .ZN(KeyArray_S10reg_gff_1_SFF_0_n2) );
  XOR2_X1 KeyArray_S10reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS11ser[0]), .B(KeyArray_outS20ser[0]), .Z(
        KeyArray_S10reg_gff_1_SFF_0_MUXInst_X) );
  AND2_X1 KeyArray_S10reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A1(KeyArray_n22), 
        .A2(KeyArray_S10reg_gff_1_SFF_0_MUXInst_X), .ZN(
        KeyArray_S10reg_gff_1_SFF_0_MUXInst_Y) );
  XOR2_X1 KeyArray_S10reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A(
        KeyArray_S10reg_gff_1_SFF_0_MUXInst_Y), .B(KeyArray_outS11ser[0]), .Z(
        KeyArray_S10reg_gff_1_SFF_0_QD) );
  INV_X1 KeyArray_S10reg_gff_1_SFF_0_Q_reg_U1 ( .A(KeyArray_outS10ser[0]), 
        .ZN(KeyArray_S10reg_gff_1_SFF_0_n10) );
  DFF_X1 KeyArray_S10reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        KeyArray_S10reg_gff_1_SFF_0_n5), .CK(clk), .Q(KeyArray_outS10ser[0]), 
        .QN() );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_1_U3 ( .A1(KeyArray_S10reg_gff_1_SFF_1_n2), .A2(KeyArray_S10reg_gff_1_SFF_1_n1), .ZN(KeyArray_S10reg_gff_1_SFF_1_n5) );
  OR2_X1 KeyArray_S10reg_gff_1_SFF_1_U2 ( .A1(KeyArray_n19), .A2(
        KeyArray_S10reg_gff_1_SFF_1_n10), .ZN(KeyArray_S10reg_gff_1_SFF_1_n1)
         );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_1_U1 ( .A1(KeyArray_S10reg_gff_1_SFF_1_QD), .A2(KeyArray_n19), .ZN(KeyArray_S10reg_gff_1_SFF_1_n2) );
  XOR2_X1 KeyArray_S10reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS11ser[1]), .B(KeyArray_outS20ser[1]), .Z(
        KeyArray_S10reg_gff_1_SFF_1_MUXInst_X) );
  AND2_X1 KeyArray_S10reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A1(KeyArray_n22), 
        .A2(KeyArray_S10reg_gff_1_SFF_1_MUXInst_X), .ZN(
        KeyArray_S10reg_gff_1_SFF_1_MUXInst_Y) );
  XOR2_X1 KeyArray_S10reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A(
        KeyArray_S10reg_gff_1_SFF_1_MUXInst_Y), .B(KeyArray_outS11ser[1]), .Z(
        KeyArray_S10reg_gff_1_SFF_1_QD) );
  INV_X1 KeyArray_S10reg_gff_1_SFF_1_Q_reg_U1 ( .A(KeyArray_outS10ser[1]), 
        .ZN(KeyArray_S10reg_gff_1_SFF_1_n10) );
  DFF_X1 KeyArray_S10reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        KeyArray_S10reg_gff_1_SFF_1_n5), .CK(clk), .Q(KeyArray_outS10ser[1]), 
        .QN() );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_2_U3 ( .A1(KeyArray_S10reg_gff_1_SFF_2_n2), .A2(KeyArray_S10reg_gff_1_SFF_2_n1), .ZN(KeyArray_S10reg_gff_1_SFF_2_n5) );
  OR2_X1 KeyArray_S10reg_gff_1_SFF_2_U2 ( .A1(KeyArray_n19), .A2(
        KeyArray_S10reg_gff_1_SFF_2_n10), .ZN(KeyArray_S10reg_gff_1_SFF_2_n1)
         );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_2_U1 ( .A1(KeyArray_S10reg_gff_1_SFF_2_QD), .A2(KeyArray_n19), .ZN(KeyArray_S10reg_gff_1_SFF_2_n2) );
  XOR2_X1 KeyArray_S10reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS11ser[2]), .B(KeyArray_outS20ser[2]), .Z(
        KeyArray_S10reg_gff_1_SFF_2_MUXInst_X) );
  AND2_X1 KeyArray_S10reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A1(KeyArray_n22), 
        .A2(KeyArray_S10reg_gff_1_SFF_2_MUXInst_X), .ZN(
        KeyArray_S10reg_gff_1_SFF_2_MUXInst_Y) );
  XOR2_X1 KeyArray_S10reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A(
        KeyArray_S10reg_gff_1_SFF_2_MUXInst_Y), .B(KeyArray_outS11ser[2]), .Z(
        KeyArray_S10reg_gff_1_SFF_2_QD) );
  INV_X1 KeyArray_S10reg_gff_1_SFF_2_Q_reg_U1 ( .A(KeyArray_outS10ser[2]), 
        .ZN(KeyArray_S10reg_gff_1_SFF_2_n10) );
  DFF_X1 KeyArray_S10reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        KeyArray_S10reg_gff_1_SFF_2_n5), .CK(clk), .Q(KeyArray_outS10ser[2]), 
        .QN() );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_3_U3 ( .A1(KeyArray_S10reg_gff_1_SFF_3_n2), .A2(KeyArray_S10reg_gff_1_SFF_3_n1), .ZN(KeyArray_S10reg_gff_1_SFF_3_n5) );
  OR2_X1 KeyArray_S10reg_gff_1_SFF_3_U2 ( .A1(KeyArray_n19), .A2(
        KeyArray_S10reg_gff_1_SFF_3_n10), .ZN(KeyArray_S10reg_gff_1_SFF_3_n1)
         );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_3_U1 ( .A1(KeyArray_S10reg_gff_1_SFF_3_QD), .A2(KeyArray_n19), .ZN(KeyArray_S10reg_gff_1_SFF_3_n2) );
  XOR2_X1 KeyArray_S10reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS11ser[3]), .B(KeyArray_outS20ser[3]), .Z(
        KeyArray_S10reg_gff_1_SFF_3_MUXInst_X) );
  AND2_X1 KeyArray_S10reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A1(KeyArray_n22), 
        .A2(KeyArray_S10reg_gff_1_SFF_3_MUXInst_X), .ZN(
        KeyArray_S10reg_gff_1_SFF_3_MUXInst_Y) );
  XOR2_X1 KeyArray_S10reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A(
        KeyArray_S10reg_gff_1_SFF_3_MUXInst_Y), .B(KeyArray_outS11ser[3]), .Z(
        KeyArray_S10reg_gff_1_SFF_3_QD) );
  INV_X1 KeyArray_S10reg_gff_1_SFF_3_Q_reg_U1 ( .A(KeyArray_outS10ser[3]), 
        .ZN(KeyArray_S10reg_gff_1_SFF_3_n10) );
  DFF_X1 KeyArray_S10reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        KeyArray_S10reg_gff_1_SFF_3_n5), .CK(clk), .Q(KeyArray_outS10ser[3]), 
        .QN() );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_4_U3 ( .A1(KeyArray_S10reg_gff_1_SFF_4_n2), .A2(KeyArray_S10reg_gff_1_SFF_4_n1), .ZN(KeyArray_S10reg_gff_1_SFF_4_n5) );
  OR2_X1 KeyArray_S10reg_gff_1_SFF_4_U2 ( .A1(KeyArray_n19), .A2(
        KeyArray_S10reg_gff_1_SFF_4_n10), .ZN(KeyArray_S10reg_gff_1_SFF_4_n1)
         );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_4_U1 ( .A1(KeyArray_S10reg_gff_1_SFF_4_QD), .A2(KeyArray_n19), .ZN(KeyArray_S10reg_gff_1_SFF_4_n2) );
  XOR2_X1 KeyArray_S10reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS11ser[4]), .B(KeyArray_outS20ser[4]), .Z(
        KeyArray_S10reg_gff_1_SFF_4_MUXInst_X) );
  AND2_X1 KeyArray_S10reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A1(KeyArray_n22), 
        .A2(KeyArray_S10reg_gff_1_SFF_4_MUXInst_X), .ZN(
        KeyArray_S10reg_gff_1_SFF_4_MUXInst_Y) );
  XOR2_X1 KeyArray_S10reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A(
        KeyArray_S10reg_gff_1_SFF_4_MUXInst_Y), .B(KeyArray_outS11ser[4]), .Z(
        KeyArray_S10reg_gff_1_SFF_4_QD) );
  INV_X1 KeyArray_S10reg_gff_1_SFF_4_Q_reg_U1 ( .A(KeyArray_outS10ser[4]), 
        .ZN(KeyArray_S10reg_gff_1_SFF_4_n10) );
  DFF_X1 KeyArray_S10reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        KeyArray_S10reg_gff_1_SFF_4_n5), .CK(clk), .Q(KeyArray_outS10ser[4]), 
        .QN() );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_5_U3 ( .A1(KeyArray_S10reg_gff_1_SFF_5_n2), .A2(KeyArray_S10reg_gff_1_SFF_5_n1), .ZN(KeyArray_S10reg_gff_1_SFF_5_n5) );
  OR2_X1 KeyArray_S10reg_gff_1_SFF_5_U2 ( .A1(KeyArray_n19), .A2(
        KeyArray_S10reg_gff_1_SFF_5_n10), .ZN(KeyArray_S10reg_gff_1_SFF_5_n1)
         );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_5_U1 ( .A1(KeyArray_S10reg_gff_1_SFF_5_QD), .A2(KeyArray_n19), .ZN(KeyArray_S10reg_gff_1_SFF_5_n2) );
  XOR2_X1 KeyArray_S10reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS11ser[5]), .B(KeyArray_outS20ser[5]), .Z(
        KeyArray_S10reg_gff_1_SFF_5_MUXInst_X) );
  AND2_X1 KeyArray_S10reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A1(KeyArray_n22), 
        .A2(KeyArray_S10reg_gff_1_SFF_5_MUXInst_X), .ZN(
        KeyArray_S10reg_gff_1_SFF_5_MUXInst_Y) );
  XOR2_X1 KeyArray_S10reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A(
        KeyArray_S10reg_gff_1_SFF_5_MUXInst_Y), .B(KeyArray_outS11ser[5]), .Z(
        KeyArray_S10reg_gff_1_SFF_5_QD) );
  INV_X1 KeyArray_S10reg_gff_1_SFF_5_Q_reg_U1 ( .A(KeyArray_outS10ser[5]), 
        .ZN(KeyArray_S10reg_gff_1_SFF_5_n10) );
  DFF_X1 KeyArray_S10reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        KeyArray_S10reg_gff_1_SFF_5_n5), .CK(clk), .Q(KeyArray_outS10ser[5]), 
        .QN() );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_6_U3 ( .A1(KeyArray_S10reg_gff_1_SFF_6_n2), .A2(KeyArray_S10reg_gff_1_SFF_6_n1), .ZN(KeyArray_S10reg_gff_1_SFF_6_n5) );
  OR2_X1 KeyArray_S10reg_gff_1_SFF_6_U2 ( .A1(KeyArray_n19), .A2(
        KeyArray_S10reg_gff_1_SFF_6_n10), .ZN(KeyArray_S10reg_gff_1_SFF_6_n1)
         );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_6_U1 ( .A1(KeyArray_S10reg_gff_1_SFF_6_QD), .A2(KeyArray_n19), .ZN(KeyArray_S10reg_gff_1_SFF_6_n2) );
  XOR2_X1 KeyArray_S10reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS11ser[6]), .B(KeyArray_outS20ser[6]), .Z(
        KeyArray_S10reg_gff_1_SFF_6_MUXInst_X) );
  AND2_X1 KeyArray_S10reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A1(KeyArray_n22), 
        .A2(KeyArray_S10reg_gff_1_SFF_6_MUXInst_X), .ZN(
        KeyArray_S10reg_gff_1_SFF_6_MUXInst_Y) );
  XOR2_X1 KeyArray_S10reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A(
        KeyArray_S10reg_gff_1_SFF_6_MUXInst_Y), .B(KeyArray_outS11ser[6]), .Z(
        KeyArray_S10reg_gff_1_SFF_6_QD) );
  INV_X1 KeyArray_S10reg_gff_1_SFF_6_Q_reg_U1 ( .A(KeyArray_outS10ser[6]), 
        .ZN(KeyArray_S10reg_gff_1_SFF_6_n10) );
  DFF_X1 KeyArray_S10reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        KeyArray_S10reg_gff_1_SFF_6_n5), .CK(clk), .Q(KeyArray_outS10ser[6]), 
        .QN() );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_7_U3 ( .A1(KeyArray_S10reg_gff_1_SFF_7_n2), .A2(KeyArray_S10reg_gff_1_SFF_7_n1), .ZN(KeyArray_S10reg_gff_1_SFF_7_n5) );
  OR2_X1 KeyArray_S10reg_gff_1_SFF_7_U2 ( .A1(KeyArray_n19), .A2(
        KeyArray_S10reg_gff_1_SFF_7_n10), .ZN(KeyArray_S10reg_gff_1_SFF_7_n1)
         );
  NAND2_X1 KeyArray_S10reg_gff_1_SFF_7_U1 ( .A1(KeyArray_S10reg_gff_1_SFF_7_QD), .A2(KeyArray_n19), .ZN(KeyArray_S10reg_gff_1_SFF_7_n2) );
  XOR2_X1 KeyArray_S10reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS11ser[7]), .B(KeyArray_outS20ser[7]), .Z(
        KeyArray_S10reg_gff_1_SFF_7_MUXInst_X) );
  AND2_X1 KeyArray_S10reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A1(KeyArray_n22), 
        .A2(KeyArray_S10reg_gff_1_SFF_7_MUXInst_X), .ZN(
        KeyArray_S10reg_gff_1_SFF_7_MUXInst_Y) );
  XOR2_X1 KeyArray_S10reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A(
        KeyArray_S10reg_gff_1_SFF_7_MUXInst_Y), .B(KeyArray_outS11ser[7]), .Z(
        KeyArray_S10reg_gff_1_SFF_7_QD) );
  INV_X1 KeyArray_S10reg_gff_1_SFF_7_Q_reg_U1 ( .A(KeyArray_outS10ser[7]), 
        .ZN(KeyArray_S10reg_gff_1_SFF_7_n10) );
  DFF_X1 KeyArray_S10reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        KeyArray_S10reg_gff_1_SFF_7_n5), .CK(clk), .Q(KeyArray_outS10ser[7]), 
        .QN() );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_0_U3 ( .A1(KeyArray_S11reg_gff_1_SFF_0_n2), .A2(KeyArray_S11reg_gff_1_SFF_0_n1), .ZN(KeyArray_S11reg_gff_1_SFF_0_n6) );
  OR2_X1 KeyArray_S11reg_gff_1_SFF_0_U2 ( .A1(KeyArray_n19), .A2(
        KeyArray_S11reg_gff_1_SFF_0_n11), .ZN(KeyArray_S11reg_gff_1_SFF_0_n1)
         );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_0_U1 ( .A1(KeyArray_S11reg_gff_1_SFF_0_QD), .A2(KeyArray_n19), .ZN(KeyArray_S11reg_gff_1_SFF_0_n2) );
  XOR2_X1 KeyArray_S11reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS12ser[0]), .B(KeyArray_outS21ser[0]), .Z(
        KeyArray_S11reg_gff_1_SFF_0_MUXInst_X) );
  AND2_X1 KeyArray_S11reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A1(KeyArray_n22), 
        .A2(KeyArray_S11reg_gff_1_SFF_0_MUXInst_X), .ZN(
        KeyArray_S11reg_gff_1_SFF_0_MUXInst_Y) );
  XOR2_X1 KeyArray_S11reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A(
        KeyArray_S11reg_gff_1_SFF_0_MUXInst_Y), .B(KeyArray_outS12ser[0]), .Z(
        KeyArray_S11reg_gff_1_SFF_0_QD) );
  INV_X1 KeyArray_S11reg_gff_1_SFF_0_Q_reg_U1 ( .A(KeyArray_outS11ser[0]), 
        .ZN(KeyArray_S11reg_gff_1_SFF_0_n11) );
  DFF_X1 KeyArray_S11reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        KeyArray_S11reg_gff_1_SFF_0_n6), .CK(clk), .Q(KeyArray_outS11ser[0]), 
        .QN() );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_1_U3 ( .A1(KeyArray_S11reg_gff_1_SFF_1_n2), .A2(KeyArray_S11reg_gff_1_SFF_1_n1), .ZN(KeyArray_S11reg_gff_1_SFF_1_n6) );
  OR2_X1 KeyArray_S11reg_gff_1_SFF_1_U2 ( .A1(KeyArray_n19), .A2(
        KeyArray_S11reg_gff_1_SFF_1_n11), .ZN(KeyArray_S11reg_gff_1_SFF_1_n1)
         );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_1_U1 ( .A1(KeyArray_S11reg_gff_1_SFF_1_QD), .A2(KeyArray_n19), .ZN(KeyArray_S11reg_gff_1_SFF_1_n2) );
  XOR2_X1 KeyArray_S11reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS12ser[1]), .B(KeyArray_outS21ser[1]), .Z(
        KeyArray_S11reg_gff_1_SFF_1_MUXInst_X) );
  AND2_X1 KeyArray_S11reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A1(KeyArray_n22), 
        .A2(KeyArray_S11reg_gff_1_SFF_1_MUXInst_X), .ZN(
        KeyArray_S11reg_gff_1_SFF_1_MUXInst_Y) );
  XOR2_X1 KeyArray_S11reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A(
        KeyArray_S11reg_gff_1_SFF_1_MUXInst_Y), .B(KeyArray_outS12ser[1]), .Z(
        KeyArray_S11reg_gff_1_SFF_1_QD) );
  INV_X1 KeyArray_S11reg_gff_1_SFF_1_Q_reg_U1 ( .A(KeyArray_outS11ser[1]), 
        .ZN(KeyArray_S11reg_gff_1_SFF_1_n11) );
  DFF_X1 KeyArray_S11reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        KeyArray_S11reg_gff_1_SFF_1_n6), .CK(clk), .Q(KeyArray_outS11ser[1]), 
        .QN() );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_2_U3 ( .A1(KeyArray_S11reg_gff_1_SFF_2_n2), .A2(KeyArray_S11reg_gff_1_SFF_2_n1), .ZN(KeyArray_S11reg_gff_1_SFF_2_n6) );
  OR2_X1 KeyArray_S11reg_gff_1_SFF_2_U2 ( .A1(KeyArray_n19), .A2(
        KeyArray_S11reg_gff_1_SFF_2_n11), .ZN(KeyArray_S11reg_gff_1_SFF_2_n1)
         );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_2_U1 ( .A1(KeyArray_S11reg_gff_1_SFF_2_QD), .A2(KeyArray_n19), .ZN(KeyArray_S11reg_gff_1_SFF_2_n2) );
  XOR2_X1 KeyArray_S11reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS12ser[2]), .B(KeyArray_outS21ser[2]), .Z(
        KeyArray_S11reg_gff_1_SFF_2_MUXInst_X) );
  AND2_X1 KeyArray_S11reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A1(KeyArray_n22), 
        .A2(KeyArray_S11reg_gff_1_SFF_2_MUXInst_X), .ZN(
        KeyArray_S11reg_gff_1_SFF_2_MUXInst_Y) );
  XOR2_X1 KeyArray_S11reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A(
        KeyArray_S11reg_gff_1_SFF_2_MUXInst_Y), .B(KeyArray_outS12ser[2]), .Z(
        KeyArray_S11reg_gff_1_SFF_2_QD) );
  INV_X1 KeyArray_S11reg_gff_1_SFF_2_Q_reg_U1 ( .A(KeyArray_outS11ser[2]), 
        .ZN(KeyArray_S11reg_gff_1_SFF_2_n11) );
  DFF_X1 KeyArray_S11reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        KeyArray_S11reg_gff_1_SFF_2_n6), .CK(clk), .Q(KeyArray_outS11ser[2]), 
        .QN() );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_3_U3 ( .A1(KeyArray_S11reg_gff_1_SFF_3_n2), .A2(KeyArray_S11reg_gff_1_SFF_3_n1), .ZN(KeyArray_S11reg_gff_1_SFF_3_n6) );
  OR2_X1 KeyArray_S11reg_gff_1_SFF_3_U2 ( .A1(KeyArray_n19), .A2(
        KeyArray_S11reg_gff_1_SFF_3_n11), .ZN(KeyArray_S11reg_gff_1_SFF_3_n1)
         );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_3_U1 ( .A1(KeyArray_S11reg_gff_1_SFF_3_QD), .A2(KeyArray_n19), .ZN(KeyArray_S11reg_gff_1_SFF_3_n2) );
  XOR2_X1 KeyArray_S11reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS12ser[3]), .B(KeyArray_outS21ser[3]), .Z(
        KeyArray_S11reg_gff_1_SFF_3_MUXInst_X) );
  AND2_X1 KeyArray_S11reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A1(KeyArray_n22), 
        .A2(KeyArray_S11reg_gff_1_SFF_3_MUXInst_X), .ZN(
        KeyArray_S11reg_gff_1_SFF_3_MUXInst_Y) );
  XOR2_X1 KeyArray_S11reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A(
        KeyArray_S11reg_gff_1_SFF_3_MUXInst_Y), .B(KeyArray_outS12ser[3]), .Z(
        KeyArray_S11reg_gff_1_SFF_3_QD) );
  INV_X1 KeyArray_S11reg_gff_1_SFF_3_Q_reg_U1 ( .A(KeyArray_outS11ser[3]), 
        .ZN(KeyArray_S11reg_gff_1_SFF_3_n11) );
  DFF_X1 KeyArray_S11reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        KeyArray_S11reg_gff_1_SFF_3_n6), .CK(clk), .Q(KeyArray_outS11ser[3]), 
        .QN() );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_4_U3 ( .A1(KeyArray_S11reg_gff_1_SFF_4_n2), .A2(KeyArray_S11reg_gff_1_SFF_4_n1), .ZN(KeyArray_S11reg_gff_1_SFF_4_n6) );
  OR2_X1 KeyArray_S11reg_gff_1_SFF_4_U2 ( .A1(KeyArray_n19), .A2(
        KeyArray_S11reg_gff_1_SFF_4_n11), .ZN(KeyArray_S11reg_gff_1_SFF_4_n1)
         );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_4_U1 ( .A1(KeyArray_S11reg_gff_1_SFF_4_QD), .A2(KeyArray_n19), .ZN(KeyArray_S11reg_gff_1_SFF_4_n2) );
  XOR2_X1 KeyArray_S11reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS12ser[4]), .B(KeyArray_outS21ser[4]), .Z(
        KeyArray_S11reg_gff_1_SFF_4_MUXInst_X) );
  AND2_X1 KeyArray_S11reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A1(KeyArray_n22), 
        .A2(KeyArray_S11reg_gff_1_SFF_4_MUXInst_X), .ZN(
        KeyArray_S11reg_gff_1_SFF_4_MUXInst_Y) );
  XOR2_X1 KeyArray_S11reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A(
        KeyArray_S11reg_gff_1_SFF_4_MUXInst_Y), .B(KeyArray_outS12ser[4]), .Z(
        KeyArray_S11reg_gff_1_SFF_4_QD) );
  INV_X1 KeyArray_S11reg_gff_1_SFF_4_Q_reg_U1 ( .A(KeyArray_outS11ser[4]), 
        .ZN(KeyArray_S11reg_gff_1_SFF_4_n11) );
  DFF_X1 KeyArray_S11reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        KeyArray_S11reg_gff_1_SFF_4_n6), .CK(clk), .Q(KeyArray_outS11ser[4]), 
        .QN() );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_5_U3 ( .A1(KeyArray_S11reg_gff_1_SFF_5_n2), .A2(KeyArray_S11reg_gff_1_SFF_5_n1), .ZN(KeyArray_S11reg_gff_1_SFF_5_n6) );
  OR2_X1 KeyArray_S11reg_gff_1_SFF_5_U2 ( .A1(KeyArray_n19), .A2(
        KeyArray_S11reg_gff_1_SFF_5_n11), .ZN(KeyArray_S11reg_gff_1_SFF_5_n1)
         );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_5_U1 ( .A1(KeyArray_S11reg_gff_1_SFF_5_QD), .A2(KeyArray_n19), .ZN(KeyArray_S11reg_gff_1_SFF_5_n2) );
  XOR2_X1 KeyArray_S11reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS12ser[5]), .B(KeyArray_outS21ser[5]), .Z(
        KeyArray_S11reg_gff_1_SFF_5_MUXInst_X) );
  AND2_X1 KeyArray_S11reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A1(KeyArray_n22), 
        .A2(KeyArray_S11reg_gff_1_SFF_5_MUXInst_X), .ZN(
        KeyArray_S11reg_gff_1_SFF_5_MUXInst_Y) );
  XOR2_X1 KeyArray_S11reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A(
        KeyArray_S11reg_gff_1_SFF_5_MUXInst_Y), .B(KeyArray_outS12ser[5]), .Z(
        KeyArray_S11reg_gff_1_SFF_5_QD) );
  INV_X1 KeyArray_S11reg_gff_1_SFF_5_Q_reg_U1 ( .A(KeyArray_outS11ser[5]), 
        .ZN(KeyArray_S11reg_gff_1_SFF_5_n11) );
  DFF_X1 KeyArray_S11reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        KeyArray_S11reg_gff_1_SFF_5_n6), .CK(clk), .Q(KeyArray_outS11ser[5]), 
        .QN() );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_6_U3 ( .A1(KeyArray_S11reg_gff_1_SFF_6_n2), .A2(KeyArray_S11reg_gff_1_SFF_6_n1), .ZN(KeyArray_S11reg_gff_1_SFF_6_n6) );
  OR2_X1 KeyArray_S11reg_gff_1_SFF_6_U2 ( .A1(KeyArray_n19), .A2(
        KeyArray_S11reg_gff_1_SFF_6_n11), .ZN(KeyArray_S11reg_gff_1_SFF_6_n1)
         );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_6_U1 ( .A1(KeyArray_S11reg_gff_1_SFF_6_QD), .A2(KeyArray_n19), .ZN(KeyArray_S11reg_gff_1_SFF_6_n2) );
  XOR2_X1 KeyArray_S11reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS12ser[6]), .B(KeyArray_outS21ser[6]), .Z(
        KeyArray_S11reg_gff_1_SFF_6_MUXInst_X) );
  AND2_X1 KeyArray_S11reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A1(KeyArray_n22), 
        .A2(KeyArray_S11reg_gff_1_SFF_6_MUXInst_X), .ZN(
        KeyArray_S11reg_gff_1_SFF_6_MUXInst_Y) );
  XOR2_X1 KeyArray_S11reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A(
        KeyArray_S11reg_gff_1_SFF_6_MUXInst_Y), .B(KeyArray_outS12ser[6]), .Z(
        KeyArray_S11reg_gff_1_SFF_6_QD) );
  INV_X1 KeyArray_S11reg_gff_1_SFF_6_Q_reg_U1 ( .A(KeyArray_outS11ser[6]), 
        .ZN(KeyArray_S11reg_gff_1_SFF_6_n11) );
  DFF_X1 KeyArray_S11reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        KeyArray_S11reg_gff_1_SFF_6_n6), .CK(clk), .Q(KeyArray_outS11ser[6]), 
        .QN() );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_7_U3 ( .A1(KeyArray_S11reg_gff_1_SFF_7_n2), .A2(KeyArray_S11reg_gff_1_SFF_7_n1), .ZN(KeyArray_S11reg_gff_1_SFF_7_n6) );
  OR2_X1 KeyArray_S11reg_gff_1_SFF_7_U2 ( .A1(KeyArray_n19), .A2(
        KeyArray_S11reg_gff_1_SFF_7_n11), .ZN(KeyArray_S11reg_gff_1_SFF_7_n1)
         );
  NAND2_X1 KeyArray_S11reg_gff_1_SFF_7_U1 ( .A1(KeyArray_S11reg_gff_1_SFF_7_QD), .A2(KeyArray_n19), .ZN(KeyArray_S11reg_gff_1_SFF_7_n2) );
  XOR2_X1 KeyArray_S11reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS12ser[7]), .B(KeyArray_outS21ser[7]), .Z(
        KeyArray_S11reg_gff_1_SFF_7_MUXInst_X) );
  AND2_X1 KeyArray_S11reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A1(KeyArray_n22), 
        .A2(KeyArray_S11reg_gff_1_SFF_7_MUXInst_X), .ZN(
        KeyArray_S11reg_gff_1_SFF_7_MUXInst_Y) );
  XOR2_X1 KeyArray_S11reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A(
        KeyArray_S11reg_gff_1_SFF_7_MUXInst_Y), .B(KeyArray_outS12ser[7]), .Z(
        KeyArray_S11reg_gff_1_SFF_7_QD) );
  INV_X1 KeyArray_S11reg_gff_1_SFF_7_Q_reg_U1 ( .A(KeyArray_outS11ser[7]), 
        .ZN(KeyArray_S11reg_gff_1_SFF_7_n11) );
  DFF_X1 KeyArray_S11reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        KeyArray_S11reg_gff_1_SFF_7_n6), .CK(clk), .Q(KeyArray_outS11ser[7]), 
        .QN() );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_0_U3 ( .A1(KeyArray_S12reg_gff_1_SFF_0_n2), .A2(KeyArray_S12reg_gff_1_SFF_0_n1), .ZN(KeyArray_S12reg_gff_1_SFF_0_n6) );
  OR2_X1 KeyArray_S12reg_gff_1_SFF_0_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S12reg_gff_1_SFF_0_n11), .ZN(KeyArray_S12reg_gff_1_SFF_0_n1)
         );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_0_U1 ( .A1(KeyArray_S12reg_gff_1_SFF_0_QD), .A2(KeyArray_n18), .ZN(KeyArray_S12reg_gff_1_SFF_0_n2) );
  XOR2_X1 KeyArray_S12reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A(keySBIn[0]), .B(
        KeyArray_outS22ser[0]), .Z(KeyArray_S12reg_gff_1_SFF_0_MUXInst_X) );
  AND2_X1 KeyArray_S12reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A1(KeyArray_n22), 
        .A2(KeyArray_S12reg_gff_1_SFF_0_MUXInst_X), .ZN(
        KeyArray_S12reg_gff_1_SFF_0_MUXInst_Y) );
  XOR2_X1 KeyArray_S12reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A(
        KeyArray_S12reg_gff_1_SFF_0_MUXInst_Y), .B(keySBIn[0]), .Z(
        KeyArray_S12reg_gff_1_SFF_0_QD) );
  INV_X1 KeyArray_S12reg_gff_1_SFF_0_Q_reg_U1 ( .A(KeyArray_outS12ser[0]), 
        .ZN(KeyArray_S12reg_gff_1_SFF_0_n11) );
  DFF_X1 KeyArray_S12reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        KeyArray_S12reg_gff_1_SFF_0_n6), .CK(clk), .Q(KeyArray_outS12ser[0]), 
        .QN() );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_1_U3 ( .A1(KeyArray_S12reg_gff_1_SFF_1_n2), .A2(KeyArray_S12reg_gff_1_SFF_1_n1), .ZN(KeyArray_S12reg_gff_1_SFF_1_n6) );
  OR2_X1 KeyArray_S12reg_gff_1_SFF_1_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S12reg_gff_1_SFF_1_n11), .ZN(KeyArray_S12reg_gff_1_SFF_1_n1)
         );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_1_U1 ( .A1(KeyArray_S12reg_gff_1_SFF_1_QD), .A2(KeyArray_n18), .ZN(KeyArray_S12reg_gff_1_SFF_1_n2) );
  XOR2_X1 KeyArray_S12reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A(keySBIn[1]), .B(
        KeyArray_outS22ser[1]), .Z(KeyArray_S12reg_gff_1_SFF_1_MUXInst_X) );
  AND2_X1 KeyArray_S12reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A1(KeyArray_n22), 
        .A2(KeyArray_S12reg_gff_1_SFF_1_MUXInst_X), .ZN(
        KeyArray_S12reg_gff_1_SFF_1_MUXInst_Y) );
  XOR2_X1 KeyArray_S12reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A(
        KeyArray_S12reg_gff_1_SFF_1_MUXInst_Y), .B(keySBIn[1]), .Z(
        KeyArray_S12reg_gff_1_SFF_1_QD) );
  INV_X1 KeyArray_S12reg_gff_1_SFF_1_Q_reg_U1 ( .A(KeyArray_outS12ser[1]), 
        .ZN(KeyArray_S12reg_gff_1_SFF_1_n11) );
  DFF_X1 KeyArray_S12reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        KeyArray_S12reg_gff_1_SFF_1_n6), .CK(clk), .Q(KeyArray_outS12ser[1]), 
        .QN() );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_2_U3 ( .A1(KeyArray_S12reg_gff_1_SFF_2_n2), .A2(KeyArray_S12reg_gff_1_SFF_2_n1), .ZN(KeyArray_S12reg_gff_1_SFF_2_n6) );
  OR2_X1 KeyArray_S12reg_gff_1_SFF_2_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S12reg_gff_1_SFF_2_n11), .ZN(KeyArray_S12reg_gff_1_SFF_2_n1)
         );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_2_U1 ( .A1(KeyArray_S12reg_gff_1_SFF_2_QD), .A2(KeyArray_n18), .ZN(KeyArray_S12reg_gff_1_SFF_2_n2) );
  XOR2_X1 KeyArray_S12reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A(keySBIn[2]), .B(
        KeyArray_outS22ser[2]), .Z(KeyArray_S12reg_gff_1_SFF_2_MUXInst_X) );
  AND2_X1 KeyArray_S12reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A1(KeyArray_n22), 
        .A2(KeyArray_S12reg_gff_1_SFF_2_MUXInst_X), .ZN(
        KeyArray_S12reg_gff_1_SFF_2_MUXInst_Y) );
  XOR2_X1 KeyArray_S12reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A(
        KeyArray_S12reg_gff_1_SFF_2_MUXInst_Y), .B(keySBIn[2]), .Z(
        KeyArray_S12reg_gff_1_SFF_2_QD) );
  INV_X1 KeyArray_S12reg_gff_1_SFF_2_Q_reg_U1 ( .A(KeyArray_outS12ser[2]), 
        .ZN(KeyArray_S12reg_gff_1_SFF_2_n11) );
  DFF_X1 KeyArray_S12reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        KeyArray_S12reg_gff_1_SFF_2_n6), .CK(clk), .Q(KeyArray_outS12ser[2]), 
        .QN() );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_3_U3 ( .A1(KeyArray_S12reg_gff_1_SFF_3_n2), .A2(KeyArray_S12reg_gff_1_SFF_3_n1), .ZN(KeyArray_S12reg_gff_1_SFF_3_n6) );
  OR2_X1 KeyArray_S12reg_gff_1_SFF_3_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S12reg_gff_1_SFF_3_n11), .ZN(KeyArray_S12reg_gff_1_SFF_3_n1)
         );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_3_U1 ( .A1(KeyArray_S12reg_gff_1_SFF_3_QD), .A2(KeyArray_n18), .ZN(KeyArray_S12reg_gff_1_SFF_3_n2) );
  XOR2_X1 KeyArray_S12reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A(keySBIn[3]), .B(
        KeyArray_outS22ser[3]), .Z(KeyArray_S12reg_gff_1_SFF_3_MUXInst_X) );
  AND2_X1 KeyArray_S12reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A1(KeyArray_n22), 
        .A2(KeyArray_S12reg_gff_1_SFF_3_MUXInst_X), .ZN(
        KeyArray_S12reg_gff_1_SFF_3_MUXInst_Y) );
  XOR2_X1 KeyArray_S12reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A(
        KeyArray_S12reg_gff_1_SFF_3_MUXInst_Y), .B(keySBIn[3]), .Z(
        KeyArray_S12reg_gff_1_SFF_3_QD) );
  INV_X1 KeyArray_S12reg_gff_1_SFF_3_Q_reg_U1 ( .A(KeyArray_outS12ser[3]), 
        .ZN(KeyArray_S12reg_gff_1_SFF_3_n11) );
  DFF_X1 KeyArray_S12reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        KeyArray_S12reg_gff_1_SFF_3_n6), .CK(clk), .Q(KeyArray_outS12ser[3]), 
        .QN() );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_4_U3 ( .A1(KeyArray_S12reg_gff_1_SFF_4_n2), .A2(KeyArray_S12reg_gff_1_SFF_4_n1), .ZN(KeyArray_S12reg_gff_1_SFF_4_n6) );
  OR2_X1 KeyArray_S12reg_gff_1_SFF_4_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S12reg_gff_1_SFF_4_n11), .ZN(KeyArray_S12reg_gff_1_SFF_4_n1)
         );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_4_U1 ( .A1(KeyArray_S12reg_gff_1_SFF_4_QD), .A2(KeyArray_n18), .ZN(KeyArray_S12reg_gff_1_SFF_4_n2) );
  XOR2_X1 KeyArray_S12reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A(keySBIn[4]), .B(
        KeyArray_outS22ser[4]), .Z(KeyArray_S12reg_gff_1_SFF_4_MUXInst_X) );
  AND2_X1 KeyArray_S12reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A1(KeyArray_n22), 
        .A2(KeyArray_S12reg_gff_1_SFF_4_MUXInst_X), .ZN(
        KeyArray_S12reg_gff_1_SFF_4_MUXInst_Y) );
  XOR2_X1 KeyArray_S12reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A(
        KeyArray_S12reg_gff_1_SFF_4_MUXInst_Y), .B(keySBIn[4]), .Z(
        KeyArray_S12reg_gff_1_SFF_4_QD) );
  INV_X1 KeyArray_S12reg_gff_1_SFF_4_Q_reg_U1 ( .A(KeyArray_outS12ser[4]), 
        .ZN(KeyArray_S12reg_gff_1_SFF_4_n11) );
  DFF_X1 KeyArray_S12reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        KeyArray_S12reg_gff_1_SFF_4_n6), .CK(clk), .Q(KeyArray_outS12ser[4]), 
        .QN() );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_5_U3 ( .A1(KeyArray_S12reg_gff_1_SFF_5_n2), .A2(KeyArray_S12reg_gff_1_SFF_5_n1), .ZN(KeyArray_S12reg_gff_1_SFF_5_n6) );
  OR2_X1 KeyArray_S12reg_gff_1_SFF_5_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S12reg_gff_1_SFF_5_n11), .ZN(KeyArray_S12reg_gff_1_SFF_5_n1)
         );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_5_U1 ( .A1(KeyArray_S12reg_gff_1_SFF_5_QD), .A2(KeyArray_n18), .ZN(KeyArray_S12reg_gff_1_SFF_5_n2) );
  XOR2_X1 KeyArray_S12reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A(keySBIn[5]), .B(
        KeyArray_outS22ser[5]), .Z(KeyArray_S12reg_gff_1_SFF_5_MUXInst_X) );
  AND2_X1 KeyArray_S12reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A1(KeyArray_n22), 
        .A2(KeyArray_S12reg_gff_1_SFF_5_MUXInst_X), .ZN(
        KeyArray_S12reg_gff_1_SFF_5_MUXInst_Y) );
  XOR2_X1 KeyArray_S12reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A(
        KeyArray_S12reg_gff_1_SFF_5_MUXInst_Y), .B(keySBIn[5]), .Z(
        KeyArray_S12reg_gff_1_SFF_5_QD) );
  INV_X1 KeyArray_S12reg_gff_1_SFF_5_Q_reg_U1 ( .A(KeyArray_outS12ser[5]), 
        .ZN(KeyArray_S12reg_gff_1_SFF_5_n11) );
  DFF_X1 KeyArray_S12reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        KeyArray_S12reg_gff_1_SFF_5_n6), .CK(clk), .Q(KeyArray_outS12ser[5]), 
        .QN() );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_6_U3 ( .A1(KeyArray_S12reg_gff_1_SFF_6_n2), .A2(KeyArray_S12reg_gff_1_SFF_6_n1), .ZN(KeyArray_S12reg_gff_1_SFF_6_n6) );
  OR2_X1 KeyArray_S12reg_gff_1_SFF_6_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S12reg_gff_1_SFF_6_n11), .ZN(KeyArray_S12reg_gff_1_SFF_6_n1)
         );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_6_U1 ( .A1(KeyArray_S12reg_gff_1_SFF_6_QD), .A2(KeyArray_n18), .ZN(KeyArray_S12reg_gff_1_SFF_6_n2) );
  XOR2_X1 KeyArray_S12reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A(keySBIn[6]), .B(
        KeyArray_outS22ser[6]), .Z(KeyArray_S12reg_gff_1_SFF_6_MUXInst_X) );
  AND2_X1 KeyArray_S12reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A1(KeyArray_n22), 
        .A2(KeyArray_S12reg_gff_1_SFF_6_MUXInst_X), .ZN(
        KeyArray_S12reg_gff_1_SFF_6_MUXInst_Y) );
  XOR2_X1 KeyArray_S12reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A(
        KeyArray_S12reg_gff_1_SFF_6_MUXInst_Y), .B(keySBIn[6]), .Z(
        KeyArray_S12reg_gff_1_SFF_6_QD) );
  INV_X1 KeyArray_S12reg_gff_1_SFF_6_Q_reg_U1 ( .A(KeyArray_outS12ser[6]), 
        .ZN(KeyArray_S12reg_gff_1_SFF_6_n11) );
  DFF_X1 KeyArray_S12reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        KeyArray_S12reg_gff_1_SFF_6_n6), .CK(clk), .Q(KeyArray_outS12ser[6]), 
        .QN() );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_7_U3 ( .A1(KeyArray_S12reg_gff_1_SFF_7_n2), .A2(KeyArray_S12reg_gff_1_SFF_7_n1), .ZN(KeyArray_S12reg_gff_1_SFF_7_n6) );
  OR2_X1 KeyArray_S12reg_gff_1_SFF_7_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S12reg_gff_1_SFF_7_n11), .ZN(KeyArray_S12reg_gff_1_SFF_7_n1)
         );
  NAND2_X1 KeyArray_S12reg_gff_1_SFF_7_U1 ( .A1(KeyArray_S12reg_gff_1_SFF_7_QD), .A2(KeyArray_n18), .ZN(KeyArray_S12reg_gff_1_SFF_7_n2) );
  XOR2_X1 KeyArray_S12reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A(keySBIn[7]), .B(
        KeyArray_outS22ser[7]), .Z(KeyArray_S12reg_gff_1_SFF_7_MUXInst_X) );
  AND2_X1 KeyArray_S12reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A1(KeyArray_n22), 
        .A2(KeyArray_S12reg_gff_1_SFF_7_MUXInst_X), .ZN(
        KeyArray_S12reg_gff_1_SFF_7_MUXInst_Y) );
  XOR2_X1 KeyArray_S12reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A(
        KeyArray_S12reg_gff_1_SFF_7_MUXInst_Y), .B(keySBIn[7]), .Z(
        KeyArray_S12reg_gff_1_SFF_7_QD) );
  INV_X1 KeyArray_S12reg_gff_1_SFF_7_Q_reg_U1 ( .A(KeyArray_outS12ser[7]), 
        .ZN(KeyArray_S12reg_gff_1_SFF_7_n11) );
  DFF_X1 KeyArray_S12reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        KeyArray_S12reg_gff_1_SFF_7_n6), .CK(clk), .Q(KeyArray_outS12ser[7]), 
        .QN() );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_0_U3 ( .A1(KeyArray_S13reg_gff_1_SFF_0_n2), .A2(KeyArray_S13reg_gff_1_SFF_0_n1), .ZN(KeyArray_S13reg_gff_1_SFF_0_n6) );
  OR2_X1 KeyArray_S13reg_gff_1_SFF_0_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S13reg_gff_1_SFF_0_n11), .ZN(KeyArray_S13reg_gff_1_SFF_0_n1)
         );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_0_U1 ( .A1(KeyArray_S13reg_gff_1_SFF_0_QD), .A2(KeyArray_n18), .ZN(KeyArray_S13reg_gff_1_SFF_0_n2) );
  XOR2_X1 KeyArray_S13reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS20ser[0]), .B(KeyArray_outS23ser[0]), .Z(
        KeyArray_S13reg_gff_1_SFF_0_MUXInst_X) );
  AND2_X1 KeyArray_S13reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A1(KeyArray_n22), 
        .A2(KeyArray_S13reg_gff_1_SFF_0_MUXInst_X), .ZN(
        KeyArray_S13reg_gff_1_SFF_0_MUXInst_Y) );
  XOR2_X1 KeyArray_S13reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A(
        KeyArray_S13reg_gff_1_SFF_0_MUXInst_Y), .B(KeyArray_outS20ser[0]), .Z(
        KeyArray_S13reg_gff_1_SFF_0_QD) );
  INV_X1 KeyArray_S13reg_gff_1_SFF_0_Q_reg_U1 ( .A(keySBIn[0]), .ZN(
        KeyArray_S13reg_gff_1_SFF_0_n11) );
  DFF_X1 KeyArray_S13reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        KeyArray_S13reg_gff_1_SFF_0_n6), .CK(clk), .Q(keySBIn[0]), .QN() );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_1_U3 ( .A1(KeyArray_S13reg_gff_1_SFF_1_n2), .A2(KeyArray_S13reg_gff_1_SFF_1_n1), .ZN(KeyArray_S13reg_gff_1_SFF_1_n6) );
  OR2_X1 KeyArray_S13reg_gff_1_SFF_1_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S13reg_gff_1_SFF_1_n11), .ZN(KeyArray_S13reg_gff_1_SFF_1_n1)
         );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_1_U1 ( .A1(KeyArray_S13reg_gff_1_SFF_1_QD), .A2(KeyArray_n18), .ZN(KeyArray_S13reg_gff_1_SFF_1_n2) );
  XOR2_X1 KeyArray_S13reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS20ser[1]), .B(KeyArray_outS23ser[1]), .Z(
        KeyArray_S13reg_gff_1_SFF_1_MUXInst_X) );
  AND2_X1 KeyArray_S13reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A1(KeyArray_n22), 
        .A2(KeyArray_S13reg_gff_1_SFF_1_MUXInst_X), .ZN(
        KeyArray_S13reg_gff_1_SFF_1_MUXInst_Y) );
  XOR2_X1 KeyArray_S13reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A(
        KeyArray_S13reg_gff_1_SFF_1_MUXInst_Y), .B(KeyArray_outS20ser[1]), .Z(
        KeyArray_S13reg_gff_1_SFF_1_QD) );
  INV_X1 KeyArray_S13reg_gff_1_SFF_1_Q_reg_U1 ( .A(keySBIn[1]), .ZN(
        KeyArray_S13reg_gff_1_SFF_1_n11) );
  DFF_X1 KeyArray_S13reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        KeyArray_S13reg_gff_1_SFF_1_n6), .CK(clk), .Q(keySBIn[1]), .QN() );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_2_U3 ( .A1(KeyArray_S13reg_gff_1_SFF_2_n2), .A2(KeyArray_S13reg_gff_1_SFF_2_n1), .ZN(KeyArray_S13reg_gff_1_SFF_2_n6) );
  OR2_X1 KeyArray_S13reg_gff_1_SFF_2_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S13reg_gff_1_SFF_2_n11), .ZN(KeyArray_S13reg_gff_1_SFF_2_n1)
         );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_2_U1 ( .A1(KeyArray_S13reg_gff_1_SFF_2_QD), .A2(KeyArray_n18), .ZN(KeyArray_S13reg_gff_1_SFF_2_n2) );
  XOR2_X1 KeyArray_S13reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS20ser[2]), .B(KeyArray_outS23ser[2]), .Z(
        KeyArray_S13reg_gff_1_SFF_2_MUXInst_X) );
  AND2_X1 KeyArray_S13reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A1(KeyArray_n22), 
        .A2(KeyArray_S13reg_gff_1_SFF_2_MUXInst_X), .ZN(
        KeyArray_S13reg_gff_1_SFF_2_MUXInst_Y) );
  XOR2_X1 KeyArray_S13reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A(
        KeyArray_S13reg_gff_1_SFF_2_MUXInst_Y), .B(KeyArray_outS20ser[2]), .Z(
        KeyArray_S13reg_gff_1_SFF_2_QD) );
  INV_X1 KeyArray_S13reg_gff_1_SFF_2_Q_reg_U1 ( .A(keySBIn[2]), .ZN(
        KeyArray_S13reg_gff_1_SFF_2_n11) );
  DFF_X1 KeyArray_S13reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        KeyArray_S13reg_gff_1_SFF_2_n6), .CK(clk), .Q(keySBIn[2]), .QN() );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_3_U3 ( .A1(KeyArray_S13reg_gff_1_SFF_3_n2), .A2(KeyArray_S13reg_gff_1_SFF_3_n1), .ZN(KeyArray_S13reg_gff_1_SFF_3_n6) );
  OR2_X1 KeyArray_S13reg_gff_1_SFF_3_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S13reg_gff_1_SFF_3_n11), .ZN(KeyArray_S13reg_gff_1_SFF_3_n1)
         );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_3_U1 ( .A1(KeyArray_S13reg_gff_1_SFF_3_QD), .A2(KeyArray_n18), .ZN(KeyArray_S13reg_gff_1_SFF_3_n2) );
  XOR2_X1 KeyArray_S13reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS20ser[3]), .B(KeyArray_outS23ser[3]), .Z(
        KeyArray_S13reg_gff_1_SFF_3_MUXInst_X) );
  AND2_X1 KeyArray_S13reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A1(KeyArray_n22), 
        .A2(KeyArray_S13reg_gff_1_SFF_3_MUXInst_X), .ZN(
        KeyArray_S13reg_gff_1_SFF_3_MUXInst_Y) );
  XOR2_X1 KeyArray_S13reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A(
        KeyArray_S13reg_gff_1_SFF_3_MUXInst_Y), .B(KeyArray_outS20ser[3]), .Z(
        KeyArray_S13reg_gff_1_SFF_3_QD) );
  INV_X1 KeyArray_S13reg_gff_1_SFF_3_Q_reg_U1 ( .A(keySBIn[3]), .ZN(
        KeyArray_S13reg_gff_1_SFF_3_n11) );
  DFF_X1 KeyArray_S13reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        KeyArray_S13reg_gff_1_SFF_3_n6), .CK(clk), .Q(keySBIn[3]), .QN() );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_4_U3 ( .A1(KeyArray_S13reg_gff_1_SFF_4_n2), .A2(KeyArray_S13reg_gff_1_SFF_4_n1), .ZN(KeyArray_S13reg_gff_1_SFF_4_n6) );
  OR2_X1 KeyArray_S13reg_gff_1_SFF_4_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S13reg_gff_1_SFF_4_n11), .ZN(KeyArray_S13reg_gff_1_SFF_4_n1)
         );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_4_U1 ( .A1(KeyArray_S13reg_gff_1_SFF_4_QD), .A2(KeyArray_n18), .ZN(KeyArray_S13reg_gff_1_SFF_4_n2) );
  XOR2_X1 KeyArray_S13reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS20ser[4]), .B(KeyArray_outS23ser[4]), .Z(
        KeyArray_S13reg_gff_1_SFF_4_MUXInst_X) );
  AND2_X1 KeyArray_S13reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A1(KeyArray_n22), 
        .A2(KeyArray_S13reg_gff_1_SFF_4_MUXInst_X), .ZN(
        KeyArray_S13reg_gff_1_SFF_4_MUXInst_Y) );
  XOR2_X1 KeyArray_S13reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A(
        KeyArray_S13reg_gff_1_SFF_4_MUXInst_Y), .B(KeyArray_outS20ser[4]), .Z(
        KeyArray_S13reg_gff_1_SFF_4_QD) );
  INV_X1 KeyArray_S13reg_gff_1_SFF_4_Q_reg_U1 ( .A(keySBIn[4]), .ZN(
        KeyArray_S13reg_gff_1_SFF_4_n11) );
  DFF_X1 KeyArray_S13reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        KeyArray_S13reg_gff_1_SFF_4_n6), .CK(clk), .Q(keySBIn[4]), .QN() );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_5_U3 ( .A1(KeyArray_S13reg_gff_1_SFF_5_n2), .A2(KeyArray_S13reg_gff_1_SFF_5_n1), .ZN(KeyArray_S13reg_gff_1_SFF_5_n5) );
  OR2_X1 KeyArray_S13reg_gff_1_SFF_5_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S13reg_gff_1_SFF_5_n10), .ZN(KeyArray_S13reg_gff_1_SFF_5_n1)
         );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_5_U1 ( .A1(KeyArray_S13reg_gff_1_SFF_5_QD), .A2(KeyArray_n18), .ZN(KeyArray_S13reg_gff_1_SFF_5_n2) );
  XOR2_X1 KeyArray_S13reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS20ser[5]), .B(KeyArray_outS23ser[5]), .Z(
        KeyArray_S13reg_gff_1_SFF_5_MUXInst_X) );
  AND2_X1 KeyArray_S13reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A1(KeyArray_n22), 
        .A2(KeyArray_S13reg_gff_1_SFF_5_MUXInst_X), .ZN(
        KeyArray_S13reg_gff_1_SFF_5_MUXInst_Y) );
  XOR2_X1 KeyArray_S13reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A(
        KeyArray_S13reg_gff_1_SFF_5_MUXInst_Y), .B(KeyArray_outS20ser[5]), .Z(
        KeyArray_S13reg_gff_1_SFF_5_QD) );
  INV_X1 KeyArray_S13reg_gff_1_SFF_5_Q_reg_U1 ( .A(keySBIn[5]), .ZN(
        KeyArray_S13reg_gff_1_SFF_5_n10) );
  DFF_X1 KeyArray_S13reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        KeyArray_S13reg_gff_1_SFF_5_n5), .CK(clk), .Q(keySBIn[5]), .QN() );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_6_U3 ( .A1(KeyArray_S13reg_gff_1_SFF_6_n2), .A2(KeyArray_S13reg_gff_1_SFF_6_n1), .ZN(KeyArray_S13reg_gff_1_SFF_6_n5) );
  OR2_X1 KeyArray_S13reg_gff_1_SFF_6_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S13reg_gff_1_SFF_6_n10), .ZN(KeyArray_S13reg_gff_1_SFF_6_n1)
         );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_6_U1 ( .A1(KeyArray_S13reg_gff_1_SFF_6_QD), .A2(KeyArray_n18), .ZN(KeyArray_S13reg_gff_1_SFF_6_n2) );
  XOR2_X1 KeyArray_S13reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS20ser[6]), .B(KeyArray_outS23ser[6]), .Z(
        KeyArray_S13reg_gff_1_SFF_6_MUXInst_X) );
  AND2_X1 KeyArray_S13reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A1(KeyArray_n22), 
        .A2(KeyArray_S13reg_gff_1_SFF_6_MUXInst_X), .ZN(
        KeyArray_S13reg_gff_1_SFF_6_MUXInst_Y) );
  XOR2_X1 KeyArray_S13reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A(
        KeyArray_S13reg_gff_1_SFF_6_MUXInst_Y), .B(KeyArray_outS20ser[6]), .Z(
        KeyArray_S13reg_gff_1_SFF_6_QD) );
  INV_X1 KeyArray_S13reg_gff_1_SFF_6_Q_reg_U1 ( .A(keySBIn[6]), .ZN(
        KeyArray_S13reg_gff_1_SFF_6_n10) );
  DFF_X1 KeyArray_S13reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        KeyArray_S13reg_gff_1_SFF_6_n5), .CK(clk), .Q(keySBIn[6]), .QN() );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_7_U3 ( .A1(KeyArray_S13reg_gff_1_SFF_7_n2), .A2(KeyArray_S13reg_gff_1_SFF_7_n1), .ZN(KeyArray_S13reg_gff_1_SFF_7_n5) );
  OR2_X1 KeyArray_S13reg_gff_1_SFF_7_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S13reg_gff_1_SFF_7_n10), .ZN(KeyArray_S13reg_gff_1_SFF_7_n1)
         );
  NAND2_X1 KeyArray_S13reg_gff_1_SFF_7_U1 ( .A1(KeyArray_S13reg_gff_1_SFF_7_QD), .A2(KeyArray_n18), .ZN(KeyArray_S13reg_gff_1_SFF_7_n2) );
  XOR2_X1 KeyArray_S13reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS20ser[7]), .B(KeyArray_outS23ser[7]), .Z(
        KeyArray_S13reg_gff_1_SFF_7_MUXInst_X) );
  AND2_X1 KeyArray_S13reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A1(KeyArray_n22), 
        .A2(KeyArray_S13reg_gff_1_SFF_7_MUXInst_X), .ZN(
        KeyArray_S13reg_gff_1_SFF_7_MUXInst_Y) );
  XOR2_X1 KeyArray_S13reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A(
        KeyArray_S13reg_gff_1_SFF_7_MUXInst_Y), .B(KeyArray_outS20ser[7]), .Z(
        KeyArray_S13reg_gff_1_SFF_7_QD) );
  INV_X1 KeyArray_S13reg_gff_1_SFF_7_Q_reg_U1 ( .A(keySBIn[7]), .ZN(
        KeyArray_S13reg_gff_1_SFF_7_n10) );
  DFF_X1 KeyArray_S13reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        KeyArray_S13reg_gff_1_SFF_7_n5), .CK(clk), .Q(keySBIn[7]), .QN() );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_0_U3 ( .A1(KeyArray_S20reg_gff_1_SFF_0_n2), .A2(KeyArray_S20reg_gff_1_SFF_0_n1), .ZN(KeyArray_S20reg_gff_1_SFF_0_n5) );
  OR2_X1 KeyArray_S20reg_gff_1_SFF_0_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S20reg_gff_1_SFF_0_n10), .ZN(KeyArray_S20reg_gff_1_SFF_0_n1)
         );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_0_U1 ( .A1(KeyArray_S20reg_gff_1_SFF_0_QD), .A2(KeyArray_n18), .ZN(KeyArray_S20reg_gff_1_SFF_0_n2) );
  XOR2_X1 KeyArray_S20reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS21ser[0]), .B(KeyArray_outS30ser[0]), .Z(
        KeyArray_S20reg_gff_1_SFF_0_MUXInst_X) );
  AND2_X1 KeyArray_S20reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A1(KeyArray_n22), 
        .A2(KeyArray_S20reg_gff_1_SFF_0_MUXInst_X), .ZN(
        KeyArray_S20reg_gff_1_SFF_0_MUXInst_Y) );
  XOR2_X1 KeyArray_S20reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A(
        KeyArray_S20reg_gff_1_SFF_0_MUXInst_Y), .B(KeyArray_outS21ser[0]), .Z(
        KeyArray_S20reg_gff_1_SFF_0_QD) );
  INV_X1 KeyArray_S20reg_gff_1_SFF_0_Q_reg_U1 ( .A(KeyArray_outS20ser[0]), 
        .ZN(KeyArray_S20reg_gff_1_SFF_0_n10) );
  DFF_X1 KeyArray_S20reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        KeyArray_S20reg_gff_1_SFF_0_n5), .CK(clk), .Q(KeyArray_outS20ser[0]), 
        .QN() );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_1_U3 ( .A1(KeyArray_S20reg_gff_1_SFF_1_n2), .A2(KeyArray_S20reg_gff_1_SFF_1_n1), .ZN(KeyArray_S20reg_gff_1_SFF_1_n5) );
  OR2_X1 KeyArray_S20reg_gff_1_SFF_1_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S20reg_gff_1_SFF_1_n10), .ZN(KeyArray_S20reg_gff_1_SFF_1_n1)
         );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_1_U1 ( .A1(KeyArray_S20reg_gff_1_SFF_1_QD), .A2(KeyArray_n18), .ZN(KeyArray_S20reg_gff_1_SFF_1_n2) );
  XOR2_X1 KeyArray_S20reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS21ser[1]), .B(KeyArray_outS30ser[1]), .Z(
        KeyArray_S20reg_gff_1_SFF_1_MUXInst_X) );
  AND2_X1 KeyArray_S20reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A1(KeyArray_n22), 
        .A2(KeyArray_S20reg_gff_1_SFF_1_MUXInst_X), .ZN(
        KeyArray_S20reg_gff_1_SFF_1_MUXInst_Y) );
  XOR2_X1 KeyArray_S20reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A(
        KeyArray_S20reg_gff_1_SFF_1_MUXInst_Y), .B(KeyArray_outS21ser[1]), .Z(
        KeyArray_S20reg_gff_1_SFF_1_QD) );
  INV_X1 KeyArray_S20reg_gff_1_SFF_1_Q_reg_U1 ( .A(KeyArray_outS20ser[1]), 
        .ZN(KeyArray_S20reg_gff_1_SFF_1_n10) );
  DFF_X1 KeyArray_S20reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        KeyArray_S20reg_gff_1_SFF_1_n5), .CK(clk), .Q(KeyArray_outS20ser[1]), 
        .QN() );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_2_U3 ( .A1(KeyArray_S20reg_gff_1_SFF_2_n2), .A2(KeyArray_S20reg_gff_1_SFF_2_n1), .ZN(KeyArray_S20reg_gff_1_SFF_2_n5) );
  OR2_X1 KeyArray_S20reg_gff_1_SFF_2_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S20reg_gff_1_SFF_2_n10), .ZN(KeyArray_S20reg_gff_1_SFF_2_n1)
         );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_2_U1 ( .A1(KeyArray_S20reg_gff_1_SFF_2_QD), .A2(KeyArray_n18), .ZN(KeyArray_S20reg_gff_1_SFF_2_n2) );
  XOR2_X1 KeyArray_S20reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS21ser[2]), .B(KeyArray_outS30ser[2]), .Z(
        KeyArray_S20reg_gff_1_SFF_2_MUXInst_X) );
  AND2_X1 KeyArray_S20reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A1(KeyArray_n22), 
        .A2(KeyArray_S20reg_gff_1_SFF_2_MUXInst_X), .ZN(
        KeyArray_S20reg_gff_1_SFF_2_MUXInst_Y) );
  XOR2_X1 KeyArray_S20reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A(
        KeyArray_S20reg_gff_1_SFF_2_MUXInst_Y), .B(KeyArray_outS21ser[2]), .Z(
        KeyArray_S20reg_gff_1_SFF_2_QD) );
  INV_X1 KeyArray_S20reg_gff_1_SFF_2_Q_reg_U1 ( .A(KeyArray_outS20ser[2]), 
        .ZN(KeyArray_S20reg_gff_1_SFF_2_n10) );
  DFF_X1 KeyArray_S20reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        KeyArray_S20reg_gff_1_SFF_2_n5), .CK(clk), .Q(KeyArray_outS20ser[2]), 
        .QN() );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_3_U3 ( .A1(KeyArray_S20reg_gff_1_SFF_3_n2), .A2(KeyArray_S20reg_gff_1_SFF_3_n1), .ZN(KeyArray_S20reg_gff_1_SFF_3_n5) );
  OR2_X1 KeyArray_S20reg_gff_1_SFF_3_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S20reg_gff_1_SFF_3_n10), .ZN(KeyArray_S20reg_gff_1_SFF_3_n1)
         );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_3_U1 ( .A1(KeyArray_S20reg_gff_1_SFF_3_QD), .A2(KeyArray_n18), .ZN(KeyArray_S20reg_gff_1_SFF_3_n2) );
  XOR2_X1 KeyArray_S20reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS21ser[3]), .B(KeyArray_outS30ser[3]), .Z(
        KeyArray_S20reg_gff_1_SFF_3_MUXInst_X) );
  AND2_X1 KeyArray_S20reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A1(KeyArray_n22), 
        .A2(KeyArray_S20reg_gff_1_SFF_3_MUXInst_X), .ZN(
        KeyArray_S20reg_gff_1_SFF_3_MUXInst_Y) );
  XOR2_X1 KeyArray_S20reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A(
        KeyArray_S20reg_gff_1_SFF_3_MUXInst_Y), .B(KeyArray_outS21ser[3]), .Z(
        KeyArray_S20reg_gff_1_SFF_3_QD) );
  INV_X1 KeyArray_S20reg_gff_1_SFF_3_Q_reg_U1 ( .A(KeyArray_outS20ser[3]), 
        .ZN(KeyArray_S20reg_gff_1_SFF_3_n10) );
  DFF_X1 KeyArray_S20reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        KeyArray_S20reg_gff_1_SFF_3_n5), .CK(clk), .Q(KeyArray_outS20ser[3]), 
        .QN() );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_4_U3 ( .A1(KeyArray_S20reg_gff_1_SFF_4_n2), .A2(KeyArray_S20reg_gff_1_SFF_4_n1), .ZN(KeyArray_S20reg_gff_1_SFF_4_n5) );
  OR2_X1 KeyArray_S20reg_gff_1_SFF_4_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S20reg_gff_1_SFF_4_n10), .ZN(KeyArray_S20reg_gff_1_SFF_4_n1)
         );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_4_U1 ( .A1(KeyArray_S20reg_gff_1_SFF_4_QD), .A2(KeyArray_n18), .ZN(KeyArray_S20reg_gff_1_SFF_4_n2) );
  XOR2_X1 KeyArray_S20reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS21ser[4]), .B(KeyArray_outS30ser[4]), .Z(
        KeyArray_S20reg_gff_1_SFF_4_MUXInst_X) );
  AND2_X1 KeyArray_S20reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A1(KeyArray_n22), 
        .A2(KeyArray_S20reg_gff_1_SFF_4_MUXInst_X), .ZN(
        KeyArray_S20reg_gff_1_SFF_4_MUXInst_Y) );
  XOR2_X1 KeyArray_S20reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A(
        KeyArray_S20reg_gff_1_SFF_4_MUXInst_Y), .B(KeyArray_outS21ser[4]), .Z(
        KeyArray_S20reg_gff_1_SFF_4_QD) );
  INV_X1 KeyArray_S20reg_gff_1_SFF_4_Q_reg_U1 ( .A(KeyArray_outS20ser[4]), 
        .ZN(KeyArray_S20reg_gff_1_SFF_4_n10) );
  DFF_X1 KeyArray_S20reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        KeyArray_S20reg_gff_1_SFF_4_n5), .CK(clk), .Q(KeyArray_outS20ser[4]), 
        .QN() );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_5_U3 ( .A1(KeyArray_S20reg_gff_1_SFF_5_n2), .A2(KeyArray_S20reg_gff_1_SFF_5_n1), .ZN(KeyArray_S20reg_gff_1_SFF_5_n5) );
  OR2_X1 KeyArray_S20reg_gff_1_SFF_5_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S20reg_gff_1_SFF_5_n10), .ZN(KeyArray_S20reg_gff_1_SFF_5_n1)
         );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_5_U1 ( .A1(KeyArray_S20reg_gff_1_SFF_5_QD), .A2(KeyArray_n18), .ZN(KeyArray_S20reg_gff_1_SFF_5_n2) );
  XOR2_X1 KeyArray_S20reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS21ser[5]), .B(KeyArray_outS30ser[5]), .Z(
        KeyArray_S20reg_gff_1_SFF_5_MUXInst_X) );
  AND2_X1 KeyArray_S20reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A1(KeyArray_n22), 
        .A2(KeyArray_S20reg_gff_1_SFF_5_MUXInst_X), .ZN(
        KeyArray_S20reg_gff_1_SFF_5_MUXInst_Y) );
  XOR2_X1 KeyArray_S20reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A(
        KeyArray_S20reg_gff_1_SFF_5_MUXInst_Y), .B(KeyArray_outS21ser[5]), .Z(
        KeyArray_S20reg_gff_1_SFF_5_QD) );
  INV_X1 KeyArray_S20reg_gff_1_SFF_5_Q_reg_U1 ( .A(KeyArray_outS20ser[5]), 
        .ZN(KeyArray_S20reg_gff_1_SFF_5_n10) );
  DFF_X1 KeyArray_S20reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        KeyArray_S20reg_gff_1_SFF_5_n5), .CK(clk), .Q(KeyArray_outS20ser[5]), 
        .QN() );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_6_U3 ( .A1(KeyArray_S20reg_gff_1_SFF_6_n2), .A2(KeyArray_S20reg_gff_1_SFF_6_n1), .ZN(KeyArray_S20reg_gff_1_SFF_6_n5) );
  OR2_X1 KeyArray_S20reg_gff_1_SFF_6_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S20reg_gff_1_SFF_6_n10), .ZN(KeyArray_S20reg_gff_1_SFF_6_n1)
         );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_6_U1 ( .A1(KeyArray_S20reg_gff_1_SFF_6_QD), .A2(KeyArray_n18), .ZN(KeyArray_S20reg_gff_1_SFF_6_n2) );
  XOR2_X1 KeyArray_S20reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS21ser[6]), .B(KeyArray_outS30ser[6]), .Z(
        KeyArray_S20reg_gff_1_SFF_6_MUXInst_X) );
  AND2_X1 KeyArray_S20reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A1(KeyArray_n22), 
        .A2(KeyArray_S20reg_gff_1_SFF_6_MUXInst_X), .ZN(
        KeyArray_S20reg_gff_1_SFF_6_MUXInst_Y) );
  XOR2_X1 KeyArray_S20reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A(
        KeyArray_S20reg_gff_1_SFF_6_MUXInst_Y), .B(KeyArray_outS21ser[6]), .Z(
        KeyArray_S20reg_gff_1_SFF_6_QD) );
  INV_X1 KeyArray_S20reg_gff_1_SFF_6_Q_reg_U1 ( .A(KeyArray_outS20ser[6]), 
        .ZN(KeyArray_S20reg_gff_1_SFF_6_n10) );
  DFF_X1 KeyArray_S20reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        KeyArray_S20reg_gff_1_SFF_6_n5), .CK(clk), .Q(KeyArray_outS20ser[6]), 
        .QN() );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_7_U3 ( .A1(KeyArray_S20reg_gff_1_SFF_7_n2), .A2(KeyArray_S20reg_gff_1_SFF_7_n1), .ZN(KeyArray_S20reg_gff_1_SFF_7_n5) );
  OR2_X1 KeyArray_S20reg_gff_1_SFF_7_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S20reg_gff_1_SFF_7_n10), .ZN(KeyArray_S20reg_gff_1_SFF_7_n1)
         );
  NAND2_X1 KeyArray_S20reg_gff_1_SFF_7_U1 ( .A1(KeyArray_S20reg_gff_1_SFF_7_QD), .A2(KeyArray_n18), .ZN(KeyArray_S20reg_gff_1_SFF_7_n2) );
  XOR2_X1 KeyArray_S20reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS21ser[7]), .B(KeyArray_outS30ser[7]), .Z(
        KeyArray_S20reg_gff_1_SFF_7_MUXInst_X) );
  AND2_X1 KeyArray_S20reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A1(KeyArray_n22), 
        .A2(KeyArray_S20reg_gff_1_SFF_7_MUXInst_X), .ZN(
        KeyArray_S20reg_gff_1_SFF_7_MUXInst_Y) );
  XOR2_X1 KeyArray_S20reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A(
        KeyArray_S20reg_gff_1_SFF_7_MUXInst_Y), .B(KeyArray_outS21ser[7]), .Z(
        KeyArray_S20reg_gff_1_SFF_7_QD) );
  INV_X1 KeyArray_S20reg_gff_1_SFF_7_Q_reg_U1 ( .A(KeyArray_outS20ser[7]), 
        .ZN(KeyArray_S20reg_gff_1_SFF_7_n10) );
  DFF_X1 KeyArray_S20reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        KeyArray_S20reg_gff_1_SFF_7_n5), .CK(clk), .Q(KeyArray_outS20ser[7]), 
        .QN() );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_0_U3 ( .A1(KeyArray_S21reg_gff_1_SFF_0_n2), .A2(KeyArray_S21reg_gff_1_SFF_0_n1), .ZN(KeyArray_S21reg_gff_1_SFF_0_n6) );
  OR2_X1 KeyArray_S21reg_gff_1_SFF_0_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S21reg_gff_1_SFF_0_n11), .ZN(KeyArray_S21reg_gff_1_SFF_0_n1)
         );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_0_U1 ( .A1(KeyArray_S21reg_gff_1_SFF_0_QD), .A2(KeyArray_n18), .ZN(KeyArray_S21reg_gff_1_SFF_0_n2) );
  XOR2_X1 KeyArray_S21reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS22ser[0]), .B(KeyArray_outS31ser[0]), .Z(
        KeyArray_S21reg_gff_1_SFF_0_MUXInst_X) );
  AND2_X1 KeyArray_S21reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A1(KeyArray_n22), 
        .A2(KeyArray_S21reg_gff_1_SFF_0_MUXInst_X), .ZN(
        KeyArray_S21reg_gff_1_SFF_0_MUXInst_Y) );
  XOR2_X1 KeyArray_S21reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A(
        KeyArray_S21reg_gff_1_SFF_0_MUXInst_Y), .B(KeyArray_outS22ser[0]), .Z(
        KeyArray_S21reg_gff_1_SFF_0_QD) );
  INV_X1 KeyArray_S21reg_gff_1_SFF_0_Q_reg_U1 ( .A(KeyArray_outS21ser[0]), 
        .ZN(KeyArray_S21reg_gff_1_SFF_0_n11) );
  DFF_X1 KeyArray_S21reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        KeyArray_S21reg_gff_1_SFF_0_n6), .CK(clk), .Q(KeyArray_outS21ser[0]), 
        .QN() );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_1_U3 ( .A1(KeyArray_S21reg_gff_1_SFF_1_n2), .A2(KeyArray_S21reg_gff_1_SFF_1_n1), .ZN(KeyArray_S21reg_gff_1_SFF_1_n6) );
  OR2_X1 KeyArray_S21reg_gff_1_SFF_1_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S21reg_gff_1_SFF_1_n11), .ZN(KeyArray_S21reg_gff_1_SFF_1_n1)
         );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_1_U1 ( .A1(KeyArray_S21reg_gff_1_SFF_1_QD), .A2(KeyArray_n18), .ZN(KeyArray_S21reg_gff_1_SFF_1_n2) );
  XOR2_X1 KeyArray_S21reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS22ser[1]), .B(KeyArray_outS31ser[1]), .Z(
        KeyArray_S21reg_gff_1_SFF_1_MUXInst_X) );
  AND2_X1 KeyArray_S21reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A1(KeyArray_n22), 
        .A2(KeyArray_S21reg_gff_1_SFF_1_MUXInst_X), .ZN(
        KeyArray_S21reg_gff_1_SFF_1_MUXInst_Y) );
  XOR2_X1 KeyArray_S21reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A(
        KeyArray_S21reg_gff_1_SFF_1_MUXInst_Y), .B(KeyArray_outS22ser[1]), .Z(
        KeyArray_S21reg_gff_1_SFF_1_QD) );
  INV_X1 KeyArray_S21reg_gff_1_SFF_1_Q_reg_U1 ( .A(KeyArray_outS21ser[1]), 
        .ZN(KeyArray_S21reg_gff_1_SFF_1_n11) );
  DFF_X1 KeyArray_S21reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        KeyArray_S21reg_gff_1_SFF_1_n6), .CK(clk), .Q(KeyArray_outS21ser[1]), 
        .QN() );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_2_U3 ( .A1(KeyArray_S21reg_gff_1_SFF_2_n2), .A2(KeyArray_S21reg_gff_1_SFF_2_n1), .ZN(KeyArray_S21reg_gff_1_SFF_2_n6) );
  OR2_X1 KeyArray_S21reg_gff_1_SFF_2_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S21reg_gff_1_SFF_2_n11), .ZN(KeyArray_S21reg_gff_1_SFF_2_n1)
         );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_2_U1 ( .A1(KeyArray_S21reg_gff_1_SFF_2_QD), .A2(KeyArray_n18), .ZN(KeyArray_S21reg_gff_1_SFF_2_n2) );
  XOR2_X1 KeyArray_S21reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS22ser[2]), .B(KeyArray_outS31ser[2]), .Z(
        KeyArray_S21reg_gff_1_SFF_2_MUXInst_X) );
  AND2_X1 KeyArray_S21reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A1(KeyArray_n22), 
        .A2(KeyArray_S21reg_gff_1_SFF_2_MUXInst_X), .ZN(
        KeyArray_S21reg_gff_1_SFF_2_MUXInst_Y) );
  XOR2_X1 KeyArray_S21reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A(
        KeyArray_S21reg_gff_1_SFF_2_MUXInst_Y), .B(KeyArray_outS22ser[2]), .Z(
        KeyArray_S21reg_gff_1_SFF_2_QD) );
  INV_X1 KeyArray_S21reg_gff_1_SFF_2_Q_reg_U1 ( .A(KeyArray_outS21ser[2]), 
        .ZN(KeyArray_S21reg_gff_1_SFF_2_n11) );
  DFF_X1 KeyArray_S21reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        KeyArray_S21reg_gff_1_SFF_2_n6), .CK(clk), .Q(KeyArray_outS21ser[2]), 
        .QN() );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_3_U3 ( .A1(KeyArray_S21reg_gff_1_SFF_3_n2), .A2(KeyArray_S21reg_gff_1_SFF_3_n1), .ZN(KeyArray_S21reg_gff_1_SFF_3_n6) );
  OR2_X1 KeyArray_S21reg_gff_1_SFF_3_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S21reg_gff_1_SFF_3_n11), .ZN(KeyArray_S21reg_gff_1_SFF_3_n1)
         );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_3_U1 ( .A1(KeyArray_S21reg_gff_1_SFF_3_QD), .A2(KeyArray_n18), .ZN(KeyArray_S21reg_gff_1_SFF_3_n2) );
  XOR2_X1 KeyArray_S21reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS22ser[3]), .B(KeyArray_outS31ser[3]), .Z(
        KeyArray_S21reg_gff_1_SFF_3_MUXInst_X) );
  AND2_X1 KeyArray_S21reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A1(KeyArray_n22), 
        .A2(KeyArray_S21reg_gff_1_SFF_3_MUXInst_X), .ZN(
        KeyArray_S21reg_gff_1_SFF_3_MUXInst_Y) );
  XOR2_X1 KeyArray_S21reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A(
        KeyArray_S21reg_gff_1_SFF_3_MUXInst_Y), .B(KeyArray_outS22ser[3]), .Z(
        KeyArray_S21reg_gff_1_SFF_3_QD) );
  INV_X1 KeyArray_S21reg_gff_1_SFF_3_Q_reg_U1 ( .A(KeyArray_outS21ser[3]), 
        .ZN(KeyArray_S21reg_gff_1_SFF_3_n11) );
  DFF_X1 KeyArray_S21reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        KeyArray_S21reg_gff_1_SFF_3_n6), .CK(clk), .Q(KeyArray_outS21ser[3]), 
        .QN() );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_4_U3 ( .A1(KeyArray_S21reg_gff_1_SFF_4_n2), .A2(KeyArray_S21reg_gff_1_SFF_4_n1), .ZN(KeyArray_S21reg_gff_1_SFF_4_n6) );
  OR2_X1 KeyArray_S21reg_gff_1_SFF_4_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S21reg_gff_1_SFF_4_n11), .ZN(KeyArray_S21reg_gff_1_SFF_4_n1)
         );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_4_U1 ( .A1(KeyArray_S21reg_gff_1_SFF_4_QD), .A2(KeyArray_n18), .ZN(KeyArray_S21reg_gff_1_SFF_4_n2) );
  XOR2_X1 KeyArray_S21reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS22ser[4]), .B(KeyArray_outS31ser[4]), .Z(
        KeyArray_S21reg_gff_1_SFF_4_MUXInst_X) );
  AND2_X1 KeyArray_S21reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A1(KeyArray_n22), 
        .A2(KeyArray_S21reg_gff_1_SFF_4_MUXInst_X), .ZN(
        KeyArray_S21reg_gff_1_SFF_4_MUXInst_Y) );
  XOR2_X1 KeyArray_S21reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A(
        KeyArray_S21reg_gff_1_SFF_4_MUXInst_Y), .B(KeyArray_outS22ser[4]), .Z(
        KeyArray_S21reg_gff_1_SFF_4_QD) );
  INV_X1 KeyArray_S21reg_gff_1_SFF_4_Q_reg_U1 ( .A(KeyArray_outS21ser[4]), 
        .ZN(KeyArray_S21reg_gff_1_SFF_4_n11) );
  DFF_X1 KeyArray_S21reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        KeyArray_S21reg_gff_1_SFF_4_n6), .CK(clk), .Q(KeyArray_outS21ser[4]), 
        .QN() );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_5_U3 ( .A1(KeyArray_S21reg_gff_1_SFF_5_n2), .A2(KeyArray_S21reg_gff_1_SFF_5_n1), .ZN(KeyArray_S21reg_gff_1_SFF_5_n6) );
  OR2_X1 KeyArray_S21reg_gff_1_SFF_5_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S21reg_gff_1_SFF_5_n11), .ZN(KeyArray_S21reg_gff_1_SFF_5_n1)
         );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_5_U1 ( .A1(KeyArray_S21reg_gff_1_SFF_5_QD), .A2(KeyArray_n18), .ZN(KeyArray_S21reg_gff_1_SFF_5_n2) );
  XOR2_X1 KeyArray_S21reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS22ser[5]), .B(KeyArray_outS31ser[5]), .Z(
        KeyArray_S21reg_gff_1_SFF_5_MUXInst_X) );
  AND2_X1 KeyArray_S21reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A1(KeyArray_n22), 
        .A2(KeyArray_S21reg_gff_1_SFF_5_MUXInst_X), .ZN(
        KeyArray_S21reg_gff_1_SFF_5_MUXInst_Y) );
  XOR2_X1 KeyArray_S21reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A(
        KeyArray_S21reg_gff_1_SFF_5_MUXInst_Y), .B(KeyArray_outS22ser[5]), .Z(
        KeyArray_S21reg_gff_1_SFF_5_QD) );
  INV_X1 KeyArray_S21reg_gff_1_SFF_5_Q_reg_U1 ( .A(KeyArray_outS21ser[5]), 
        .ZN(KeyArray_S21reg_gff_1_SFF_5_n11) );
  DFF_X1 KeyArray_S21reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        KeyArray_S21reg_gff_1_SFF_5_n6), .CK(clk), .Q(KeyArray_outS21ser[5]), 
        .QN() );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_6_U3 ( .A1(KeyArray_S21reg_gff_1_SFF_6_n2), .A2(KeyArray_S21reg_gff_1_SFF_6_n1), .ZN(KeyArray_S21reg_gff_1_SFF_6_n6) );
  OR2_X1 KeyArray_S21reg_gff_1_SFF_6_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S21reg_gff_1_SFF_6_n11), .ZN(KeyArray_S21reg_gff_1_SFF_6_n1)
         );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_6_U1 ( .A1(KeyArray_S21reg_gff_1_SFF_6_QD), .A2(KeyArray_n18), .ZN(KeyArray_S21reg_gff_1_SFF_6_n2) );
  XOR2_X1 KeyArray_S21reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS22ser[6]), .B(KeyArray_outS31ser[6]), .Z(
        KeyArray_S21reg_gff_1_SFF_6_MUXInst_X) );
  AND2_X1 KeyArray_S21reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A1(KeyArray_n22), 
        .A2(KeyArray_S21reg_gff_1_SFF_6_MUXInst_X), .ZN(
        KeyArray_S21reg_gff_1_SFF_6_MUXInst_Y) );
  XOR2_X1 KeyArray_S21reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A(
        KeyArray_S21reg_gff_1_SFF_6_MUXInst_Y), .B(KeyArray_outS22ser[6]), .Z(
        KeyArray_S21reg_gff_1_SFF_6_QD) );
  INV_X1 KeyArray_S21reg_gff_1_SFF_6_Q_reg_U1 ( .A(KeyArray_outS21ser[6]), 
        .ZN(KeyArray_S21reg_gff_1_SFF_6_n11) );
  DFF_X1 KeyArray_S21reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        KeyArray_S21reg_gff_1_SFF_6_n6), .CK(clk), .Q(KeyArray_outS21ser[6]), 
        .QN() );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_7_U3 ( .A1(KeyArray_S21reg_gff_1_SFF_7_n2), .A2(KeyArray_S21reg_gff_1_SFF_7_n1), .ZN(KeyArray_S21reg_gff_1_SFF_7_n6) );
  OR2_X1 KeyArray_S21reg_gff_1_SFF_7_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S21reg_gff_1_SFF_7_n11), .ZN(KeyArray_S21reg_gff_1_SFF_7_n1)
         );
  NAND2_X1 KeyArray_S21reg_gff_1_SFF_7_U1 ( .A1(KeyArray_S21reg_gff_1_SFF_7_QD), .A2(KeyArray_n18), .ZN(KeyArray_S21reg_gff_1_SFF_7_n2) );
  XOR2_X1 KeyArray_S21reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS22ser[7]), .B(KeyArray_outS31ser[7]), .Z(
        KeyArray_S21reg_gff_1_SFF_7_MUXInst_X) );
  AND2_X1 KeyArray_S21reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A1(KeyArray_n22), 
        .A2(KeyArray_S21reg_gff_1_SFF_7_MUXInst_X), .ZN(
        KeyArray_S21reg_gff_1_SFF_7_MUXInst_Y) );
  XOR2_X1 KeyArray_S21reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A(
        KeyArray_S21reg_gff_1_SFF_7_MUXInst_Y), .B(KeyArray_outS22ser[7]), .Z(
        KeyArray_S21reg_gff_1_SFF_7_QD) );
  INV_X1 KeyArray_S21reg_gff_1_SFF_7_Q_reg_U1 ( .A(KeyArray_outS21ser[7]), 
        .ZN(KeyArray_S21reg_gff_1_SFF_7_n11) );
  DFF_X1 KeyArray_S21reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        KeyArray_S21reg_gff_1_SFF_7_n6), .CK(clk), .Q(KeyArray_outS21ser[7]), 
        .QN() );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_0_U3 ( .A1(KeyArray_S22reg_gff_1_SFF_0_n2), .A2(KeyArray_S22reg_gff_1_SFF_0_n1), .ZN(KeyArray_S22reg_gff_1_SFF_0_n6) );
  OR2_X1 KeyArray_S22reg_gff_1_SFF_0_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S22reg_gff_1_SFF_0_n11), .ZN(KeyArray_S22reg_gff_1_SFF_0_n1)
         );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_0_U1 ( .A1(KeyArray_S22reg_gff_1_SFF_0_QD), .A2(KeyArray_n18), .ZN(KeyArray_S22reg_gff_1_SFF_0_n2) );
  XOR2_X1 KeyArray_S22reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS23ser[0]), .B(KeyArray_outS32ser[0]), .Z(
        KeyArray_S22reg_gff_1_SFF_0_MUXInst_X) );
  AND2_X1 KeyArray_S22reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A1(KeyArray_n21), 
        .A2(KeyArray_S22reg_gff_1_SFF_0_MUXInst_X), .ZN(
        KeyArray_S22reg_gff_1_SFF_0_MUXInst_Y) );
  XOR2_X1 KeyArray_S22reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A(
        KeyArray_S22reg_gff_1_SFF_0_MUXInst_Y), .B(KeyArray_outS23ser[0]), .Z(
        KeyArray_S22reg_gff_1_SFF_0_QD) );
  INV_X1 KeyArray_S22reg_gff_1_SFF_0_Q_reg_U1 ( .A(KeyArray_outS22ser[0]), 
        .ZN(KeyArray_S22reg_gff_1_SFF_0_n11) );
  DFF_X1 KeyArray_S22reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        KeyArray_S22reg_gff_1_SFF_0_n6), .CK(clk), .Q(KeyArray_outS22ser[0]), 
        .QN() );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_1_U3 ( .A1(KeyArray_S22reg_gff_1_SFF_1_n2), .A2(KeyArray_S22reg_gff_1_SFF_1_n1), .ZN(KeyArray_S22reg_gff_1_SFF_1_n6) );
  OR2_X1 KeyArray_S22reg_gff_1_SFF_1_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S22reg_gff_1_SFF_1_n11), .ZN(KeyArray_S22reg_gff_1_SFF_1_n1)
         );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_1_U1 ( .A1(KeyArray_S22reg_gff_1_SFF_1_QD), .A2(KeyArray_n18), .ZN(KeyArray_S22reg_gff_1_SFF_1_n2) );
  XOR2_X1 KeyArray_S22reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS23ser[1]), .B(KeyArray_outS32ser[1]), .Z(
        KeyArray_S22reg_gff_1_SFF_1_MUXInst_X) );
  AND2_X1 KeyArray_S22reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A1(KeyArray_n21), 
        .A2(KeyArray_S22reg_gff_1_SFF_1_MUXInst_X), .ZN(
        KeyArray_S22reg_gff_1_SFF_1_MUXInst_Y) );
  XOR2_X1 KeyArray_S22reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A(
        KeyArray_S22reg_gff_1_SFF_1_MUXInst_Y), .B(KeyArray_outS23ser[1]), .Z(
        KeyArray_S22reg_gff_1_SFF_1_QD) );
  INV_X1 KeyArray_S22reg_gff_1_SFF_1_Q_reg_U1 ( .A(KeyArray_outS22ser[1]), 
        .ZN(KeyArray_S22reg_gff_1_SFF_1_n11) );
  DFF_X1 KeyArray_S22reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        KeyArray_S22reg_gff_1_SFF_1_n6), .CK(clk), .Q(KeyArray_outS22ser[1]), 
        .QN() );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_2_U3 ( .A1(KeyArray_S22reg_gff_1_SFF_2_n2), .A2(KeyArray_S22reg_gff_1_SFF_2_n1), .ZN(KeyArray_S22reg_gff_1_SFF_2_n6) );
  OR2_X1 KeyArray_S22reg_gff_1_SFF_2_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S22reg_gff_1_SFF_2_n11), .ZN(KeyArray_S22reg_gff_1_SFF_2_n1)
         );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_2_U1 ( .A1(KeyArray_S22reg_gff_1_SFF_2_QD), .A2(KeyArray_n18), .ZN(KeyArray_S22reg_gff_1_SFF_2_n2) );
  XOR2_X1 KeyArray_S22reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS23ser[2]), .B(KeyArray_outS32ser[2]), .Z(
        KeyArray_S22reg_gff_1_SFF_2_MUXInst_X) );
  AND2_X1 KeyArray_S22reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A1(KeyArray_n21), 
        .A2(KeyArray_S22reg_gff_1_SFF_2_MUXInst_X), .ZN(
        KeyArray_S22reg_gff_1_SFF_2_MUXInst_Y) );
  XOR2_X1 KeyArray_S22reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A(
        KeyArray_S22reg_gff_1_SFF_2_MUXInst_Y), .B(KeyArray_outS23ser[2]), .Z(
        KeyArray_S22reg_gff_1_SFF_2_QD) );
  INV_X1 KeyArray_S22reg_gff_1_SFF_2_Q_reg_U1 ( .A(KeyArray_outS22ser[2]), 
        .ZN(KeyArray_S22reg_gff_1_SFF_2_n11) );
  DFF_X1 KeyArray_S22reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        KeyArray_S22reg_gff_1_SFF_2_n6), .CK(clk), .Q(KeyArray_outS22ser[2]), 
        .QN() );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_3_U3 ( .A1(KeyArray_S22reg_gff_1_SFF_3_n2), .A2(KeyArray_S22reg_gff_1_SFF_3_n1), .ZN(KeyArray_S22reg_gff_1_SFF_3_n6) );
  OR2_X1 KeyArray_S22reg_gff_1_SFF_3_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S22reg_gff_1_SFF_3_n11), .ZN(KeyArray_S22reg_gff_1_SFF_3_n1)
         );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_3_U1 ( .A1(KeyArray_S22reg_gff_1_SFF_3_QD), .A2(KeyArray_n18), .ZN(KeyArray_S22reg_gff_1_SFF_3_n2) );
  XOR2_X1 KeyArray_S22reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS23ser[3]), .B(KeyArray_outS32ser[3]), .Z(
        KeyArray_S22reg_gff_1_SFF_3_MUXInst_X) );
  AND2_X1 KeyArray_S22reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A1(KeyArray_n21), 
        .A2(KeyArray_S22reg_gff_1_SFF_3_MUXInst_X), .ZN(
        KeyArray_S22reg_gff_1_SFF_3_MUXInst_Y) );
  XOR2_X1 KeyArray_S22reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A(
        KeyArray_S22reg_gff_1_SFF_3_MUXInst_Y), .B(KeyArray_outS23ser[3]), .Z(
        KeyArray_S22reg_gff_1_SFF_3_QD) );
  INV_X1 KeyArray_S22reg_gff_1_SFF_3_Q_reg_U1 ( .A(KeyArray_outS22ser[3]), 
        .ZN(KeyArray_S22reg_gff_1_SFF_3_n11) );
  DFF_X1 KeyArray_S22reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        KeyArray_S22reg_gff_1_SFF_3_n6), .CK(clk), .Q(KeyArray_outS22ser[3]), 
        .QN() );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_4_U3 ( .A1(KeyArray_S22reg_gff_1_SFF_4_n2), .A2(KeyArray_S22reg_gff_1_SFF_4_n1), .ZN(KeyArray_S22reg_gff_1_SFF_4_n6) );
  OR2_X1 KeyArray_S22reg_gff_1_SFF_4_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S22reg_gff_1_SFF_4_n11), .ZN(KeyArray_S22reg_gff_1_SFF_4_n1)
         );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_4_U1 ( .A1(KeyArray_S22reg_gff_1_SFF_4_QD), .A2(KeyArray_n18), .ZN(KeyArray_S22reg_gff_1_SFF_4_n2) );
  XOR2_X1 KeyArray_S22reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS23ser[4]), .B(KeyArray_outS32ser[4]), .Z(
        KeyArray_S22reg_gff_1_SFF_4_MUXInst_X) );
  AND2_X1 KeyArray_S22reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A1(KeyArray_n21), 
        .A2(KeyArray_S22reg_gff_1_SFF_4_MUXInst_X), .ZN(
        KeyArray_S22reg_gff_1_SFF_4_MUXInst_Y) );
  XOR2_X1 KeyArray_S22reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A(
        KeyArray_S22reg_gff_1_SFF_4_MUXInst_Y), .B(KeyArray_outS23ser[4]), .Z(
        KeyArray_S22reg_gff_1_SFF_4_QD) );
  INV_X1 KeyArray_S22reg_gff_1_SFF_4_Q_reg_U1 ( .A(KeyArray_outS22ser[4]), 
        .ZN(KeyArray_S22reg_gff_1_SFF_4_n11) );
  DFF_X1 KeyArray_S22reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        KeyArray_S22reg_gff_1_SFF_4_n6), .CK(clk), .Q(KeyArray_outS22ser[4]), 
        .QN() );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_5_U3 ( .A1(KeyArray_S22reg_gff_1_SFF_5_n2), .A2(KeyArray_S22reg_gff_1_SFF_5_n1), .ZN(KeyArray_S22reg_gff_1_SFF_5_n6) );
  OR2_X1 KeyArray_S22reg_gff_1_SFF_5_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S22reg_gff_1_SFF_5_n11), .ZN(KeyArray_S22reg_gff_1_SFF_5_n1)
         );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_5_U1 ( .A1(KeyArray_S22reg_gff_1_SFF_5_QD), .A2(KeyArray_n18), .ZN(KeyArray_S22reg_gff_1_SFF_5_n2) );
  XOR2_X1 KeyArray_S22reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS23ser[5]), .B(KeyArray_outS32ser[5]), .Z(
        KeyArray_S22reg_gff_1_SFF_5_MUXInst_X) );
  AND2_X1 KeyArray_S22reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A1(KeyArray_n21), 
        .A2(KeyArray_S22reg_gff_1_SFF_5_MUXInst_X), .ZN(
        KeyArray_S22reg_gff_1_SFF_5_MUXInst_Y) );
  XOR2_X1 KeyArray_S22reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A(
        KeyArray_S22reg_gff_1_SFF_5_MUXInst_Y), .B(KeyArray_outS23ser[5]), .Z(
        KeyArray_S22reg_gff_1_SFF_5_QD) );
  INV_X1 KeyArray_S22reg_gff_1_SFF_5_Q_reg_U1 ( .A(KeyArray_outS22ser[5]), 
        .ZN(KeyArray_S22reg_gff_1_SFF_5_n11) );
  DFF_X1 KeyArray_S22reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        KeyArray_S22reg_gff_1_SFF_5_n6), .CK(clk), .Q(KeyArray_outS22ser[5]), 
        .QN() );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_6_U3 ( .A1(KeyArray_S22reg_gff_1_SFF_6_n2), .A2(KeyArray_S22reg_gff_1_SFF_6_n1), .ZN(KeyArray_S22reg_gff_1_SFF_6_n6) );
  OR2_X1 KeyArray_S22reg_gff_1_SFF_6_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S22reg_gff_1_SFF_6_n11), .ZN(KeyArray_S22reg_gff_1_SFF_6_n1)
         );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_6_U1 ( .A1(KeyArray_S22reg_gff_1_SFF_6_QD), .A2(KeyArray_n18), .ZN(KeyArray_S22reg_gff_1_SFF_6_n2) );
  XOR2_X1 KeyArray_S22reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS23ser[6]), .B(KeyArray_outS32ser[6]), .Z(
        KeyArray_S22reg_gff_1_SFF_6_MUXInst_X) );
  AND2_X1 KeyArray_S22reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A1(KeyArray_n21), 
        .A2(KeyArray_S22reg_gff_1_SFF_6_MUXInst_X), .ZN(
        KeyArray_S22reg_gff_1_SFF_6_MUXInst_Y) );
  XOR2_X1 KeyArray_S22reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A(
        KeyArray_S22reg_gff_1_SFF_6_MUXInst_Y), .B(KeyArray_outS23ser[6]), .Z(
        KeyArray_S22reg_gff_1_SFF_6_QD) );
  INV_X1 KeyArray_S22reg_gff_1_SFF_6_Q_reg_U1 ( .A(KeyArray_outS22ser[6]), 
        .ZN(KeyArray_S22reg_gff_1_SFF_6_n11) );
  DFF_X1 KeyArray_S22reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        KeyArray_S22reg_gff_1_SFF_6_n6), .CK(clk), .Q(KeyArray_outS22ser[6]), 
        .QN() );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_7_U3 ( .A1(KeyArray_S22reg_gff_1_SFF_7_n2), .A2(KeyArray_S22reg_gff_1_SFF_7_n1), .ZN(KeyArray_S22reg_gff_1_SFF_7_n6) );
  OR2_X1 KeyArray_S22reg_gff_1_SFF_7_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S22reg_gff_1_SFF_7_n11), .ZN(KeyArray_S22reg_gff_1_SFF_7_n1)
         );
  NAND2_X1 KeyArray_S22reg_gff_1_SFF_7_U1 ( .A1(KeyArray_S22reg_gff_1_SFF_7_QD), .A2(KeyArray_n18), .ZN(KeyArray_S22reg_gff_1_SFF_7_n2) );
  XOR2_X1 KeyArray_S22reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS23ser[7]), .B(KeyArray_outS32ser[7]), .Z(
        KeyArray_S22reg_gff_1_SFF_7_MUXInst_X) );
  AND2_X1 KeyArray_S22reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A1(KeyArray_n21), 
        .A2(KeyArray_S22reg_gff_1_SFF_7_MUXInst_X), .ZN(
        KeyArray_S22reg_gff_1_SFF_7_MUXInst_Y) );
  XOR2_X1 KeyArray_S22reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A(
        KeyArray_S22reg_gff_1_SFF_7_MUXInst_Y), .B(KeyArray_outS23ser[7]), .Z(
        KeyArray_S22reg_gff_1_SFF_7_QD) );
  INV_X1 KeyArray_S22reg_gff_1_SFF_7_Q_reg_U1 ( .A(KeyArray_outS22ser[7]), 
        .ZN(KeyArray_S22reg_gff_1_SFF_7_n11) );
  DFF_X1 KeyArray_S22reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        KeyArray_S22reg_gff_1_SFF_7_n6), .CK(clk), .Q(KeyArray_outS22ser[7]), 
        .QN() );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_0_U3 ( .A1(KeyArray_S23reg_gff_1_SFF_0_n2), .A2(KeyArray_S23reg_gff_1_SFF_0_n1), .ZN(KeyArray_S23reg_gff_1_SFF_0_n6) );
  OR2_X1 KeyArray_S23reg_gff_1_SFF_0_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S23reg_gff_1_SFF_0_n11), .ZN(KeyArray_S23reg_gff_1_SFF_0_n1)
         );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_0_U1 ( .A1(KeyArray_S23reg_gff_1_SFF_0_QD), .A2(KeyArray_n18), .ZN(KeyArray_S23reg_gff_1_SFF_0_n2) );
  XOR2_X1 KeyArray_S23reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS30ser[0]), .B(KeyArray_outS33ser[0]), .Z(
        KeyArray_S23reg_gff_1_SFF_0_MUXInst_X) );
  AND2_X1 KeyArray_S23reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A1(KeyArray_n21), 
        .A2(KeyArray_S23reg_gff_1_SFF_0_MUXInst_X), .ZN(
        KeyArray_S23reg_gff_1_SFF_0_MUXInst_Y) );
  XOR2_X1 KeyArray_S23reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A(
        KeyArray_S23reg_gff_1_SFF_0_MUXInst_Y), .B(KeyArray_outS30ser[0]), .Z(
        KeyArray_S23reg_gff_1_SFF_0_QD) );
  INV_X1 KeyArray_S23reg_gff_1_SFF_0_Q_reg_U1 ( .A(KeyArray_outS23ser[0]), 
        .ZN(KeyArray_S23reg_gff_1_SFF_0_n11) );
  DFF_X1 KeyArray_S23reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        KeyArray_S23reg_gff_1_SFF_0_n6), .CK(clk), .Q(KeyArray_outS23ser[0]), 
        .QN() );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_1_U3 ( .A1(KeyArray_S23reg_gff_1_SFF_1_n2), .A2(KeyArray_S23reg_gff_1_SFF_1_n1), .ZN(KeyArray_S23reg_gff_1_SFF_1_n6) );
  OR2_X1 KeyArray_S23reg_gff_1_SFF_1_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S23reg_gff_1_SFF_1_n11), .ZN(KeyArray_S23reg_gff_1_SFF_1_n1)
         );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_1_U1 ( .A1(KeyArray_S23reg_gff_1_SFF_1_QD), .A2(KeyArray_n18), .ZN(KeyArray_S23reg_gff_1_SFF_1_n2) );
  XOR2_X1 KeyArray_S23reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS30ser[1]), .B(KeyArray_outS33ser[1]), .Z(
        KeyArray_S23reg_gff_1_SFF_1_MUXInst_X) );
  AND2_X1 KeyArray_S23reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A1(KeyArray_n21), 
        .A2(KeyArray_S23reg_gff_1_SFF_1_MUXInst_X), .ZN(
        KeyArray_S23reg_gff_1_SFF_1_MUXInst_Y) );
  XOR2_X1 KeyArray_S23reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A(
        KeyArray_S23reg_gff_1_SFF_1_MUXInst_Y), .B(KeyArray_outS30ser[1]), .Z(
        KeyArray_S23reg_gff_1_SFF_1_QD) );
  INV_X1 KeyArray_S23reg_gff_1_SFF_1_Q_reg_U1 ( .A(KeyArray_outS23ser[1]), 
        .ZN(KeyArray_S23reg_gff_1_SFF_1_n11) );
  DFF_X1 KeyArray_S23reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        KeyArray_S23reg_gff_1_SFF_1_n6), .CK(clk), .Q(KeyArray_outS23ser[1]), 
        .QN() );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_2_U3 ( .A1(KeyArray_S23reg_gff_1_SFF_2_n2), .A2(KeyArray_S23reg_gff_1_SFF_2_n1), .ZN(KeyArray_S23reg_gff_1_SFF_2_n6) );
  OR2_X1 KeyArray_S23reg_gff_1_SFF_2_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S23reg_gff_1_SFF_2_n11), .ZN(KeyArray_S23reg_gff_1_SFF_2_n1)
         );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_2_U1 ( .A1(KeyArray_S23reg_gff_1_SFF_2_QD), .A2(KeyArray_n18), .ZN(KeyArray_S23reg_gff_1_SFF_2_n2) );
  XOR2_X1 KeyArray_S23reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS30ser[2]), .B(KeyArray_outS33ser[2]), .Z(
        KeyArray_S23reg_gff_1_SFF_2_MUXInst_X) );
  AND2_X1 KeyArray_S23reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A1(KeyArray_n21), 
        .A2(KeyArray_S23reg_gff_1_SFF_2_MUXInst_X), .ZN(
        KeyArray_S23reg_gff_1_SFF_2_MUXInst_Y) );
  XOR2_X1 KeyArray_S23reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A(
        KeyArray_S23reg_gff_1_SFF_2_MUXInst_Y), .B(KeyArray_outS30ser[2]), .Z(
        KeyArray_S23reg_gff_1_SFF_2_QD) );
  INV_X1 KeyArray_S23reg_gff_1_SFF_2_Q_reg_U1 ( .A(KeyArray_outS23ser[2]), 
        .ZN(KeyArray_S23reg_gff_1_SFF_2_n11) );
  DFF_X1 KeyArray_S23reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        KeyArray_S23reg_gff_1_SFF_2_n6), .CK(clk), .Q(KeyArray_outS23ser[2]), 
        .QN() );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_3_U3 ( .A1(KeyArray_S23reg_gff_1_SFF_3_n2), .A2(KeyArray_S23reg_gff_1_SFF_3_n1), .ZN(KeyArray_S23reg_gff_1_SFF_3_n6) );
  OR2_X1 KeyArray_S23reg_gff_1_SFF_3_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S23reg_gff_1_SFF_3_n11), .ZN(KeyArray_S23reg_gff_1_SFF_3_n1)
         );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_3_U1 ( .A1(KeyArray_S23reg_gff_1_SFF_3_QD), .A2(KeyArray_n18), .ZN(KeyArray_S23reg_gff_1_SFF_3_n2) );
  XOR2_X1 KeyArray_S23reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS30ser[3]), .B(KeyArray_outS33ser[3]), .Z(
        KeyArray_S23reg_gff_1_SFF_3_MUXInst_X) );
  AND2_X1 KeyArray_S23reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A1(KeyArray_n21), 
        .A2(KeyArray_S23reg_gff_1_SFF_3_MUXInst_X), .ZN(
        KeyArray_S23reg_gff_1_SFF_3_MUXInst_Y) );
  XOR2_X1 KeyArray_S23reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A(
        KeyArray_S23reg_gff_1_SFF_3_MUXInst_Y), .B(KeyArray_outS30ser[3]), .Z(
        KeyArray_S23reg_gff_1_SFF_3_QD) );
  INV_X1 KeyArray_S23reg_gff_1_SFF_3_Q_reg_U1 ( .A(KeyArray_outS23ser[3]), 
        .ZN(KeyArray_S23reg_gff_1_SFF_3_n11) );
  DFF_X1 KeyArray_S23reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        KeyArray_S23reg_gff_1_SFF_3_n6), .CK(clk), .Q(KeyArray_outS23ser[3]), 
        .QN() );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_4_U3 ( .A1(KeyArray_S23reg_gff_1_SFF_4_n2), .A2(KeyArray_S23reg_gff_1_SFF_4_n1), .ZN(KeyArray_S23reg_gff_1_SFF_4_n6) );
  OR2_X1 KeyArray_S23reg_gff_1_SFF_4_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S23reg_gff_1_SFF_4_n11), .ZN(KeyArray_S23reg_gff_1_SFF_4_n1)
         );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_4_U1 ( .A1(KeyArray_S23reg_gff_1_SFF_4_QD), .A2(KeyArray_n18), .ZN(KeyArray_S23reg_gff_1_SFF_4_n2) );
  XOR2_X1 KeyArray_S23reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS30ser[4]), .B(KeyArray_outS33ser[4]), .Z(
        KeyArray_S23reg_gff_1_SFF_4_MUXInst_X) );
  AND2_X1 KeyArray_S23reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A1(KeyArray_n21), 
        .A2(KeyArray_S23reg_gff_1_SFF_4_MUXInst_X), .ZN(
        KeyArray_S23reg_gff_1_SFF_4_MUXInst_Y) );
  XOR2_X1 KeyArray_S23reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A(
        KeyArray_S23reg_gff_1_SFF_4_MUXInst_Y), .B(KeyArray_outS30ser[4]), .Z(
        KeyArray_S23reg_gff_1_SFF_4_QD) );
  INV_X1 KeyArray_S23reg_gff_1_SFF_4_Q_reg_U1 ( .A(KeyArray_outS23ser[4]), 
        .ZN(KeyArray_S23reg_gff_1_SFF_4_n11) );
  DFF_X1 KeyArray_S23reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        KeyArray_S23reg_gff_1_SFF_4_n6), .CK(clk), .Q(KeyArray_outS23ser[4]), 
        .QN() );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_5_U3 ( .A1(KeyArray_S23reg_gff_1_SFF_5_n2), .A2(KeyArray_S23reg_gff_1_SFF_5_n1), .ZN(KeyArray_S23reg_gff_1_SFF_5_n5) );
  OR2_X1 KeyArray_S23reg_gff_1_SFF_5_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S23reg_gff_1_SFF_5_n10), .ZN(KeyArray_S23reg_gff_1_SFF_5_n1)
         );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_5_U1 ( .A1(KeyArray_S23reg_gff_1_SFF_5_QD), .A2(KeyArray_n18), .ZN(KeyArray_S23reg_gff_1_SFF_5_n2) );
  XOR2_X1 KeyArray_S23reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS30ser[5]), .B(KeyArray_outS33ser[5]), .Z(
        KeyArray_S23reg_gff_1_SFF_5_MUXInst_X) );
  AND2_X1 KeyArray_S23reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A1(KeyArray_n21), 
        .A2(KeyArray_S23reg_gff_1_SFF_5_MUXInst_X), .ZN(
        KeyArray_S23reg_gff_1_SFF_5_MUXInst_Y) );
  XOR2_X1 KeyArray_S23reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A(
        KeyArray_S23reg_gff_1_SFF_5_MUXInst_Y), .B(KeyArray_outS30ser[5]), .Z(
        KeyArray_S23reg_gff_1_SFF_5_QD) );
  INV_X1 KeyArray_S23reg_gff_1_SFF_5_Q_reg_U1 ( .A(KeyArray_outS23ser[5]), 
        .ZN(KeyArray_S23reg_gff_1_SFF_5_n10) );
  DFF_X1 KeyArray_S23reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        KeyArray_S23reg_gff_1_SFF_5_n5), .CK(clk), .Q(KeyArray_outS23ser[5]), 
        .QN() );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_6_U3 ( .A1(KeyArray_S23reg_gff_1_SFF_6_n2), .A2(KeyArray_S23reg_gff_1_SFF_6_n1), .ZN(KeyArray_S23reg_gff_1_SFF_6_n5) );
  OR2_X1 KeyArray_S23reg_gff_1_SFF_6_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S23reg_gff_1_SFF_6_n10), .ZN(KeyArray_S23reg_gff_1_SFF_6_n1)
         );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_6_U1 ( .A1(KeyArray_S23reg_gff_1_SFF_6_QD), .A2(KeyArray_n18), .ZN(KeyArray_S23reg_gff_1_SFF_6_n2) );
  XOR2_X1 KeyArray_S23reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS30ser[6]), .B(KeyArray_outS33ser[6]), .Z(
        KeyArray_S23reg_gff_1_SFF_6_MUXInst_X) );
  AND2_X1 KeyArray_S23reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A1(KeyArray_n21), 
        .A2(KeyArray_S23reg_gff_1_SFF_6_MUXInst_X), .ZN(
        KeyArray_S23reg_gff_1_SFF_6_MUXInst_Y) );
  XOR2_X1 KeyArray_S23reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A(
        KeyArray_S23reg_gff_1_SFF_6_MUXInst_Y), .B(KeyArray_outS30ser[6]), .Z(
        KeyArray_S23reg_gff_1_SFF_6_QD) );
  INV_X1 KeyArray_S23reg_gff_1_SFF_6_Q_reg_U1 ( .A(KeyArray_outS23ser[6]), 
        .ZN(KeyArray_S23reg_gff_1_SFF_6_n10) );
  DFF_X1 KeyArray_S23reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        KeyArray_S23reg_gff_1_SFF_6_n5), .CK(clk), .Q(KeyArray_outS23ser[6]), 
        .QN() );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_7_U3 ( .A1(KeyArray_S23reg_gff_1_SFF_7_n2), .A2(KeyArray_S23reg_gff_1_SFF_7_n1), .ZN(KeyArray_S23reg_gff_1_SFF_7_n5) );
  OR2_X1 KeyArray_S23reg_gff_1_SFF_7_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S23reg_gff_1_SFF_7_n10), .ZN(KeyArray_S23reg_gff_1_SFF_7_n1)
         );
  NAND2_X1 KeyArray_S23reg_gff_1_SFF_7_U1 ( .A1(KeyArray_S23reg_gff_1_SFF_7_QD), .A2(KeyArray_n18), .ZN(KeyArray_S23reg_gff_1_SFF_7_n2) );
  XOR2_X1 KeyArray_S23reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS30ser[7]), .B(KeyArray_outS33ser[7]), .Z(
        KeyArray_S23reg_gff_1_SFF_7_MUXInst_X) );
  AND2_X1 KeyArray_S23reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A1(KeyArray_n21), 
        .A2(KeyArray_S23reg_gff_1_SFF_7_MUXInst_X), .ZN(
        KeyArray_S23reg_gff_1_SFF_7_MUXInst_Y) );
  XOR2_X1 KeyArray_S23reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A(
        KeyArray_S23reg_gff_1_SFF_7_MUXInst_Y), .B(KeyArray_outS30ser[7]), .Z(
        KeyArray_S23reg_gff_1_SFF_7_QD) );
  INV_X1 KeyArray_S23reg_gff_1_SFF_7_Q_reg_U1 ( .A(KeyArray_outS23ser[7]), 
        .ZN(KeyArray_S23reg_gff_1_SFF_7_n10) );
  DFF_X1 KeyArray_S23reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        KeyArray_S23reg_gff_1_SFF_7_n5), .CK(clk), .Q(KeyArray_outS23ser[7]), 
        .QN() );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_0_U3 ( .A1(KeyArray_S30reg_gff_1_SFF_0_n2), .A2(KeyArray_S30reg_gff_1_SFF_0_n1), .ZN(KeyArray_S30reg_gff_1_SFF_0_n5) );
  OR2_X1 KeyArray_S30reg_gff_1_SFF_0_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S30reg_gff_1_SFF_0_n10), .ZN(KeyArray_S30reg_gff_1_SFF_0_n1)
         );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_0_U1 ( .A1(KeyArray_S30reg_gff_1_SFF_0_QD), .A2(KeyArray_n18), .ZN(KeyArray_S30reg_gff_1_SFF_0_n2) );
  XOR2_X1 KeyArray_S30reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS31ser[0]), .B(KeyArray_inS30par[0]), .Z(
        KeyArray_S30reg_gff_1_SFF_0_MUXInst_X) );
  AND2_X1 KeyArray_S30reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A1(KeyArray_n21), 
        .A2(KeyArray_S30reg_gff_1_SFF_0_MUXInst_X), .ZN(
        KeyArray_S30reg_gff_1_SFF_0_MUXInst_Y) );
  XOR2_X1 KeyArray_S30reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A(
        KeyArray_S30reg_gff_1_SFF_0_MUXInst_Y), .B(KeyArray_outS31ser[0]), .Z(
        KeyArray_S30reg_gff_1_SFF_0_QD) );
  INV_X1 KeyArray_S30reg_gff_1_SFF_0_Q_reg_U1 ( .A(KeyArray_outS30ser[0]), 
        .ZN(KeyArray_S30reg_gff_1_SFF_0_n10) );
  DFF_X1 KeyArray_S30reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        KeyArray_S30reg_gff_1_SFF_0_n5), .CK(clk), .Q(KeyArray_outS30ser[0]), 
        .QN() );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_1_U3 ( .A1(KeyArray_S30reg_gff_1_SFF_1_n2), .A2(KeyArray_S30reg_gff_1_SFF_1_n1), .ZN(KeyArray_S30reg_gff_1_SFF_1_n5) );
  OR2_X1 KeyArray_S30reg_gff_1_SFF_1_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S30reg_gff_1_SFF_1_n10), .ZN(KeyArray_S30reg_gff_1_SFF_1_n1)
         );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_1_U1 ( .A1(KeyArray_S30reg_gff_1_SFF_1_QD), .A2(KeyArray_n18), .ZN(KeyArray_S30reg_gff_1_SFF_1_n2) );
  XOR2_X1 KeyArray_S30reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS31ser[1]), .B(KeyArray_inS30par[1]), .Z(
        KeyArray_S30reg_gff_1_SFF_1_MUXInst_X) );
  AND2_X1 KeyArray_S30reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A1(KeyArray_n21), 
        .A2(KeyArray_S30reg_gff_1_SFF_1_MUXInst_X), .ZN(
        KeyArray_S30reg_gff_1_SFF_1_MUXInst_Y) );
  XOR2_X1 KeyArray_S30reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A(
        KeyArray_S30reg_gff_1_SFF_1_MUXInst_Y), .B(KeyArray_outS31ser[1]), .Z(
        KeyArray_S30reg_gff_1_SFF_1_QD) );
  INV_X1 KeyArray_S30reg_gff_1_SFF_1_Q_reg_U1 ( .A(KeyArray_outS30ser[1]), 
        .ZN(KeyArray_S30reg_gff_1_SFF_1_n10) );
  DFF_X1 KeyArray_S30reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        KeyArray_S30reg_gff_1_SFF_1_n5), .CK(clk), .Q(KeyArray_outS30ser[1]), 
        .QN() );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_2_U3 ( .A1(KeyArray_S30reg_gff_1_SFF_2_n2), .A2(KeyArray_S30reg_gff_1_SFF_2_n1), .ZN(KeyArray_S30reg_gff_1_SFF_2_n5) );
  OR2_X1 KeyArray_S30reg_gff_1_SFF_2_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S30reg_gff_1_SFF_2_n10), .ZN(KeyArray_S30reg_gff_1_SFF_2_n1)
         );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_2_U1 ( .A1(KeyArray_S30reg_gff_1_SFF_2_QD), .A2(KeyArray_n18), .ZN(KeyArray_S30reg_gff_1_SFF_2_n2) );
  XOR2_X1 KeyArray_S30reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS31ser[2]), .B(KeyArray_inS30par[2]), .Z(
        KeyArray_S30reg_gff_1_SFF_2_MUXInst_X) );
  AND2_X1 KeyArray_S30reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A1(KeyArray_n21), 
        .A2(KeyArray_S30reg_gff_1_SFF_2_MUXInst_X), .ZN(
        KeyArray_S30reg_gff_1_SFF_2_MUXInst_Y) );
  XOR2_X1 KeyArray_S30reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A(
        KeyArray_S30reg_gff_1_SFF_2_MUXInst_Y), .B(KeyArray_outS31ser[2]), .Z(
        KeyArray_S30reg_gff_1_SFF_2_QD) );
  INV_X1 KeyArray_S30reg_gff_1_SFF_2_Q_reg_U1 ( .A(KeyArray_outS30ser[2]), 
        .ZN(KeyArray_S30reg_gff_1_SFF_2_n10) );
  DFF_X1 KeyArray_S30reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        KeyArray_S30reg_gff_1_SFF_2_n5), .CK(clk), .Q(KeyArray_outS30ser[2]), 
        .QN() );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_3_U3 ( .A1(KeyArray_S30reg_gff_1_SFF_3_n2), .A2(KeyArray_S30reg_gff_1_SFF_3_n1), .ZN(KeyArray_S30reg_gff_1_SFF_3_n5) );
  OR2_X1 KeyArray_S30reg_gff_1_SFF_3_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S30reg_gff_1_SFF_3_n10), .ZN(KeyArray_S30reg_gff_1_SFF_3_n1)
         );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_3_U1 ( .A1(KeyArray_S30reg_gff_1_SFF_3_QD), .A2(KeyArray_n18), .ZN(KeyArray_S30reg_gff_1_SFF_3_n2) );
  XOR2_X1 KeyArray_S30reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS31ser[3]), .B(KeyArray_inS30par[3]), .Z(
        KeyArray_S30reg_gff_1_SFF_3_MUXInst_X) );
  AND2_X1 KeyArray_S30reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A1(KeyArray_n21), 
        .A2(KeyArray_S30reg_gff_1_SFF_3_MUXInst_X), .ZN(
        KeyArray_S30reg_gff_1_SFF_3_MUXInst_Y) );
  XOR2_X1 KeyArray_S30reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A(
        KeyArray_S30reg_gff_1_SFF_3_MUXInst_Y), .B(KeyArray_outS31ser[3]), .Z(
        KeyArray_S30reg_gff_1_SFF_3_QD) );
  INV_X1 KeyArray_S30reg_gff_1_SFF_3_Q_reg_U1 ( .A(KeyArray_outS30ser[3]), 
        .ZN(KeyArray_S30reg_gff_1_SFF_3_n10) );
  DFF_X1 KeyArray_S30reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        KeyArray_S30reg_gff_1_SFF_3_n5), .CK(clk), .Q(KeyArray_outS30ser[3]), 
        .QN() );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_4_U3 ( .A1(KeyArray_S30reg_gff_1_SFF_4_n2), .A2(KeyArray_S30reg_gff_1_SFF_4_n1), .ZN(KeyArray_S30reg_gff_1_SFF_4_n5) );
  OR2_X1 KeyArray_S30reg_gff_1_SFF_4_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S30reg_gff_1_SFF_4_n10), .ZN(KeyArray_S30reg_gff_1_SFF_4_n1)
         );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_4_U1 ( .A1(KeyArray_S30reg_gff_1_SFF_4_QD), .A2(KeyArray_n18), .ZN(KeyArray_S30reg_gff_1_SFF_4_n2) );
  XOR2_X1 KeyArray_S30reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS31ser[4]), .B(KeyArray_inS30par[4]), .Z(
        KeyArray_S30reg_gff_1_SFF_4_MUXInst_X) );
  AND2_X1 KeyArray_S30reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A1(KeyArray_n21), 
        .A2(KeyArray_S30reg_gff_1_SFF_4_MUXInst_X), .ZN(
        KeyArray_S30reg_gff_1_SFF_4_MUXInst_Y) );
  XOR2_X1 KeyArray_S30reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A(
        KeyArray_S30reg_gff_1_SFF_4_MUXInst_Y), .B(KeyArray_outS31ser[4]), .Z(
        KeyArray_S30reg_gff_1_SFF_4_QD) );
  INV_X1 KeyArray_S30reg_gff_1_SFF_4_Q_reg_U1 ( .A(KeyArray_outS30ser[4]), 
        .ZN(KeyArray_S30reg_gff_1_SFF_4_n10) );
  DFF_X1 KeyArray_S30reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        KeyArray_S30reg_gff_1_SFF_4_n5), .CK(clk), .Q(KeyArray_outS30ser[4]), 
        .QN() );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_5_U3 ( .A1(KeyArray_S30reg_gff_1_SFF_5_n2), .A2(KeyArray_S30reg_gff_1_SFF_5_n1), .ZN(KeyArray_S30reg_gff_1_SFF_5_n5) );
  OR2_X1 KeyArray_S30reg_gff_1_SFF_5_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S30reg_gff_1_SFF_5_n10), .ZN(KeyArray_S30reg_gff_1_SFF_5_n1)
         );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_5_U1 ( .A1(KeyArray_S30reg_gff_1_SFF_5_QD), .A2(KeyArray_n18), .ZN(KeyArray_S30reg_gff_1_SFF_5_n2) );
  XOR2_X1 KeyArray_S30reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS31ser[5]), .B(KeyArray_inS30par[5]), .Z(
        KeyArray_S30reg_gff_1_SFF_5_MUXInst_X) );
  AND2_X1 KeyArray_S30reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A1(KeyArray_n21), 
        .A2(KeyArray_S30reg_gff_1_SFF_5_MUXInst_X), .ZN(
        KeyArray_S30reg_gff_1_SFF_5_MUXInst_Y) );
  XOR2_X1 KeyArray_S30reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A(
        KeyArray_S30reg_gff_1_SFF_5_MUXInst_Y), .B(KeyArray_outS31ser[5]), .Z(
        KeyArray_S30reg_gff_1_SFF_5_QD) );
  INV_X1 KeyArray_S30reg_gff_1_SFF_5_Q_reg_U1 ( .A(KeyArray_outS30ser[5]), 
        .ZN(KeyArray_S30reg_gff_1_SFF_5_n10) );
  DFF_X1 KeyArray_S30reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        KeyArray_S30reg_gff_1_SFF_5_n5), .CK(clk), .Q(KeyArray_outS30ser[5]), 
        .QN() );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_6_U3 ( .A1(KeyArray_S30reg_gff_1_SFF_6_n2), .A2(KeyArray_S30reg_gff_1_SFF_6_n1), .ZN(KeyArray_S30reg_gff_1_SFF_6_n5) );
  OR2_X1 KeyArray_S30reg_gff_1_SFF_6_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S30reg_gff_1_SFF_6_n10), .ZN(KeyArray_S30reg_gff_1_SFF_6_n1)
         );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_6_U1 ( .A1(KeyArray_S30reg_gff_1_SFF_6_QD), .A2(KeyArray_n18), .ZN(KeyArray_S30reg_gff_1_SFF_6_n2) );
  XOR2_X1 KeyArray_S30reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS31ser[6]), .B(KeyArray_inS30par[6]), .Z(
        KeyArray_S30reg_gff_1_SFF_6_MUXInst_X) );
  AND2_X1 KeyArray_S30reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A1(KeyArray_n21), 
        .A2(KeyArray_S30reg_gff_1_SFF_6_MUXInst_X), .ZN(
        KeyArray_S30reg_gff_1_SFF_6_MUXInst_Y) );
  XOR2_X1 KeyArray_S30reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A(
        KeyArray_S30reg_gff_1_SFF_6_MUXInst_Y), .B(KeyArray_outS31ser[6]), .Z(
        KeyArray_S30reg_gff_1_SFF_6_QD) );
  INV_X1 KeyArray_S30reg_gff_1_SFF_6_Q_reg_U1 ( .A(KeyArray_outS30ser[6]), 
        .ZN(KeyArray_S30reg_gff_1_SFF_6_n10) );
  DFF_X1 KeyArray_S30reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        KeyArray_S30reg_gff_1_SFF_6_n5), .CK(clk), .Q(KeyArray_outS30ser[6]), 
        .QN() );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_7_U3 ( .A1(KeyArray_S30reg_gff_1_SFF_7_n2), .A2(KeyArray_S30reg_gff_1_SFF_7_n1), .ZN(KeyArray_S30reg_gff_1_SFF_7_n5) );
  OR2_X1 KeyArray_S30reg_gff_1_SFF_7_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S30reg_gff_1_SFF_7_n10), .ZN(KeyArray_S30reg_gff_1_SFF_7_n1)
         );
  NAND2_X1 KeyArray_S30reg_gff_1_SFF_7_U1 ( .A1(KeyArray_S30reg_gff_1_SFF_7_QD), .A2(KeyArray_n18), .ZN(KeyArray_S30reg_gff_1_SFF_7_n2) );
  XOR2_X1 KeyArray_S30reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS31ser[7]), .B(KeyArray_inS30par[7]), .Z(
        KeyArray_S30reg_gff_1_SFF_7_MUXInst_X) );
  AND2_X1 KeyArray_S30reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A1(KeyArray_n21), 
        .A2(KeyArray_S30reg_gff_1_SFF_7_MUXInst_X), .ZN(
        KeyArray_S30reg_gff_1_SFF_7_MUXInst_Y) );
  XOR2_X1 KeyArray_S30reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A(
        KeyArray_S30reg_gff_1_SFF_7_MUXInst_Y), .B(KeyArray_outS31ser[7]), .Z(
        KeyArray_S30reg_gff_1_SFF_7_QD) );
  INV_X1 KeyArray_S30reg_gff_1_SFF_7_Q_reg_U1 ( .A(KeyArray_outS30ser[7]), 
        .ZN(KeyArray_S30reg_gff_1_SFF_7_n10) );
  DFF_X1 KeyArray_S30reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        KeyArray_S30reg_gff_1_SFF_7_n5), .CK(clk), .Q(KeyArray_outS30ser[7]), 
        .QN() );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_0_U3 ( .A1(KeyArray_S31reg_gff_1_SFF_0_n2), .A2(KeyArray_S31reg_gff_1_SFF_0_n1), .ZN(KeyArray_S31reg_gff_1_SFF_0_n6) );
  OR2_X1 KeyArray_S31reg_gff_1_SFF_0_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S31reg_gff_1_SFF_0_n11), .ZN(KeyArray_S31reg_gff_1_SFF_0_n1)
         );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_0_U1 ( .A1(KeyArray_S31reg_gff_1_SFF_0_QD), .A2(KeyArray_n18), .ZN(KeyArray_S31reg_gff_1_SFF_0_n2) );
  XOR2_X1 KeyArray_S31reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS32ser[0]), .B(KeyArray_outS01ser_0_), .Z(
        KeyArray_S31reg_gff_1_SFF_0_MUXInst_X) );
  AND2_X1 KeyArray_S31reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A1(KeyArray_n21), 
        .A2(KeyArray_S31reg_gff_1_SFF_0_MUXInst_X), .ZN(
        KeyArray_S31reg_gff_1_SFF_0_MUXInst_Y) );
  XOR2_X1 KeyArray_S31reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A(
        KeyArray_S31reg_gff_1_SFF_0_MUXInst_Y), .B(KeyArray_outS32ser[0]), .Z(
        KeyArray_S31reg_gff_1_SFF_0_QD) );
  INV_X1 KeyArray_S31reg_gff_1_SFF_0_Q_reg_U1 ( .A(KeyArray_outS31ser[0]), 
        .ZN(KeyArray_S31reg_gff_1_SFF_0_n11) );
  DFF_X1 KeyArray_S31reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        KeyArray_S31reg_gff_1_SFF_0_n6), .CK(clk), .Q(KeyArray_outS31ser[0]), 
        .QN() );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_1_U3 ( .A1(KeyArray_S31reg_gff_1_SFF_1_n2), .A2(KeyArray_S31reg_gff_1_SFF_1_n1), .ZN(KeyArray_S31reg_gff_1_SFF_1_n6) );
  OR2_X1 KeyArray_S31reg_gff_1_SFF_1_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S31reg_gff_1_SFF_1_n11), .ZN(KeyArray_S31reg_gff_1_SFF_1_n1)
         );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_1_U1 ( .A1(KeyArray_S31reg_gff_1_SFF_1_QD), .A2(KeyArray_n18), .ZN(KeyArray_S31reg_gff_1_SFF_1_n2) );
  XOR2_X1 KeyArray_S31reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS32ser[1]), .B(KeyArray_outS01ser_1_), .Z(
        KeyArray_S31reg_gff_1_SFF_1_MUXInst_X) );
  AND2_X1 KeyArray_S31reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A1(KeyArray_n21), 
        .A2(KeyArray_S31reg_gff_1_SFF_1_MUXInst_X), .ZN(
        KeyArray_S31reg_gff_1_SFF_1_MUXInst_Y) );
  XOR2_X1 KeyArray_S31reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A(
        KeyArray_S31reg_gff_1_SFF_1_MUXInst_Y), .B(KeyArray_outS32ser[1]), .Z(
        KeyArray_S31reg_gff_1_SFF_1_QD) );
  INV_X1 KeyArray_S31reg_gff_1_SFF_1_Q_reg_U1 ( .A(KeyArray_outS31ser[1]), 
        .ZN(KeyArray_S31reg_gff_1_SFF_1_n11) );
  DFF_X1 KeyArray_S31reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        KeyArray_S31reg_gff_1_SFF_1_n6), .CK(clk), .Q(KeyArray_outS31ser[1]), 
        .QN() );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_2_U3 ( .A1(KeyArray_S31reg_gff_1_SFF_2_n2), .A2(KeyArray_S31reg_gff_1_SFF_2_n1), .ZN(KeyArray_S31reg_gff_1_SFF_2_n6) );
  OR2_X1 KeyArray_S31reg_gff_1_SFF_2_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S31reg_gff_1_SFF_2_n11), .ZN(KeyArray_S31reg_gff_1_SFF_2_n1)
         );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_2_U1 ( .A1(KeyArray_S31reg_gff_1_SFF_2_QD), .A2(KeyArray_n18), .ZN(KeyArray_S31reg_gff_1_SFF_2_n2) );
  XOR2_X1 KeyArray_S31reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS32ser[2]), .B(KeyArray_outS01ser_2_), .Z(
        KeyArray_S31reg_gff_1_SFF_2_MUXInst_X) );
  AND2_X1 KeyArray_S31reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A1(KeyArray_n21), 
        .A2(KeyArray_S31reg_gff_1_SFF_2_MUXInst_X), .ZN(
        KeyArray_S31reg_gff_1_SFF_2_MUXInst_Y) );
  XOR2_X1 KeyArray_S31reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A(
        KeyArray_S31reg_gff_1_SFF_2_MUXInst_Y), .B(KeyArray_outS32ser[2]), .Z(
        KeyArray_S31reg_gff_1_SFF_2_QD) );
  INV_X1 KeyArray_S31reg_gff_1_SFF_2_Q_reg_U1 ( .A(KeyArray_outS31ser[2]), 
        .ZN(KeyArray_S31reg_gff_1_SFF_2_n11) );
  DFF_X1 KeyArray_S31reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        KeyArray_S31reg_gff_1_SFF_2_n6), .CK(clk), .Q(KeyArray_outS31ser[2]), 
        .QN() );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_3_U3 ( .A1(KeyArray_S31reg_gff_1_SFF_3_n2), .A2(KeyArray_S31reg_gff_1_SFF_3_n1), .ZN(KeyArray_S31reg_gff_1_SFF_3_n6) );
  OR2_X1 KeyArray_S31reg_gff_1_SFF_3_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S31reg_gff_1_SFF_3_n11), .ZN(KeyArray_S31reg_gff_1_SFF_3_n1)
         );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_3_U1 ( .A1(KeyArray_S31reg_gff_1_SFF_3_QD), .A2(KeyArray_n18), .ZN(KeyArray_S31reg_gff_1_SFF_3_n2) );
  XOR2_X1 KeyArray_S31reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS32ser[3]), .B(KeyArray_outS01ser_3_), .Z(
        KeyArray_S31reg_gff_1_SFF_3_MUXInst_X) );
  AND2_X1 KeyArray_S31reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A1(KeyArray_n21), 
        .A2(KeyArray_S31reg_gff_1_SFF_3_MUXInst_X), .ZN(
        KeyArray_S31reg_gff_1_SFF_3_MUXInst_Y) );
  XOR2_X1 KeyArray_S31reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A(
        KeyArray_S31reg_gff_1_SFF_3_MUXInst_Y), .B(KeyArray_outS32ser[3]), .Z(
        KeyArray_S31reg_gff_1_SFF_3_QD) );
  INV_X1 KeyArray_S31reg_gff_1_SFF_3_Q_reg_U1 ( .A(KeyArray_outS31ser[3]), 
        .ZN(KeyArray_S31reg_gff_1_SFF_3_n11) );
  DFF_X1 KeyArray_S31reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        KeyArray_S31reg_gff_1_SFF_3_n6), .CK(clk), .Q(KeyArray_outS31ser[3]), 
        .QN() );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_4_U3 ( .A1(KeyArray_S31reg_gff_1_SFF_4_n2), .A2(KeyArray_S31reg_gff_1_SFF_4_n1), .ZN(KeyArray_S31reg_gff_1_SFF_4_n6) );
  OR2_X1 KeyArray_S31reg_gff_1_SFF_4_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S31reg_gff_1_SFF_4_n11), .ZN(KeyArray_S31reg_gff_1_SFF_4_n1)
         );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_4_U1 ( .A1(KeyArray_S31reg_gff_1_SFF_4_QD), .A2(KeyArray_n18), .ZN(KeyArray_S31reg_gff_1_SFF_4_n2) );
  XOR2_X1 KeyArray_S31reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS32ser[4]), .B(KeyArray_outS01ser_4_), .Z(
        KeyArray_S31reg_gff_1_SFF_4_MUXInst_X) );
  AND2_X1 KeyArray_S31reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A1(KeyArray_n21), 
        .A2(KeyArray_S31reg_gff_1_SFF_4_MUXInst_X), .ZN(
        KeyArray_S31reg_gff_1_SFF_4_MUXInst_Y) );
  XOR2_X1 KeyArray_S31reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A(
        KeyArray_S31reg_gff_1_SFF_4_MUXInst_Y), .B(KeyArray_outS32ser[4]), .Z(
        KeyArray_S31reg_gff_1_SFF_4_QD) );
  INV_X1 KeyArray_S31reg_gff_1_SFF_4_Q_reg_U1 ( .A(KeyArray_outS31ser[4]), 
        .ZN(KeyArray_S31reg_gff_1_SFF_4_n11) );
  DFF_X1 KeyArray_S31reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        KeyArray_S31reg_gff_1_SFF_4_n6), .CK(clk), .Q(KeyArray_outS31ser[4]), 
        .QN() );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_5_U3 ( .A1(KeyArray_S31reg_gff_1_SFF_5_n2), .A2(KeyArray_S31reg_gff_1_SFF_5_n1), .ZN(KeyArray_S31reg_gff_1_SFF_5_n6) );
  OR2_X1 KeyArray_S31reg_gff_1_SFF_5_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S31reg_gff_1_SFF_5_n11), .ZN(KeyArray_S31reg_gff_1_SFF_5_n1)
         );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_5_U1 ( .A1(KeyArray_S31reg_gff_1_SFF_5_QD), .A2(KeyArray_n18), .ZN(KeyArray_S31reg_gff_1_SFF_5_n2) );
  XOR2_X1 KeyArray_S31reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS32ser[5]), .B(KeyArray_outS01ser_5_), .Z(
        KeyArray_S31reg_gff_1_SFF_5_MUXInst_X) );
  AND2_X1 KeyArray_S31reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A1(KeyArray_n21), 
        .A2(KeyArray_S31reg_gff_1_SFF_5_MUXInst_X), .ZN(
        KeyArray_S31reg_gff_1_SFF_5_MUXInst_Y) );
  XOR2_X1 KeyArray_S31reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A(
        KeyArray_S31reg_gff_1_SFF_5_MUXInst_Y), .B(KeyArray_outS32ser[5]), .Z(
        KeyArray_S31reg_gff_1_SFF_5_QD) );
  INV_X1 KeyArray_S31reg_gff_1_SFF_5_Q_reg_U1 ( .A(KeyArray_outS31ser[5]), 
        .ZN(KeyArray_S31reg_gff_1_SFF_5_n11) );
  DFF_X1 KeyArray_S31reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        KeyArray_S31reg_gff_1_SFF_5_n6), .CK(clk), .Q(KeyArray_outS31ser[5]), 
        .QN() );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_6_U3 ( .A1(KeyArray_S31reg_gff_1_SFF_6_n2), .A2(KeyArray_S31reg_gff_1_SFF_6_n1), .ZN(KeyArray_S31reg_gff_1_SFF_6_n6) );
  OR2_X1 KeyArray_S31reg_gff_1_SFF_6_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S31reg_gff_1_SFF_6_n11), .ZN(KeyArray_S31reg_gff_1_SFF_6_n1)
         );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_6_U1 ( .A1(KeyArray_S31reg_gff_1_SFF_6_QD), .A2(KeyArray_n18), .ZN(KeyArray_S31reg_gff_1_SFF_6_n2) );
  XOR2_X1 KeyArray_S31reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS32ser[6]), .B(KeyArray_outS01ser_6_), .Z(
        KeyArray_S31reg_gff_1_SFF_6_MUXInst_X) );
  AND2_X1 KeyArray_S31reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A1(KeyArray_n21), 
        .A2(KeyArray_S31reg_gff_1_SFF_6_MUXInst_X), .ZN(
        KeyArray_S31reg_gff_1_SFF_6_MUXInst_Y) );
  XOR2_X1 KeyArray_S31reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A(
        KeyArray_S31reg_gff_1_SFF_6_MUXInst_Y), .B(KeyArray_outS32ser[6]), .Z(
        KeyArray_S31reg_gff_1_SFF_6_QD) );
  INV_X1 KeyArray_S31reg_gff_1_SFF_6_Q_reg_U1 ( .A(KeyArray_outS31ser[6]), 
        .ZN(KeyArray_S31reg_gff_1_SFF_6_n11) );
  DFF_X1 KeyArray_S31reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        KeyArray_S31reg_gff_1_SFF_6_n6), .CK(clk), .Q(KeyArray_outS31ser[6]), 
        .QN() );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_7_U3 ( .A1(KeyArray_S31reg_gff_1_SFF_7_n2), .A2(KeyArray_S31reg_gff_1_SFF_7_n1), .ZN(KeyArray_S31reg_gff_1_SFF_7_n6) );
  OR2_X1 KeyArray_S31reg_gff_1_SFF_7_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S31reg_gff_1_SFF_7_n11), .ZN(KeyArray_S31reg_gff_1_SFF_7_n1)
         );
  NAND2_X1 KeyArray_S31reg_gff_1_SFF_7_U1 ( .A1(KeyArray_S31reg_gff_1_SFF_7_QD), .A2(KeyArray_n18), .ZN(KeyArray_S31reg_gff_1_SFF_7_n2) );
  XOR2_X1 KeyArray_S31reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS32ser[7]), .B(KeyArray_outS01ser_7_), .Z(
        KeyArray_S31reg_gff_1_SFF_7_MUXInst_X) );
  AND2_X1 KeyArray_S31reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A1(KeyArray_n21), 
        .A2(KeyArray_S31reg_gff_1_SFF_7_MUXInst_X), .ZN(
        KeyArray_S31reg_gff_1_SFF_7_MUXInst_Y) );
  XOR2_X1 KeyArray_S31reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A(
        KeyArray_S31reg_gff_1_SFF_7_MUXInst_Y), .B(KeyArray_outS32ser[7]), .Z(
        KeyArray_S31reg_gff_1_SFF_7_QD) );
  INV_X1 KeyArray_S31reg_gff_1_SFF_7_Q_reg_U1 ( .A(KeyArray_outS31ser[7]), 
        .ZN(KeyArray_S31reg_gff_1_SFF_7_n11) );
  DFF_X1 KeyArray_S31reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        KeyArray_S31reg_gff_1_SFF_7_n6), .CK(clk), .Q(KeyArray_outS31ser[7]), 
        .QN() );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_0_U3 ( .A1(KeyArray_S32reg_gff_1_SFF_0_n2), .A2(KeyArray_S32reg_gff_1_SFF_0_n1), .ZN(KeyArray_S32reg_gff_1_SFF_0_n6) );
  OR2_X1 KeyArray_S32reg_gff_1_SFF_0_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S32reg_gff_1_SFF_0_n11), .ZN(KeyArray_S32reg_gff_1_SFF_0_n1)
         );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_0_U1 ( .A1(KeyArray_S32reg_gff_1_SFF_0_QD), .A2(KeyArray_n18), .ZN(KeyArray_S32reg_gff_1_SFF_0_n2) );
  XOR2_X1 KeyArray_S32reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS33ser[0]), .B(KeyArray_outS02ser[0]), .Z(
        KeyArray_S32reg_gff_1_SFF_0_MUXInst_X) );
  AND2_X1 KeyArray_S32reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A1(KeyArray_n21), 
        .A2(KeyArray_S32reg_gff_1_SFF_0_MUXInst_X), .ZN(
        KeyArray_S32reg_gff_1_SFF_0_MUXInst_Y) );
  XOR2_X1 KeyArray_S32reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A(
        KeyArray_S32reg_gff_1_SFF_0_MUXInst_Y), .B(KeyArray_outS33ser[0]), .Z(
        KeyArray_S32reg_gff_1_SFF_0_QD) );
  INV_X1 KeyArray_S32reg_gff_1_SFF_0_Q_reg_U1 ( .A(KeyArray_outS32ser[0]), 
        .ZN(KeyArray_S32reg_gff_1_SFF_0_n11) );
  DFF_X1 KeyArray_S32reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        KeyArray_S32reg_gff_1_SFF_0_n6), .CK(clk), .Q(KeyArray_outS32ser[0]), 
        .QN() );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_1_U3 ( .A1(KeyArray_S32reg_gff_1_SFF_1_n2), .A2(KeyArray_S32reg_gff_1_SFF_1_n1), .ZN(KeyArray_S32reg_gff_1_SFF_1_n6) );
  OR2_X1 KeyArray_S32reg_gff_1_SFF_1_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S32reg_gff_1_SFF_1_n11), .ZN(KeyArray_S32reg_gff_1_SFF_1_n1)
         );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_1_U1 ( .A1(KeyArray_S32reg_gff_1_SFF_1_QD), .A2(KeyArray_n18), .ZN(KeyArray_S32reg_gff_1_SFF_1_n2) );
  XOR2_X1 KeyArray_S32reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS33ser[1]), .B(KeyArray_outS02ser[1]), .Z(
        KeyArray_S32reg_gff_1_SFF_1_MUXInst_X) );
  AND2_X1 KeyArray_S32reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A1(KeyArray_n21), 
        .A2(KeyArray_S32reg_gff_1_SFF_1_MUXInst_X), .ZN(
        KeyArray_S32reg_gff_1_SFF_1_MUXInst_Y) );
  XOR2_X1 KeyArray_S32reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A(
        KeyArray_S32reg_gff_1_SFF_1_MUXInst_Y), .B(KeyArray_outS33ser[1]), .Z(
        KeyArray_S32reg_gff_1_SFF_1_QD) );
  INV_X1 KeyArray_S32reg_gff_1_SFF_1_Q_reg_U1 ( .A(KeyArray_outS32ser[1]), 
        .ZN(KeyArray_S32reg_gff_1_SFF_1_n11) );
  DFF_X1 KeyArray_S32reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        KeyArray_S32reg_gff_1_SFF_1_n6), .CK(clk), .Q(KeyArray_outS32ser[1]), 
        .QN() );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_2_U3 ( .A1(KeyArray_S32reg_gff_1_SFF_2_n2), .A2(KeyArray_S32reg_gff_1_SFF_2_n1), .ZN(KeyArray_S32reg_gff_1_SFF_2_n6) );
  OR2_X1 KeyArray_S32reg_gff_1_SFF_2_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S32reg_gff_1_SFF_2_n11), .ZN(KeyArray_S32reg_gff_1_SFF_2_n1)
         );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_2_U1 ( .A1(KeyArray_S32reg_gff_1_SFF_2_QD), .A2(KeyArray_n18), .ZN(KeyArray_S32reg_gff_1_SFF_2_n2) );
  XOR2_X1 KeyArray_S32reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS33ser[2]), .B(KeyArray_outS02ser[2]), .Z(
        KeyArray_S32reg_gff_1_SFF_2_MUXInst_X) );
  AND2_X1 KeyArray_S32reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A1(KeyArray_n21), 
        .A2(KeyArray_S32reg_gff_1_SFF_2_MUXInst_X), .ZN(
        KeyArray_S32reg_gff_1_SFF_2_MUXInst_Y) );
  XOR2_X1 KeyArray_S32reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A(
        KeyArray_S32reg_gff_1_SFF_2_MUXInst_Y), .B(KeyArray_outS33ser[2]), .Z(
        KeyArray_S32reg_gff_1_SFF_2_QD) );
  INV_X1 KeyArray_S32reg_gff_1_SFF_2_Q_reg_U1 ( .A(KeyArray_outS32ser[2]), 
        .ZN(KeyArray_S32reg_gff_1_SFF_2_n11) );
  DFF_X1 KeyArray_S32reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        KeyArray_S32reg_gff_1_SFF_2_n6), .CK(clk), .Q(KeyArray_outS32ser[2]), 
        .QN() );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_3_U3 ( .A1(KeyArray_S32reg_gff_1_SFF_3_n2), .A2(KeyArray_S32reg_gff_1_SFF_3_n1), .ZN(KeyArray_S32reg_gff_1_SFF_3_n6) );
  OR2_X1 KeyArray_S32reg_gff_1_SFF_3_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S32reg_gff_1_SFF_3_n11), .ZN(KeyArray_S32reg_gff_1_SFF_3_n1)
         );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_3_U1 ( .A1(KeyArray_S32reg_gff_1_SFF_3_QD), .A2(KeyArray_n18), .ZN(KeyArray_S32reg_gff_1_SFF_3_n2) );
  XOR2_X1 KeyArray_S32reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS33ser[3]), .B(KeyArray_outS02ser[3]), .Z(
        KeyArray_S32reg_gff_1_SFF_3_MUXInst_X) );
  AND2_X1 KeyArray_S32reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A1(KeyArray_n21), 
        .A2(KeyArray_S32reg_gff_1_SFF_3_MUXInst_X), .ZN(
        KeyArray_S32reg_gff_1_SFF_3_MUXInst_Y) );
  XOR2_X1 KeyArray_S32reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A(
        KeyArray_S32reg_gff_1_SFF_3_MUXInst_Y), .B(KeyArray_outS33ser[3]), .Z(
        KeyArray_S32reg_gff_1_SFF_3_QD) );
  INV_X1 KeyArray_S32reg_gff_1_SFF_3_Q_reg_U1 ( .A(KeyArray_outS32ser[3]), 
        .ZN(KeyArray_S32reg_gff_1_SFF_3_n11) );
  DFF_X1 KeyArray_S32reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        KeyArray_S32reg_gff_1_SFF_3_n6), .CK(clk), .Q(KeyArray_outS32ser[3]), 
        .QN() );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_4_U3 ( .A1(KeyArray_S32reg_gff_1_SFF_4_n2), .A2(KeyArray_S32reg_gff_1_SFF_4_n1), .ZN(KeyArray_S32reg_gff_1_SFF_4_n6) );
  OR2_X1 KeyArray_S32reg_gff_1_SFF_4_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S32reg_gff_1_SFF_4_n11), .ZN(KeyArray_S32reg_gff_1_SFF_4_n1)
         );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_4_U1 ( .A1(KeyArray_S32reg_gff_1_SFF_4_QD), .A2(KeyArray_n18), .ZN(KeyArray_S32reg_gff_1_SFF_4_n2) );
  XOR2_X1 KeyArray_S32reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS33ser[4]), .B(KeyArray_outS02ser[4]), .Z(
        KeyArray_S32reg_gff_1_SFF_4_MUXInst_X) );
  AND2_X1 KeyArray_S32reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A1(KeyArray_n21), 
        .A2(KeyArray_S32reg_gff_1_SFF_4_MUXInst_X), .ZN(
        KeyArray_S32reg_gff_1_SFF_4_MUXInst_Y) );
  XOR2_X1 KeyArray_S32reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A(
        KeyArray_S32reg_gff_1_SFF_4_MUXInst_Y), .B(KeyArray_outS33ser[4]), .Z(
        KeyArray_S32reg_gff_1_SFF_4_QD) );
  INV_X1 KeyArray_S32reg_gff_1_SFF_4_Q_reg_U1 ( .A(KeyArray_outS32ser[4]), 
        .ZN(KeyArray_S32reg_gff_1_SFF_4_n11) );
  DFF_X1 KeyArray_S32reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        KeyArray_S32reg_gff_1_SFF_4_n6), .CK(clk), .Q(KeyArray_outS32ser[4]), 
        .QN() );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_5_U3 ( .A1(KeyArray_S32reg_gff_1_SFF_5_n2), .A2(KeyArray_S32reg_gff_1_SFF_5_n1), .ZN(KeyArray_S32reg_gff_1_SFF_5_n5) );
  OR2_X1 KeyArray_S32reg_gff_1_SFF_5_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S32reg_gff_1_SFF_5_n10), .ZN(KeyArray_S32reg_gff_1_SFF_5_n1)
         );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_5_U1 ( .A1(KeyArray_S32reg_gff_1_SFF_5_QD), .A2(KeyArray_n18), .ZN(KeyArray_S32reg_gff_1_SFF_5_n2) );
  XOR2_X1 KeyArray_S32reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS33ser[5]), .B(KeyArray_outS02ser[5]), .Z(
        KeyArray_S32reg_gff_1_SFF_5_MUXInst_X) );
  AND2_X1 KeyArray_S32reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A1(KeyArray_n21), 
        .A2(KeyArray_S32reg_gff_1_SFF_5_MUXInst_X), .ZN(
        KeyArray_S32reg_gff_1_SFF_5_MUXInst_Y) );
  XOR2_X1 KeyArray_S32reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A(
        KeyArray_S32reg_gff_1_SFF_5_MUXInst_Y), .B(KeyArray_outS33ser[5]), .Z(
        KeyArray_S32reg_gff_1_SFF_5_QD) );
  INV_X1 KeyArray_S32reg_gff_1_SFF_5_Q_reg_U1 ( .A(KeyArray_outS32ser[5]), 
        .ZN(KeyArray_S32reg_gff_1_SFF_5_n10) );
  DFF_X1 KeyArray_S32reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        KeyArray_S32reg_gff_1_SFF_5_n5), .CK(clk), .Q(KeyArray_outS32ser[5]), 
        .QN() );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_6_U3 ( .A1(KeyArray_S32reg_gff_1_SFF_6_n2), .A2(KeyArray_S32reg_gff_1_SFF_6_n1), .ZN(KeyArray_S32reg_gff_1_SFF_6_n5) );
  OR2_X1 KeyArray_S32reg_gff_1_SFF_6_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S32reg_gff_1_SFF_6_n10), .ZN(KeyArray_S32reg_gff_1_SFF_6_n1)
         );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_6_U1 ( .A1(KeyArray_S32reg_gff_1_SFF_6_QD), .A2(KeyArray_n18), .ZN(KeyArray_S32reg_gff_1_SFF_6_n2) );
  XOR2_X1 KeyArray_S32reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS33ser[6]), .B(KeyArray_outS02ser[6]), .Z(
        KeyArray_S32reg_gff_1_SFF_6_MUXInst_X) );
  AND2_X1 KeyArray_S32reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A1(KeyArray_n21), 
        .A2(KeyArray_S32reg_gff_1_SFF_6_MUXInst_X), .ZN(
        KeyArray_S32reg_gff_1_SFF_6_MUXInst_Y) );
  XOR2_X1 KeyArray_S32reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A(
        KeyArray_S32reg_gff_1_SFF_6_MUXInst_Y), .B(KeyArray_outS33ser[6]), .Z(
        KeyArray_S32reg_gff_1_SFF_6_QD) );
  INV_X1 KeyArray_S32reg_gff_1_SFF_6_Q_reg_U1 ( .A(KeyArray_outS32ser[6]), 
        .ZN(KeyArray_S32reg_gff_1_SFF_6_n10) );
  DFF_X1 KeyArray_S32reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        KeyArray_S32reg_gff_1_SFF_6_n5), .CK(clk), .Q(KeyArray_outS32ser[6]), 
        .QN() );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_7_U3 ( .A1(KeyArray_S32reg_gff_1_SFF_7_n2), .A2(KeyArray_S32reg_gff_1_SFF_7_n1), .ZN(KeyArray_S32reg_gff_1_SFF_7_n5) );
  OR2_X1 KeyArray_S32reg_gff_1_SFF_7_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S32reg_gff_1_SFF_7_n10), .ZN(KeyArray_S32reg_gff_1_SFF_7_n1)
         );
  NAND2_X1 KeyArray_S32reg_gff_1_SFF_7_U1 ( .A1(KeyArray_S32reg_gff_1_SFF_7_QD), .A2(KeyArray_n18), .ZN(KeyArray_S32reg_gff_1_SFF_7_n2) );
  XOR2_X1 KeyArray_S32reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A(
        KeyArray_outS33ser[7]), .B(KeyArray_outS02ser[7]), .Z(
        KeyArray_S32reg_gff_1_SFF_7_MUXInst_X) );
  AND2_X1 KeyArray_S32reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A1(KeyArray_n21), 
        .A2(KeyArray_S32reg_gff_1_SFF_7_MUXInst_X), .ZN(
        KeyArray_S32reg_gff_1_SFF_7_MUXInst_Y) );
  XOR2_X1 KeyArray_S32reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A(
        KeyArray_S32reg_gff_1_SFF_7_MUXInst_Y), .B(KeyArray_outS33ser[7]), .Z(
        KeyArray_S32reg_gff_1_SFF_7_QD) );
  INV_X1 KeyArray_S32reg_gff_1_SFF_7_Q_reg_U1 ( .A(KeyArray_outS32ser[7]), 
        .ZN(KeyArray_S32reg_gff_1_SFF_7_n10) );
  DFF_X1 KeyArray_S32reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        KeyArray_S32reg_gff_1_SFF_7_n5), .CK(clk), .Q(KeyArray_outS32ser[7]), 
        .QN() );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_0_U3 ( .A1(KeyArray_S33reg_gff_1_SFF_0_n2), .A2(KeyArray_S33reg_gff_1_SFF_0_n1), .ZN(KeyArray_S33reg_gff_1_SFF_0_n5) );
  OR2_X1 KeyArray_S33reg_gff_1_SFF_0_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S33reg_gff_1_SFF_0_n10), .ZN(KeyArray_S33reg_gff_1_SFF_0_n1)
         );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_0_U1 ( .A1(KeyArray_S33reg_gff_1_SFF_0_QD), .A2(KeyArray_n18), .ZN(KeyArray_S33reg_gff_1_SFF_0_n2) );
  XOR2_X1 KeyArray_S33reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A(
        KeyArray_inS33ser[0]), .B(KeyArray_outS03ser[0]), .Z(
        KeyArray_S33reg_gff_1_SFF_0_MUXInst_X) );
  AND2_X1 KeyArray_S33reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A1(KeyArray_n21), 
        .A2(KeyArray_S33reg_gff_1_SFF_0_MUXInst_X), .ZN(
        KeyArray_S33reg_gff_1_SFF_0_MUXInst_Y) );
  XOR2_X1 KeyArray_S33reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A(
        KeyArray_S33reg_gff_1_SFF_0_MUXInst_Y), .B(KeyArray_inS33ser[0]), .Z(
        KeyArray_S33reg_gff_1_SFF_0_QD) );
  INV_X1 KeyArray_S33reg_gff_1_SFF_0_Q_reg_U1 ( .A(KeyArray_outS33ser[0]), 
        .ZN(KeyArray_S33reg_gff_1_SFF_0_n10) );
  DFF_X1 KeyArray_S33reg_gff_1_SFF_0_Q_reg_FF_FF ( .D(
        KeyArray_S33reg_gff_1_SFF_0_n5), .CK(clk), .Q(KeyArray_outS33ser[0]), 
        .QN() );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_1_U3 ( .A1(KeyArray_S33reg_gff_1_SFF_1_n2), .A2(KeyArray_S33reg_gff_1_SFF_1_n1), .ZN(KeyArray_S33reg_gff_1_SFF_1_n5) );
  OR2_X1 KeyArray_S33reg_gff_1_SFF_1_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S33reg_gff_1_SFF_1_n10), .ZN(KeyArray_S33reg_gff_1_SFF_1_n1)
         );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_1_U1 ( .A1(KeyArray_S33reg_gff_1_SFF_1_QD), .A2(KeyArray_n18), .ZN(KeyArray_S33reg_gff_1_SFF_1_n2) );
  XOR2_X1 KeyArray_S33reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A(
        KeyArray_inS33ser[1]), .B(KeyArray_outS03ser[1]), .Z(
        KeyArray_S33reg_gff_1_SFF_1_MUXInst_X) );
  AND2_X1 KeyArray_S33reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A1(KeyArray_n21), 
        .A2(KeyArray_S33reg_gff_1_SFF_1_MUXInst_X), .ZN(
        KeyArray_S33reg_gff_1_SFF_1_MUXInst_Y) );
  XOR2_X1 KeyArray_S33reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A(
        KeyArray_S33reg_gff_1_SFF_1_MUXInst_Y), .B(KeyArray_inS33ser[1]), .Z(
        KeyArray_S33reg_gff_1_SFF_1_QD) );
  INV_X1 KeyArray_S33reg_gff_1_SFF_1_Q_reg_U1 ( .A(KeyArray_outS33ser[1]), 
        .ZN(KeyArray_S33reg_gff_1_SFF_1_n10) );
  DFF_X1 KeyArray_S33reg_gff_1_SFF_1_Q_reg_FF_FF ( .D(
        KeyArray_S33reg_gff_1_SFF_1_n5), .CK(clk), .Q(KeyArray_outS33ser[1]), 
        .QN() );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_2_U3 ( .A1(KeyArray_S33reg_gff_1_SFF_2_n2), .A2(KeyArray_S33reg_gff_1_SFF_2_n1), .ZN(KeyArray_S33reg_gff_1_SFF_2_n5) );
  OR2_X1 KeyArray_S33reg_gff_1_SFF_2_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S33reg_gff_1_SFF_2_n10), .ZN(KeyArray_S33reg_gff_1_SFF_2_n1)
         );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_2_U1 ( .A1(KeyArray_S33reg_gff_1_SFF_2_QD), .A2(KeyArray_n18), .ZN(KeyArray_S33reg_gff_1_SFF_2_n2) );
  XOR2_X1 KeyArray_S33reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A(
        KeyArray_inS33ser[2]), .B(KeyArray_outS03ser[2]), .Z(
        KeyArray_S33reg_gff_1_SFF_2_MUXInst_X) );
  AND2_X1 KeyArray_S33reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A1(KeyArray_n21), 
        .A2(KeyArray_S33reg_gff_1_SFF_2_MUXInst_X), .ZN(
        KeyArray_S33reg_gff_1_SFF_2_MUXInst_Y) );
  XOR2_X1 KeyArray_S33reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A(
        KeyArray_S33reg_gff_1_SFF_2_MUXInst_Y), .B(KeyArray_inS33ser[2]), .Z(
        KeyArray_S33reg_gff_1_SFF_2_QD) );
  INV_X1 KeyArray_S33reg_gff_1_SFF_2_Q_reg_U1 ( .A(KeyArray_outS33ser[2]), 
        .ZN(KeyArray_S33reg_gff_1_SFF_2_n10) );
  DFF_X1 KeyArray_S33reg_gff_1_SFF_2_Q_reg_FF_FF ( .D(
        KeyArray_S33reg_gff_1_SFF_2_n5), .CK(clk), .Q(KeyArray_outS33ser[2]), 
        .QN() );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_3_U3 ( .A1(KeyArray_S33reg_gff_1_SFF_3_n2), .A2(KeyArray_S33reg_gff_1_SFF_3_n1), .ZN(KeyArray_S33reg_gff_1_SFF_3_n5) );
  OR2_X1 KeyArray_S33reg_gff_1_SFF_3_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S33reg_gff_1_SFF_3_n10), .ZN(KeyArray_S33reg_gff_1_SFF_3_n1)
         );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_3_U1 ( .A1(KeyArray_S33reg_gff_1_SFF_3_QD), .A2(KeyArray_n18), .ZN(KeyArray_S33reg_gff_1_SFF_3_n2) );
  XOR2_X1 KeyArray_S33reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A(
        KeyArray_inS33ser[3]), .B(KeyArray_outS03ser[3]), .Z(
        KeyArray_S33reg_gff_1_SFF_3_MUXInst_X) );
  AND2_X1 KeyArray_S33reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A1(KeyArray_n21), 
        .A2(KeyArray_S33reg_gff_1_SFF_3_MUXInst_X), .ZN(
        KeyArray_S33reg_gff_1_SFF_3_MUXInst_Y) );
  XOR2_X1 KeyArray_S33reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A(
        KeyArray_S33reg_gff_1_SFF_3_MUXInst_Y), .B(KeyArray_inS33ser[3]), .Z(
        KeyArray_S33reg_gff_1_SFF_3_QD) );
  INV_X1 KeyArray_S33reg_gff_1_SFF_3_Q_reg_U1 ( .A(KeyArray_outS33ser[3]), 
        .ZN(KeyArray_S33reg_gff_1_SFF_3_n10) );
  DFF_X1 KeyArray_S33reg_gff_1_SFF_3_Q_reg_FF_FF ( .D(
        KeyArray_S33reg_gff_1_SFF_3_n5), .CK(clk), .Q(KeyArray_outS33ser[3]), 
        .QN() );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_4_U3 ( .A1(KeyArray_S33reg_gff_1_SFF_4_n2), .A2(KeyArray_S33reg_gff_1_SFF_4_n1), .ZN(KeyArray_S33reg_gff_1_SFF_4_n5) );
  OR2_X1 KeyArray_S33reg_gff_1_SFF_4_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S33reg_gff_1_SFF_4_n10), .ZN(KeyArray_S33reg_gff_1_SFF_4_n1)
         );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_4_U1 ( .A1(KeyArray_S33reg_gff_1_SFF_4_QD), .A2(KeyArray_n18), .ZN(KeyArray_S33reg_gff_1_SFF_4_n2) );
  XOR2_X1 KeyArray_S33reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A(
        KeyArray_inS33ser[4]), .B(KeyArray_outS03ser[4]), .Z(
        KeyArray_S33reg_gff_1_SFF_4_MUXInst_X) );
  AND2_X1 KeyArray_S33reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A1(KeyArray_n21), 
        .A2(KeyArray_S33reg_gff_1_SFF_4_MUXInst_X), .ZN(
        KeyArray_S33reg_gff_1_SFF_4_MUXInst_Y) );
  XOR2_X1 KeyArray_S33reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A(
        KeyArray_S33reg_gff_1_SFF_4_MUXInst_Y), .B(KeyArray_inS33ser[4]), .Z(
        KeyArray_S33reg_gff_1_SFF_4_QD) );
  INV_X1 KeyArray_S33reg_gff_1_SFF_4_Q_reg_U1 ( .A(KeyArray_outS33ser[4]), 
        .ZN(KeyArray_S33reg_gff_1_SFF_4_n10) );
  DFF_X1 KeyArray_S33reg_gff_1_SFF_4_Q_reg_FF_FF ( .D(
        KeyArray_S33reg_gff_1_SFF_4_n5), .CK(clk), .Q(KeyArray_outS33ser[4]), 
        .QN() );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_5_U3 ( .A1(KeyArray_S33reg_gff_1_SFF_5_n2), .A2(KeyArray_S33reg_gff_1_SFF_5_n1), .ZN(KeyArray_S33reg_gff_1_SFF_5_n5) );
  OR2_X1 KeyArray_S33reg_gff_1_SFF_5_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S33reg_gff_1_SFF_5_n10), .ZN(KeyArray_S33reg_gff_1_SFF_5_n1)
         );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_5_U1 ( .A1(KeyArray_S33reg_gff_1_SFF_5_QD), .A2(KeyArray_n18), .ZN(KeyArray_S33reg_gff_1_SFF_5_n2) );
  XOR2_X1 KeyArray_S33reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A(
        KeyArray_inS33ser[5]), .B(KeyArray_outS03ser[5]), .Z(
        KeyArray_S33reg_gff_1_SFF_5_MUXInst_X) );
  AND2_X1 KeyArray_S33reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A1(KeyArray_n21), 
        .A2(KeyArray_S33reg_gff_1_SFF_5_MUXInst_X), .ZN(
        KeyArray_S33reg_gff_1_SFF_5_MUXInst_Y) );
  XOR2_X1 KeyArray_S33reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A(
        KeyArray_S33reg_gff_1_SFF_5_MUXInst_Y), .B(KeyArray_inS33ser[5]), .Z(
        KeyArray_S33reg_gff_1_SFF_5_QD) );
  INV_X1 KeyArray_S33reg_gff_1_SFF_5_Q_reg_U1 ( .A(KeyArray_outS33ser[5]), 
        .ZN(KeyArray_S33reg_gff_1_SFF_5_n10) );
  DFF_X1 KeyArray_S33reg_gff_1_SFF_5_Q_reg_FF_FF ( .D(
        KeyArray_S33reg_gff_1_SFF_5_n5), .CK(clk), .Q(KeyArray_outS33ser[5]), 
        .QN() );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_6_U3 ( .A1(KeyArray_S33reg_gff_1_SFF_6_n2), .A2(KeyArray_S33reg_gff_1_SFF_6_n1), .ZN(KeyArray_S33reg_gff_1_SFF_6_n5) );
  OR2_X1 KeyArray_S33reg_gff_1_SFF_6_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S33reg_gff_1_SFF_6_n10), .ZN(KeyArray_S33reg_gff_1_SFF_6_n1)
         );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_6_U1 ( .A1(KeyArray_S33reg_gff_1_SFF_6_QD), .A2(KeyArray_n18), .ZN(KeyArray_S33reg_gff_1_SFF_6_n2) );
  XOR2_X1 KeyArray_S33reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A(
        KeyArray_inS33ser[6]), .B(KeyArray_outS03ser[6]), .Z(
        KeyArray_S33reg_gff_1_SFF_6_MUXInst_X) );
  AND2_X1 KeyArray_S33reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A1(KeyArray_n21), 
        .A2(KeyArray_S33reg_gff_1_SFF_6_MUXInst_X), .ZN(
        KeyArray_S33reg_gff_1_SFF_6_MUXInst_Y) );
  XOR2_X1 KeyArray_S33reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A(
        KeyArray_S33reg_gff_1_SFF_6_MUXInst_Y), .B(KeyArray_inS33ser[6]), .Z(
        KeyArray_S33reg_gff_1_SFF_6_QD) );
  INV_X1 KeyArray_S33reg_gff_1_SFF_6_Q_reg_U1 ( .A(KeyArray_outS33ser[6]), 
        .ZN(KeyArray_S33reg_gff_1_SFF_6_n10) );
  DFF_X1 KeyArray_S33reg_gff_1_SFF_6_Q_reg_FF_FF ( .D(
        KeyArray_S33reg_gff_1_SFF_6_n5), .CK(clk), .Q(KeyArray_outS33ser[6]), 
        .QN() );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_7_U3 ( .A1(KeyArray_S33reg_gff_1_SFF_7_n2), .A2(KeyArray_S33reg_gff_1_SFF_7_n1), .ZN(KeyArray_S33reg_gff_1_SFF_7_n5) );
  OR2_X1 KeyArray_S33reg_gff_1_SFF_7_U2 ( .A1(KeyArray_n18), .A2(
        KeyArray_S33reg_gff_1_SFF_7_n10), .ZN(KeyArray_S33reg_gff_1_SFF_7_n1)
         );
  NAND2_X1 KeyArray_S33reg_gff_1_SFF_7_U1 ( .A1(KeyArray_S33reg_gff_1_SFF_7_QD), .A2(KeyArray_n18), .ZN(KeyArray_S33reg_gff_1_SFF_7_n2) );
  XOR2_X1 KeyArray_S33reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A(
        KeyArray_inS33ser[7]), .B(KeyArray_outS03ser[7]), .Z(
        KeyArray_S33reg_gff_1_SFF_7_MUXInst_X) );
  AND2_X1 KeyArray_S33reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A1(KeyArray_n21), 
        .A2(KeyArray_S33reg_gff_1_SFF_7_MUXInst_X), .ZN(
        KeyArray_S33reg_gff_1_SFF_7_MUXInst_Y) );
  XOR2_X1 KeyArray_S33reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A(
        KeyArray_S33reg_gff_1_SFF_7_MUXInst_Y), .B(KeyArray_inS33ser[7]), .Z(
        KeyArray_S33reg_gff_1_SFF_7_QD) );
  INV_X1 KeyArray_S33reg_gff_1_SFF_7_Q_reg_U1 ( .A(KeyArray_outS33ser[7]), 
        .ZN(KeyArray_S33reg_gff_1_SFF_7_n10) );
  DFF_X1 KeyArray_S33reg_gff_1_SFF_7_Q_reg_FF_FF ( .D(
        KeyArray_S33reg_gff_1_SFF_7_n5), .CK(clk), .Q(KeyArray_outS33ser[7]), 
        .QN() );
  XOR2_X1 KeyArray_MUX_inS00ser_mux_inst_0_XOR1_U1 ( .A(KeyArray_outS01ser_0_), 
        .B(KeyArray_outS01ser_XOR_00[0]), .Z(
        KeyArray_MUX_inS00ser_mux_inst_0_X) );
  AND2_X1 KeyArray_MUX_inS00ser_mux_inst_0_AND1_U1 ( .A1(
        KeyArray_nReset_selXOR), .A2(KeyArray_MUX_inS00ser_mux_inst_0_X), .ZN(
        KeyArray_MUX_inS00ser_mux_inst_0_Y) );
  XOR2_X1 KeyArray_MUX_inS00ser_mux_inst_0_XOR2_U1 ( .A(
        KeyArray_MUX_inS00ser_mux_inst_0_Y), .B(KeyArray_outS01ser_0_), .Z(
        KeyArray_inS00ser[0]) );
  XOR2_X1 KeyArray_MUX_inS00ser_mux_inst_1_XOR1_U1 ( .A(KeyArray_outS01ser_1_), 
        .B(KeyArray_outS01ser_XOR_00[1]), .Z(
        KeyArray_MUX_inS00ser_mux_inst_1_X) );
  AND2_X1 KeyArray_MUX_inS00ser_mux_inst_1_AND1_U1 ( .A1(
        KeyArray_nReset_selXOR), .A2(KeyArray_MUX_inS00ser_mux_inst_1_X), .ZN(
        KeyArray_MUX_inS00ser_mux_inst_1_Y) );
  XOR2_X1 KeyArray_MUX_inS00ser_mux_inst_1_XOR2_U1 ( .A(
        KeyArray_MUX_inS00ser_mux_inst_1_Y), .B(KeyArray_outS01ser_1_), .Z(
        KeyArray_inS00ser[1]) );
  XOR2_X1 KeyArray_MUX_inS00ser_mux_inst_2_XOR1_U1 ( .A(KeyArray_outS01ser_2_), 
        .B(KeyArray_outS01ser_XOR_00[2]), .Z(
        KeyArray_MUX_inS00ser_mux_inst_2_X) );
  AND2_X1 KeyArray_MUX_inS00ser_mux_inst_2_AND1_U1 ( .A1(
        KeyArray_nReset_selXOR), .A2(KeyArray_MUX_inS00ser_mux_inst_2_X), .ZN(
        KeyArray_MUX_inS00ser_mux_inst_2_Y) );
  XOR2_X1 KeyArray_MUX_inS00ser_mux_inst_2_XOR2_U1 ( .A(
        KeyArray_MUX_inS00ser_mux_inst_2_Y), .B(KeyArray_outS01ser_2_), .Z(
        KeyArray_inS00ser[2]) );
  XOR2_X1 KeyArray_MUX_inS00ser_mux_inst_3_XOR1_U1 ( .A(KeyArray_outS01ser_3_), 
        .B(KeyArray_outS01ser_XOR_00[3]), .Z(
        KeyArray_MUX_inS00ser_mux_inst_3_X) );
  AND2_X1 KeyArray_MUX_inS00ser_mux_inst_3_AND1_U1 ( .A1(
        KeyArray_nReset_selXOR), .A2(KeyArray_MUX_inS00ser_mux_inst_3_X), .ZN(
        KeyArray_MUX_inS00ser_mux_inst_3_Y) );
  XOR2_X1 KeyArray_MUX_inS00ser_mux_inst_3_XOR2_U1 ( .A(
        KeyArray_MUX_inS00ser_mux_inst_3_Y), .B(KeyArray_outS01ser_3_), .Z(
        KeyArray_inS00ser[3]) );
  XOR2_X1 KeyArray_MUX_inS00ser_mux_inst_4_XOR1_U1 ( .A(KeyArray_outS01ser_4_), 
        .B(KeyArray_outS01ser_XOR_00[4]), .Z(
        KeyArray_MUX_inS00ser_mux_inst_4_X) );
  AND2_X1 KeyArray_MUX_inS00ser_mux_inst_4_AND1_U1 ( .A1(
        KeyArray_nReset_selXOR), .A2(KeyArray_MUX_inS00ser_mux_inst_4_X), .ZN(
        KeyArray_MUX_inS00ser_mux_inst_4_Y) );
  XOR2_X1 KeyArray_MUX_inS00ser_mux_inst_4_XOR2_U1 ( .A(
        KeyArray_MUX_inS00ser_mux_inst_4_Y), .B(KeyArray_outS01ser_4_), .Z(
        KeyArray_inS00ser[4]) );
  XOR2_X1 KeyArray_MUX_inS00ser_mux_inst_5_XOR1_U1 ( .A(KeyArray_outS01ser_5_), 
        .B(KeyArray_outS01ser_XOR_00[5]), .Z(
        KeyArray_MUX_inS00ser_mux_inst_5_X) );
  AND2_X1 KeyArray_MUX_inS00ser_mux_inst_5_AND1_U1 ( .A1(
        KeyArray_nReset_selXOR), .A2(KeyArray_MUX_inS00ser_mux_inst_5_X), .ZN(
        KeyArray_MUX_inS00ser_mux_inst_5_Y) );
  XOR2_X1 KeyArray_MUX_inS00ser_mux_inst_5_XOR2_U1 ( .A(
        KeyArray_MUX_inS00ser_mux_inst_5_Y), .B(KeyArray_outS01ser_5_), .Z(
        KeyArray_inS00ser[5]) );
  XOR2_X1 KeyArray_MUX_inS00ser_mux_inst_6_XOR1_U1 ( .A(KeyArray_outS01ser_6_), 
        .B(KeyArray_outS01ser_XOR_00[6]), .Z(
        KeyArray_MUX_inS00ser_mux_inst_6_X) );
  AND2_X1 KeyArray_MUX_inS00ser_mux_inst_6_AND1_U1 ( .A1(
        KeyArray_nReset_selXOR), .A2(KeyArray_MUX_inS00ser_mux_inst_6_X), .ZN(
        KeyArray_MUX_inS00ser_mux_inst_6_Y) );
  XOR2_X1 KeyArray_MUX_inS00ser_mux_inst_6_XOR2_U1 ( .A(
        KeyArray_MUX_inS00ser_mux_inst_6_Y), .B(KeyArray_outS01ser_6_), .Z(
        KeyArray_inS00ser[6]) );
  XOR2_X1 KeyArray_MUX_inS00ser_mux_inst_7_XOR1_U1 ( .A(KeyArray_outS01ser_7_), 
        .B(KeyArray_outS01ser_XOR_00[7]), .Z(
        KeyArray_MUX_inS00ser_mux_inst_7_X) );
  AND2_X1 KeyArray_MUX_inS00ser_mux_inst_7_AND1_U1 ( .A1(
        KeyArray_nReset_selXOR), .A2(KeyArray_MUX_inS00ser_mux_inst_7_X), .ZN(
        KeyArray_MUX_inS00ser_mux_inst_7_Y) );
  XOR2_X1 KeyArray_MUX_inS00ser_mux_inst_7_XOR2_U1 ( .A(
        KeyArray_MUX_inS00ser_mux_inst_7_Y), .B(KeyArray_outS01ser_7_), .Z(
        KeyArray_inS00ser[7]) );
  XOR2_X1 KeyArray_MUX_inS33ser_mux_inst_0_XOR1_U1 ( .A(port_out[0]), .B(
        keyStateIn[0]), .Z(KeyArray_MUX_inS33ser_mux_inst_0_X) );
  AND2_X1 KeyArray_MUX_inS33ser_mux_inst_0_AND1_U1 ( .A1(n2), .A2(
        KeyArray_MUX_inS33ser_mux_inst_0_X), .ZN(
        KeyArray_MUX_inS33ser_mux_inst_0_Y) );
  XOR2_X1 KeyArray_MUX_inS33ser_mux_inst_0_XOR2_U1 ( .A(
        KeyArray_MUX_inS33ser_mux_inst_0_Y), .B(port_out[0]), .Z(
        KeyArray_inS33ser[0]) );
  XOR2_X1 KeyArray_MUX_inS33ser_mux_inst_1_XOR1_U1 ( .A(port_out[1]), .B(
        keyStateIn[1]), .Z(KeyArray_MUX_inS33ser_mux_inst_1_X) );
  AND2_X1 KeyArray_MUX_inS33ser_mux_inst_1_AND1_U1 ( .A1(n2), .A2(
        KeyArray_MUX_inS33ser_mux_inst_1_X), .ZN(
        KeyArray_MUX_inS33ser_mux_inst_1_Y) );
  XOR2_X1 KeyArray_MUX_inS33ser_mux_inst_1_XOR2_U1 ( .A(
        KeyArray_MUX_inS33ser_mux_inst_1_Y), .B(port_out[1]), .Z(
        KeyArray_inS33ser[1]) );
  XOR2_X1 KeyArray_MUX_inS33ser_mux_inst_2_XOR1_U1 ( .A(port_out[2]), .B(
        keyStateIn[2]), .Z(KeyArray_MUX_inS33ser_mux_inst_2_X) );
  AND2_X1 KeyArray_MUX_inS33ser_mux_inst_2_AND1_U1 ( .A1(n2), .A2(
        KeyArray_MUX_inS33ser_mux_inst_2_X), .ZN(
        KeyArray_MUX_inS33ser_mux_inst_2_Y) );
  XOR2_X1 KeyArray_MUX_inS33ser_mux_inst_2_XOR2_U1 ( .A(
        KeyArray_MUX_inS33ser_mux_inst_2_Y), .B(port_out[2]), .Z(
        KeyArray_inS33ser[2]) );
  XOR2_X1 KeyArray_MUX_inS33ser_mux_inst_3_XOR1_U1 ( .A(port_out[3]), .B(
        keyStateIn[3]), .Z(KeyArray_MUX_inS33ser_mux_inst_3_X) );
  AND2_X1 KeyArray_MUX_inS33ser_mux_inst_3_AND1_U1 ( .A1(n2), .A2(
        KeyArray_MUX_inS33ser_mux_inst_3_X), .ZN(
        KeyArray_MUX_inS33ser_mux_inst_3_Y) );
  XOR2_X1 KeyArray_MUX_inS33ser_mux_inst_3_XOR2_U1 ( .A(
        KeyArray_MUX_inS33ser_mux_inst_3_Y), .B(port_out[3]), .Z(
        KeyArray_inS33ser[3]) );
  XOR2_X1 KeyArray_MUX_inS33ser_mux_inst_4_XOR1_U1 ( .A(port_out[4]), .B(
        keyStateIn[4]), .Z(KeyArray_MUX_inS33ser_mux_inst_4_X) );
  AND2_X1 KeyArray_MUX_inS33ser_mux_inst_4_AND1_U1 ( .A1(n2), .A2(
        KeyArray_MUX_inS33ser_mux_inst_4_X), .ZN(
        KeyArray_MUX_inS33ser_mux_inst_4_Y) );
  XOR2_X1 KeyArray_MUX_inS33ser_mux_inst_4_XOR2_U1 ( .A(
        KeyArray_MUX_inS33ser_mux_inst_4_Y), .B(port_out[4]), .Z(
        KeyArray_inS33ser[4]) );
  XOR2_X1 KeyArray_MUX_inS33ser_mux_inst_5_XOR1_U1 ( .A(port_out[5]), .B(
        keyStateIn[5]), .Z(KeyArray_MUX_inS33ser_mux_inst_5_X) );
  AND2_X1 KeyArray_MUX_inS33ser_mux_inst_5_AND1_U1 ( .A1(n2), .A2(
        KeyArray_MUX_inS33ser_mux_inst_5_X), .ZN(
        KeyArray_MUX_inS33ser_mux_inst_5_Y) );
  XOR2_X1 KeyArray_MUX_inS33ser_mux_inst_5_XOR2_U1 ( .A(
        KeyArray_MUX_inS33ser_mux_inst_5_Y), .B(port_out[5]), .Z(
        KeyArray_inS33ser[5]) );
  XOR2_X1 KeyArray_MUX_inS33ser_mux_inst_6_XOR1_U1 ( .A(port_out[6]), .B(
        keyStateIn[6]), .Z(KeyArray_MUX_inS33ser_mux_inst_6_X) );
  AND2_X1 KeyArray_MUX_inS33ser_mux_inst_6_AND1_U1 ( .A1(n2), .A2(
        KeyArray_MUX_inS33ser_mux_inst_6_X), .ZN(
        KeyArray_MUX_inS33ser_mux_inst_6_Y) );
  XOR2_X1 KeyArray_MUX_inS33ser_mux_inst_6_XOR2_U1 ( .A(
        KeyArray_MUX_inS33ser_mux_inst_6_Y), .B(port_out[6]), .Z(
        KeyArray_inS33ser[6]) );
  XOR2_X1 KeyArray_MUX_inS33ser_mux_inst_7_XOR1_U1 ( .A(port_out[7]), .B(
        keyStateIn[7]), .Z(KeyArray_MUX_inS33ser_mux_inst_7_X) );
  AND2_X1 KeyArray_MUX_inS33ser_mux_inst_7_AND1_U1 ( .A1(n2), .A2(
        KeyArray_MUX_inS33ser_mux_inst_7_X), .ZN(
        KeyArray_MUX_inS33ser_mux_inst_7_Y) );
  XOR2_X1 KeyArray_MUX_inS33ser_mux_inst_7_XOR2_U1 ( .A(
        KeyArray_MUX_inS33ser_mux_inst_7_Y), .B(port_out[7]), .Z(
        KeyArray_inS33ser[7]) );
  XNOR2_X1 MixColumns_line0_U24 ( .A(MixColumns_line0_n16), .B(
        MixColumns_line0_n15), .ZN(MCout[31]) );
  XNOR2_X1 MixColumns_line0_U23 ( .A(MixColumns_line2_S02[0]), .B(
        MixColumns_line3_S02[0]), .ZN(MixColumns_line0_n15) );
  XOR2_X1 MixColumns_line0_U22 ( .A(port_out[6]), .B(MixColumns_line0_S13[7]), 
        .Z(MixColumns_line0_n16) );
  XNOR2_X1 MixColumns_line0_U21 ( .A(MixColumns_line0_n14), .B(
        MixColumns_line0_n13), .ZN(MCout[30]) );
  XNOR2_X1 MixColumns_line0_U20 ( .A(MixColumns_line2_S02[7]), .B(
        MixColumns_line3_S02[7]), .ZN(MixColumns_line0_n13) );
  XOR2_X1 MixColumns_line0_U19 ( .A(port_out[5]), .B(MixColumns_line0_S13[6]), 
        .Z(MixColumns_line0_n14) );
  XNOR2_X1 MixColumns_line0_U18 ( .A(MixColumns_line0_n12), .B(
        MixColumns_line0_n11), .ZN(MCout[29]) );
  XNOR2_X1 MixColumns_line0_U17 ( .A(MixColumns_line2_S02[6]), .B(
        MixColumns_line3_S02[6]), .ZN(MixColumns_line0_n11) );
  XOR2_X1 MixColumns_line0_U16 ( .A(port_out[4]), .B(MixColumns_line0_S13[5]), 
        .Z(MixColumns_line0_n12) );
  XNOR2_X1 MixColumns_line0_U15 ( .A(MixColumns_line0_n10), .B(
        MixColumns_line0_n9), .ZN(MCout[28]) );
  XNOR2_X1 MixColumns_line0_U14 ( .A(MixColumns_line2_S02[5]), .B(
        MixColumns_line3_S02[5]), .ZN(MixColumns_line0_n9) );
  XOR2_X1 MixColumns_line0_U13 ( .A(MixColumns_line0_S02[4]), .B(
        MixColumns_line0_S13[4]), .Z(MixColumns_line0_n10) );
  XNOR2_X1 MixColumns_line0_U12 ( .A(MixColumns_line0_n8), .B(
        MixColumns_line0_n7), .ZN(MCout[27]) );
  XNOR2_X1 MixColumns_line0_U11 ( .A(MCin[11]), .B(MCin[3]), .ZN(
        MixColumns_line0_n7) );
  XOR2_X1 MixColumns_line0_U10 ( .A(MixColumns_line0_S02[3]), .B(
        MixColumns_line0_S13[3]), .Z(MixColumns_line0_n8) );
  XNOR2_X1 MixColumns_line0_U9 ( .A(MixColumns_line0_n6), .B(
        MixColumns_line0_n5), .ZN(MCout[26]) );
  XNOR2_X1 MixColumns_line0_U8 ( .A(MCin[10]), .B(MCin[2]), .ZN(
        MixColumns_line0_n5) );
  XOR2_X1 MixColumns_line0_U7 ( .A(port_out[1]), .B(MixColumns_line0_S13[2]), 
        .Z(MixColumns_line0_n6) );
  XNOR2_X1 MixColumns_line0_U6 ( .A(MixColumns_line0_n4), .B(
        MixColumns_line0_n3), .ZN(MCout[25]) );
  XNOR2_X1 MixColumns_line0_U5 ( .A(MixColumns_line3_S02[2]), .B(
        MixColumns_line2_S02[2]), .ZN(MixColumns_line0_n3) );
  XOR2_X1 MixColumns_line0_U4 ( .A(MixColumns_line0_S02[1]), .B(
        MixColumns_line0_S13[1]), .Z(MixColumns_line0_n4) );
  XNOR2_X1 MixColumns_line0_U3 ( .A(MixColumns_line0_n2), .B(
        MixColumns_line0_n1), .ZN(MCout[24]) );
  XNOR2_X1 MixColumns_line0_U2 ( .A(MCin[0]), .B(MCin[8]), .ZN(
        MixColumns_line0_n1) );
  XOR2_X1 MixColumns_line0_U1 ( .A(port_out[7]), .B(MixColumns_line0_S13[0]), 
        .Z(MixColumns_line0_n2) );
  XOR2_X1 MixColumns_line0_timesTWO_U3 ( .A(port_out[7]), .B(port_out[3]), .Z(
        MixColumns_line0_S02[4]) );
  XOR2_X1 MixColumns_line0_timesTWO_U2 ( .A(port_out[7]), .B(port_out[2]), .Z(
        MixColumns_line0_S02[3]) );
  XOR2_X1 MixColumns_line0_timesTWO_U1 ( .A(port_out[7]), .B(port_out[0]), .Z(
        MixColumns_line0_S02[1]) );
  XOR2_X1 MixColumns_line0_timesTHREE_U8 ( .A(MixColumns_line1_S02[0]), .B(
        MixColumns_line1_S02[7]), .Z(MixColumns_line0_S13[7]) );
  XOR2_X1 MixColumns_line0_timesTHREE_U7 ( .A(MixColumns_line1_S02[7]), .B(
        MixColumns_line1_S02[6]), .Z(MixColumns_line0_S13[6]) );
  XOR2_X1 MixColumns_line0_timesTHREE_U6 ( .A(MixColumns_line1_S02[6]), .B(
        MixColumns_line1_S02[5]), .Z(MixColumns_line0_S13[5]) );
  XOR2_X1 MixColumns_line0_timesTHREE_U5 ( .A(MixColumns_line1_S02[5]), .B(
        MixColumns_line0_timesTHREE_input2[4]), .Z(MixColumns_line0_S13[4]) );
  XOR2_X1 MixColumns_line0_timesTHREE_U4 ( .A(MCin[19]), .B(
        MixColumns_line0_timesTHREE_input2[3]), .Z(MixColumns_line0_S13[3]) );
  XOR2_X1 MixColumns_line0_timesTHREE_U3 ( .A(MCin[18]), .B(
        MixColumns_line1_S02[2]), .Z(MixColumns_line0_S13[2]) );
  XOR2_X1 MixColumns_line0_timesTHREE_U2 ( .A(MixColumns_line1_S02[2]), .B(
        MixColumns_line0_timesTHREE_input2[1]), .Z(MixColumns_line0_S13[1]) );
  XOR2_X1 MixColumns_line0_timesTHREE_U1 ( .A(MCin[16]), .B(
        MixColumns_line1_S02[0]), .Z(MixColumns_line0_S13[0]) );
  XOR2_X1 MixColumns_line0_timesTHREE_timesTWO_U3 ( .A(MixColumns_line1_S02[0]), .B(MCin[19]), .Z(MixColumns_line0_timesTHREE_input2[4]) );
  XOR2_X1 MixColumns_line0_timesTHREE_timesTWO_U2 ( .A(MixColumns_line1_S02[0]), .B(MCin[18]), .Z(MixColumns_line0_timesTHREE_input2[3]) );
  XOR2_X1 MixColumns_line0_timesTHREE_timesTWO_U1 ( .A(MixColumns_line1_S02[0]), .B(MCin[16]), .Z(MixColumns_line0_timesTHREE_input2[1]) );
  XNOR2_X1 MixColumns_line1_U24 ( .A(MixColumns_line1_n16), .B(
        MixColumns_line1_n15), .ZN(MCout[23]) );
  XNOR2_X1 MixColumns_line1_U23 ( .A(MixColumns_line3_S02[0]), .B(port_out[7]), 
        .ZN(MixColumns_line1_n15) );
  XOR2_X1 MixColumns_line1_U22 ( .A(MixColumns_line1_S02[7]), .B(
        MixColumns_line1_S13[7]), .Z(MixColumns_line1_n16) );
  XNOR2_X1 MixColumns_line1_U21 ( .A(MixColumns_line1_n14), .B(
        MixColumns_line1_n13), .ZN(MCout[22]) );
  XNOR2_X1 MixColumns_line1_U20 ( .A(MixColumns_line3_S02[7]), .B(port_out[6]), 
        .ZN(MixColumns_line1_n13) );
  XOR2_X1 MixColumns_line1_U19 ( .A(MixColumns_line1_S02[6]), .B(
        MixColumns_line1_S13[6]), .Z(MixColumns_line1_n14) );
  XNOR2_X1 MixColumns_line1_U18 ( .A(MixColumns_line1_n12), .B(
        MixColumns_line1_n11), .ZN(MCout[21]) );
  XNOR2_X1 MixColumns_line1_U17 ( .A(MixColumns_line3_S02[6]), .B(port_out[5]), 
        .ZN(MixColumns_line1_n11) );
  XOR2_X1 MixColumns_line1_U16 ( .A(MixColumns_line1_S02[5]), .B(
        MixColumns_line1_S13[5]), .Z(MixColumns_line1_n12) );
  XNOR2_X1 MixColumns_line1_U15 ( .A(MixColumns_line1_n10), .B(
        MixColumns_line1_n9), .ZN(MCout[20]) );
  XNOR2_X1 MixColumns_line1_U14 ( .A(MixColumns_line3_S02[5]), .B(port_out[4]), 
        .ZN(MixColumns_line1_n9) );
  XOR2_X1 MixColumns_line1_U13 ( .A(MixColumns_line1_S02[4]), .B(
        MixColumns_line1_S13[4]), .Z(MixColumns_line1_n10) );
  XNOR2_X1 MixColumns_line1_U12 ( .A(MixColumns_line1_n8), .B(
        MixColumns_line1_n7), .ZN(MCout[19]) );
  XNOR2_X1 MixColumns_line1_U11 ( .A(MCin[3]), .B(port_out[3]), .ZN(
        MixColumns_line1_n7) );
  XOR2_X1 MixColumns_line1_U10 ( .A(MixColumns_line1_S02[3]), .B(
        MixColumns_line1_S13[3]), .Z(MixColumns_line1_n8) );
  XNOR2_X1 MixColumns_line1_U9 ( .A(MixColumns_line1_n6), .B(
        MixColumns_line1_n5), .ZN(MCout[18]) );
  XNOR2_X1 MixColumns_line1_U8 ( .A(MCin[2]), .B(port_out[2]), .ZN(
        MixColumns_line1_n5) );
  XOR2_X1 MixColumns_line1_U7 ( .A(MixColumns_line1_S02[2]), .B(
        MixColumns_line1_S13[2]), .Z(MixColumns_line1_n6) );
  XNOR2_X1 MixColumns_line1_U6 ( .A(MixColumns_line1_n4), .B(
        MixColumns_line1_n3), .ZN(MCout[17]) );
  XNOR2_X1 MixColumns_line1_U5 ( .A(port_out[1]), .B(MixColumns_line3_S02[2]), 
        .ZN(MixColumns_line1_n3) );
  XOR2_X1 MixColumns_line1_U4 ( .A(MixColumns_line1_S02[1]), .B(
        MixColumns_line1_S13[1]), .Z(MixColumns_line1_n4) );
  XNOR2_X1 MixColumns_line1_U3 ( .A(MixColumns_line1_n2), .B(
        MixColumns_line1_n1), .ZN(MCout[16]) );
  XNOR2_X1 MixColumns_line1_U2 ( .A(port_out[0]), .B(MCin[0]), .ZN(
        MixColumns_line1_n1) );
  XOR2_X1 MixColumns_line1_U1 ( .A(MixColumns_line1_S02[0]), .B(
        MixColumns_line1_S13[0]), .Z(MixColumns_line1_n2) );
  XOR2_X1 MixColumns_line1_timesTWO_U3 ( .A(MixColumns_line1_S02[0]), .B(
        MCin[19]), .Z(MixColumns_line1_S02[4]) );
  XOR2_X1 MixColumns_line1_timesTWO_U2 ( .A(MixColumns_line1_S02[0]), .B(
        MCin[18]), .Z(MixColumns_line1_S02[3]) );
  XOR2_X1 MixColumns_line1_timesTWO_U1 ( .A(MixColumns_line1_S02[0]), .B(
        MCin[16]), .Z(MixColumns_line1_S02[1]) );
  XOR2_X1 MixColumns_line1_timesTHREE_U8 ( .A(MixColumns_line2_S02[0]), .B(
        MixColumns_line2_S02[7]), .Z(MixColumns_line1_S13[7]) );
  XOR2_X1 MixColumns_line1_timesTHREE_U7 ( .A(MixColumns_line2_S02[7]), .B(
        MixColumns_line2_S02[6]), .Z(MixColumns_line1_S13[6]) );
  XOR2_X1 MixColumns_line1_timesTHREE_U6 ( .A(MixColumns_line2_S02[6]), .B(
        MixColumns_line2_S02[5]), .Z(MixColumns_line1_S13[5]) );
  XOR2_X1 MixColumns_line1_timesTHREE_U5 ( .A(MixColumns_line2_S02[5]), .B(
        MixColumns_line1_timesTHREE_input2[4]), .Z(MixColumns_line1_S13[4]) );
  XOR2_X1 MixColumns_line1_timesTHREE_U4 ( .A(MCin[11]), .B(
        MixColumns_line1_timesTHREE_input2[3]), .Z(MixColumns_line1_S13[3]) );
  XOR2_X1 MixColumns_line1_timesTHREE_U3 ( .A(MCin[10]), .B(
        MixColumns_line2_S02[2]), .Z(MixColumns_line1_S13[2]) );
  XOR2_X1 MixColumns_line1_timesTHREE_U2 ( .A(MixColumns_line2_S02[2]), .B(
        MixColumns_line1_timesTHREE_input2[1]), .Z(MixColumns_line1_S13[1]) );
  XOR2_X1 MixColumns_line1_timesTHREE_U1 ( .A(MCin[8]), .B(
        MixColumns_line2_S02[0]), .Z(MixColumns_line1_S13[0]) );
  XOR2_X1 MixColumns_line1_timesTHREE_timesTWO_U3 ( .A(MixColumns_line2_S02[0]), .B(MCin[11]), .Z(MixColumns_line1_timesTHREE_input2[4]) );
  XOR2_X1 MixColumns_line1_timesTHREE_timesTWO_U2 ( .A(MixColumns_line2_S02[0]), .B(MCin[10]), .Z(MixColumns_line1_timesTHREE_input2[3]) );
  XOR2_X1 MixColumns_line1_timesTHREE_timesTWO_U1 ( .A(MixColumns_line2_S02[0]), .B(MCin[8]), .Z(MixColumns_line1_timesTHREE_input2[1]) );
  XNOR2_X1 MixColumns_line2_U24 ( .A(MixColumns_line2_n16), .B(
        MixColumns_line2_n15), .ZN(MCout[15]) );
  XNOR2_X1 MixColumns_line2_U23 ( .A(port_out[7]), .B(MixColumns_line1_S02[0]), 
        .ZN(MixColumns_line2_n15) );
  XOR2_X1 MixColumns_line2_U22 ( .A(MixColumns_line2_S02[7]), .B(
        MixColumns_line2_S13[7]), .Z(MixColumns_line2_n16) );
  XNOR2_X1 MixColumns_line2_U21 ( .A(MixColumns_line2_n14), .B(
        MixColumns_line2_n13), .ZN(MCout[14]) );
  XNOR2_X1 MixColumns_line2_U20 ( .A(port_out[6]), .B(MixColumns_line1_S02[7]), 
        .ZN(MixColumns_line2_n13) );
  XOR2_X1 MixColumns_line2_U19 ( .A(MixColumns_line2_S02[6]), .B(
        MixColumns_line2_S13[6]), .Z(MixColumns_line2_n14) );
  XNOR2_X1 MixColumns_line2_U18 ( .A(MixColumns_line2_n12), .B(
        MixColumns_line2_n11), .ZN(MCout[13]) );
  XNOR2_X1 MixColumns_line2_U17 ( .A(port_out[5]), .B(MixColumns_line1_S02[6]), 
        .ZN(MixColumns_line2_n11) );
  XOR2_X1 MixColumns_line2_U16 ( .A(MixColumns_line2_S02[5]), .B(
        MixColumns_line2_S13[5]), .Z(MixColumns_line2_n12) );
  XNOR2_X1 MixColumns_line2_U15 ( .A(MixColumns_line2_n10), .B(
        MixColumns_line2_n9), .ZN(MCout[12]) );
  XNOR2_X1 MixColumns_line2_U14 ( .A(port_out[4]), .B(MixColumns_line1_S02[5]), 
        .ZN(MixColumns_line2_n9) );
  XOR2_X1 MixColumns_line2_U13 ( .A(MixColumns_line2_S02[4]), .B(
        MixColumns_line2_S13[4]), .Z(MixColumns_line2_n10) );
  XNOR2_X1 MixColumns_line2_U12 ( .A(MixColumns_line2_n8), .B(
        MixColumns_line2_n7), .ZN(MCout[11]) );
  XNOR2_X1 MixColumns_line2_U11 ( .A(port_out[3]), .B(MCin[19]), .ZN(
        MixColumns_line2_n7) );
  XOR2_X1 MixColumns_line2_U10 ( .A(MixColumns_line2_S02[3]), .B(
        MixColumns_line2_S13[3]), .Z(MixColumns_line2_n8) );
  XNOR2_X1 MixColumns_line2_U9 ( .A(MixColumns_line2_n6), .B(
        MixColumns_line2_n5), .ZN(MCout[10]) );
  XNOR2_X1 MixColumns_line2_U8 ( .A(port_out[2]), .B(MCin[18]), .ZN(
        MixColumns_line2_n5) );
  XOR2_X1 MixColumns_line2_U7 ( .A(MixColumns_line2_S02[2]), .B(
        MixColumns_line2_S13[2]), .Z(MixColumns_line2_n6) );
  XNOR2_X1 MixColumns_line2_U6 ( .A(MixColumns_line2_n4), .B(
        MixColumns_line2_n3), .ZN(MCout[9]) );
  XNOR2_X1 MixColumns_line2_U5 ( .A(MixColumns_line1_S02[2]), .B(port_out[1]), 
        .ZN(MixColumns_line2_n3) );
  XOR2_X1 MixColumns_line2_U4 ( .A(MixColumns_line2_S02[1]), .B(
        MixColumns_line2_S13[1]), .Z(MixColumns_line2_n4) );
  XNOR2_X1 MixColumns_line2_U3 ( .A(MixColumns_line2_n2), .B(
        MixColumns_line2_n1), .ZN(MCout[8]) );
  XNOR2_X1 MixColumns_line2_U2 ( .A(MCin[16]), .B(port_out[0]), .ZN(
        MixColumns_line2_n1) );
  XOR2_X1 MixColumns_line2_U1 ( .A(MixColumns_line2_S02[0]), .B(
        MixColumns_line2_S13[0]), .Z(MixColumns_line2_n2) );
  XOR2_X1 MixColumns_line2_timesTWO_U3 ( .A(MixColumns_line2_S02[0]), .B(
        MCin[11]), .Z(MixColumns_line2_S02[4]) );
  XOR2_X1 MixColumns_line2_timesTWO_U2 ( .A(MixColumns_line2_S02[0]), .B(
        MCin[10]), .Z(MixColumns_line2_S02[3]) );
  XOR2_X1 MixColumns_line2_timesTWO_U1 ( .A(MixColumns_line2_S02[0]), .B(
        MCin[8]), .Z(MixColumns_line2_S02[1]) );
  XOR2_X1 MixColumns_line2_timesTHREE_U8 ( .A(MixColumns_line3_S02[0]), .B(
        MixColumns_line3_S02[7]), .Z(MixColumns_line2_S13[7]) );
  XOR2_X1 MixColumns_line2_timesTHREE_U7 ( .A(MixColumns_line3_S02[7]), .B(
        MixColumns_line3_S02[6]), .Z(MixColumns_line2_S13[6]) );
  XOR2_X1 MixColumns_line2_timesTHREE_U6 ( .A(MixColumns_line3_S02[6]), .B(
        MixColumns_line3_S02[5]), .Z(MixColumns_line2_S13[5]) );
  XOR2_X1 MixColumns_line2_timesTHREE_U5 ( .A(MixColumns_line3_S02[5]), .B(
        MixColumns_line2_timesTHREE_input2[4]), .Z(MixColumns_line2_S13[4]) );
  XOR2_X1 MixColumns_line2_timesTHREE_U4 ( .A(MCin[3]), .B(
        MixColumns_line2_timesTHREE_input2[3]), .Z(MixColumns_line2_S13[3]) );
  XOR2_X1 MixColumns_line2_timesTHREE_U3 ( .A(MCin[2]), .B(
        MixColumns_line3_S02[2]), .Z(MixColumns_line2_S13[2]) );
  XOR2_X1 MixColumns_line2_timesTHREE_U2 ( .A(MixColumns_line3_S02[2]), .B(
        MixColumns_line2_timesTHREE_input2[1]), .Z(MixColumns_line2_S13[1]) );
  XOR2_X1 MixColumns_line2_timesTHREE_U1 ( .A(MCin[0]), .B(
        MixColumns_line3_S02[0]), .Z(MixColumns_line2_S13[0]) );
  XOR2_X1 MixColumns_line2_timesTHREE_timesTWO_U3 ( .A(MixColumns_line3_S02[0]), .B(MCin[3]), .Z(MixColumns_line2_timesTHREE_input2[4]) );
  XOR2_X1 MixColumns_line2_timesTHREE_timesTWO_U2 ( .A(MixColumns_line3_S02[0]), .B(MCin[2]), .Z(MixColumns_line2_timesTHREE_input2[3]) );
  XOR2_X1 MixColumns_line2_timesTHREE_timesTWO_U1 ( .A(MixColumns_line3_S02[0]), .B(MCin[0]), .Z(MixColumns_line2_timesTHREE_input2[1]) );
  XNOR2_X1 MixColumns_line3_U24 ( .A(MixColumns_line3_n16), .B(
        MixColumns_line3_n15), .ZN(MCout[7]) );
  XNOR2_X1 MixColumns_line3_U23 ( .A(MixColumns_line1_S02[0]), .B(
        MixColumns_line2_S02[0]), .ZN(MixColumns_line3_n15) );
  XOR2_X1 MixColumns_line3_U22 ( .A(MixColumns_line3_S02[7]), .B(
        MixColumns_line3_S13[7]), .Z(MixColumns_line3_n16) );
  XNOR2_X1 MixColumns_line3_U21 ( .A(MixColumns_line3_n14), .B(
        MixColumns_line3_n13), .ZN(MCout[6]) );
  XNOR2_X1 MixColumns_line3_U20 ( .A(MixColumns_line1_S02[7]), .B(
        MixColumns_line2_S02[7]), .ZN(MixColumns_line3_n13) );
  XOR2_X1 MixColumns_line3_U19 ( .A(MixColumns_line3_S02[6]), .B(
        MixColumns_line3_S13[6]), .Z(MixColumns_line3_n14) );
  XNOR2_X1 MixColumns_line3_U18 ( .A(MixColumns_line3_n12), .B(
        MixColumns_line3_n11), .ZN(MCout[5]) );
  XNOR2_X1 MixColumns_line3_U17 ( .A(MixColumns_line1_S02[6]), .B(
        MixColumns_line2_S02[6]), .ZN(MixColumns_line3_n11) );
  XOR2_X1 MixColumns_line3_U16 ( .A(MixColumns_line3_S02[5]), .B(
        MixColumns_line3_S13[5]), .Z(MixColumns_line3_n12) );
  XNOR2_X1 MixColumns_line3_U15 ( .A(MixColumns_line3_n10), .B(
        MixColumns_line3_n9), .ZN(MCout[4]) );
  XNOR2_X1 MixColumns_line3_U14 ( .A(MixColumns_line1_S02[5]), .B(
        MixColumns_line2_S02[5]), .ZN(MixColumns_line3_n9) );
  XOR2_X1 MixColumns_line3_U13 ( .A(MixColumns_line3_S02[4]), .B(
        MixColumns_line3_S13[4]), .Z(MixColumns_line3_n10) );
  XNOR2_X1 MixColumns_line3_U12 ( .A(MixColumns_line3_n8), .B(
        MixColumns_line3_n7), .ZN(MCout[3]) );
  XNOR2_X1 MixColumns_line3_U11 ( .A(MCin[19]), .B(MCin[11]), .ZN(
        MixColumns_line3_n7) );
  XOR2_X1 MixColumns_line3_U10 ( .A(MixColumns_line3_S02[3]), .B(
        MixColumns_line3_S13[3]), .Z(MixColumns_line3_n8) );
  XNOR2_X1 MixColumns_line3_U9 ( .A(MixColumns_line3_n6), .B(
        MixColumns_line3_n5), .ZN(MCout[2]) );
  XNOR2_X1 MixColumns_line3_U8 ( .A(MCin[18]), .B(MCin[10]), .ZN(
        MixColumns_line3_n5) );
  XOR2_X1 MixColumns_line3_U7 ( .A(MixColumns_line3_S02[2]), .B(
        MixColumns_line3_S13[2]), .Z(MixColumns_line3_n6) );
  XNOR2_X1 MixColumns_line3_U6 ( .A(MixColumns_line3_n4), .B(
        MixColumns_line3_n3), .ZN(MCout[1]) );
  XNOR2_X1 MixColumns_line3_U5 ( .A(MixColumns_line2_S02[2]), .B(
        MixColumns_line1_S02[2]), .ZN(MixColumns_line3_n3) );
  XOR2_X1 MixColumns_line3_U4 ( .A(MixColumns_line3_S02[1]), .B(
        MixColumns_line3_S13[1]), .Z(MixColumns_line3_n4) );
  XNOR2_X1 MixColumns_line3_U3 ( .A(MixColumns_line3_n2), .B(
        MixColumns_line3_n1), .ZN(MCout[0]) );
  XNOR2_X1 MixColumns_line3_U2 ( .A(MCin[8]), .B(MCin[16]), .ZN(
        MixColumns_line3_n1) );
  XOR2_X1 MixColumns_line3_U1 ( .A(MixColumns_line3_S02[0]), .B(
        MixColumns_line3_S13[0]), .Z(MixColumns_line3_n2) );
  XOR2_X1 MixColumns_line3_timesTWO_U3 ( .A(MixColumns_line3_S02[0]), .B(
        MCin[3]), .Z(MixColumns_line3_S02[4]) );
  XOR2_X1 MixColumns_line3_timesTWO_U2 ( .A(MixColumns_line3_S02[0]), .B(
        MCin[2]), .Z(MixColumns_line3_S02[3]) );
  XOR2_X1 MixColumns_line3_timesTWO_U1 ( .A(MixColumns_line3_S02[0]), .B(
        MCin[0]), .Z(MixColumns_line3_S02[1]) );
  XOR2_X1 MixColumns_line3_timesTHREE_U8 ( .A(port_out[7]), .B(port_out[6]), 
        .Z(MixColumns_line3_S13[7]) );
  XOR2_X1 MixColumns_line3_timesTHREE_U7 ( .A(port_out[6]), .B(port_out[5]), 
        .Z(MixColumns_line3_S13[6]) );
  XOR2_X1 MixColumns_line3_timesTHREE_U6 ( .A(port_out[5]), .B(port_out[4]), 
        .Z(MixColumns_line3_S13[5]) );
  XOR2_X1 MixColumns_line3_timesTHREE_U5 ( .A(port_out[4]), .B(
        MixColumns_line3_timesTHREE_input2_4_), .Z(MixColumns_line3_S13[4]) );
  XOR2_X1 MixColumns_line3_timesTHREE_U4 ( .A(port_out[3]), .B(
        MixColumns_line3_timesTHREE_input2_3_), .Z(MixColumns_line3_S13[3]) );
  XOR2_X1 MixColumns_line3_timesTHREE_U3 ( .A(port_out[2]), .B(port_out[1]), 
        .Z(MixColumns_line3_S13[2]) );
  XOR2_X1 MixColumns_line3_timesTHREE_U2 ( .A(port_out[1]), .B(
        MixColumns_line3_timesTHREE_input2_1_), .Z(MixColumns_line3_S13[1]) );
  XOR2_X1 MixColumns_line3_timesTHREE_U1 ( .A(port_out[0]), .B(port_out[7]), 
        .Z(MixColumns_line3_S13[0]) );
  XOR2_X1 MixColumns_line3_timesTHREE_timesTWO_U3 ( .A(port_out[7]), .B(
        port_out[3]), .Z(MixColumns_line3_timesTHREE_input2_4_) );
  XOR2_X1 MixColumns_line3_timesTHREE_timesTWO_U2 ( .A(port_out[7]), .B(
        port_out[2]), .Z(MixColumns_line3_timesTHREE_input2_3_) );
  XOR2_X1 MixColumns_line3_timesTHREE_timesTWO_U1 ( .A(port_out[7]), .B(
        port_out[0]), .Z(MixColumns_line3_timesTHREE_input2_1_) );
  NOR2_X1 calcRCon_U53 ( .A1(calcRCon_n10), .A2(calcRCon_n43), .ZN(
        roundConstant[7]) );
  NOR2_X1 calcRCon_U52 ( .A1(calcRCon_n2), .A2(calcRCon_n43), .ZN(
        roundConstant[6]) );
  NOR2_X1 calcRCon_U51 ( .A1(calcRCon_n4), .A2(calcRCon_n43), .ZN(
        roundConstant[5]) );
  NOR2_X1 calcRCon_U50 ( .A1(calcRCon_n3), .A2(calcRCon_n43), .ZN(
        roundConstant[4]) );
  AND2_X1 calcRCon_U49 ( .A1(calcRCon_s_current_state_3_), .A2(enRCon), .ZN(
        roundConstant[3]) );
  NOR2_X1 calcRCon_U48 ( .A1(calcRCon_n11), .A2(calcRCon_n43), .ZN(
        roundConstant[2]) );
  NOR2_X1 calcRCon_U47 ( .A1(calcRCon_n1), .A2(calcRCon_n43), .ZN(
        roundConstant[1]) );
  NOR2_X1 calcRCon_U46 ( .A1(calcRCon_n12), .A2(calcRCon_n43), .ZN(
        roundConstant[0]) );
  INV_X1 calcRCon_U45 ( .A(enRCon), .ZN(calcRCon_n43) );
  NAND2_X1 calcRCon_U44 ( .A1(calcRCon_n42), .A2(calcRCon_n41), .ZN(notFirst)
         );
  NOR2_X1 calcRCon_U43 ( .A1(calcRCon_n40), .A2(calcRCon_n39), .ZN(
        calcRCon_n41) );
  NAND2_X1 calcRCon_U42 ( .A1(calcRCon_n2), .A2(calcRCon_n4), .ZN(calcRCon_n39) );
  NAND2_X1 calcRCon_U41 ( .A1(calcRCon_s_current_state_3_), .A2(
        calcRCon_s_current_state_7_), .ZN(calcRCon_n40) );
  NOR2_X1 calcRCon_U40 ( .A1(calcRCon_n38), .A2(calcRCon_n37), .ZN(
        calcRCon_n42) );
  NAND2_X1 calcRCon_U39 ( .A1(calcRCon_s_current_state_2_), .A2(
        calcRCon_s_current_state_0_), .ZN(calcRCon_n37) );
  NAND2_X1 calcRCon_U38 ( .A1(calcRCon_n1), .A2(calcRCon_n3), .ZN(calcRCon_n38) );
  NAND2_X1 calcRCon_U37 ( .A1(calcRCon_n36), .A2(calcRCon_n35), .ZN(
        calcRCon_n51) );
  NAND2_X1 calcRCon_U36 ( .A1(calcRCon_n34), .A2(calcRCon_s_current_state_0_), 
        .ZN(calcRCon_n35) );
  NOR2_X1 calcRCon_U35 ( .A1(calcRCon_n6), .A2(calcRCon_n33), .ZN(calcRCon_n36) );
  NOR2_X1 calcRCon_U34 ( .A1(calcRCon_n34), .A2(calcRCon_n10), .ZN(
        calcRCon_n33) );
  NAND2_X1 calcRCon_U33 ( .A1(calcRCon_n32), .A2(calcRCon_n31), .ZN(
        calcRCon_n50) );
  NAND2_X1 calcRCon_U32 ( .A1(calcRCon_n34), .A2(calcRCon_s_current_state_1_), 
        .ZN(calcRCon_n31) );
  NAND2_X1 calcRCon_U31 ( .A1(calcRCon_n30), .A2(calcRCon_n29), .ZN(
        calcRCon_n32) );
  XOR2_X1 calcRCon_U30 ( .A(calcRCon_s_current_state_0_), .B(
        calcRCon_s_current_state_7_), .Z(calcRCon_n30) );
  NAND2_X1 calcRCon_U29 ( .A1(n2), .A2(calcRCon_n28), .ZN(calcRCon_n49) );
  NOR2_X1 calcRCon_U28 ( .A1(calcRCon_n27), .A2(calcRCon_n26), .ZN(
        calcRCon_n28) );
  NOR2_X1 calcRCon_U27 ( .A1(selSR), .A2(calcRCon_n11), .ZN(calcRCon_n26) );
  NOR2_X1 calcRCon_U26 ( .A1(calcRCon_n34), .A2(calcRCon_n1), .ZN(calcRCon_n27) );
  NAND2_X1 calcRCon_U25 ( .A1(calcRCon_n25), .A2(calcRCon_n24), .ZN(
        calcRCon_n48) );
  NAND2_X1 calcRCon_U24 ( .A1(calcRCon_n34), .A2(calcRCon_s_current_state_3_), 
        .ZN(calcRCon_n24) );
  NOR2_X1 calcRCon_U23 ( .A1(calcRCon_n23), .A2(calcRCon_n6), .ZN(calcRCon_n25) );
  NOR2_X1 calcRCon_U22 ( .A1(calcRCon_n34), .A2(calcRCon_n22), .ZN(
        calcRCon_n23) );
  XOR2_X1 calcRCon_U21 ( .A(calcRCon_n11), .B(calcRCon_s_current_state_7_), 
        .Z(calcRCon_n22) );
  NAND2_X1 calcRCon_U20 ( .A1(calcRCon_n21), .A2(calcRCon_n20), .ZN(
        calcRCon_n47) );
  NAND2_X1 calcRCon_U19 ( .A1(calcRCon_n34), .A2(calcRCon_s_current_state_4_), 
        .ZN(calcRCon_n20) );
  NAND2_X1 calcRCon_U18 ( .A1(calcRCon_n19), .A2(calcRCon_n29), .ZN(
        calcRCon_n21) );
  XOR2_X1 calcRCon_U17 ( .A(calcRCon_s_current_state_3_), .B(
        calcRCon_s_current_state_7_), .Z(calcRCon_n19) );
  NAND2_X1 calcRCon_U16 ( .A1(calcRCon_n18), .A2(calcRCon_n17), .ZN(
        calcRCon_n46) );
  NAND2_X1 calcRCon_U15 ( .A1(calcRCon_s_current_state_5_), .A2(calcRCon_n34), 
        .ZN(calcRCon_n17) );
  NAND2_X1 calcRCon_U14 ( .A1(calcRCon_s_current_state_4_), .A2(calcRCon_n29), 
        .ZN(calcRCon_n18) );
  NAND2_X1 calcRCon_U13 ( .A1(calcRCon_n16), .A2(calcRCon_n15), .ZN(
        calcRCon_n45) );
  NAND2_X1 calcRCon_U12 ( .A1(calcRCon_s_current_state_6_), .A2(calcRCon_n34), 
        .ZN(calcRCon_n15) );
  NAND2_X1 calcRCon_U11 ( .A1(calcRCon_s_current_state_5_), .A2(calcRCon_n29), 
        .ZN(calcRCon_n16) );
  NOR2_X1 calcRCon_U10 ( .A1(calcRCon_n34), .A2(calcRCon_n6), .ZN(calcRCon_n29) );
  NAND2_X1 calcRCon_U9 ( .A1(n2), .A2(calcRCon_n14), .ZN(calcRCon_n44) );
  NOR2_X1 calcRCon_U8 ( .A1(calcRCon_n13), .A2(calcRCon_n9), .ZN(calcRCon_n14)
         );
  NOR2_X1 calcRCon_U7 ( .A1(selSR), .A2(calcRCon_n10), .ZN(calcRCon_n9) );
  NOR2_X1 calcRCon_U6 ( .A1(calcRCon_n34), .A2(calcRCon_n2), .ZN(calcRCon_n13)
         );
  NAND2_X1 calcRCon_U5 ( .A1(calcRCon_s_current_state_5_), .A2(
        calcRCon_s_current_state_4_), .ZN(calcRCon_n7) );
  NAND2_X1 calcRCon_U4 ( .A1(calcRCon_s_current_state_1_), .A2(
        calcRCon_s_current_state_2_), .ZN(calcRCon_n8) );
  INV_X1 calcRCon_U3 ( .A(n2), .ZN(calcRCon_n6) );
  NOR2_X1 calcRCon_U2 ( .A1(selSR), .A2(calcRCon_n6), .ZN(calcRCon_n34) );
  NOR2_X1 calcRCon_U1 ( .A1(calcRCon_n8), .A2(calcRCon_n7), .ZN(intFinal) );
  INV_X1 calcRCon_s_current_state_reg_0__U1 ( .A(calcRCon_s_current_state_0_), 
        .ZN(calcRCon_n12) );
  DFF_X1 calcRCon_s_current_state_reg_0__FF_FF ( .D(calcRCon_n51), .CK(clk), 
        .Q(calcRCon_s_current_state_0_), .QN() );
  INV_X1 calcRCon_s_current_state_reg_1__U1 ( .A(calcRCon_s_current_state_1_), 
        .ZN(calcRCon_n1) );
  DFF_X1 calcRCon_s_current_state_reg_1__FF_FF ( .D(calcRCon_n50), .CK(clk), 
        .Q(calcRCon_s_current_state_1_), .QN() );
  INV_X1 calcRCon_s_current_state_reg_2__U1 ( .A(calcRCon_s_current_state_2_), 
        .ZN(calcRCon_n11) );
  DFF_X1 calcRCon_s_current_state_reg_2__FF_FF ( .D(calcRCon_n49), .CK(clk), 
        .Q(calcRCon_s_current_state_2_), .QN() );
  INV_X1 calcRCon_s_current_state_reg_3__U1 ( .A(calcRCon_s_current_state_3_), 
        .ZN(calcRCon_s_current_state_reg_3__QN) );
  DFF_X1 calcRCon_s_current_state_reg_3__FF_FF ( .D(calcRCon_n48), .CK(clk), 
        .Q(calcRCon_s_current_state_3_), .QN() );
  INV_X1 calcRCon_s_current_state_reg_4__U1 ( .A(calcRCon_s_current_state_4_), 
        .ZN(calcRCon_n3) );
  DFF_X1 calcRCon_s_current_state_reg_4__FF_FF ( .D(calcRCon_n47), .CK(clk), 
        .Q(calcRCon_s_current_state_4_), .QN() );
  INV_X1 calcRCon_s_current_state_reg_5__U1 ( .A(calcRCon_s_current_state_5_), 
        .ZN(calcRCon_n4) );
  DFF_X1 calcRCon_s_current_state_reg_5__FF_FF ( .D(calcRCon_n46), .CK(clk), 
        .Q(calcRCon_s_current_state_5_), .QN() );
  INV_X1 calcRCon_s_current_state_reg_6__U1 ( .A(calcRCon_s_current_state_6_), 
        .ZN(calcRCon_n2) );
  DFF_X1 calcRCon_s_current_state_reg_6__FF_FF ( .D(calcRCon_n45), .CK(clk), 
        .Q(calcRCon_s_current_state_6_), .QN() );
  INV_X1 calcRCon_s_current_state_reg_7__U1 ( .A(calcRCon_s_current_state_7_), 
        .ZN(calcRCon_n10) );
  DFF_X1 calcRCon_s_current_state_reg_7__FF_FF ( .D(calcRCon_n44), .CK(clk), 
        .Q(calcRCon_s_current_state_7_), .QN() );
  XOR2_X1 MUX_SboxIn_mux_inst_0_XOR1_U1 ( .A(StateOutXORroundKey[0]), .B(
        keySBIn[0]), .Z(MUX_SboxIn_mux_inst_0_X) );
  AND2_X1 MUX_SboxIn_mux_inst_0_AND1_U1 ( .A1(selMC), .A2(
        MUX_SboxIn_mux_inst_0_X), .ZN(MUX_SboxIn_mux_inst_0_Y) );
  XOR2_X1 MUX_SboxIn_mux_inst_0_XOR2_U1 ( .A(MUX_SboxIn_mux_inst_0_Y), .B(
        StateOutXORroundKey[0]), .Z(SboxIn[0]) );
  XOR2_X1 MUX_SboxIn_mux_inst_1_XOR1_U1 ( .A(StateOutXORroundKey[1]), .B(
        keySBIn[1]), .Z(MUX_SboxIn_mux_inst_1_X) );
  AND2_X1 MUX_SboxIn_mux_inst_1_AND1_U1 ( .A1(selMC), .A2(
        MUX_SboxIn_mux_inst_1_X), .ZN(MUX_SboxIn_mux_inst_1_Y) );
  XOR2_X1 MUX_SboxIn_mux_inst_1_XOR2_U1 ( .A(MUX_SboxIn_mux_inst_1_Y), .B(
        StateOutXORroundKey[1]), .Z(SboxIn[1]) );
  XOR2_X1 MUX_SboxIn_mux_inst_2_XOR1_U1 ( .A(StateOutXORroundKey[2]), .B(
        keySBIn[2]), .Z(MUX_SboxIn_mux_inst_2_X) );
  AND2_X1 MUX_SboxIn_mux_inst_2_AND1_U1 ( .A1(selMC), .A2(
        MUX_SboxIn_mux_inst_2_X), .ZN(MUX_SboxIn_mux_inst_2_Y) );
  XOR2_X1 MUX_SboxIn_mux_inst_2_XOR2_U1 ( .A(MUX_SboxIn_mux_inst_2_Y), .B(
        StateOutXORroundKey[2]), .Z(SboxIn[2]) );
  XOR2_X1 MUX_SboxIn_mux_inst_3_XOR1_U1 ( .A(StateOutXORroundKey[3]), .B(
        keySBIn[3]), .Z(MUX_SboxIn_mux_inst_3_X) );
  AND2_X1 MUX_SboxIn_mux_inst_3_AND1_U1 ( .A1(selMC), .A2(
        MUX_SboxIn_mux_inst_3_X), .ZN(MUX_SboxIn_mux_inst_3_Y) );
  XOR2_X1 MUX_SboxIn_mux_inst_3_XOR2_U1 ( .A(MUX_SboxIn_mux_inst_3_Y), .B(
        StateOutXORroundKey[3]), .Z(SboxIn[3]) );
  XOR2_X1 MUX_SboxIn_mux_inst_4_XOR1_U1 ( .A(StateOutXORroundKey[4]), .B(
        keySBIn[4]), .Z(MUX_SboxIn_mux_inst_4_X) );
  AND2_X1 MUX_SboxIn_mux_inst_4_AND1_U1 ( .A1(selMC), .A2(
        MUX_SboxIn_mux_inst_4_X), .ZN(MUX_SboxIn_mux_inst_4_Y) );
  XOR2_X1 MUX_SboxIn_mux_inst_4_XOR2_U1 ( .A(MUX_SboxIn_mux_inst_4_Y), .B(
        StateOutXORroundKey[4]), .Z(SboxIn[4]) );
  XOR2_X1 MUX_SboxIn_mux_inst_5_XOR1_U1 ( .A(StateOutXORroundKey[5]), .B(
        keySBIn[5]), .Z(MUX_SboxIn_mux_inst_5_X) );
  AND2_X1 MUX_SboxIn_mux_inst_5_AND1_U1 ( .A1(selMC), .A2(
        MUX_SboxIn_mux_inst_5_X), .ZN(MUX_SboxIn_mux_inst_5_Y) );
  XOR2_X1 MUX_SboxIn_mux_inst_5_XOR2_U1 ( .A(MUX_SboxIn_mux_inst_5_Y), .B(
        StateOutXORroundKey[5]), .Z(SboxIn[5]) );
  XOR2_X1 MUX_SboxIn_mux_inst_6_XOR1_U1 ( .A(StateOutXORroundKey[6]), .B(
        keySBIn[6]), .Z(MUX_SboxIn_mux_inst_6_X) );
  AND2_X1 MUX_SboxIn_mux_inst_6_AND1_U1 ( .A1(selMC), .A2(
        MUX_SboxIn_mux_inst_6_X), .ZN(MUX_SboxIn_mux_inst_6_Y) );
  XOR2_X1 MUX_SboxIn_mux_inst_6_XOR2_U1 ( .A(MUX_SboxIn_mux_inst_6_Y), .B(
        StateOutXORroundKey[6]), .Z(SboxIn[6]) );
  XOR2_X1 MUX_SboxIn_mux_inst_7_XOR1_U1 ( .A(StateOutXORroundKey[7]), .B(
        keySBIn[7]), .Z(MUX_SboxIn_mux_inst_7_X) );
  AND2_X1 MUX_SboxIn_mux_inst_7_AND1_U1 ( .A1(selMC), .A2(
        MUX_SboxIn_mux_inst_7_X), .ZN(MUX_SboxIn_mux_inst_7_Y) );
  XOR2_X1 MUX_SboxIn_mux_inst_7_XOR2_U1 ( .A(MUX_SboxIn_mux_inst_7_Y), .B(
        StateOutXORroundKey[7]), .Z(SboxIn[7]) );
  XOR2_X1 Inst_bSbox_XOR_T1_U1 ( .A(SboxIn[7]), .B(SboxIn[4]), .Z(
        Inst_bSbox_T1) );
  XOR2_X1 Inst_bSbox_XOR_T2_U1 ( .A(SboxIn[7]), .B(SboxIn[2]), .Z(
        Inst_bSbox_T2) );
  XOR2_X1 Inst_bSbox_XOR_T3_U1 ( .A(SboxIn[7]), .B(SboxIn[1]), .Z(
        Inst_bSbox_T3) );
  XOR2_X1 Inst_bSbox_XOR_T4_U1 ( .A(SboxIn[4]), .B(SboxIn[2]), .Z(
        Inst_bSbox_T4) );
  XOR2_X1 Inst_bSbox_XOR_T5_U1 ( .A(SboxIn[3]), .B(SboxIn[1]), .Z(
        Inst_bSbox_T5) );
  XOR2_X1 Inst_bSbox_XOR_T6_U1 ( .A(Inst_bSbox_T1), .B(Inst_bSbox_T5), .Z(
        Inst_bSbox_T6) );
  XOR2_X1 Inst_bSbox_XOR_T7_U1 ( .A(SboxIn[6]), .B(SboxIn[5]), .Z(
        Inst_bSbox_T7) );
  XOR2_X1 Inst_bSbox_XOR_T8_U1 ( .A(SboxIn[0]), .B(Inst_bSbox_T6), .Z(
        Inst_bSbox_T8) );
  XOR2_X1 Inst_bSbox_XOR_T9_U1 ( .A(SboxIn[0]), .B(Inst_bSbox_T7), .Z(
        Inst_bSbox_T9) );
  XOR2_X1 Inst_bSbox_XOR_T10_U1 ( .A(Inst_bSbox_T6), .B(Inst_bSbox_T7), .Z(
        Inst_bSbox_T10) );
  XOR2_X1 Inst_bSbox_XOR_T11_U1 ( .A(SboxIn[6]), .B(SboxIn[2]), .Z(
        Inst_bSbox_T11) );
  XOR2_X1 Inst_bSbox_XOR_T12_U1 ( .A(SboxIn[5]), .B(SboxIn[2]), .Z(
        Inst_bSbox_T12) );
  XOR2_X1 Inst_bSbox_XOR_T13_U1 ( .A(Inst_bSbox_T3), .B(Inst_bSbox_T4), .Z(
        Inst_bSbox_T13) );
  XOR2_X1 Inst_bSbox_XOR_T14_U1 ( .A(Inst_bSbox_T6), .B(Inst_bSbox_T11), .Z(
        Inst_bSbox_T14) );
  XOR2_X1 Inst_bSbox_XOR_T15_U1 ( .A(Inst_bSbox_T5), .B(Inst_bSbox_T11), .Z(
        Inst_bSbox_T15) );
  XOR2_X1 Inst_bSbox_XOR_T16_U1 ( .A(Inst_bSbox_T5), .B(Inst_bSbox_T12), .Z(
        Inst_bSbox_T16) );
  XOR2_X1 Inst_bSbox_XOR_T17_U1 ( .A(Inst_bSbox_T9), .B(Inst_bSbox_T16), .Z(
        Inst_bSbox_T17) );
  XOR2_X1 Inst_bSbox_XOR_T18_U1 ( .A(SboxIn[4]), .B(SboxIn[0]), .Z(
        Inst_bSbox_T18) );
  XOR2_X1 Inst_bSbox_XOR_T19_U1 ( .A(Inst_bSbox_T7), .B(Inst_bSbox_T18), .Z(
        Inst_bSbox_T19) );
  XOR2_X1 Inst_bSbox_XOR_T20_U1 ( .A(Inst_bSbox_T1), .B(Inst_bSbox_T19), .Z(
        Inst_bSbox_T20) );
  XOR2_X1 Inst_bSbox_XOR_T21_U1 ( .A(SboxIn[1]), .B(SboxIn[0]), .Z(
        Inst_bSbox_T21) );
  XOR2_X1 Inst_bSbox_XOR_T22_U1 ( .A(Inst_bSbox_T7), .B(Inst_bSbox_T21), .Z(
        Inst_bSbox_T22) );
  XOR2_X1 Inst_bSbox_XOR_T23_U1 ( .A(Inst_bSbox_T2), .B(Inst_bSbox_T22), .Z(
        Inst_bSbox_T23) );
  XOR2_X1 Inst_bSbox_XOR_T24_U1 ( .A(Inst_bSbox_T2), .B(Inst_bSbox_T10), .Z(
        Inst_bSbox_T24) );
  XOR2_X1 Inst_bSbox_XOR_T25_U1 ( .A(Inst_bSbox_T20), .B(Inst_bSbox_T17), .Z(
        Inst_bSbox_T25) );
  XOR2_X1 Inst_bSbox_XOR_T26_U1 ( .A(Inst_bSbox_T3), .B(Inst_bSbox_T16), .Z(
        Inst_bSbox_T26) );
  XOR2_X1 Inst_bSbox_XOR_T27_U1 ( .A(Inst_bSbox_T1), .B(Inst_bSbox_T12), .Z(
        Inst_bSbox_T27) );
  AND2_X1 Inst_bSbox_AND_M1_U1 ( .A1(Inst_bSbox_T13), .A2(Inst_bSbox_T6), .ZN(
        Inst_bSbox_M1) );
  AND2_X1 Inst_bSbox_AND_M2_U1 ( .A1(Inst_bSbox_T23), .A2(Inst_bSbox_T8), .ZN(
        Inst_bSbox_M2) );
  XOR2_X1 Inst_bSbox_XOR_M3_U1 ( .A(Inst_bSbox_T14), .B(Inst_bSbox_M1), .Z(
        Inst_bSbox_M3) );
  AND2_X1 Inst_bSbox_AND_M4_U1 ( .A1(Inst_bSbox_T19), .A2(SboxIn[0]), .ZN(
        Inst_bSbox_M4) );
  XOR2_X1 Inst_bSbox_XOR_M5_U1 ( .A(Inst_bSbox_M4), .B(Inst_bSbox_M1), .Z(
        Inst_bSbox_M5) );
  AND2_X1 Inst_bSbox_AND_M6_U1 ( .A1(Inst_bSbox_T3), .A2(Inst_bSbox_T16), .ZN(
        Inst_bSbox_M6) );
  AND2_X1 Inst_bSbox_AND_M7_U1 ( .A1(Inst_bSbox_T22), .A2(Inst_bSbox_T9), .ZN(
        Inst_bSbox_M7) );
  XOR2_X1 Inst_bSbox_XOR_M8_U1 ( .A(Inst_bSbox_T26), .B(Inst_bSbox_M6), .Z(
        Inst_bSbox_M8) );
  AND2_X1 Inst_bSbox_AND_M9_U1 ( .A1(Inst_bSbox_T20), .A2(Inst_bSbox_T17), 
        .ZN(Inst_bSbox_M9) );
  XOR2_X1 Inst_bSbox_XOR_M10_U1 ( .A(Inst_bSbox_M9), .B(Inst_bSbox_M6), .Z(
        Inst_bSbox_M10) );
  AND2_X1 Inst_bSbox_AND_M11_U1 ( .A1(Inst_bSbox_T1), .A2(Inst_bSbox_T15), 
        .ZN(Inst_bSbox_M11) );
  AND2_X1 Inst_bSbox_AND_M12_U1 ( .A1(Inst_bSbox_T4), .A2(Inst_bSbox_T27), 
        .ZN(Inst_bSbox_M12) );
  XOR2_X1 Inst_bSbox_XOR_M13_U1 ( .A(Inst_bSbox_M12), .B(Inst_bSbox_M11), .Z(
        Inst_bSbox_M13) );
  AND2_X1 Inst_bSbox_AND_M14_U1 ( .A1(Inst_bSbox_T2), .A2(Inst_bSbox_T10), 
        .ZN(Inst_bSbox_M14) );
  XOR2_X1 Inst_bSbox_XOR_M15_U1 ( .A(Inst_bSbox_M14), .B(Inst_bSbox_M11), .Z(
        Inst_bSbox_M15) );
  XOR2_X1 Inst_bSbox_XOR_M16_U1 ( .A(Inst_bSbox_M3), .B(Inst_bSbox_M2), .Z(
        Inst_bSbox_M16) );
  XOR2_X1 Inst_bSbox_XOR_M17_U1 ( .A(Inst_bSbox_M5), .B(Inst_bSbox_T24), .Z(
        Inst_bSbox_M17) );
  XOR2_X1 Inst_bSbox_XOR_M18_U1 ( .A(Inst_bSbox_M8), .B(Inst_bSbox_M7), .Z(
        Inst_bSbox_M18) );
  XOR2_X1 Inst_bSbox_XOR_M19_U1 ( .A(Inst_bSbox_M10), .B(Inst_bSbox_M15), .Z(
        Inst_bSbox_M19) );
  XOR2_X1 Inst_bSbox_XOR_M20_U1 ( .A(Inst_bSbox_M16), .B(Inst_bSbox_M13), .Z(
        Inst_bSbox_M20) );
  XOR2_X1 Inst_bSbox_XOR_M21_U1 ( .A(Inst_bSbox_M17), .B(Inst_bSbox_M15), .Z(
        Inst_bSbox_M21) );
  XOR2_X1 Inst_bSbox_XOR_M22_U1 ( .A(Inst_bSbox_M18), .B(Inst_bSbox_M13), .Z(
        Inst_bSbox_M22) );
  XOR2_X1 Inst_bSbox_XOR_M23_U1 ( .A(Inst_bSbox_M19), .B(Inst_bSbox_T25), .Z(
        Inst_bSbox_M23) );
  XOR2_X1 Inst_bSbox_XOR_M24_U1 ( .A(Inst_bSbox_M22), .B(Inst_bSbox_M23), .Z(
        Inst_bSbox_M24) );
  AND2_X1 Inst_bSbox_AND_M25_U1 ( .A1(Inst_bSbox_M22), .A2(Inst_bSbox_M20), 
        .ZN(Inst_bSbox_M25) );
  XOR2_X1 Inst_bSbox_XOR_M26_U1 ( .A(Inst_bSbox_M21), .B(Inst_bSbox_M25), .Z(
        Inst_bSbox_M26) );
  XOR2_X1 Inst_bSbox_XOR_M27_U1 ( .A(Inst_bSbox_M20), .B(Inst_bSbox_M21), .Z(
        Inst_bSbox_M27) );
  XOR2_X1 Inst_bSbox_XOR_M28_U1 ( .A(Inst_bSbox_M23), .B(Inst_bSbox_M25), .Z(
        Inst_bSbox_M28) );
  AND2_X1 Inst_bSbox_AND_M29_U1 ( .A1(Inst_bSbox_M28), .A2(Inst_bSbox_M27), 
        .ZN(Inst_bSbox_M29) );
  AND2_X1 Inst_bSbox_AND_M30_U1 ( .A1(Inst_bSbox_M26), .A2(Inst_bSbox_M24), 
        .ZN(Inst_bSbox_M30) );
  AND2_X1 Inst_bSbox_AND_M31_U1 ( .A1(Inst_bSbox_M20), .A2(Inst_bSbox_M23), 
        .ZN(Inst_bSbox_M31) );
  AND2_X1 Inst_bSbox_AND_M32_U1 ( .A1(Inst_bSbox_M27), .A2(Inst_bSbox_M31), 
        .ZN(Inst_bSbox_M32) );
  XOR2_X1 Inst_bSbox_XOR_M33_U1 ( .A(Inst_bSbox_M27), .B(Inst_bSbox_M25), .Z(
        Inst_bSbox_M33) );
  AND2_X1 Inst_bSbox_AND_M34_U1 ( .A1(Inst_bSbox_M21), .A2(Inst_bSbox_M22), 
        .ZN(Inst_bSbox_M34) );
  AND2_X1 Inst_bSbox_AND_M35_U1 ( .A1(Inst_bSbox_M24), .A2(Inst_bSbox_M34), 
        .ZN(Inst_bSbox_M35) );
  XOR2_X1 Inst_bSbox_XOR_M36_U1 ( .A(Inst_bSbox_M24), .B(Inst_bSbox_M25), .Z(
        Inst_bSbox_M36) );
  XOR2_X1 Inst_bSbox_XOR_M37_U1 ( .A(Inst_bSbox_M21), .B(Inst_bSbox_M29), .Z(
        Inst_bSbox_M37) );
  XOR2_X1 Inst_bSbox_XOR_M38_U1 ( .A(Inst_bSbox_M32), .B(Inst_bSbox_M33), .Z(
        Inst_bSbox_M38) );
  XOR2_X1 Inst_bSbox_XOR_M39_U1 ( .A(Inst_bSbox_M23), .B(Inst_bSbox_M30), .Z(
        Inst_bSbox_M39) );
  XOR2_X1 Inst_bSbox_XOR_M40_U1 ( .A(Inst_bSbox_M35), .B(Inst_bSbox_M36), .Z(
        Inst_bSbox_M40) );
  XOR2_X1 Inst_bSbox_XOR_M41_U1 ( .A(Inst_bSbox_M38), .B(Inst_bSbox_M40), .Z(
        Inst_bSbox_M41) );
  XOR2_X1 Inst_bSbox_XOR_M42_U1 ( .A(Inst_bSbox_M37), .B(Inst_bSbox_M39), .Z(
        Inst_bSbox_M42) );
  XOR2_X1 Inst_bSbox_XOR_M43_U1 ( .A(Inst_bSbox_M37), .B(Inst_bSbox_M38), .Z(
        Inst_bSbox_M43) );
  XOR2_X1 Inst_bSbox_XOR_M44_U1 ( .A(Inst_bSbox_M39), .B(Inst_bSbox_M40), .Z(
        Inst_bSbox_M44) );
  XOR2_X1 Inst_bSbox_XOR_M45_U1 ( .A(Inst_bSbox_M42), .B(Inst_bSbox_M41), .Z(
        Inst_bSbox_M45) );
  AND2_X1 Inst_bSbox_AND_M46_U1 ( .A1(Inst_bSbox_M44), .A2(Inst_bSbox_T6), 
        .ZN(Inst_bSbox_M46) );
  AND2_X1 Inst_bSbox_AND_M47_U1 ( .A1(Inst_bSbox_M40), .A2(Inst_bSbox_T8), 
        .ZN(Inst_bSbox_M47) );
  AND2_X1 Inst_bSbox_AND_M48_U1 ( .A1(Inst_bSbox_M39), .A2(SboxIn[0]), .ZN(
        Inst_bSbox_M48) );
  AND2_X1 Inst_bSbox_AND_M49_U1 ( .A1(Inst_bSbox_M43), .A2(Inst_bSbox_T16), 
        .ZN(Inst_bSbox_M49) );
  AND2_X1 Inst_bSbox_AND_M50_U1 ( .A1(Inst_bSbox_M38), .A2(Inst_bSbox_T9), 
        .ZN(Inst_bSbox_M50) );
  AND2_X1 Inst_bSbox_AND_M51_U1 ( .A1(Inst_bSbox_M37), .A2(Inst_bSbox_T17), 
        .ZN(Inst_bSbox_M51) );
  AND2_X1 Inst_bSbox_AND_M52_U1 ( .A1(Inst_bSbox_M42), .A2(Inst_bSbox_T15), 
        .ZN(Inst_bSbox_M52) );
  AND2_X1 Inst_bSbox_AND_M53_U1 ( .A1(Inst_bSbox_M45), .A2(Inst_bSbox_T27), 
        .ZN(Inst_bSbox_M53) );
  AND2_X1 Inst_bSbox_AND_M54_U1 ( .A1(Inst_bSbox_M41), .A2(Inst_bSbox_T10), 
        .ZN(Inst_bSbox_M54) );
  AND2_X1 Inst_bSbox_AND_M55_U1 ( .A1(Inst_bSbox_M44), .A2(Inst_bSbox_T13), 
        .ZN(Inst_bSbox_M55) );
  AND2_X1 Inst_bSbox_AND_M56_U1 ( .A1(Inst_bSbox_M40), .A2(Inst_bSbox_T23), 
        .ZN(Inst_bSbox_M56) );
  AND2_X1 Inst_bSbox_AND_M57_U1 ( .A1(Inst_bSbox_M39), .A2(Inst_bSbox_T19), 
        .ZN(Inst_bSbox_M57) );
  AND2_X1 Inst_bSbox_AND_M58_U1 ( .A1(Inst_bSbox_M43), .A2(Inst_bSbox_T3), 
        .ZN(Inst_bSbox_M58) );
  AND2_X1 Inst_bSbox_AND_M59_U1 ( .A1(Inst_bSbox_M38), .A2(Inst_bSbox_T22), 
        .ZN(Inst_bSbox_M59) );
  AND2_X1 Inst_bSbox_AND_M60_U1 ( .A1(Inst_bSbox_M37), .A2(Inst_bSbox_T20), 
        .ZN(Inst_bSbox_M60) );
  AND2_X1 Inst_bSbox_AND_M61_U1 ( .A1(Inst_bSbox_M42), .A2(Inst_bSbox_T1), 
        .ZN(Inst_bSbox_M61) );
  AND2_X1 Inst_bSbox_AND_M62_U1 ( .A1(Inst_bSbox_M45), .A2(Inst_bSbox_T4), 
        .ZN(Inst_bSbox_M62) );
  AND2_X1 Inst_bSbox_AND_M63_U1 ( .A1(Inst_bSbox_M41), .A2(Inst_bSbox_T2), 
        .ZN(Inst_bSbox_M63) );
  XOR2_X1 Inst_bSbox_XOR_L0_U1 ( .A(Inst_bSbox_M61), .B(Inst_bSbox_M62), .Z(
        Inst_bSbox_L0) );
  XOR2_X1 Inst_bSbox_XOR_L1_U1 ( .A(Inst_bSbox_M50), .B(Inst_bSbox_M56), .Z(
        Inst_bSbox_L1) );
  XOR2_X1 Inst_bSbox_XOR_L2_U1 ( .A(Inst_bSbox_M46), .B(Inst_bSbox_M48), .Z(
        Inst_bSbox_L2) );
  XOR2_X1 Inst_bSbox_XOR_L3_U1 ( .A(Inst_bSbox_M47), .B(Inst_bSbox_M55), .Z(
        Inst_bSbox_L3) );
  XOR2_X1 Inst_bSbox_XOR_L4_U1 ( .A(Inst_bSbox_M54), .B(Inst_bSbox_M58), .Z(
        Inst_bSbox_L4) );
  XOR2_X1 Inst_bSbox_XOR_L5_U1 ( .A(Inst_bSbox_M49), .B(Inst_bSbox_M61), .Z(
        Inst_bSbox_L5) );
  XOR2_X1 Inst_bSbox_XOR_L6_U1 ( .A(Inst_bSbox_M62), .B(Inst_bSbox_L5), .Z(
        Inst_bSbox_L6) );
  XOR2_X1 Inst_bSbox_XOR_L7_U1 ( .A(Inst_bSbox_M46), .B(Inst_bSbox_L3), .Z(
        Inst_bSbox_L7) );
  XOR2_X1 Inst_bSbox_XOR_L8_U1 ( .A(Inst_bSbox_M51), .B(Inst_bSbox_M59), .Z(
        Inst_bSbox_L8) );
  XOR2_X1 Inst_bSbox_XOR_L9_U1 ( .A(Inst_bSbox_M52), .B(Inst_bSbox_M53), .Z(
        Inst_bSbox_L9) );
  XOR2_X1 Inst_bSbox_XOR_L10_U1 ( .A(Inst_bSbox_M53), .B(Inst_bSbox_L4), .Z(
        Inst_bSbox_L10) );
  XOR2_X1 Inst_bSbox_XOR_L11_U1 ( .A(Inst_bSbox_M60), .B(Inst_bSbox_L2), .Z(
        Inst_bSbox_L11) );
  XOR2_X1 Inst_bSbox_XOR_L12_U1 ( .A(Inst_bSbox_M48), .B(Inst_bSbox_M51), .Z(
        Inst_bSbox_L12) );
  XOR2_X1 Inst_bSbox_XOR_L13_U1 ( .A(Inst_bSbox_M50), .B(Inst_bSbox_L0), .Z(
        Inst_bSbox_L13) );
  XOR2_X1 Inst_bSbox_XOR_L14_U1 ( .A(Inst_bSbox_M52), .B(Inst_bSbox_M61), .Z(
        Inst_bSbox_L14) );
  XOR2_X1 Inst_bSbox_XOR_L15_U1 ( .A(Inst_bSbox_M55), .B(Inst_bSbox_L1), .Z(
        Inst_bSbox_L15) );
  XOR2_X1 Inst_bSbox_XOR_L16_U1 ( .A(Inst_bSbox_M56), .B(Inst_bSbox_L0), .Z(
        Inst_bSbox_L16) );
  XOR2_X1 Inst_bSbox_XOR_L17_U1 ( .A(Inst_bSbox_M57), .B(Inst_bSbox_L1), .Z(
        Inst_bSbox_L17) );
  XOR2_X1 Inst_bSbox_XOR_L18_U1 ( .A(Inst_bSbox_M58), .B(Inst_bSbox_L8), .Z(
        Inst_bSbox_L18) );
  XOR2_X1 Inst_bSbox_XOR_L19_U1 ( .A(Inst_bSbox_M63), .B(Inst_bSbox_L4), .Z(
        Inst_bSbox_L19) );
  XOR2_X1 Inst_bSbox_XOR_L20_U1 ( .A(Inst_bSbox_L0), .B(Inst_bSbox_L1), .Z(
        Inst_bSbox_L20) );
  XOR2_X1 Inst_bSbox_XOR_L21_U1 ( .A(Inst_bSbox_L1), .B(Inst_bSbox_L7), .Z(
        Inst_bSbox_L21) );
  XOR2_X1 Inst_bSbox_XOR_L22_U1 ( .A(Inst_bSbox_L3), .B(Inst_bSbox_L12), .Z(
        Inst_bSbox_L22) );
  XOR2_X1 Inst_bSbox_XOR_L23_U1 ( .A(Inst_bSbox_L18), .B(Inst_bSbox_L2), .Z(
        Inst_bSbox_L23) );
  XOR2_X1 Inst_bSbox_XOR_L24_U1 ( .A(Inst_bSbox_L15), .B(Inst_bSbox_L9), .Z(
        Inst_bSbox_L24) );
  XOR2_X1 Inst_bSbox_XOR_L25_U1 ( .A(Inst_bSbox_L6), .B(Inst_bSbox_L10), .Z(
        Inst_bSbox_L25) );
  XOR2_X1 Inst_bSbox_XOR_L26_U1 ( .A(Inst_bSbox_L7), .B(Inst_bSbox_L9), .Z(
        Inst_bSbox_L26) );
  XOR2_X1 Inst_bSbox_XOR_L27_U1 ( .A(Inst_bSbox_L8), .B(Inst_bSbox_L10), .Z(
        Inst_bSbox_L27) );
  XOR2_X1 Inst_bSbox_XOR_L28_U1 ( .A(Inst_bSbox_L11), .B(Inst_bSbox_L14), .Z(
        Inst_bSbox_L28) );
  XOR2_X1 Inst_bSbox_XOR_L29_U1 ( .A(Inst_bSbox_L11), .B(Inst_bSbox_L17), .Z(
        Inst_bSbox_L29) );
  XOR2_X1 Inst_bSbox_XOR_S0_U1 ( .A(Inst_bSbox_L6), .B(Inst_bSbox_L24), .Z(
        SboxOut[7]) );
  XNOR2_X1 Inst_bSbox_XOR_S1_U1 ( .A(Inst_bSbox_L16), .B(Inst_bSbox_L26), .ZN(
        SboxOut[6]) );
  XNOR2_X1 Inst_bSbox_XOR_S2_U1 ( .A(Inst_bSbox_L19), .B(Inst_bSbox_L28), .ZN(
        SboxOut[5]) );
  XOR2_X1 Inst_bSbox_XOR_S3_U1 ( .A(Inst_bSbox_L6), .B(Inst_bSbox_L21), .Z(
        SboxOut[4]) );
  XOR2_X1 Inst_bSbox_XOR_S4_U1 ( .A(Inst_bSbox_L20), .B(Inst_bSbox_L22), .Z(
        SboxOut[3]) );
  XOR2_X1 Inst_bSbox_XOR_S5_U1 ( .A(Inst_bSbox_L25), .B(Inst_bSbox_L29), .Z(
        SboxOut[2]) );
  XNOR2_X1 Inst_bSbox_XOR_S6_U1 ( .A(Inst_bSbox_L13), .B(Inst_bSbox_L27), .ZN(
        SboxOut[1]) );
  XNOR2_X1 Inst_bSbox_XOR_S7_U1 ( .A(Inst_bSbox_L6), .B(Inst_bSbox_L23), .ZN(
        SboxOut[0]) );
endmodule

