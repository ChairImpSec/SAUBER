module eFPGA
    #(
        parameter MaxFramesPerCol=20,
        parameter FrameBitsPerRow=32,
        parameter NoConfigBits=0
    )
    (
        input Tile_X0Y1_A_O_top_0_t, //EXTERNAL
        input Tile_X0Y1_A_O_top_0_f, //EXTERNAL
        input Tile_X0Y1_A_O_top_1_t, //EXTERNAL
        input Tile_X0Y1_A_O_top_1_f, //EXTERNAL
        input Tile_X0Y1_A_prech1, //EXTERNAL
        input Tile_X0Y1_A_prech2, //EXTERNAL
        input Tile_X0Y1_A_DR_fault, //EXTERNAL
        output Tile_X0Y1_A_I_top_0_t, //EXTERNAL
        output Tile_X0Y1_A_I_top_0_f, //EXTERNAL
        output Tile_X0Y1_A_I_top_1_t, //EXTERNAL
        output Tile_X0Y1_A_I_top_1_f, //EXTERNAL
        output Tile_X0Y1_A_T_top, //EXTERNAL
        output Tile_X0Y1_A_F_masked1, //EXTERNAL
        output Tile_X0Y1_A_F_masked2, //EXTERNAL
        output Tile_X0Y1_A_config_C_bit0, //EXTERNAL
        output Tile_X0Y1_A_config_C_bit1, //EXTERNAL
        output Tile_X0Y1_A_config_C_bit2, //EXTERNAL
        output Tile_X0Y1_A_config_C_bit3, //EXTERNAL
        output Tile_X0Y1_B_config_C_bit0, //EXTERNAL
        output Tile_X0Y1_B_config_C_bit1, //EXTERNAL
        output Tile_X0Y1_B_config_C_bit2, //EXTERNAL
        output Tile_X0Y1_B_config_C_bit3, //EXTERNAL
        output Tile_X1Y1_F_masked1, //EXTERNAL
        output Tile_X1Y1_F_masked2, //EXTERNAL
        output Tile_X2Y1_F_masked1, //EXTERNAL
        output Tile_X2Y1_F_masked2, //EXTERNAL
        input Tile_X3Y1_R_t, //EXTERNAL
        input Tile_X3Y1_R_f, //EXTERNAL
        output Tile_X3Y1_F_masked1, //EXTERNAL
        output Tile_X3Y1_F_masked2, //EXTERNAL
        output Tile_X4Y1_F_masked1, //EXTERNAL
        output Tile_X4Y1_F_masked2, //EXTERNAL
        output Tile_X5Y1_F_masked1, //EXTERNAL
        output Tile_X5Y1_F_masked2, //EXTERNAL
        input Tile_X6Y1_R_t, //EXTERNAL
        input Tile_X6Y1_R_f, //EXTERNAL
        output Tile_X6Y1_F_masked1, //EXTERNAL
        output Tile_X6Y1_F_masked2, //EXTERNAL
        output Tile_X7Y1_F_masked1, //EXTERNAL
        output Tile_X7Y1_F_masked2, //EXTERNAL
        output Tile_X9Y1_F_ctrl, //EXTERNAL
        input Tile_X10Y1_A_O_top_0_t, //EXTERNAL
        input Tile_X10Y1_A_O_top_0_f, //EXTERNAL
        input Tile_X10Y1_A_prech2, //EXTERNAL
        input Tile_X10Y1_A_DR_fault, //EXTERNAL
        output Tile_X10Y1_A_I_top_0_t, //EXTERNAL
        output Tile_X10Y1_A_I_top_0_f, //EXTERNAL
        output Tile_X10Y1_A_T_top, //EXTERNAL
        output Tile_X10Y1_A_F_ctrl, //EXTERNAL
        input Tile_X0Y2_A_O_top_0_t, //EXTERNAL
        input Tile_X0Y2_A_O_top_0_f, //EXTERNAL
        input Tile_X0Y2_A_O_top_1_t, //EXTERNAL
        input Tile_X0Y2_A_O_top_1_f, //EXTERNAL
        input Tile_X0Y2_A_prech1, //EXTERNAL
        input Tile_X0Y2_A_prech2, //EXTERNAL
        input Tile_X0Y2_A_DR_fault, //EXTERNAL
        output Tile_X0Y2_A_I_top_0_t, //EXTERNAL
        output Tile_X0Y2_A_I_top_0_f, //EXTERNAL
        output Tile_X0Y2_A_I_top_1_t, //EXTERNAL
        output Tile_X0Y2_A_I_top_1_f, //EXTERNAL
        output Tile_X0Y2_A_T_top, //EXTERNAL
        output Tile_X0Y2_A_F_masked1, //EXTERNAL
        output Tile_X0Y2_A_F_masked2, //EXTERNAL
        output Tile_X0Y2_A_config_C_bit0, //EXTERNAL
        output Tile_X0Y2_A_config_C_bit1, //EXTERNAL
        output Tile_X0Y2_A_config_C_bit2, //EXTERNAL
        output Tile_X0Y2_A_config_C_bit3, //EXTERNAL
        output Tile_X0Y2_B_config_C_bit0, //EXTERNAL
        output Tile_X0Y2_B_config_C_bit1, //EXTERNAL
        output Tile_X0Y2_B_config_C_bit2, //EXTERNAL
        output Tile_X0Y2_B_config_C_bit3, //EXTERNAL
        output Tile_X1Y2_F_masked1, //EXTERNAL
        output Tile_X1Y2_F_masked2, //EXTERNAL
        output Tile_X2Y2_F_masked1, //EXTERNAL
        output Tile_X2Y2_F_masked2, //EXTERNAL
        input Tile_X3Y2_R_t, //EXTERNAL
        input Tile_X3Y2_R_f, //EXTERNAL
        output Tile_X3Y2_F_masked1, //EXTERNAL
        output Tile_X3Y2_F_masked2, //EXTERNAL
        output Tile_X4Y2_F_masked1, //EXTERNAL
        output Tile_X4Y2_F_masked2, //EXTERNAL
        output Tile_X5Y2_F_masked1, //EXTERNAL
        output Tile_X5Y2_F_masked2, //EXTERNAL
        input Tile_X6Y2_R_t, //EXTERNAL
        input Tile_X6Y2_R_f, //EXTERNAL
        output Tile_X6Y2_F_masked1, //EXTERNAL
        output Tile_X6Y2_F_masked2, //EXTERNAL
        output Tile_X7Y2_F_masked1, //EXTERNAL
        output Tile_X7Y2_F_masked2, //EXTERNAL
        output Tile_X9Y2_F_ctrl, //EXTERNAL
        input Tile_X10Y2_A_O_top_0_t, //EXTERNAL
        input Tile_X10Y2_A_O_top_0_f, //EXTERNAL
        input Tile_X10Y2_A_prech2, //EXTERNAL
        input Tile_X10Y2_A_DR_fault, //EXTERNAL
        output Tile_X10Y2_A_I_top_0_t, //EXTERNAL
        output Tile_X10Y2_A_I_top_0_f, //EXTERNAL
        output Tile_X10Y2_A_T_top, //EXTERNAL
        output Tile_X10Y2_A_F_ctrl, //EXTERNAL
        input Tile_X0Y3_A_O_top_0_t, //EXTERNAL
        input Tile_X0Y3_A_O_top_0_f, //EXTERNAL
        input Tile_X0Y3_A_O_top_1_t, //EXTERNAL
        input Tile_X0Y3_A_O_top_1_f, //EXTERNAL
        input Tile_X0Y3_A_prech1, //EXTERNAL
        input Tile_X0Y3_A_prech2, //EXTERNAL
        input Tile_X0Y3_A_DR_fault, //EXTERNAL
        output Tile_X0Y3_A_I_top_0_t, //EXTERNAL
        output Tile_X0Y3_A_I_top_0_f, //EXTERNAL
        output Tile_X0Y3_A_I_top_1_t, //EXTERNAL
        output Tile_X0Y3_A_I_top_1_f, //EXTERNAL
        output Tile_X0Y3_A_T_top, //EXTERNAL
        output Tile_X0Y3_A_F_masked1, //EXTERNAL
        output Tile_X0Y3_A_F_masked2, //EXTERNAL
        output Tile_X0Y3_A_config_C_bit0, //EXTERNAL
        output Tile_X0Y3_A_config_C_bit1, //EXTERNAL
        output Tile_X0Y3_A_config_C_bit2, //EXTERNAL
        output Tile_X0Y3_A_config_C_bit3, //EXTERNAL
        output Tile_X0Y3_B_config_C_bit0, //EXTERNAL
        output Tile_X0Y3_B_config_C_bit1, //EXTERNAL
        output Tile_X0Y3_B_config_C_bit2, //EXTERNAL
        output Tile_X0Y3_B_config_C_bit3, //EXTERNAL
        output Tile_X1Y3_F_masked1, //EXTERNAL
        output Tile_X1Y3_F_masked2, //EXTERNAL
        output Tile_X2Y3_F_masked1, //EXTERNAL
        output Tile_X2Y3_F_masked2, //EXTERNAL
        input Tile_X3Y3_R_t, //EXTERNAL
        input Tile_X3Y3_R_f, //EXTERNAL
        output Tile_X3Y3_F_masked1, //EXTERNAL
        output Tile_X3Y3_F_masked2, //EXTERNAL
        output Tile_X4Y3_F_masked1, //EXTERNAL
        output Tile_X4Y3_F_masked2, //EXTERNAL
        output Tile_X5Y3_F_masked1, //EXTERNAL
        output Tile_X5Y3_F_masked2, //EXTERNAL
        input Tile_X6Y3_R_t, //EXTERNAL
        input Tile_X6Y3_R_f, //EXTERNAL
        output Tile_X6Y3_F_masked1, //EXTERNAL
        output Tile_X6Y3_F_masked2, //EXTERNAL
        output Tile_X7Y3_F_masked1, //EXTERNAL
        output Tile_X7Y3_F_masked2, //EXTERNAL
        output Tile_X9Y3_F_ctrl, //EXTERNAL
        input Tile_X10Y3_A_O_top_0_t, //EXTERNAL
        input Tile_X10Y3_A_O_top_0_f, //EXTERNAL
        input Tile_X10Y3_A_prech2, //EXTERNAL
        input Tile_X10Y3_A_DR_fault, //EXTERNAL
        output Tile_X10Y3_A_I_top_0_t, //EXTERNAL
        output Tile_X10Y3_A_I_top_0_f, //EXTERNAL
        output Tile_X10Y3_A_T_top, //EXTERNAL
        output Tile_X10Y3_A_F_ctrl, //EXTERNAL
        input Tile_X0Y4_A_O_top_0_t, //EXTERNAL
        input Tile_X0Y4_A_O_top_0_f, //EXTERNAL
        input Tile_X0Y4_A_O_top_1_t, //EXTERNAL
        input Tile_X0Y4_A_O_top_1_f, //EXTERNAL
        input Tile_X0Y4_A_prech1, //EXTERNAL
        input Tile_X0Y4_A_prech2, //EXTERNAL
        input Tile_X0Y4_A_DR_fault, //EXTERNAL
        output Tile_X0Y4_A_I_top_0_t, //EXTERNAL
        output Tile_X0Y4_A_I_top_0_f, //EXTERNAL
        output Tile_X0Y4_A_I_top_1_t, //EXTERNAL
        output Tile_X0Y4_A_I_top_1_f, //EXTERNAL
        output Tile_X0Y4_A_T_top, //EXTERNAL
        output Tile_X0Y4_A_F_masked1, //EXTERNAL
        output Tile_X0Y4_A_F_masked2, //EXTERNAL
        output Tile_X0Y4_A_config_C_bit0, //EXTERNAL
        output Tile_X0Y4_A_config_C_bit1, //EXTERNAL
        output Tile_X0Y4_A_config_C_bit2, //EXTERNAL
        output Tile_X0Y4_A_config_C_bit3, //EXTERNAL
        output Tile_X0Y4_B_config_C_bit0, //EXTERNAL
        output Tile_X0Y4_B_config_C_bit1, //EXTERNAL
        output Tile_X0Y4_B_config_C_bit2, //EXTERNAL
        output Tile_X0Y4_B_config_C_bit3, //EXTERNAL
        output Tile_X1Y4_F_masked1, //EXTERNAL
        output Tile_X1Y4_F_masked2, //EXTERNAL
        output Tile_X2Y4_F_masked1, //EXTERNAL
        output Tile_X2Y4_F_masked2, //EXTERNAL
        input Tile_X3Y4_R_t, //EXTERNAL
        input Tile_X3Y4_R_f, //EXTERNAL
        output Tile_X3Y4_F_masked1, //EXTERNAL
        output Tile_X3Y4_F_masked2, //EXTERNAL
        output Tile_X4Y4_F_masked1, //EXTERNAL
        output Tile_X4Y4_F_masked2, //EXTERNAL
        output Tile_X5Y4_F_masked1, //EXTERNAL
        output Tile_X5Y4_F_masked2, //EXTERNAL
        input Tile_X6Y4_R_t, //EXTERNAL
        input Tile_X6Y4_R_f, //EXTERNAL
        output Tile_X6Y4_F_masked1, //EXTERNAL
        output Tile_X6Y4_F_masked2, //EXTERNAL
        output Tile_X7Y4_F_masked1, //EXTERNAL
        output Tile_X7Y4_F_masked2, //EXTERNAL
        output Tile_X9Y4_F_ctrl, //EXTERNAL
        input Tile_X10Y4_A_O_top_0_t, //EXTERNAL
        input Tile_X10Y4_A_O_top_0_f, //EXTERNAL
        input Tile_X10Y4_A_prech2, //EXTERNAL
        input Tile_X10Y4_A_DR_fault, //EXTERNAL
        output Tile_X10Y4_A_I_top_0_t, //EXTERNAL
        output Tile_X10Y4_A_I_top_0_f, //EXTERNAL
        output Tile_X10Y4_A_T_top, //EXTERNAL
        output Tile_X10Y4_A_F_ctrl, //EXTERNAL
        input Tile_X0Y5_A_O_top_0_t, //EXTERNAL
        input Tile_X0Y5_A_O_top_0_f, //EXTERNAL
        input Tile_X0Y5_A_O_top_1_t, //EXTERNAL
        input Tile_X0Y5_A_O_top_1_f, //EXTERNAL
        input Tile_X0Y5_A_prech1, //EXTERNAL
        input Tile_X0Y5_A_prech2, //EXTERNAL
        input Tile_X0Y5_A_DR_fault, //EXTERNAL
        output Tile_X0Y5_A_I_top_0_t, //EXTERNAL
        output Tile_X0Y5_A_I_top_0_f, //EXTERNAL
        output Tile_X0Y5_A_I_top_1_t, //EXTERNAL
        output Tile_X0Y5_A_I_top_1_f, //EXTERNAL
        output Tile_X0Y5_A_T_top, //EXTERNAL
        output Tile_X0Y5_A_F_masked1, //EXTERNAL
        output Tile_X0Y5_A_F_masked2, //EXTERNAL
        output Tile_X0Y5_A_config_C_bit0, //EXTERNAL
        output Tile_X0Y5_A_config_C_bit1, //EXTERNAL
        output Tile_X0Y5_A_config_C_bit2, //EXTERNAL
        output Tile_X0Y5_A_config_C_bit3, //EXTERNAL
        output Tile_X0Y5_B_config_C_bit0, //EXTERNAL
        output Tile_X0Y5_B_config_C_bit1, //EXTERNAL
        output Tile_X0Y5_B_config_C_bit2, //EXTERNAL
        output Tile_X0Y5_B_config_C_bit3, //EXTERNAL
        output Tile_X1Y5_F_masked1, //EXTERNAL
        output Tile_X1Y5_F_masked2, //EXTERNAL
        output Tile_X2Y5_F_masked1, //EXTERNAL
        output Tile_X2Y5_F_masked2, //EXTERNAL
        input Tile_X3Y5_R_t, //EXTERNAL
        input Tile_X3Y5_R_f, //EXTERNAL
        output Tile_X3Y5_F_masked1, //EXTERNAL
        output Tile_X3Y5_F_masked2, //EXTERNAL
        output Tile_X4Y5_F_masked1, //EXTERNAL
        output Tile_X4Y5_F_masked2, //EXTERNAL
        output Tile_X5Y5_F_masked1, //EXTERNAL
        output Tile_X5Y5_F_masked2, //EXTERNAL
        input Tile_X6Y5_R_t, //EXTERNAL
        input Tile_X6Y5_R_f, //EXTERNAL
        output Tile_X6Y5_F_masked1, //EXTERNAL
        output Tile_X6Y5_F_masked2, //EXTERNAL
        output Tile_X7Y5_F_masked1, //EXTERNAL
        output Tile_X7Y5_F_masked2, //EXTERNAL
        output Tile_X9Y5_F_ctrl, //EXTERNAL
        input Tile_X10Y5_A_O_top_0_t, //EXTERNAL
        input Tile_X10Y5_A_O_top_0_f, //EXTERNAL
        input Tile_X10Y5_A_prech2, //EXTERNAL
        input Tile_X10Y5_A_DR_fault, //EXTERNAL
        output Tile_X10Y5_A_I_top_0_t, //EXTERNAL
        output Tile_X10Y5_A_I_top_0_f, //EXTERNAL
        output Tile_X10Y5_A_T_top, //EXTERNAL
        output Tile_X10Y5_A_F_ctrl, //EXTERNAL
        input Tile_X0Y6_A_O_top_0_t, //EXTERNAL
        input Tile_X0Y6_A_O_top_0_f, //EXTERNAL
        input Tile_X0Y6_A_O_top_1_t, //EXTERNAL
        input Tile_X0Y6_A_O_top_1_f, //EXTERNAL
        input Tile_X0Y6_A_prech1, //EXTERNAL
        input Tile_X0Y6_A_prech2, //EXTERNAL
        input Tile_X0Y6_A_DR_fault, //EXTERNAL
        output Tile_X0Y6_A_I_top_0_t, //EXTERNAL
        output Tile_X0Y6_A_I_top_0_f, //EXTERNAL
        output Tile_X0Y6_A_I_top_1_t, //EXTERNAL
        output Tile_X0Y6_A_I_top_1_f, //EXTERNAL
        output Tile_X0Y6_A_T_top, //EXTERNAL
        output Tile_X0Y6_A_F_masked1, //EXTERNAL
        output Tile_X0Y6_A_F_masked2, //EXTERNAL
        output Tile_X0Y6_A_config_C_bit0, //EXTERNAL
        output Tile_X0Y6_A_config_C_bit1, //EXTERNAL
        output Tile_X0Y6_A_config_C_bit2, //EXTERNAL
        output Tile_X0Y6_A_config_C_bit3, //EXTERNAL
        output Tile_X0Y6_B_config_C_bit0, //EXTERNAL
        output Tile_X0Y6_B_config_C_bit1, //EXTERNAL
        output Tile_X0Y6_B_config_C_bit2, //EXTERNAL
        output Tile_X0Y6_B_config_C_bit3, //EXTERNAL
        output Tile_X1Y6_F_masked1, //EXTERNAL
        output Tile_X1Y6_F_masked2, //EXTERNAL
        output Tile_X2Y6_F_masked1, //EXTERNAL
        output Tile_X2Y6_F_masked2, //EXTERNAL
        input Tile_X3Y6_R_t, //EXTERNAL
        input Tile_X3Y6_R_f, //EXTERNAL
        output Tile_X3Y6_F_masked1, //EXTERNAL
        output Tile_X3Y6_F_masked2, //EXTERNAL
        output Tile_X4Y6_F_masked1, //EXTERNAL
        output Tile_X4Y6_F_masked2, //EXTERNAL
        output Tile_X5Y6_F_masked1, //EXTERNAL
        output Tile_X5Y6_F_masked2, //EXTERNAL
        input Tile_X6Y6_R_t, //EXTERNAL
        input Tile_X6Y6_R_f, //EXTERNAL
        output Tile_X6Y6_F_masked1, //EXTERNAL
        output Tile_X6Y6_F_masked2, //EXTERNAL
        output Tile_X7Y6_F_masked1, //EXTERNAL
        output Tile_X7Y6_F_masked2, //EXTERNAL
        output Tile_X9Y6_F_ctrl, //EXTERNAL
        input Tile_X10Y6_A_O_top_0_t, //EXTERNAL
        input Tile_X10Y6_A_O_top_0_f, //EXTERNAL
        input Tile_X10Y6_A_prech2, //EXTERNAL
        input Tile_X10Y6_A_DR_fault, //EXTERNAL
        output Tile_X10Y6_A_I_top_0_t, //EXTERNAL
        output Tile_X10Y6_A_I_top_0_f, //EXTERNAL
        output Tile_X10Y6_A_T_top, //EXTERNAL
        output Tile_X10Y6_A_F_ctrl, //EXTERNAL
        input Tile_X0Y7_A_O_top_0_t, //EXTERNAL
        input Tile_X0Y7_A_O_top_0_f, //EXTERNAL
        input Tile_X0Y7_A_O_top_1_t, //EXTERNAL
        input Tile_X0Y7_A_O_top_1_f, //EXTERNAL
        input Tile_X0Y7_A_prech1, //EXTERNAL
        input Tile_X0Y7_A_prech2, //EXTERNAL
        input Tile_X0Y7_A_DR_fault, //EXTERNAL
        output Tile_X0Y7_A_I_top_0_t, //EXTERNAL
        output Tile_X0Y7_A_I_top_0_f, //EXTERNAL
        output Tile_X0Y7_A_I_top_1_t, //EXTERNAL
        output Tile_X0Y7_A_I_top_1_f, //EXTERNAL
        output Tile_X0Y7_A_T_top, //EXTERNAL
        output Tile_X0Y7_A_F_masked1, //EXTERNAL
        output Tile_X0Y7_A_F_masked2, //EXTERNAL
        output Tile_X0Y7_A_config_C_bit0, //EXTERNAL
        output Tile_X0Y7_A_config_C_bit1, //EXTERNAL
        output Tile_X0Y7_A_config_C_bit2, //EXTERNAL
        output Tile_X0Y7_A_config_C_bit3, //EXTERNAL
        output Tile_X0Y7_B_config_C_bit0, //EXTERNAL
        output Tile_X0Y7_B_config_C_bit1, //EXTERNAL
        output Tile_X0Y7_B_config_C_bit2, //EXTERNAL
        output Tile_X0Y7_B_config_C_bit3, //EXTERNAL
        output Tile_X1Y7_F_masked1, //EXTERNAL
        output Tile_X1Y7_F_masked2, //EXTERNAL
        output Tile_X2Y7_F_masked1, //EXTERNAL
        output Tile_X2Y7_F_masked2, //EXTERNAL
        input Tile_X3Y7_R_t, //EXTERNAL
        input Tile_X3Y7_R_f, //EXTERNAL
        output Tile_X3Y7_F_masked1, //EXTERNAL
        output Tile_X3Y7_F_masked2, //EXTERNAL
        output Tile_X4Y7_F_masked1, //EXTERNAL
        output Tile_X4Y7_F_masked2, //EXTERNAL
        output Tile_X5Y7_F_masked1, //EXTERNAL
        output Tile_X5Y7_F_masked2, //EXTERNAL
        input Tile_X6Y7_R_t, //EXTERNAL
        input Tile_X6Y7_R_f, //EXTERNAL
        output Tile_X6Y7_F_masked1, //EXTERNAL
        output Tile_X6Y7_F_masked2, //EXTERNAL
        output Tile_X7Y7_F_masked1, //EXTERNAL
        output Tile_X7Y7_F_masked2, //EXTERNAL
        output Tile_X9Y7_F_ctrl, //EXTERNAL
        input Tile_X10Y7_A_O_top_0_t, //EXTERNAL
        input Tile_X10Y7_A_O_top_0_f, //EXTERNAL
        input Tile_X10Y7_A_prech2, //EXTERNAL
        input Tile_X10Y7_A_DR_fault, //EXTERNAL
        output Tile_X10Y7_A_I_top_0_t, //EXTERNAL
        output Tile_X10Y7_A_I_top_0_f, //EXTERNAL
        output Tile_X10Y7_A_T_top, //EXTERNAL
        output Tile_X10Y7_A_F_ctrl, //EXTERNAL
        input Tile_X0Y8_A_O_top_0_t, //EXTERNAL
        input Tile_X0Y8_A_O_top_0_f, //EXTERNAL
        input Tile_X0Y8_A_O_top_1_t, //EXTERNAL
        input Tile_X0Y8_A_O_top_1_f, //EXTERNAL
        input Tile_X0Y8_A_prech1, //EXTERNAL
        input Tile_X0Y8_A_prech2, //EXTERNAL
        input Tile_X0Y8_A_DR_fault, //EXTERNAL
        output Tile_X0Y8_A_I_top_0_t, //EXTERNAL
        output Tile_X0Y8_A_I_top_0_f, //EXTERNAL
        output Tile_X0Y8_A_I_top_1_t, //EXTERNAL
        output Tile_X0Y8_A_I_top_1_f, //EXTERNAL
        output Tile_X0Y8_A_T_top, //EXTERNAL
        output Tile_X0Y8_A_F_masked1, //EXTERNAL
        output Tile_X0Y8_A_F_masked2, //EXTERNAL
        output Tile_X0Y8_A_config_C_bit0, //EXTERNAL
        output Tile_X0Y8_A_config_C_bit1, //EXTERNAL
        output Tile_X0Y8_A_config_C_bit2, //EXTERNAL
        output Tile_X0Y8_A_config_C_bit3, //EXTERNAL
        output Tile_X0Y8_B_config_C_bit0, //EXTERNAL
        output Tile_X0Y8_B_config_C_bit1, //EXTERNAL
        output Tile_X0Y8_B_config_C_bit2, //EXTERNAL
        output Tile_X0Y8_B_config_C_bit3, //EXTERNAL
        output Tile_X1Y8_F_masked1, //EXTERNAL
        output Tile_X1Y8_F_masked2, //EXTERNAL
        output Tile_X2Y8_F_masked1, //EXTERNAL
        output Tile_X2Y8_F_masked2, //EXTERNAL
        input Tile_X3Y8_R_t, //EXTERNAL
        input Tile_X3Y8_R_f, //EXTERNAL
        output Tile_X3Y8_F_masked1, //EXTERNAL
        output Tile_X3Y8_F_masked2, //EXTERNAL
        output Tile_X4Y8_F_masked1, //EXTERNAL
        output Tile_X4Y8_F_masked2, //EXTERNAL
        output Tile_X5Y8_F_masked1, //EXTERNAL
        output Tile_X5Y8_F_masked2, //EXTERNAL
        input Tile_X6Y8_R_t, //EXTERNAL
        input Tile_X6Y8_R_f, //EXTERNAL
        output Tile_X6Y8_F_masked1, //EXTERNAL
        output Tile_X6Y8_F_masked2, //EXTERNAL
        output Tile_X7Y8_F_masked1, //EXTERNAL
        output Tile_X7Y8_F_masked2, //EXTERNAL
        output Tile_X9Y8_F_ctrl, //EXTERNAL
        input Tile_X10Y8_A_O_top_0_t, //EXTERNAL
        input Tile_X10Y8_A_O_top_0_f, //EXTERNAL
        input Tile_X10Y8_A_prech2, //EXTERNAL
        input Tile_X10Y8_A_DR_fault, //EXTERNAL
        output Tile_X10Y8_A_I_top_0_t, //EXTERNAL
        output Tile_X10Y8_A_I_top_0_f, //EXTERNAL
        output Tile_X10Y8_A_T_top, //EXTERNAL
        output Tile_X10Y8_A_F_ctrl, //EXTERNAL
        input Tile_X0Y9_A_O_top_0_t, //EXTERNAL
        input Tile_X0Y9_A_O_top_0_f, //EXTERNAL
        input Tile_X0Y9_A_O_top_1_t, //EXTERNAL
        input Tile_X0Y9_A_O_top_1_f, //EXTERNAL
        input Tile_X0Y9_A_prech1, //EXTERNAL
        input Tile_X0Y9_A_prech2, //EXTERNAL
        input Tile_X0Y9_A_DR_fault, //EXTERNAL
        output Tile_X0Y9_A_I_top_0_t, //EXTERNAL
        output Tile_X0Y9_A_I_top_0_f, //EXTERNAL
        output Tile_X0Y9_A_I_top_1_t, //EXTERNAL
        output Tile_X0Y9_A_I_top_1_f, //EXTERNAL
        output Tile_X0Y9_A_T_top, //EXTERNAL
        output Tile_X0Y9_A_F_masked1, //EXTERNAL
        output Tile_X0Y9_A_F_masked2, //EXTERNAL
        output Tile_X0Y9_A_config_C_bit0, //EXTERNAL
        output Tile_X0Y9_A_config_C_bit1, //EXTERNAL
        output Tile_X0Y9_A_config_C_bit2, //EXTERNAL
        output Tile_X0Y9_A_config_C_bit3, //EXTERNAL
        output Tile_X0Y9_B_config_C_bit0, //EXTERNAL
        output Tile_X0Y9_B_config_C_bit1, //EXTERNAL
        output Tile_X0Y9_B_config_C_bit2, //EXTERNAL
        output Tile_X0Y9_B_config_C_bit3, //EXTERNAL
        output Tile_X1Y9_F_masked1, //EXTERNAL
        output Tile_X1Y9_F_masked2, //EXTERNAL
        output Tile_X2Y9_F_masked1, //EXTERNAL
        output Tile_X2Y9_F_masked2, //EXTERNAL
        input Tile_X3Y9_R_t, //EXTERNAL
        input Tile_X3Y9_R_f, //EXTERNAL
        output Tile_X3Y9_F_masked1, //EXTERNAL
        output Tile_X3Y9_F_masked2, //EXTERNAL
        output Tile_X4Y9_F_masked1, //EXTERNAL
        output Tile_X4Y9_F_masked2, //EXTERNAL
        output Tile_X5Y9_F_masked1, //EXTERNAL
        output Tile_X5Y9_F_masked2, //EXTERNAL
        input Tile_X6Y9_R_t, //EXTERNAL
        input Tile_X6Y9_R_f, //EXTERNAL
        output Tile_X6Y9_F_masked1, //EXTERNAL
        output Tile_X6Y9_F_masked2, //EXTERNAL
        output Tile_X7Y9_F_masked1, //EXTERNAL
        output Tile_X7Y9_F_masked2, //EXTERNAL
        output Tile_X9Y9_F_ctrl, //EXTERNAL
        input Tile_X10Y9_A_O_top_0_t, //EXTERNAL
        input Tile_X10Y9_A_O_top_0_f, //EXTERNAL
        input Tile_X10Y9_A_prech2, //EXTERNAL
        input Tile_X10Y9_A_DR_fault, //EXTERNAL
        output Tile_X10Y9_A_I_top_0_t, //EXTERNAL
        output Tile_X10Y9_A_I_top_0_f, //EXTERNAL
        output Tile_X10Y9_A_T_top, //EXTERNAL
        output Tile_X10Y9_A_F_ctrl, //EXTERNAL
        input Tile_X0Y10_A_O_top_0_t, //EXTERNAL
        input Tile_X0Y10_A_O_top_0_f, //EXTERNAL
        input Tile_X0Y10_A_O_top_1_t, //EXTERNAL
        input Tile_X0Y10_A_O_top_1_f, //EXTERNAL
        input Tile_X0Y10_A_prech1, //EXTERNAL
        input Tile_X0Y10_A_prech2, //EXTERNAL
        input Tile_X0Y10_A_DR_fault, //EXTERNAL
        output Tile_X0Y10_A_I_top_0_t, //EXTERNAL
        output Tile_X0Y10_A_I_top_0_f, //EXTERNAL
        output Tile_X0Y10_A_I_top_1_t, //EXTERNAL
        output Tile_X0Y10_A_I_top_1_f, //EXTERNAL
        output Tile_X0Y10_A_T_top, //EXTERNAL
        output Tile_X0Y10_A_F_masked1, //EXTERNAL
        output Tile_X0Y10_A_F_masked2, //EXTERNAL
        output Tile_X0Y10_A_config_C_bit0, //EXTERNAL
        output Tile_X0Y10_A_config_C_bit1, //EXTERNAL
        output Tile_X0Y10_A_config_C_bit2, //EXTERNAL
        output Tile_X0Y10_A_config_C_bit3, //EXTERNAL
        output Tile_X0Y10_B_config_C_bit0, //EXTERNAL
        output Tile_X0Y10_B_config_C_bit1, //EXTERNAL
        output Tile_X0Y10_B_config_C_bit2, //EXTERNAL
        output Tile_X0Y10_B_config_C_bit3, //EXTERNAL
        output Tile_X1Y10_F_masked1, //EXTERNAL
        output Tile_X1Y10_F_masked2, //EXTERNAL
        output Tile_X2Y10_F_masked1, //EXTERNAL
        output Tile_X2Y10_F_masked2, //EXTERNAL
        input Tile_X3Y10_R_t, //EXTERNAL
        input Tile_X3Y10_R_f, //EXTERNAL
        output Tile_X3Y10_F_masked1, //EXTERNAL
        output Tile_X3Y10_F_masked2, //EXTERNAL
        output Tile_X4Y10_F_masked1, //EXTERNAL
        output Tile_X4Y10_F_masked2, //EXTERNAL
        output Tile_X5Y10_F_masked1, //EXTERNAL
        output Tile_X5Y10_F_masked2, //EXTERNAL
        input Tile_X6Y10_R_t, //EXTERNAL
        input Tile_X6Y10_R_f, //EXTERNAL
        output Tile_X6Y10_F_masked1, //EXTERNAL
        output Tile_X6Y10_F_masked2, //EXTERNAL
        output Tile_X7Y10_F_masked1, //EXTERNAL
        output Tile_X7Y10_F_masked2, //EXTERNAL
        output Tile_X9Y10_F_ctrl, //EXTERNAL
        input Tile_X10Y10_A_O_top_0_t, //EXTERNAL
        input Tile_X10Y10_A_O_top_0_f, //EXTERNAL
        input Tile_X10Y10_A_prech2, //EXTERNAL
        input Tile_X10Y10_A_DR_fault, //EXTERNAL
        output Tile_X10Y10_A_I_top_0_t, //EXTERNAL
        output Tile_X10Y10_A_I_top_0_f, //EXTERNAL
        output Tile_X10Y10_A_T_top, //EXTERNAL
        output Tile_X10Y10_A_F_ctrl, //EXTERNAL
        input Tile_X0Y11_A_O_top_0_t, //EXTERNAL
        input Tile_X0Y11_A_O_top_0_f, //EXTERNAL
        input Tile_X0Y11_A_O_top_1_t, //EXTERNAL
        input Tile_X0Y11_A_O_top_1_f, //EXTERNAL
        input Tile_X0Y11_A_prech1, //EXTERNAL
        input Tile_X0Y11_A_prech2, //EXTERNAL
        input Tile_X0Y11_A_DR_fault, //EXTERNAL
        output Tile_X0Y11_A_I_top_0_t, //EXTERNAL
        output Tile_X0Y11_A_I_top_0_f, //EXTERNAL
        output Tile_X0Y11_A_I_top_1_t, //EXTERNAL
        output Tile_X0Y11_A_I_top_1_f, //EXTERNAL
        output Tile_X0Y11_A_T_top, //EXTERNAL
        output Tile_X0Y11_A_F_masked1, //EXTERNAL
        output Tile_X0Y11_A_F_masked2, //EXTERNAL
        output Tile_X0Y11_A_config_C_bit0, //EXTERNAL
        output Tile_X0Y11_A_config_C_bit1, //EXTERNAL
        output Tile_X0Y11_A_config_C_bit2, //EXTERNAL
        output Tile_X0Y11_A_config_C_bit3, //EXTERNAL
        output Tile_X0Y11_B_config_C_bit0, //EXTERNAL
        output Tile_X0Y11_B_config_C_bit1, //EXTERNAL
        output Tile_X0Y11_B_config_C_bit2, //EXTERNAL
        output Tile_X0Y11_B_config_C_bit3, //EXTERNAL
        output Tile_X1Y11_F_masked1, //EXTERNAL
        output Tile_X1Y11_F_masked2, //EXTERNAL
        output Tile_X2Y11_F_masked1, //EXTERNAL
        output Tile_X2Y11_F_masked2, //EXTERNAL
        input Tile_X3Y11_R_t, //EXTERNAL
        input Tile_X3Y11_R_f, //EXTERNAL
        output Tile_X3Y11_F_masked1, //EXTERNAL
        output Tile_X3Y11_F_masked2, //EXTERNAL
        output Tile_X4Y11_F_masked1, //EXTERNAL
        output Tile_X4Y11_F_masked2, //EXTERNAL
        output Tile_X5Y11_F_masked1, //EXTERNAL
        output Tile_X5Y11_F_masked2, //EXTERNAL
        input Tile_X6Y11_R_t, //EXTERNAL
        input Tile_X6Y11_R_f, //EXTERNAL
        output Tile_X6Y11_F_masked1, //EXTERNAL
        output Tile_X6Y11_F_masked2, //EXTERNAL
        output Tile_X7Y11_F_masked1, //EXTERNAL
        output Tile_X7Y11_F_masked2, //EXTERNAL
        output Tile_X9Y11_F_ctrl, //EXTERNAL
        input Tile_X10Y11_A_O_top_0_t, //EXTERNAL
        input Tile_X10Y11_A_O_top_0_f, //EXTERNAL
        input Tile_X10Y11_A_prech2, //EXTERNAL
        input Tile_X10Y11_A_DR_fault, //EXTERNAL
        output Tile_X10Y11_A_I_top_0_t, //EXTERNAL
        output Tile_X10Y11_A_I_top_0_f, //EXTERNAL
        output Tile_X10Y11_A_T_top, //EXTERNAL
        output Tile_X10Y11_A_F_ctrl, //EXTERNAL
        input Tile_X0Y12_A_O_top_0_t, //EXTERNAL
        input Tile_X0Y12_A_O_top_0_f, //EXTERNAL
        input Tile_X0Y12_A_O_top_1_t, //EXTERNAL
        input Tile_X0Y12_A_O_top_1_f, //EXTERNAL
        input Tile_X0Y12_A_prech1, //EXTERNAL
        input Tile_X0Y12_A_prech2, //EXTERNAL
        input Tile_X0Y12_A_DR_fault, //EXTERNAL
        output Tile_X0Y12_A_I_top_0_t, //EXTERNAL
        output Tile_X0Y12_A_I_top_0_f, //EXTERNAL
        output Tile_X0Y12_A_I_top_1_t, //EXTERNAL
        output Tile_X0Y12_A_I_top_1_f, //EXTERNAL
        output Tile_X0Y12_A_T_top, //EXTERNAL
        output Tile_X0Y12_A_F_masked1, //EXTERNAL
        output Tile_X0Y12_A_F_masked2, //EXTERNAL
        output Tile_X0Y12_A_config_C_bit0, //EXTERNAL
        output Tile_X0Y12_A_config_C_bit1, //EXTERNAL
        output Tile_X0Y12_A_config_C_bit2, //EXTERNAL
        output Tile_X0Y12_A_config_C_bit3, //EXTERNAL
        output Tile_X0Y12_B_config_C_bit0, //EXTERNAL
        output Tile_X0Y12_B_config_C_bit1, //EXTERNAL
        output Tile_X0Y12_B_config_C_bit2, //EXTERNAL
        output Tile_X0Y12_B_config_C_bit3, //EXTERNAL
        output Tile_X1Y12_F_masked1, //EXTERNAL
        output Tile_X1Y12_F_masked2, //EXTERNAL
        output Tile_X2Y12_F_masked1, //EXTERNAL
        output Tile_X2Y12_F_masked2, //EXTERNAL
        input Tile_X3Y12_R_t, //EXTERNAL
        input Tile_X3Y12_R_f, //EXTERNAL
        output Tile_X3Y12_F_masked1, //EXTERNAL
        output Tile_X3Y12_F_masked2, //EXTERNAL
        output Tile_X4Y12_F_masked1, //EXTERNAL
        output Tile_X4Y12_F_masked2, //EXTERNAL
        output Tile_X5Y12_F_masked1, //EXTERNAL
        output Tile_X5Y12_F_masked2, //EXTERNAL
        input Tile_X6Y12_R_t, //EXTERNAL
        input Tile_X6Y12_R_f, //EXTERNAL
        output Tile_X6Y12_F_masked1, //EXTERNAL
        output Tile_X6Y12_F_masked2, //EXTERNAL
        output Tile_X7Y12_F_masked1, //EXTERNAL
        output Tile_X7Y12_F_masked2, //EXTERNAL
        output Tile_X9Y12_F_ctrl, //EXTERNAL
        input Tile_X10Y12_A_O_top_0_t, //EXTERNAL
        input Tile_X10Y12_A_O_top_0_f, //EXTERNAL
        input Tile_X10Y12_A_prech2, //EXTERNAL
        input Tile_X10Y12_A_DR_fault, //EXTERNAL
        output Tile_X10Y12_A_I_top_0_t, //EXTERNAL
        output Tile_X10Y12_A_I_top_0_f, //EXTERNAL
        output Tile_X10Y12_A_T_top, //EXTERNAL
        output Tile_X10Y12_A_F_ctrl, //EXTERNAL
        input Tile_X0Y13_A_O_top_0_t, //EXTERNAL
        input Tile_X0Y13_A_O_top_0_f, //EXTERNAL
        input Tile_X0Y13_A_O_top_1_t, //EXTERNAL
        input Tile_X0Y13_A_O_top_1_f, //EXTERNAL
        input Tile_X0Y13_A_prech1, //EXTERNAL
        input Tile_X0Y13_A_prech2, //EXTERNAL
        input Tile_X0Y13_A_DR_fault, //EXTERNAL
        output Tile_X0Y13_A_I_top_0_t, //EXTERNAL
        output Tile_X0Y13_A_I_top_0_f, //EXTERNAL
        output Tile_X0Y13_A_I_top_1_t, //EXTERNAL
        output Tile_X0Y13_A_I_top_1_f, //EXTERNAL
        output Tile_X0Y13_A_T_top, //EXTERNAL
        output Tile_X0Y13_A_F_masked1, //EXTERNAL
        output Tile_X0Y13_A_F_masked2, //EXTERNAL
        output Tile_X0Y13_A_config_C_bit0, //EXTERNAL
        output Tile_X0Y13_A_config_C_bit1, //EXTERNAL
        output Tile_X0Y13_A_config_C_bit2, //EXTERNAL
        output Tile_X0Y13_A_config_C_bit3, //EXTERNAL
        output Tile_X0Y13_B_config_C_bit0, //EXTERNAL
        output Tile_X0Y13_B_config_C_bit1, //EXTERNAL
        output Tile_X0Y13_B_config_C_bit2, //EXTERNAL
        output Tile_X0Y13_B_config_C_bit3, //EXTERNAL
        output Tile_X1Y13_F_masked1, //EXTERNAL
        output Tile_X1Y13_F_masked2, //EXTERNAL
        output Tile_X2Y13_F_masked1, //EXTERNAL
        output Tile_X2Y13_F_masked2, //EXTERNAL
        input Tile_X3Y13_R_t, //EXTERNAL
        input Tile_X3Y13_R_f, //EXTERNAL
        output Tile_X3Y13_F_masked1, //EXTERNAL
        output Tile_X3Y13_F_masked2, //EXTERNAL
        output Tile_X4Y13_F_masked1, //EXTERNAL
        output Tile_X4Y13_F_masked2, //EXTERNAL
        output Tile_X5Y13_F_masked1, //EXTERNAL
        output Tile_X5Y13_F_masked2, //EXTERNAL
        input Tile_X6Y13_R_t, //EXTERNAL
        input Tile_X6Y13_R_f, //EXTERNAL
        output Tile_X6Y13_F_masked1, //EXTERNAL
        output Tile_X6Y13_F_masked2, //EXTERNAL
        output Tile_X7Y13_F_masked1, //EXTERNAL
        output Tile_X7Y13_F_masked2, //EXTERNAL
        output Tile_X9Y13_F_ctrl, //EXTERNAL
        input Tile_X10Y13_A_O_top_0_t, //EXTERNAL
        input Tile_X10Y13_A_O_top_0_f, //EXTERNAL
        input Tile_X10Y13_A_prech2, //EXTERNAL
        input Tile_X10Y13_A_DR_fault, //EXTERNAL
        output Tile_X10Y13_A_I_top_0_t, //EXTERNAL
        output Tile_X10Y13_A_I_top_0_f, //EXTERNAL
        output Tile_X10Y13_A_T_top, //EXTERNAL
        output Tile_X10Y13_A_F_ctrl, //EXTERNAL
        input Tile_X0Y14_A_O_top_0_t, //EXTERNAL
        input Tile_X0Y14_A_O_top_0_f, //EXTERNAL
        input Tile_X0Y14_A_O_top_1_t, //EXTERNAL
        input Tile_X0Y14_A_O_top_1_f, //EXTERNAL
        input Tile_X0Y14_A_prech1, //EXTERNAL
        input Tile_X0Y14_A_prech2, //EXTERNAL
        input Tile_X0Y14_A_DR_fault, //EXTERNAL
        output Tile_X0Y14_A_I_top_0_t, //EXTERNAL
        output Tile_X0Y14_A_I_top_0_f, //EXTERNAL
        output Tile_X0Y14_A_I_top_1_t, //EXTERNAL
        output Tile_X0Y14_A_I_top_1_f, //EXTERNAL
        output Tile_X0Y14_A_T_top, //EXTERNAL
        output Tile_X0Y14_A_F_masked1, //EXTERNAL
        output Tile_X0Y14_A_F_masked2, //EXTERNAL
        output Tile_X0Y14_A_config_C_bit0, //EXTERNAL
        output Tile_X0Y14_A_config_C_bit1, //EXTERNAL
        output Tile_X0Y14_A_config_C_bit2, //EXTERNAL
        output Tile_X0Y14_A_config_C_bit3, //EXTERNAL
        output Tile_X0Y14_B_config_C_bit0, //EXTERNAL
        output Tile_X0Y14_B_config_C_bit1, //EXTERNAL
        output Tile_X0Y14_B_config_C_bit2, //EXTERNAL
        output Tile_X0Y14_B_config_C_bit3, //EXTERNAL
        output Tile_X1Y14_F_masked1, //EXTERNAL
        output Tile_X1Y14_F_masked2, //EXTERNAL
        output Tile_X2Y14_F_masked1, //EXTERNAL
        output Tile_X2Y14_F_masked2, //EXTERNAL
        input Tile_X3Y14_R_t, //EXTERNAL
        input Tile_X3Y14_R_f, //EXTERNAL
        output Tile_X3Y14_F_masked1, //EXTERNAL
        output Tile_X3Y14_F_masked2, //EXTERNAL
        output Tile_X4Y14_F_masked1, //EXTERNAL
        output Tile_X4Y14_F_masked2, //EXTERNAL
        output Tile_X5Y14_F_masked1, //EXTERNAL
        output Tile_X5Y14_F_masked2, //EXTERNAL
        input Tile_X6Y14_R_t, //EXTERNAL
        input Tile_X6Y14_R_f, //EXTERNAL
        output Tile_X6Y14_F_masked1, //EXTERNAL
        output Tile_X6Y14_F_masked2, //EXTERNAL
        output Tile_X7Y14_F_masked1, //EXTERNAL
        output Tile_X7Y14_F_masked2, //EXTERNAL
        output Tile_X9Y14_F_ctrl, //EXTERNAL
        input Tile_X10Y14_A_O_top_0_t, //EXTERNAL
        input Tile_X10Y14_A_O_top_0_f, //EXTERNAL
        input Tile_X10Y14_A_prech2, //EXTERNAL
        input Tile_X10Y14_A_DR_fault, //EXTERNAL
        output Tile_X10Y14_A_I_top_0_t, //EXTERNAL
        output Tile_X10Y14_A_I_top_0_f, //EXTERNAL
        output Tile_X10Y14_A_T_top, //EXTERNAL
        output Tile_X10Y14_A_F_ctrl, //EXTERNAL
        input Tile_X0Y15_A_O_top_0_t, //EXTERNAL
        input Tile_X0Y15_A_O_top_0_f, //EXTERNAL
        input Tile_X0Y15_A_O_top_1_t, //EXTERNAL
        input Tile_X0Y15_A_O_top_1_f, //EXTERNAL
        input Tile_X0Y15_A_prech1, //EXTERNAL
        input Tile_X0Y15_A_prech2, //EXTERNAL
        input Tile_X0Y15_A_DR_fault, //EXTERNAL
        output Tile_X0Y15_A_I_top_0_t, //EXTERNAL
        output Tile_X0Y15_A_I_top_0_f, //EXTERNAL
        output Tile_X0Y15_A_I_top_1_t, //EXTERNAL
        output Tile_X0Y15_A_I_top_1_f, //EXTERNAL
        output Tile_X0Y15_A_T_top, //EXTERNAL
        output Tile_X0Y15_A_F_masked1, //EXTERNAL
        output Tile_X0Y15_A_F_masked2, //EXTERNAL
        output Tile_X0Y15_A_config_C_bit0, //EXTERNAL
        output Tile_X0Y15_A_config_C_bit1, //EXTERNAL
        output Tile_X0Y15_A_config_C_bit2, //EXTERNAL
        output Tile_X0Y15_A_config_C_bit3, //EXTERNAL
        output Tile_X0Y15_B_config_C_bit0, //EXTERNAL
        output Tile_X0Y15_B_config_C_bit1, //EXTERNAL
        output Tile_X0Y15_B_config_C_bit2, //EXTERNAL
        output Tile_X0Y15_B_config_C_bit3, //EXTERNAL
        output Tile_X1Y15_F_masked1, //EXTERNAL
        output Tile_X1Y15_F_masked2, //EXTERNAL
        output Tile_X2Y15_F_masked1, //EXTERNAL
        output Tile_X2Y15_F_masked2, //EXTERNAL
        input Tile_X3Y15_R_t, //EXTERNAL
        input Tile_X3Y15_R_f, //EXTERNAL
        output Tile_X3Y15_F_masked1, //EXTERNAL
        output Tile_X3Y15_F_masked2, //EXTERNAL
        output Tile_X4Y15_F_masked1, //EXTERNAL
        output Tile_X4Y15_F_masked2, //EXTERNAL
        output Tile_X5Y15_F_masked1, //EXTERNAL
        output Tile_X5Y15_F_masked2, //EXTERNAL
        input Tile_X6Y15_R_t, //EXTERNAL
        input Tile_X6Y15_R_f, //EXTERNAL
        output Tile_X6Y15_F_masked1, //EXTERNAL
        output Tile_X6Y15_F_masked2, //EXTERNAL
        output Tile_X7Y15_F_masked1, //EXTERNAL
        output Tile_X7Y15_F_masked2, //EXTERNAL
        output Tile_X9Y15_F_ctrl, //EXTERNAL
        input Tile_X10Y15_A_O_top_0_t, //EXTERNAL
        input Tile_X10Y15_A_O_top_0_f, //EXTERNAL
        input Tile_X10Y15_A_prech2, //EXTERNAL
        input Tile_X10Y15_A_DR_fault, //EXTERNAL
        output Tile_X10Y15_A_I_top_0_t, //EXTERNAL
        output Tile_X10Y15_A_I_top_0_f, //EXTERNAL
        output Tile_X10Y15_A_T_top, //EXTERNAL
        output Tile_X10Y15_A_F_ctrl, //EXTERNAL
        input Tile_X0Y16_A_O_top_0_t, //EXTERNAL
        input Tile_X0Y16_A_O_top_0_f, //EXTERNAL
        input Tile_X0Y16_A_O_top_1_t, //EXTERNAL
        input Tile_X0Y16_A_O_top_1_f, //EXTERNAL
        input Tile_X0Y16_A_prech1, //EXTERNAL
        input Tile_X0Y16_A_prech2, //EXTERNAL
        input Tile_X0Y16_A_DR_fault, //EXTERNAL
        output Tile_X0Y16_A_I_top_0_t, //EXTERNAL
        output Tile_X0Y16_A_I_top_0_f, //EXTERNAL
        output Tile_X0Y16_A_I_top_1_t, //EXTERNAL
        output Tile_X0Y16_A_I_top_1_f, //EXTERNAL
        output Tile_X0Y16_A_T_top, //EXTERNAL
        output Tile_X0Y16_A_F_masked1, //EXTERNAL
        output Tile_X0Y16_A_F_masked2, //EXTERNAL
        output Tile_X0Y16_A_config_C_bit0, //EXTERNAL
        output Tile_X0Y16_A_config_C_bit1, //EXTERNAL
        output Tile_X0Y16_A_config_C_bit2, //EXTERNAL
        output Tile_X0Y16_A_config_C_bit3, //EXTERNAL
        output Tile_X0Y16_B_config_C_bit0, //EXTERNAL
        output Tile_X0Y16_B_config_C_bit1, //EXTERNAL
        output Tile_X0Y16_B_config_C_bit2, //EXTERNAL
        output Tile_X0Y16_B_config_C_bit3, //EXTERNAL
        output Tile_X1Y16_F_masked1, //EXTERNAL
        output Tile_X1Y16_F_masked2, //EXTERNAL
        output Tile_X2Y16_F_masked1, //EXTERNAL
        output Tile_X2Y16_F_masked2, //EXTERNAL
        input Tile_X3Y16_R_t, //EXTERNAL
        input Tile_X3Y16_R_f, //EXTERNAL
        output Tile_X3Y16_F_masked1, //EXTERNAL
        output Tile_X3Y16_F_masked2, //EXTERNAL
        output Tile_X4Y16_F_masked1, //EXTERNAL
        output Tile_X4Y16_F_masked2, //EXTERNAL
        output Tile_X5Y16_F_masked1, //EXTERNAL
        output Tile_X5Y16_F_masked2, //EXTERNAL
        input Tile_X6Y16_R_t, //EXTERNAL
        input Tile_X6Y16_R_f, //EXTERNAL
        output Tile_X6Y16_F_masked1, //EXTERNAL
        output Tile_X6Y16_F_masked2, //EXTERNAL
        output Tile_X7Y16_F_masked1, //EXTERNAL
        output Tile_X7Y16_F_masked2, //EXTERNAL
        output Tile_X9Y16_F_ctrl, //EXTERNAL
        input Tile_X10Y16_A_O_top_0_t, //EXTERNAL
        input Tile_X10Y16_A_O_top_0_f, //EXTERNAL
        input Tile_X10Y16_A_prech2, //EXTERNAL
        input Tile_X10Y16_A_DR_fault, //EXTERNAL
        output Tile_X10Y16_A_I_top_0_t, //EXTERNAL
        output Tile_X10Y16_A_I_top_0_f, //EXTERNAL
        output Tile_X10Y16_A_T_top, //EXTERNAL
        output Tile_X10Y16_A_F_ctrl, //EXTERNAL
        input Tile_X0Y17_A_O_top_0_t, //EXTERNAL
        input Tile_X0Y17_A_O_top_0_f, //EXTERNAL
        input Tile_X0Y17_A_O_top_1_t, //EXTERNAL
        input Tile_X0Y17_A_O_top_1_f, //EXTERNAL
        input Tile_X0Y17_A_prech1, //EXTERNAL
        input Tile_X0Y17_A_prech2, //EXTERNAL
        input Tile_X0Y17_A_DR_fault, //EXTERNAL
        output Tile_X0Y17_A_I_top_0_t, //EXTERNAL
        output Tile_X0Y17_A_I_top_0_f, //EXTERNAL
        output Tile_X0Y17_A_I_top_1_t, //EXTERNAL
        output Tile_X0Y17_A_I_top_1_f, //EXTERNAL
        output Tile_X0Y17_A_T_top, //EXTERNAL
        output Tile_X0Y17_A_F_masked1, //EXTERNAL
        output Tile_X0Y17_A_F_masked2, //EXTERNAL
        output Tile_X0Y17_A_config_C_bit0, //EXTERNAL
        output Tile_X0Y17_A_config_C_bit1, //EXTERNAL
        output Tile_X0Y17_A_config_C_bit2, //EXTERNAL
        output Tile_X0Y17_A_config_C_bit3, //EXTERNAL
        output Tile_X0Y17_B_config_C_bit0, //EXTERNAL
        output Tile_X0Y17_B_config_C_bit1, //EXTERNAL
        output Tile_X0Y17_B_config_C_bit2, //EXTERNAL
        output Tile_X0Y17_B_config_C_bit3, //EXTERNAL
        output Tile_X1Y17_F_masked1, //EXTERNAL
        output Tile_X1Y17_F_masked2, //EXTERNAL
        output Tile_X2Y17_F_masked1, //EXTERNAL
        output Tile_X2Y17_F_masked2, //EXTERNAL
        input Tile_X3Y17_R_t, //EXTERNAL
        input Tile_X3Y17_R_f, //EXTERNAL
        output Tile_X3Y17_F_masked1, //EXTERNAL
        output Tile_X3Y17_F_masked2, //EXTERNAL
        output Tile_X4Y17_F_masked1, //EXTERNAL
        output Tile_X4Y17_F_masked2, //EXTERNAL
        output Tile_X5Y17_F_masked1, //EXTERNAL
        output Tile_X5Y17_F_masked2, //EXTERNAL
        input Tile_X6Y17_R_t, //EXTERNAL
        input Tile_X6Y17_R_f, //EXTERNAL
        output Tile_X6Y17_F_masked1, //EXTERNAL
        output Tile_X6Y17_F_masked2, //EXTERNAL
        output Tile_X7Y17_F_masked1, //EXTERNAL
        output Tile_X7Y17_F_masked2, //EXTERNAL
        output Tile_X9Y17_F_ctrl, //EXTERNAL
        input Tile_X10Y17_A_O_top_0_t, //EXTERNAL
        input Tile_X10Y17_A_O_top_0_f, //EXTERNAL
        input Tile_X10Y17_A_prech2, //EXTERNAL
        input Tile_X10Y17_A_DR_fault, //EXTERNAL
        output Tile_X10Y17_A_I_top_0_t, //EXTERNAL
        output Tile_X10Y17_A_I_top_0_f, //EXTERNAL
        output Tile_X10Y17_A_T_top, //EXTERNAL
        output Tile_X10Y17_A_F_ctrl, //EXTERNAL
        input Tile_X0Y18_A_O_top_0_t, //EXTERNAL
        input Tile_X0Y18_A_O_top_0_f, //EXTERNAL
        input Tile_X0Y18_A_O_top_1_t, //EXTERNAL
        input Tile_X0Y18_A_O_top_1_f, //EXTERNAL
        input Tile_X0Y18_A_prech1, //EXTERNAL
        input Tile_X0Y18_A_prech2, //EXTERNAL
        input Tile_X0Y18_A_DR_fault, //EXTERNAL
        output Tile_X0Y18_A_I_top_0_t, //EXTERNAL
        output Tile_X0Y18_A_I_top_0_f, //EXTERNAL
        output Tile_X0Y18_A_I_top_1_t, //EXTERNAL
        output Tile_X0Y18_A_I_top_1_f, //EXTERNAL
        output Tile_X0Y18_A_T_top, //EXTERNAL
        output Tile_X0Y18_A_F_masked1, //EXTERNAL
        output Tile_X0Y18_A_F_masked2, //EXTERNAL
        output Tile_X0Y18_A_config_C_bit0, //EXTERNAL
        output Tile_X0Y18_A_config_C_bit1, //EXTERNAL
        output Tile_X0Y18_A_config_C_bit2, //EXTERNAL
        output Tile_X0Y18_A_config_C_bit3, //EXTERNAL
        output Tile_X0Y18_B_config_C_bit0, //EXTERNAL
        output Tile_X0Y18_B_config_C_bit1, //EXTERNAL
        output Tile_X0Y18_B_config_C_bit2, //EXTERNAL
        output Tile_X0Y18_B_config_C_bit3, //EXTERNAL
        output Tile_X1Y18_F_masked1, //EXTERNAL
        output Tile_X1Y18_F_masked2, //EXTERNAL
        output Tile_X2Y18_F_masked1, //EXTERNAL
        output Tile_X2Y18_F_masked2, //EXTERNAL
        input Tile_X3Y18_R_t, //EXTERNAL
        input Tile_X3Y18_R_f, //EXTERNAL
        output Tile_X3Y18_F_masked1, //EXTERNAL
        output Tile_X3Y18_F_masked2, //EXTERNAL
        output Tile_X4Y18_F_masked1, //EXTERNAL
        output Tile_X4Y18_F_masked2, //EXTERNAL
        output Tile_X5Y18_F_masked1, //EXTERNAL
        output Tile_X5Y18_F_masked2, //EXTERNAL
        input Tile_X6Y18_R_t, //EXTERNAL
        input Tile_X6Y18_R_f, //EXTERNAL
        output Tile_X6Y18_F_masked1, //EXTERNAL
        output Tile_X6Y18_F_masked2, //EXTERNAL
        output Tile_X7Y18_F_masked1, //EXTERNAL
        output Tile_X7Y18_F_masked2, //EXTERNAL
        output Tile_X9Y18_F_ctrl, //EXTERNAL
        input Tile_X10Y18_A_O_top_0_t, //EXTERNAL
        input Tile_X10Y18_A_O_top_0_f, //EXTERNAL
        input Tile_X10Y18_A_prech2, //EXTERNAL
        input Tile_X10Y18_A_DR_fault, //EXTERNAL
        output Tile_X10Y18_A_I_top_0_t, //EXTERNAL
        output Tile_X10Y18_A_I_top_0_f, //EXTERNAL
        output Tile_X10Y18_A_T_top, //EXTERNAL
        output Tile_X10Y18_A_F_ctrl, //EXTERNAL
        input Tile_X0Y19_A_O_top_0_t, //EXTERNAL
        input Tile_X0Y19_A_O_top_0_f, //EXTERNAL
        input Tile_X0Y19_A_O_top_1_t, //EXTERNAL
        input Tile_X0Y19_A_O_top_1_f, //EXTERNAL
        input Tile_X0Y19_A_prech1, //EXTERNAL
        input Tile_X0Y19_A_prech2, //EXTERNAL
        input Tile_X0Y19_A_DR_fault, //EXTERNAL
        output Tile_X0Y19_A_I_top_0_t, //EXTERNAL
        output Tile_X0Y19_A_I_top_0_f, //EXTERNAL
        output Tile_X0Y19_A_I_top_1_t, //EXTERNAL
        output Tile_X0Y19_A_I_top_1_f, //EXTERNAL
        output Tile_X0Y19_A_T_top, //EXTERNAL
        output Tile_X0Y19_A_F_masked1, //EXTERNAL
        output Tile_X0Y19_A_F_masked2, //EXTERNAL
        output Tile_X0Y19_A_config_C_bit0, //EXTERNAL
        output Tile_X0Y19_A_config_C_bit1, //EXTERNAL
        output Tile_X0Y19_A_config_C_bit2, //EXTERNAL
        output Tile_X0Y19_A_config_C_bit3, //EXTERNAL
        output Tile_X0Y19_B_config_C_bit0, //EXTERNAL
        output Tile_X0Y19_B_config_C_bit1, //EXTERNAL
        output Tile_X0Y19_B_config_C_bit2, //EXTERNAL
        output Tile_X0Y19_B_config_C_bit3, //EXTERNAL
        output Tile_X1Y19_F_masked1, //EXTERNAL
        output Tile_X1Y19_F_masked2, //EXTERNAL
        output Tile_X2Y19_F_masked1, //EXTERNAL
        output Tile_X2Y19_F_masked2, //EXTERNAL
        input Tile_X3Y19_R_t, //EXTERNAL
        input Tile_X3Y19_R_f, //EXTERNAL
        output Tile_X3Y19_F_masked1, //EXTERNAL
        output Tile_X3Y19_F_masked2, //EXTERNAL
        output Tile_X4Y19_F_masked1, //EXTERNAL
        output Tile_X4Y19_F_masked2, //EXTERNAL
        output Tile_X5Y19_F_masked1, //EXTERNAL
        output Tile_X5Y19_F_masked2, //EXTERNAL
        input Tile_X6Y19_R_t, //EXTERNAL
        input Tile_X6Y19_R_f, //EXTERNAL
        output Tile_X6Y19_F_masked1, //EXTERNAL
        output Tile_X6Y19_F_masked2, //EXTERNAL
        output Tile_X7Y19_F_masked1, //EXTERNAL
        output Tile_X7Y19_F_masked2, //EXTERNAL
        output Tile_X9Y19_F_ctrl, //EXTERNAL
        input Tile_X10Y19_A_O_top_0_t, //EXTERNAL
        input Tile_X10Y19_A_O_top_0_f, //EXTERNAL
        input Tile_X10Y19_A_prech2, //EXTERNAL
        input Tile_X10Y19_A_DR_fault, //EXTERNAL
        output Tile_X10Y19_A_I_top_0_t, //EXTERNAL
        output Tile_X10Y19_A_I_top_0_f, //EXTERNAL
        output Tile_X10Y19_A_T_top, //EXTERNAL
        output Tile_X10Y19_A_F_ctrl, //EXTERNAL
        input Tile_X0Y20_A_O_top_0_t, //EXTERNAL
        input Tile_X0Y20_A_O_top_0_f, //EXTERNAL
        input Tile_X0Y20_A_O_top_1_t, //EXTERNAL
        input Tile_X0Y20_A_O_top_1_f, //EXTERNAL
        input Tile_X0Y20_A_prech1, //EXTERNAL
        input Tile_X0Y20_A_prech2, //EXTERNAL
        input Tile_X0Y20_A_DR_fault, //EXTERNAL
        output Tile_X0Y20_A_I_top_0_t, //EXTERNAL
        output Tile_X0Y20_A_I_top_0_f, //EXTERNAL
        output Tile_X0Y20_A_I_top_1_t, //EXTERNAL
        output Tile_X0Y20_A_I_top_1_f, //EXTERNAL
        output Tile_X0Y20_A_T_top, //EXTERNAL
        output Tile_X0Y20_A_F_masked1, //EXTERNAL
        output Tile_X0Y20_A_F_masked2, //EXTERNAL
        output Tile_X0Y20_A_config_C_bit0, //EXTERNAL
        output Tile_X0Y20_A_config_C_bit1, //EXTERNAL
        output Tile_X0Y20_A_config_C_bit2, //EXTERNAL
        output Tile_X0Y20_A_config_C_bit3, //EXTERNAL
        output Tile_X0Y20_B_config_C_bit0, //EXTERNAL
        output Tile_X0Y20_B_config_C_bit1, //EXTERNAL
        output Tile_X0Y20_B_config_C_bit2, //EXTERNAL
        output Tile_X0Y20_B_config_C_bit3, //EXTERNAL
        output Tile_X1Y20_F_masked1, //EXTERNAL
        output Tile_X1Y20_F_masked2, //EXTERNAL
        output Tile_X2Y20_F_masked1, //EXTERNAL
        output Tile_X2Y20_F_masked2, //EXTERNAL
        input Tile_X3Y20_R_t, //EXTERNAL
        input Tile_X3Y20_R_f, //EXTERNAL
        output Tile_X3Y20_F_masked1, //EXTERNAL
        output Tile_X3Y20_F_masked2, //EXTERNAL
        output Tile_X4Y20_F_masked1, //EXTERNAL
        output Tile_X4Y20_F_masked2, //EXTERNAL
        output Tile_X5Y20_F_masked1, //EXTERNAL
        output Tile_X5Y20_F_masked2, //EXTERNAL
        input Tile_X6Y20_R_t, //EXTERNAL
        input Tile_X6Y20_R_f, //EXTERNAL
        output Tile_X6Y20_F_masked1, //EXTERNAL
        output Tile_X6Y20_F_masked2, //EXTERNAL
        output Tile_X7Y20_F_masked1, //EXTERNAL
        output Tile_X7Y20_F_masked2, //EXTERNAL
        output Tile_X9Y20_F_ctrl, //EXTERNAL
        input Tile_X10Y20_A_O_top_0_t, //EXTERNAL
        input Tile_X10Y20_A_O_top_0_f, //EXTERNAL
        input Tile_X10Y20_A_prech2, //EXTERNAL
        input Tile_X10Y20_A_DR_fault, //EXTERNAL
        output Tile_X10Y20_A_I_top_0_t, //EXTERNAL
        output Tile_X10Y20_A_I_top_0_f, //EXTERNAL
        output Tile_X10Y20_A_T_top, //EXTERNAL
        output Tile_X10Y20_A_F_ctrl, //EXTERNAL
        input Tile_X0Y21_A_O_top_0_t, //EXTERNAL
        input Tile_X0Y21_A_O_top_0_f, //EXTERNAL
        input Tile_X0Y21_A_O_top_1_t, //EXTERNAL
        input Tile_X0Y21_A_O_top_1_f, //EXTERNAL
        input Tile_X0Y21_A_prech1, //EXTERNAL
        input Tile_X0Y21_A_prech2, //EXTERNAL
        input Tile_X0Y21_A_DR_fault, //EXTERNAL
        output Tile_X0Y21_A_I_top_0_t, //EXTERNAL
        output Tile_X0Y21_A_I_top_0_f, //EXTERNAL
        output Tile_X0Y21_A_I_top_1_t, //EXTERNAL
        output Tile_X0Y21_A_I_top_1_f, //EXTERNAL
        output Tile_X0Y21_A_T_top, //EXTERNAL
        output Tile_X0Y21_A_F_masked1, //EXTERNAL
        output Tile_X0Y21_A_F_masked2, //EXTERNAL
        output Tile_X0Y21_A_config_C_bit0, //EXTERNAL
        output Tile_X0Y21_A_config_C_bit1, //EXTERNAL
        output Tile_X0Y21_A_config_C_bit2, //EXTERNAL
        output Tile_X0Y21_A_config_C_bit3, //EXTERNAL
        output Tile_X0Y21_B_config_C_bit0, //EXTERNAL
        output Tile_X0Y21_B_config_C_bit1, //EXTERNAL
        output Tile_X0Y21_B_config_C_bit2, //EXTERNAL
        output Tile_X0Y21_B_config_C_bit3, //EXTERNAL
        output Tile_X1Y21_F_masked1, //EXTERNAL
        output Tile_X1Y21_F_masked2, //EXTERNAL
        output Tile_X2Y21_F_masked1, //EXTERNAL
        output Tile_X2Y21_F_masked2, //EXTERNAL
        input Tile_X3Y21_R_t, //EXTERNAL
        input Tile_X3Y21_R_f, //EXTERNAL
        output Tile_X3Y21_F_masked1, //EXTERNAL
        output Tile_X3Y21_F_masked2, //EXTERNAL
        output Tile_X4Y21_F_masked1, //EXTERNAL
        output Tile_X4Y21_F_masked2, //EXTERNAL
        output Tile_X5Y21_F_masked1, //EXTERNAL
        output Tile_X5Y21_F_masked2, //EXTERNAL
        input Tile_X6Y21_R_t, //EXTERNAL
        input Tile_X6Y21_R_f, //EXTERNAL
        output Tile_X6Y21_F_masked1, //EXTERNAL
        output Tile_X6Y21_F_masked2, //EXTERNAL
        output Tile_X7Y21_F_masked1, //EXTERNAL
        output Tile_X7Y21_F_masked2, //EXTERNAL
        output Tile_X9Y21_F_ctrl, //EXTERNAL
        input Tile_X10Y21_A_O_top_0_t, //EXTERNAL
        input Tile_X10Y21_A_O_top_0_f, //EXTERNAL
        input Tile_X10Y21_A_prech2, //EXTERNAL
        input Tile_X10Y21_A_DR_fault, //EXTERNAL
        output Tile_X10Y21_A_I_top_0_t, //EXTERNAL
        output Tile_X10Y21_A_I_top_0_f, //EXTERNAL
        output Tile_X10Y21_A_T_top, //EXTERNAL
        output Tile_X10Y21_A_F_ctrl, //EXTERNAL
        input Tile_X0Y22_A_O_top_0_t, //EXTERNAL
        input Tile_X0Y22_A_O_top_0_f, //EXTERNAL
        input Tile_X0Y22_A_O_top_1_t, //EXTERNAL
        input Tile_X0Y22_A_O_top_1_f, //EXTERNAL
        input Tile_X0Y22_A_prech1, //EXTERNAL
        input Tile_X0Y22_A_prech2, //EXTERNAL
        input Tile_X0Y22_A_DR_fault, //EXTERNAL
        output Tile_X0Y22_A_I_top_0_t, //EXTERNAL
        output Tile_X0Y22_A_I_top_0_f, //EXTERNAL
        output Tile_X0Y22_A_I_top_1_t, //EXTERNAL
        output Tile_X0Y22_A_I_top_1_f, //EXTERNAL
        output Tile_X0Y22_A_T_top, //EXTERNAL
        output Tile_X0Y22_A_F_masked1, //EXTERNAL
        output Tile_X0Y22_A_F_masked2, //EXTERNAL
        output Tile_X0Y22_A_config_C_bit0, //EXTERNAL
        output Tile_X0Y22_A_config_C_bit1, //EXTERNAL
        output Tile_X0Y22_A_config_C_bit2, //EXTERNAL
        output Tile_X0Y22_A_config_C_bit3, //EXTERNAL
        output Tile_X0Y22_B_config_C_bit0, //EXTERNAL
        output Tile_X0Y22_B_config_C_bit1, //EXTERNAL
        output Tile_X0Y22_B_config_C_bit2, //EXTERNAL
        output Tile_X0Y22_B_config_C_bit3, //EXTERNAL
        output Tile_X1Y22_F_masked1, //EXTERNAL
        output Tile_X1Y22_F_masked2, //EXTERNAL
        output Tile_X2Y22_F_masked1, //EXTERNAL
        output Tile_X2Y22_F_masked2, //EXTERNAL
        input Tile_X3Y22_R_t, //EXTERNAL
        input Tile_X3Y22_R_f, //EXTERNAL
        output Tile_X3Y22_F_masked1, //EXTERNAL
        output Tile_X3Y22_F_masked2, //EXTERNAL
        output Tile_X4Y22_F_masked1, //EXTERNAL
        output Tile_X4Y22_F_masked2, //EXTERNAL
        output Tile_X5Y22_F_masked1, //EXTERNAL
        output Tile_X5Y22_F_masked2, //EXTERNAL
        input Tile_X6Y22_R_t, //EXTERNAL
        input Tile_X6Y22_R_f, //EXTERNAL
        output Tile_X6Y22_F_masked1, //EXTERNAL
        output Tile_X6Y22_F_masked2, //EXTERNAL
        output Tile_X7Y22_F_masked1, //EXTERNAL
        output Tile_X7Y22_F_masked2, //EXTERNAL
        output Tile_X9Y22_F_ctrl, //EXTERNAL
        input Tile_X10Y22_A_O_top_0_t, //EXTERNAL
        input Tile_X10Y22_A_O_top_0_f, //EXTERNAL
        input Tile_X10Y22_A_prech2, //EXTERNAL
        input Tile_X10Y22_A_DR_fault, //EXTERNAL
        output Tile_X10Y22_A_I_top_0_t, //EXTERNAL
        output Tile_X10Y22_A_I_top_0_f, //EXTERNAL
        output Tile_X10Y22_A_T_top, //EXTERNAL
        output Tile_X10Y22_A_F_ctrl, //EXTERNAL
        input Tile_X0Y23_A_O_top_0_t, //EXTERNAL
        input Tile_X0Y23_A_O_top_0_f, //EXTERNAL
        input Tile_X0Y23_A_O_top_1_t, //EXTERNAL
        input Tile_X0Y23_A_O_top_1_f, //EXTERNAL
        input Tile_X0Y23_A_prech1, //EXTERNAL
        input Tile_X0Y23_A_prech2, //EXTERNAL
        input Tile_X0Y23_A_DR_fault, //EXTERNAL
        output Tile_X0Y23_A_I_top_0_t, //EXTERNAL
        output Tile_X0Y23_A_I_top_0_f, //EXTERNAL
        output Tile_X0Y23_A_I_top_1_t, //EXTERNAL
        output Tile_X0Y23_A_I_top_1_f, //EXTERNAL
        output Tile_X0Y23_A_T_top, //EXTERNAL
        output Tile_X0Y23_A_F_masked1, //EXTERNAL
        output Tile_X0Y23_A_F_masked2, //EXTERNAL
        output Tile_X0Y23_A_config_C_bit0, //EXTERNAL
        output Tile_X0Y23_A_config_C_bit1, //EXTERNAL
        output Tile_X0Y23_A_config_C_bit2, //EXTERNAL
        output Tile_X0Y23_A_config_C_bit3, //EXTERNAL
        output Tile_X0Y23_B_config_C_bit0, //EXTERNAL
        output Tile_X0Y23_B_config_C_bit1, //EXTERNAL
        output Tile_X0Y23_B_config_C_bit2, //EXTERNAL
        output Tile_X0Y23_B_config_C_bit3, //EXTERNAL
        output Tile_X1Y23_F_masked1, //EXTERNAL
        output Tile_X1Y23_F_masked2, //EXTERNAL
        output Tile_X2Y23_F_masked1, //EXTERNAL
        output Tile_X2Y23_F_masked2, //EXTERNAL
        input Tile_X3Y23_R_t, //EXTERNAL
        input Tile_X3Y23_R_f, //EXTERNAL
        output Tile_X3Y23_F_masked1, //EXTERNAL
        output Tile_X3Y23_F_masked2, //EXTERNAL
        output Tile_X4Y23_F_masked1, //EXTERNAL
        output Tile_X4Y23_F_masked2, //EXTERNAL
        output Tile_X5Y23_F_masked1, //EXTERNAL
        output Tile_X5Y23_F_masked2, //EXTERNAL
        input Tile_X6Y23_R_t, //EXTERNAL
        input Tile_X6Y23_R_f, //EXTERNAL
        output Tile_X6Y23_F_masked1, //EXTERNAL
        output Tile_X6Y23_F_masked2, //EXTERNAL
        output Tile_X7Y23_F_masked1, //EXTERNAL
        output Tile_X7Y23_F_masked2, //EXTERNAL
        output Tile_X9Y23_F_ctrl, //EXTERNAL
        input Tile_X10Y23_A_O_top_0_t, //EXTERNAL
        input Tile_X10Y23_A_O_top_0_f, //EXTERNAL
        input Tile_X10Y23_A_prech2, //EXTERNAL
        input Tile_X10Y23_A_DR_fault, //EXTERNAL
        output Tile_X10Y23_A_I_top_0_t, //EXTERNAL
        output Tile_X10Y23_A_I_top_0_f, //EXTERNAL
        output Tile_X10Y23_A_T_top, //EXTERNAL
        output Tile_X10Y23_A_F_ctrl, //EXTERNAL
        input [(FrameBitsPerRow*25)-1:0] FrameData, //CONFIG_PORT
        input [(MaxFramesPerCol*11)-1:0] FrameStrobe, //CONFIG_PORT
        input UserCLK,
        input rst
);

 //signal declarations

wire Tile_X0Y0_UserCLKo;
wire Tile_X0Y0_rsto;
wire Tile_X1Y0_UserCLKo;
wire Tile_X1Y0_rsto;
wire Tile_X2Y0_UserCLKo;
wire Tile_X2Y0_rsto;
wire Tile_X3Y0_UserCLKo;
wire Tile_X3Y0_rsto;
wire Tile_X4Y0_UserCLKo;
wire Tile_X4Y0_rsto;
wire Tile_X5Y0_UserCLKo;
wire Tile_X5Y0_rsto;
wire Tile_X6Y0_UserCLKo;
wire Tile_X6Y0_rsto;
wire Tile_X7Y0_UserCLKo;
wire Tile_X7Y0_rsto;
wire Tile_X8Y0_UserCLKo;
wire Tile_X8Y0_rsto;
wire Tile_X9Y0_UserCLKo;
wire Tile_X9Y0_rsto;
wire Tile_X10Y0_UserCLKo;
wire Tile_X10Y0_rsto;
wire Tile_X0Y1_UserCLKo;
wire Tile_X0Y1_rsto;
wire Tile_X1Y1_UserCLKo;
wire Tile_X1Y1_rsto;
wire Tile_X2Y1_UserCLKo;
wire Tile_X2Y1_rsto;
wire Tile_X3Y1_UserCLKo;
wire Tile_X3Y1_rsto;
wire Tile_X4Y1_UserCLKo;
wire Tile_X4Y1_rsto;
wire Tile_X5Y1_UserCLKo;
wire Tile_X5Y1_rsto;
wire Tile_X6Y1_UserCLKo;
wire Tile_X6Y1_rsto;
wire Tile_X7Y1_UserCLKo;
wire Tile_X7Y1_rsto;
wire Tile_X8Y1_UserCLKo;
wire Tile_X8Y1_rsto;
wire Tile_X9Y1_UserCLKo;
wire Tile_X9Y1_rsto;
wire Tile_X10Y1_UserCLKo;
wire Tile_X10Y1_rsto;
wire Tile_X0Y2_UserCLKo;
wire Tile_X0Y2_rsto;
wire Tile_X1Y2_UserCLKo;
wire Tile_X1Y2_rsto;
wire Tile_X2Y2_UserCLKo;
wire Tile_X2Y2_rsto;
wire Tile_X3Y2_UserCLKo;
wire Tile_X3Y2_rsto;
wire Tile_X4Y2_UserCLKo;
wire Tile_X4Y2_rsto;
wire Tile_X5Y2_UserCLKo;
wire Tile_X5Y2_rsto;
wire Tile_X6Y2_UserCLKo;
wire Tile_X6Y2_rsto;
wire Tile_X7Y2_UserCLKo;
wire Tile_X7Y2_rsto;
wire Tile_X8Y2_UserCLKo;
wire Tile_X8Y2_rsto;
wire Tile_X9Y2_UserCLKo;
wire Tile_X9Y2_rsto;
wire Tile_X10Y2_UserCLKo;
wire Tile_X10Y2_rsto;
wire Tile_X0Y3_UserCLKo;
wire Tile_X0Y3_rsto;
wire Tile_X1Y3_UserCLKo;
wire Tile_X1Y3_rsto;
wire Tile_X2Y3_UserCLKo;
wire Tile_X2Y3_rsto;
wire Tile_X3Y3_UserCLKo;
wire Tile_X3Y3_rsto;
wire Tile_X4Y3_UserCLKo;
wire Tile_X4Y3_rsto;
wire Tile_X5Y3_UserCLKo;
wire Tile_X5Y3_rsto;
wire Tile_X6Y3_UserCLKo;
wire Tile_X6Y3_rsto;
wire Tile_X7Y3_UserCLKo;
wire Tile_X7Y3_rsto;
wire Tile_X8Y3_UserCLKo;
wire Tile_X8Y3_rsto;
wire Tile_X9Y3_UserCLKo;
wire Tile_X9Y3_rsto;
wire Tile_X10Y3_UserCLKo;
wire Tile_X10Y3_rsto;
wire Tile_X0Y4_UserCLKo;
wire Tile_X0Y4_rsto;
wire Tile_X1Y4_UserCLKo;
wire Tile_X1Y4_rsto;
wire Tile_X2Y4_UserCLKo;
wire Tile_X2Y4_rsto;
wire Tile_X3Y4_UserCLKo;
wire Tile_X3Y4_rsto;
wire Tile_X4Y4_UserCLKo;
wire Tile_X4Y4_rsto;
wire Tile_X5Y4_UserCLKo;
wire Tile_X5Y4_rsto;
wire Tile_X6Y4_UserCLKo;
wire Tile_X6Y4_rsto;
wire Tile_X7Y4_UserCLKo;
wire Tile_X7Y4_rsto;
wire Tile_X8Y4_UserCLKo;
wire Tile_X8Y4_rsto;
wire Tile_X9Y4_UserCLKo;
wire Tile_X9Y4_rsto;
wire Tile_X10Y4_UserCLKo;
wire Tile_X10Y4_rsto;
wire Tile_X0Y5_UserCLKo;
wire Tile_X0Y5_rsto;
wire Tile_X1Y5_UserCLKo;
wire Tile_X1Y5_rsto;
wire Tile_X2Y5_UserCLKo;
wire Tile_X2Y5_rsto;
wire Tile_X3Y5_UserCLKo;
wire Tile_X3Y5_rsto;
wire Tile_X4Y5_UserCLKo;
wire Tile_X4Y5_rsto;
wire Tile_X5Y5_UserCLKo;
wire Tile_X5Y5_rsto;
wire Tile_X6Y5_UserCLKo;
wire Tile_X6Y5_rsto;
wire Tile_X7Y5_UserCLKo;
wire Tile_X7Y5_rsto;
wire Tile_X8Y5_UserCLKo;
wire Tile_X8Y5_rsto;
wire Tile_X9Y5_UserCLKo;
wire Tile_X9Y5_rsto;
wire Tile_X10Y5_UserCLKo;
wire Tile_X10Y5_rsto;
wire Tile_X0Y6_UserCLKo;
wire Tile_X0Y6_rsto;
wire Tile_X1Y6_UserCLKo;
wire Tile_X1Y6_rsto;
wire Tile_X2Y6_UserCLKo;
wire Tile_X2Y6_rsto;
wire Tile_X3Y6_UserCLKo;
wire Tile_X3Y6_rsto;
wire Tile_X4Y6_UserCLKo;
wire Tile_X4Y6_rsto;
wire Tile_X5Y6_UserCLKo;
wire Tile_X5Y6_rsto;
wire Tile_X6Y6_UserCLKo;
wire Tile_X6Y6_rsto;
wire Tile_X7Y6_UserCLKo;
wire Tile_X7Y6_rsto;
wire Tile_X8Y6_UserCLKo;
wire Tile_X8Y6_rsto;
wire Tile_X9Y6_UserCLKo;
wire Tile_X9Y6_rsto;
wire Tile_X10Y6_UserCLKo;
wire Tile_X10Y6_rsto;
wire Tile_X0Y7_UserCLKo;
wire Tile_X0Y7_rsto;
wire Tile_X1Y7_UserCLKo;
wire Tile_X1Y7_rsto;
wire Tile_X2Y7_UserCLKo;
wire Tile_X2Y7_rsto;
wire Tile_X3Y7_UserCLKo;
wire Tile_X3Y7_rsto;
wire Tile_X4Y7_UserCLKo;
wire Tile_X4Y7_rsto;
wire Tile_X5Y7_UserCLKo;
wire Tile_X5Y7_rsto;
wire Tile_X6Y7_UserCLKo;
wire Tile_X6Y7_rsto;
wire Tile_X7Y7_UserCLKo;
wire Tile_X7Y7_rsto;
wire Tile_X8Y7_UserCLKo;
wire Tile_X8Y7_rsto;
wire Tile_X9Y7_UserCLKo;
wire Tile_X9Y7_rsto;
wire Tile_X10Y7_UserCLKo;
wire Tile_X10Y7_rsto;
wire Tile_X0Y8_UserCLKo;
wire Tile_X0Y8_rsto;
wire Tile_X1Y8_UserCLKo;
wire Tile_X1Y8_rsto;
wire Tile_X2Y8_UserCLKo;
wire Tile_X2Y8_rsto;
wire Tile_X3Y8_UserCLKo;
wire Tile_X3Y8_rsto;
wire Tile_X4Y8_UserCLKo;
wire Tile_X4Y8_rsto;
wire Tile_X5Y8_UserCLKo;
wire Tile_X5Y8_rsto;
wire Tile_X6Y8_UserCLKo;
wire Tile_X6Y8_rsto;
wire Tile_X7Y8_UserCLKo;
wire Tile_X7Y8_rsto;
wire Tile_X8Y8_UserCLKo;
wire Tile_X8Y8_rsto;
wire Tile_X9Y8_UserCLKo;
wire Tile_X9Y8_rsto;
wire Tile_X10Y8_UserCLKo;
wire Tile_X10Y8_rsto;
wire Tile_X0Y9_UserCLKo;
wire Tile_X0Y9_rsto;
wire Tile_X1Y9_UserCLKo;
wire Tile_X1Y9_rsto;
wire Tile_X2Y9_UserCLKo;
wire Tile_X2Y9_rsto;
wire Tile_X3Y9_UserCLKo;
wire Tile_X3Y9_rsto;
wire Tile_X4Y9_UserCLKo;
wire Tile_X4Y9_rsto;
wire Tile_X5Y9_UserCLKo;
wire Tile_X5Y9_rsto;
wire Tile_X6Y9_UserCLKo;
wire Tile_X6Y9_rsto;
wire Tile_X7Y9_UserCLKo;
wire Tile_X7Y9_rsto;
wire Tile_X8Y9_UserCLKo;
wire Tile_X8Y9_rsto;
wire Tile_X9Y9_UserCLKo;
wire Tile_X9Y9_rsto;
wire Tile_X10Y9_UserCLKo;
wire Tile_X10Y9_rsto;
wire Tile_X0Y10_UserCLKo;
wire Tile_X0Y10_rsto;
wire Tile_X1Y10_UserCLKo;
wire Tile_X1Y10_rsto;
wire Tile_X2Y10_UserCLKo;
wire Tile_X2Y10_rsto;
wire Tile_X3Y10_UserCLKo;
wire Tile_X3Y10_rsto;
wire Tile_X4Y10_UserCLKo;
wire Tile_X4Y10_rsto;
wire Tile_X5Y10_UserCLKo;
wire Tile_X5Y10_rsto;
wire Tile_X6Y10_UserCLKo;
wire Tile_X6Y10_rsto;
wire Tile_X7Y10_UserCLKo;
wire Tile_X7Y10_rsto;
wire Tile_X8Y10_UserCLKo;
wire Tile_X8Y10_rsto;
wire Tile_X9Y10_UserCLKo;
wire Tile_X9Y10_rsto;
wire Tile_X10Y10_UserCLKo;
wire Tile_X10Y10_rsto;
wire Tile_X0Y11_UserCLKo;
wire Tile_X0Y11_rsto;
wire Tile_X1Y11_UserCLKo;
wire Tile_X1Y11_rsto;
wire Tile_X2Y11_UserCLKo;
wire Tile_X2Y11_rsto;
wire Tile_X3Y11_UserCLKo;
wire Tile_X3Y11_rsto;
wire Tile_X4Y11_UserCLKo;
wire Tile_X4Y11_rsto;
wire Tile_X5Y11_UserCLKo;
wire Tile_X5Y11_rsto;
wire Tile_X6Y11_UserCLKo;
wire Tile_X6Y11_rsto;
wire Tile_X7Y11_UserCLKo;
wire Tile_X7Y11_rsto;
wire Tile_X8Y11_UserCLKo;
wire Tile_X8Y11_rsto;
wire Tile_X9Y11_UserCLKo;
wire Tile_X9Y11_rsto;
wire Tile_X10Y11_UserCLKo;
wire Tile_X10Y11_rsto;
wire Tile_X0Y12_UserCLKo;
wire Tile_X0Y12_rsto;
wire Tile_X1Y12_UserCLKo;
wire Tile_X1Y12_rsto;
wire Tile_X2Y12_UserCLKo;
wire Tile_X2Y12_rsto;
wire Tile_X3Y12_UserCLKo;
wire Tile_X3Y12_rsto;
wire Tile_X4Y12_UserCLKo;
wire Tile_X4Y12_rsto;
wire Tile_X5Y12_UserCLKo;
wire Tile_X5Y12_rsto;
wire Tile_X6Y12_UserCLKo;
wire Tile_X6Y12_rsto;
wire Tile_X7Y12_UserCLKo;
wire Tile_X7Y12_rsto;
wire Tile_X8Y12_UserCLKo;
wire Tile_X8Y12_rsto;
wire Tile_X9Y12_UserCLKo;
wire Tile_X9Y12_rsto;
wire Tile_X10Y12_UserCLKo;
wire Tile_X10Y12_rsto;
wire Tile_X0Y13_UserCLKo;
wire Tile_X0Y13_rsto;
wire Tile_X1Y13_UserCLKo;
wire Tile_X1Y13_rsto;
wire Tile_X2Y13_UserCLKo;
wire Tile_X2Y13_rsto;
wire Tile_X3Y13_UserCLKo;
wire Tile_X3Y13_rsto;
wire Tile_X4Y13_UserCLKo;
wire Tile_X4Y13_rsto;
wire Tile_X5Y13_UserCLKo;
wire Tile_X5Y13_rsto;
wire Tile_X6Y13_UserCLKo;
wire Tile_X6Y13_rsto;
wire Tile_X7Y13_UserCLKo;
wire Tile_X7Y13_rsto;
wire Tile_X8Y13_UserCLKo;
wire Tile_X8Y13_rsto;
wire Tile_X9Y13_UserCLKo;
wire Tile_X9Y13_rsto;
wire Tile_X10Y13_UserCLKo;
wire Tile_X10Y13_rsto;
wire Tile_X0Y14_UserCLKo;
wire Tile_X0Y14_rsto;
wire Tile_X1Y14_UserCLKo;
wire Tile_X1Y14_rsto;
wire Tile_X2Y14_UserCLKo;
wire Tile_X2Y14_rsto;
wire Tile_X3Y14_UserCLKo;
wire Tile_X3Y14_rsto;
wire Tile_X4Y14_UserCLKo;
wire Tile_X4Y14_rsto;
wire Tile_X5Y14_UserCLKo;
wire Tile_X5Y14_rsto;
wire Tile_X6Y14_UserCLKo;
wire Tile_X6Y14_rsto;
wire Tile_X7Y14_UserCLKo;
wire Tile_X7Y14_rsto;
wire Tile_X8Y14_UserCLKo;
wire Tile_X8Y14_rsto;
wire Tile_X9Y14_UserCLKo;
wire Tile_X9Y14_rsto;
wire Tile_X10Y14_UserCLKo;
wire Tile_X10Y14_rsto;
wire Tile_X0Y15_UserCLKo;
wire Tile_X0Y15_rsto;
wire Tile_X1Y15_UserCLKo;
wire Tile_X1Y15_rsto;
wire Tile_X2Y15_UserCLKo;
wire Tile_X2Y15_rsto;
wire Tile_X3Y15_UserCLKo;
wire Tile_X3Y15_rsto;
wire Tile_X4Y15_UserCLKo;
wire Tile_X4Y15_rsto;
wire Tile_X5Y15_UserCLKo;
wire Tile_X5Y15_rsto;
wire Tile_X6Y15_UserCLKo;
wire Tile_X6Y15_rsto;
wire Tile_X7Y15_UserCLKo;
wire Tile_X7Y15_rsto;
wire Tile_X8Y15_UserCLKo;
wire Tile_X8Y15_rsto;
wire Tile_X9Y15_UserCLKo;
wire Tile_X9Y15_rsto;
wire Tile_X10Y15_UserCLKo;
wire Tile_X10Y15_rsto;
wire Tile_X0Y16_UserCLKo;
wire Tile_X0Y16_rsto;
wire Tile_X1Y16_UserCLKo;
wire Tile_X1Y16_rsto;
wire Tile_X2Y16_UserCLKo;
wire Tile_X2Y16_rsto;
wire Tile_X3Y16_UserCLKo;
wire Tile_X3Y16_rsto;
wire Tile_X4Y16_UserCLKo;
wire Tile_X4Y16_rsto;
wire Tile_X5Y16_UserCLKo;
wire Tile_X5Y16_rsto;
wire Tile_X6Y16_UserCLKo;
wire Tile_X6Y16_rsto;
wire Tile_X7Y16_UserCLKo;
wire Tile_X7Y16_rsto;
wire Tile_X8Y16_UserCLKo;
wire Tile_X8Y16_rsto;
wire Tile_X9Y16_UserCLKo;
wire Tile_X9Y16_rsto;
wire Tile_X10Y16_UserCLKo;
wire Tile_X10Y16_rsto;
wire Tile_X0Y17_UserCLKo;
wire Tile_X0Y17_rsto;
wire Tile_X1Y17_UserCLKo;
wire Tile_X1Y17_rsto;
wire Tile_X2Y17_UserCLKo;
wire Tile_X2Y17_rsto;
wire Tile_X3Y17_UserCLKo;
wire Tile_X3Y17_rsto;
wire Tile_X4Y17_UserCLKo;
wire Tile_X4Y17_rsto;
wire Tile_X5Y17_UserCLKo;
wire Tile_X5Y17_rsto;
wire Tile_X6Y17_UserCLKo;
wire Tile_X6Y17_rsto;
wire Tile_X7Y17_UserCLKo;
wire Tile_X7Y17_rsto;
wire Tile_X8Y17_UserCLKo;
wire Tile_X8Y17_rsto;
wire Tile_X9Y17_UserCLKo;
wire Tile_X9Y17_rsto;
wire Tile_X10Y17_UserCLKo;
wire Tile_X10Y17_rsto;
wire Tile_X0Y18_UserCLKo;
wire Tile_X0Y18_rsto;
wire Tile_X1Y18_UserCLKo;
wire Tile_X1Y18_rsto;
wire Tile_X2Y18_UserCLKo;
wire Tile_X2Y18_rsto;
wire Tile_X3Y18_UserCLKo;
wire Tile_X3Y18_rsto;
wire Tile_X4Y18_UserCLKo;
wire Tile_X4Y18_rsto;
wire Tile_X5Y18_UserCLKo;
wire Tile_X5Y18_rsto;
wire Tile_X6Y18_UserCLKo;
wire Tile_X6Y18_rsto;
wire Tile_X7Y18_UserCLKo;
wire Tile_X7Y18_rsto;
wire Tile_X8Y18_UserCLKo;
wire Tile_X8Y18_rsto;
wire Tile_X9Y18_UserCLKo;
wire Tile_X9Y18_rsto;
wire Tile_X10Y18_UserCLKo;
wire Tile_X10Y18_rsto;
wire Tile_X0Y19_UserCLKo;
wire Tile_X0Y19_rsto;
wire Tile_X1Y19_UserCLKo;
wire Tile_X1Y19_rsto;
wire Tile_X2Y19_UserCLKo;
wire Tile_X2Y19_rsto;
wire Tile_X3Y19_UserCLKo;
wire Tile_X3Y19_rsto;
wire Tile_X4Y19_UserCLKo;
wire Tile_X4Y19_rsto;
wire Tile_X5Y19_UserCLKo;
wire Tile_X5Y19_rsto;
wire Tile_X6Y19_UserCLKo;
wire Tile_X6Y19_rsto;
wire Tile_X7Y19_UserCLKo;
wire Tile_X7Y19_rsto;
wire Tile_X8Y19_UserCLKo;
wire Tile_X8Y19_rsto;
wire Tile_X9Y19_UserCLKo;
wire Tile_X9Y19_rsto;
wire Tile_X10Y19_UserCLKo;
wire Tile_X10Y19_rsto;
wire Tile_X0Y20_UserCLKo;
wire Tile_X0Y20_rsto;
wire Tile_X1Y20_UserCLKo;
wire Tile_X1Y20_rsto;
wire Tile_X2Y20_UserCLKo;
wire Tile_X2Y20_rsto;
wire Tile_X3Y20_UserCLKo;
wire Tile_X3Y20_rsto;
wire Tile_X4Y20_UserCLKo;
wire Tile_X4Y20_rsto;
wire Tile_X5Y20_UserCLKo;
wire Tile_X5Y20_rsto;
wire Tile_X6Y20_UserCLKo;
wire Tile_X6Y20_rsto;
wire Tile_X7Y20_UserCLKo;
wire Tile_X7Y20_rsto;
wire Tile_X8Y20_UserCLKo;
wire Tile_X8Y20_rsto;
wire Tile_X9Y20_UserCLKo;
wire Tile_X9Y20_rsto;
wire Tile_X10Y20_UserCLKo;
wire Tile_X10Y20_rsto;
wire Tile_X0Y21_UserCLKo;
wire Tile_X0Y21_rsto;
wire Tile_X1Y21_UserCLKo;
wire Tile_X1Y21_rsto;
wire Tile_X2Y21_UserCLKo;
wire Tile_X2Y21_rsto;
wire Tile_X3Y21_UserCLKo;
wire Tile_X3Y21_rsto;
wire Tile_X4Y21_UserCLKo;
wire Tile_X4Y21_rsto;
wire Tile_X5Y21_UserCLKo;
wire Tile_X5Y21_rsto;
wire Tile_X6Y21_UserCLKo;
wire Tile_X6Y21_rsto;
wire Tile_X7Y21_UserCLKo;
wire Tile_X7Y21_rsto;
wire Tile_X8Y21_UserCLKo;
wire Tile_X8Y21_rsto;
wire Tile_X9Y21_UserCLKo;
wire Tile_X9Y21_rsto;
wire Tile_X10Y21_UserCLKo;
wire Tile_X10Y21_rsto;
wire Tile_X0Y22_UserCLKo;
wire Tile_X0Y22_rsto;
wire Tile_X1Y22_UserCLKo;
wire Tile_X1Y22_rsto;
wire Tile_X2Y22_UserCLKo;
wire Tile_X2Y22_rsto;
wire Tile_X3Y22_UserCLKo;
wire Tile_X3Y22_rsto;
wire Tile_X4Y22_UserCLKo;
wire Tile_X4Y22_rsto;
wire Tile_X5Y22_UserCLKo;
wire Tile_X5Y22_rsto;
wire Tile_X6Y22_UserCLKo;
wire Tile_X6Y22_rsto;
wire Tile_X7Y22_UserCLKo;
wire Tile_X7Y22_rsto;
wire Tile_X8Y22_UserCLKo;
wire Tile_X8Y22_rsto;
wire Tile_X9Y22_UserCLKo;
wire Tile_X9Y22_rsto;
wire Tile_X10Y22_UserCLKo;
wire Tile_X10Y22_rsto;
wire Tile_X0Y23_UserCLKo;
wire Tile_X0Y23_rsto;
wire Tile_X1Y23_UserCLKo;
wire Tile_X1Y23_rsto;
wire Tile_X2Y23_UserCLKo;
wire Tile_X2Y23_rsto;
wire Tile_X3Y23_UserCLKo;
wire Tile_X3Y23_rsto;
wire Tile_X4Y23_UserCLKo;
wire Tile_X4Y23_rsto;
wire Tile_X5Y23_UserCLKo;
wire Tile_X5Y23_rsto;
wire Tile_X6Y23_UserCLKo;
wire Tile_X6Y23_rsto;
wire Tile_X7Y23_UserCLKo;
wire Tile_X7Y23_rsto;
wire Tile_X8Y23_UserCLKo;
wire Tile_X8Y23_rsto;
wire Tile_X9Y23_UserCLKo;
wire Tile_X9Y23_rsto;
wire Tile_X10Y23_UserCLKo;
wire Tile_X10Y23_rsto;
wire Tile_X0Y24_UserCLKo;
wire Tile_X0Y24_rsto;
wire Tile_X1Y24_UserCLKo;
wire Tile_X1Y24_rsto;
wire Tile_X2Y24_UserCLKo;
wire Tile_X2Y24_rsto;
wire Tile_X3Y24_UserCLKo;
wire Tile_X3Y24_rsto;
wire Tile_X4Y24_UserCLKo;
wire Tile_X4Y24_rsto;
wire Tile_X5Y24_UserCLKo;
wire Tile_X5Y24_rsto;
wire Tile_X6Y24_UserCLKo;
wire Tile_X6Y24_rsto;
wire Tile_X7Y24_UserCLKo;
wire Tile_X7Y24_rsto;
wire Tile_X8Y24_UserCLKo;
wire Tile_X8Y24_rsto;
wire Tile_X9Y24_UserCLKo;
wire Tile_X9Y24_rsto;
wire Tile_X10Y24_UserCLKo;
wire Tile_X10Y24_rsto;
 //configuration signal declarations

wire[FrameBitsPerRow -1:0] Tile_Y0_FrameData;
wire[FrameBitsPerRow -1:0] Tile_Y1_FrameData;
wire[FrameBitsPerRow -1:0] Tile_Y2_FrameData;
wire[FrameBitsPerRow -1:0] Tile_Y3_FrameData;
wire[FrameBitsPerRow -1:0] Tile_Y4_FrameData;
wire[FrameBitsPerRow -1:0] Tile_Y5_FrameData;
wire[FrameBitsPerRow -1:0] Tile_Y6_FrameData;
wire[FrameBitsPerRow -1:0] Tile_Y7_FrameData;
wire[FrameBitsPerRow -1:0] Tile_Y8_FrameData;
wire[FrameBitsPerRow -1:0] Tile_Y9_FrameData;
wire[FrameBitsPerRow -1:0] Tile_Y10_FrameData;
wire[FrameBitsPerRow -1:0] Tile_Y11_FrameData;
wire[FrameBitsPerRow -1:0] Tile_Y12_FrameData;
wire[FrameBitsPerRow -1:0] Tile_Y13_FrameData;
wire[FrameBitsPerRow -1:0] Tile_Y14_FrameData;
wire[FrameBitsPerRow -1:0] Tile_Y15_FrameData;
wire[FrameBitsPerRow -1:0] Tile_Y16_FrameData;
wire[FrameBitsPerRow -1:0] Tile_Y17_FrameData;
wire[FrameBitsPerRow -1:0] Tile_Y18_FrameData;
wire[FrameBitsPerRow -1:0] Tile_Y19_FrameData;
wire[FrameBitsPerRow -1:0] Tile_Y20_FrameData;
wire[FrameBitsPerRow -1:0] Tile_Y21_FrameData;
wire[FrameBitsPerRow -1:0] Tile_Y22_FrameData;
wire[FrameBitsPerRow -1:0] Tile_Y23_FrameData;
wire[FrameBitsPerRow -1:0] Tile_Y24_FrameData;
wire[MaxFramesPerCol - 1:0] Tile_X0_FrameStrobe;
wire[MaxFramesPerCol - 1:0] Tile_X1_FrameStrobe;
wire[MaxFramesPerCol - 1:0] Tile_X2_FrameStrobe;
wire[MaxFramesPerCol - 1:0] Tile_X3_FrameStrobe;
wire[MaxFramesPerCol - 1:0] Tile_X4_FrameStrobe;
wire[MaxFramesPerCol - 1:0] Tile_X5_FrameStrobe;
wire[MaxFramesPerCol - 1:0] Tile_X6_FrameStrobe;
wire[MaxFramesPerCol - 1:0] Tile_X7_FrameStrobe;
wire[MaxFramesPerCol - 1:0] Tile_X8_FrameStrobe;
wire[MaxFramesPerCol - 1:0] Tile_X9_FrameStrobe;
wire[MaxFramesPerCol - 1:0] Tile_X10_FrameStrobe;
wire[FrameBitsPerRow - 1:0] Tile_X0Y0_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X1Y0_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X2Y0_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X3Y0_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X4Y0_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X5Y0_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X6Y0_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X7Y0_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X8Y0_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X9Y0_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X10Y0_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X0Y1_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X1Y1_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X2Y1_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X3Y1_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X4Y1_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X5Y1_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X6Y1_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X7Y1_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X8Y1_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X9Y1_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X10Y1_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X0Y2_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X1Y2_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X2Y2_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X3Y2_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X4Y2_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X5Y2_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X6Y2_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X7Y2_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X8Y2_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X9Y2_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X10Y2_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X0Y3_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X1Y3_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X2Y3_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X3Y3_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X4Y3_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X5Y3_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X6Y3_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X7Y3_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X8Y3_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X9Y3_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X10Y3_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X0Y4_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X1Y4_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X2Y4_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X3Y4_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X4Y4_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X5Y4_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X6Y4_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X7Y4_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X8Y4_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X9Y4_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X10Y4_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X0Y5_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X1Y5_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X2Y5_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X3Y5_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X4Y5_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X5Y5_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X6Y5_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X7Y5_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X8Y5_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X9Y5_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X10Y5_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X0Y6_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X1Y6_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X2Y6_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X3Y6_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X4Y6_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X5Y6_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X6Y6_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X7Y6_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X8Y6_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X9Y6_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X10Y6_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X0Y7_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X1Y7_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X2Y7_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X3Y7_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X4Y7_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X5Y7_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X6Y7_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X7Y7_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X8Y7_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X9Y7_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X10Y7_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X0Y8_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X1Y8_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X2Y8_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X3Y8_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X4Y8_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X5Y8_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X6Y8_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X7Y8_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X8Y8_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X9Y8_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X10Y8_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X0Y9_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X1Y9_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X2Y9_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X3Y9_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X4Y9_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X5Y9_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X6Y9_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X7Y9_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X8Y9_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X9Y9_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X10Y9_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X0Y10_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X1Y10_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X2Y10_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X3Y10_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X4Y10_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X5Y10_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X6Y10_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X7Y10_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X8Y10_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X9Y10_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X10Y10_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X0Y11_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X1Y11_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X2Y11_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X3Y11_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X4Y11_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X5Y11_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X6Y11_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X7Y11_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X8Y11_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X9Y11_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X10Y11_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X0Y12_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X1Y12_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X2Y12_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X3Y12_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X4Y12_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X5Y12_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X6Y12_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X7Y12_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X8Y12_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X9Y12_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X10Y12_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X0Y13_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X1Y13_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X2Y13_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X3Y13_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X4Y13_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X5Y13_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X6Y13_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X7Y13_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X8Y13_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X9Y13_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X10Y13_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X0Y14_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X1Y14_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X2Y14_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X3Y14_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X4Y14_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X5Y14_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X6Y14_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X7Y14_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X8Y14_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X9Y14_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X10Y14_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X0Y15_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X1Y15_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X2Y15_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X3Y15_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X4Y15_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X5Y15_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X6Y15_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X7Y15_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X8Y15_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X9Y15_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X10Y15_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X0Y16_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X1Y16_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X2Y16_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X3Y16_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X4Y16_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X5Y16_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X6Y16_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X7Y16_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X8Y16_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X9Y16_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X10Y16_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X0Y17_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X1Y17_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X2Y17_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X3Y17_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X4Y17_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X5Y17_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X6Y17_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X7Y17_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X8Y17_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X9Y17_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X10Y17_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X0Y18_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X1Y18_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X2Y18_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X3Y18_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X4Y18_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X5Y18_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X6Y18_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X7Y18_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X8Y18_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X9Y18_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X10Y18_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X0Y19_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X1Y19_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X2Y19_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X3Y19_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X4Y19_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X5Y19_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X6Y19_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X7Y19_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X8Y19_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X9Y19_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X10Y19_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X0Y20_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X1Y20_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X2Y20_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X3Y20_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X4Y20_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X5Y20_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X6Y20_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X7Y20_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X8Y20_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X9Y20_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X10Y20_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X0Y21_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X1Y21_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X2Y21_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X3Y21_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X4Y21_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X5Y21_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X6Y21_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X7Y21_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X8Y21_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X9Y21_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X10Y21_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X0Y22_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X1Y22_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X2Y22_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X3Y22_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X4Y22_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X5Y22_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X6Y22_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X7Y22_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X8Y22_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X9Y22_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X10Y22_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X0Y23_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X1Y23_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X2Y23_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X3Y23_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X4Y23_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X5Y23_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X6Y23_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X7Y23_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X8Y23_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X9Y23_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X10Y23_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X0Y24_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X1Y24_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X2Y24_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X3Y24_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X4Y24_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X5Y24_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X6Y24_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X7Y24_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X8Y24_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X9Y24_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X10Y24_FrameData_O;
wire[MaxFramesPerCol - 1:0] Tile_X0Y0_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X1Y0_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X2Y0_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X3Y0_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X4Y0_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X5Y0_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X6Y0_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X7Y0_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X8Y0_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X9Y0_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X10Y0_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X0Y1_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X1Y1_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X2Y1_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X3Y1_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X4Y1_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X5Y1_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X6Y1_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X7Y1_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X8Y1_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X9Y1_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X10Y1_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X0Y2_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X1Y2_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X2Y2_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X3Y2_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X4Y2_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X5Y2_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X6Y2_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X7Y2_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X8Y2_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X9Y2_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X10Y2_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X0Y3_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X1Y3_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X2Y3_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X3Y3_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X4Y3_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X5Y3_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X6Y3_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X7Y3_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X8Y3_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X9Y3_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X10Y3_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X0Y4_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X1Y4_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X2Y4_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X3Y4_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X4Y4_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X5Y4_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X6Y4_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X7Y4_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X8Y4_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X9Y4_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X10Y4_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X0Y5_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X1Y5_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X2Y5_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X3Y5_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X4Y5_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X5Y5_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X6Y5_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X7Y5_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X8Y5_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X9Y5_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X10Y5_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X0Y6_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X1Y6_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X2Y6_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X3Y6_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X4Y6_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X5Y6_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X6Y6_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X7Y6_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X8Y6_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X9Y6_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X10Y6_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X0Y7_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X1Y7_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X2Y7_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X3Y7_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X4Y7_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X5Y7_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X6Y7_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X7Y7_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X8Y7_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X9Y7_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X10Y7_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X0Y8_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X1Y8_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X2Y8_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X3Y8_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X4Y8_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X5Y8_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X6Y8_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X7Y8_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X8Y8_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X9Y8_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X10Y8_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X0Y9_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X1Y9_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X2Y9_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X3Y9_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X4Y9_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X5Y9_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X6Y9_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X7Y9_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X8Y9_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X9Y9_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X10Y9_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X0Y10_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X1Y10_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X2Y10_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X3Y10_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X4Y10_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X5Y10_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X6Y10_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X7Y10_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X8Y10_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X9Y10_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X10Y10_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X0Y11_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X1Y11_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X2Y11_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X3Y11_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X4Y11_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X5Y11_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X6Y11_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X7Y11_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X8Y11_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X9Y11_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X10Y11_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X0Y12_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X1Y12_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X2Y12_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X3Y12_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X4Y12_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X5Y12_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X6Y12_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X7Y12_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X8Y12_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X9Y12_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X10Y12_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X0Y13_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X1Y13_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X2Y13_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X3Y13_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X4Y13_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X5Y13_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X6Y13_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X7Y13_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X8Y13_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X9Y13_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X10Y13_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X0Y14_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X1Y14_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X2Y14_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X3Y14_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X4Y14_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X5Y14_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X6Y14_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X7Y14_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X8Y14_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X9Y14_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X10Y14_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X0Y15_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X1Y15_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X2Y15_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X3Y15_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X4Y15_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X5Y15_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X6Y15_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X7Y15_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X8Y15_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X9Y15_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X10Y15_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X0Y16_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X1Y16_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X2Y16_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X3Y16_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X4Y16_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X5Y16_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X6Y16_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X7Y16_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X8Y16_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X9Y16_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X10Y16_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X0Y17_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X1Y17_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X2Y17_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X3Y17_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X4Y17_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X5Y17_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X6Y17_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X7Y17_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X8Y17_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X9Y17_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X10Y17_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X0Y18_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X1Y18_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X2Y18_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X3Y18_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X4Y18_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X5Y18_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X6Y18_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X7Y18_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X8Y18_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X9Y18_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X10Y18_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X0Y19_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X1Y19_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X2Y19_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X3Y19_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X4Y19_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X5Y19_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X6Y19_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X7Y19_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X8Y19_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X9Y19_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X10Y19_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X0Y20_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X1Y20_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X2Y20_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X3Y20_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X4Y20_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X5Y20_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X6Y20_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X7Y20_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X8Y20_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X9Y20_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X10Y20_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X0Y21_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X1Y21_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X2Y21_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X3Y21_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X4Y21_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X5Y21_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X6Y21_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X7Y21_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X8Y21_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X9Y21_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X10Y21_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X0Y22_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X1Y22_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X2Y22_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X3Y22_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X4Y22_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X5Y22_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X6Y22_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X7Y22_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X8Y22_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X9Y22_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X10Y22_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X0Y23_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X1Y23_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X2Y23_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X3Y23_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X4Y23_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X5Y23_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X6Y23_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X7Y23_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X8Y23_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X9Y23_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X10Y23_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X0Y24_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X1Y24_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X2Y24_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X3Y24_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X4Y24_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X5Y24_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X6Y24_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X7Y24_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X8Y24_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X9Y24_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X10Y24_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X0Y25_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X1Y25_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X2Y25_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X3Y25_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X4Y25_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X5Y25_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X6Y25_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X7Y25_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X8Y25_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X9Y25_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X10Y25_FrameStrobe_O;
 //tile-to-tile signal declarations
wire[3:0] Tile_X0Y0_to_SA;
wire[3:0] Tile_X0Y0_to_SB;
wire[3:0] Tile_X0Y0_to_SC;
wire[3:0] Tile_X0Y0_to_SD;
wire[3:0] Tile_X0Y0_to_SF;
wire[7:0] Tile_X0Y0_to_SG;
wire[7:0] Tile_X0Y0_to_SH;
wire[11:0] Tile_X0Y0_to_SI;
wire[3:0] Tile_X1Y0_to_SA;
wire[3:0] Tile_X1Y0_to_SB;
wire[3:0] Tile_X1Y0_to_SC;
wire[3:0] Tile_X1Y0_to_SD;
wire[3:0] Tile_X1Y0_to_SF;
wire[7:0] Tile_X1Y0_to_SG;
wire[7:0] Tile_X1Y0_to_SH;
wire[11:0] Tile_X1Y0_to_SI;
wire[3:0] Tile_X2Y0_to_SA;
wire[3:0] Tile_X2Y0_to_SB;
wire[3:0] Tile_X2Y0_to_SC;
wire[3:0] Tile_X2Y0_to_SD;
wire[3:0] Tile_X2Y0_to_SF;
wire[7:0] Tile_X2Y0_to_SG;
wire[7:0] Tile_X2Y0_to_SH;
wire[11:0] Tile_X2Y0_to_SI;
wire[3:0] Tile_X3Y0_to_SA;
wire[3:0] Tile_X3Y0_to_SB;
wire[3:0] Tile_X3Y0_to_SC;
wire[3:0] Tile_X3Y0_to_SD;
wire[3:0] Tile_X3Y0_to_SF;
wire[7:0] Tile_X3Y0_to_SG;
wire[7:0] Tile_X3Y0_to_SH;
wire[11:0] Tile_X3Y0_to_SI;
wire[3:0] Tile_X4Y0_to_SA;
wire[3:0] Tile_X4Y0_to_SB;
wire[3:0] Tile_X4Y0_to_SC;
wire[3:0] Tile_X4Y0_to_SD;
wire[3:0] Tile_X4Y0_to_SF;
wire[7:0] Tile_X4Y0_to_SG;
wire[7:0] Tile_X4Y0_to_SH;
wire[11:0] Tile_X4Y0_to_SI;
wire[3:0] Tile_X5Y0_to_SA;
wire[3:0] Tile_X5Y0_to_SB;
wire[3:0] Tile_X5Y0_to_SC;
wire[3:0] Tile_X5Y0_to_SD;
wire[3:0] Tile_X5Y0_to_SF;
wire[7:0] Tile_X5Y0_to_SG;
wire[7:0] Tile_X5Y0_to_SH;
wire[11:0] Tile_X5Y0_to_SI;
wire[3:0] Tile_X6Y0_to_SA;
wire[3:0] Tile_X6Y0_to_SB;
wire[3:0] Tile_X6Y0_to_SC;
wire[3:0] Tile_X6Y0_to_SD;
wire[3:0] Tile_X6Y0_to_SF;
wire[7:0] Tile_X6Y0_to_SG;
wire[7:0] Tile_X6Y0_to_SH;
wire[11:0] Tile_X6Y0_to_SI;
wire[3:0] Tile_X7Y0_to_SA;
wire[3:0] Tile_X7Y0_to_SB;
wire[3:0] Tile_X7Y0_to_SC;
wire[3:0] Tile_X7Y0_to_SD;
wire[3:0] Tile_X7Y0_to_SF;
wire[7:0] Tile_X7Y0_to_SG;
wire[7:0] Tile_X7Y0_to_SH;
wire[11:0] Tile_X7Y0_to_SI;
wire[3:0] Tile_X8Y0_to_SA;
wire[3:0] Tile_X8Y0_to_SB;
wire[3:0] Tile_X8Y0_to_SC;
wire[3:0] Tile_X8Y0_to_SD;
wire[3:0] Tile_X8Y0_to_SF;
wire[7:0] Tile_X8Y0_to_SG;
wire[7:0] Tile_X8Y0_to_SH;
wire[11:0] Tile_X8Y0_to_SI;
wire[1:0] Tile_X9Y0_to_SA_1s;
wire[1:0] Tile_X9Y0_to_SB_1s;
wire[1:0] Tile_X9Y0_to_SC_1s;
wire[1:0] Tile_X9Y0_to_SD_1s;
wire[1:0] Tile_X9Y0_to_SF_1s;
wire[1:0] Tile_X9Y0_to_SG_1s;
wire[1:0] Tile_X9Y0_to_SH_1s;
wire[1:0] Tile_X9Y0_to_SI_1s;
wire[1:0] Tile_X10Y0_to_SA_1s;
wire[1:0] Tile_X10Y0_to_SB_1s;
wire[1:0] Tile_X10Y0_to_SC_1s;
wire[1:0] Tile_X10Y0_to_SD_1s;
wire[1:0] Tile_X10Y0_to_SF_1s;
wire[1:0] Tile_X10Y0_to_SG_1s;
wire[1:0] Tile_X10Y0_to_SH_1s;
wire[1:0] Tile_X10Y0_to_SI_1s;
wire[3:0] Tile_X0Y1_to_EA;
wire[3:0] Tile_X0Y1_to_EB;
wire[3:0] Tile_X0Y1_to_EC;
wire[3:0] Tile_X0Y1_to_ED;
wire[3:0] Tile_X0Y1_to_EF;
wire[7:0] Tile_X0Y1_to_EG;
wire[7:0] Tile_X0Y1_to_EH;
wire[11:0] Tile_X0Y1_to_EI;
wire[3:0] Tile_X0Y1_to_NA;
wire[3:0] Tile_X0Y1_to_NB;
wire[3:0] Tile_X0Y1_to_NC;
wire[3:0] Tile_X0Y1_to_ND;
wire[3:0] Tile_X0Y1_to_NF;
wire[7:0] Tile_X0Y1_to_NG;
wire[7:0] Tile_X0Y1_to_NH;
wire[11:0] Tile_X0Y1_to_NI;
wire[3:0] Tile_X0Y1_to_SA;
wire[3:0] Tile_X0Y1_to_SB;
wire[3:0] Tile_X0Y1_to_SC;
wire[3:0] Tile_X0Y1_to_SD;
wire[3:0] Tile_X0Y1_to_SF;
wire[7:0] Tile_X0Y1_to_SG;
wire[7:0] Tile_X0Y1_to_SH;
wire[11:0] Tile_X0Y1_to_SI;
wire[3:0] Tile_X1Y1_to_EA;
wire[3:0] Tile_X1Y1_to_EB;
wire[3:0] Tile_X1Y1_to_EC;
wire[3:0] Tile_X1Y1_to_ED;
wire[3:0] Tile_X1Y1_to_EF;
wire[7:0] Tile_X1Y1_to_EG;
wire[7:0] Tile_X1Y1_to_EH;
wire[11:0] Tile_X1Y1_to_EI;
wire[3:0] Tile_X1Y1_to_WA;
wire[3:0] Tile_X1Y1_to_WB;
wire[3:0] Tile_X1Y1_to_WC;
wire[3:0] Tile_X1Y1_to_WD;
wire[3:0] Tile_X1Y1_to_WF;
wire[7:0] Tile_X1Y1_to_WG;
wire[7:0] Tile_X1Y1_to_WH;
wire[11:0] Tile_X1Y1_to_WI;
wire[3:0] Tile_X1Y1_to_NA;
wire[3:0] Tile_X1Y1_to_NB;
wire[3:0] Tile_X1Y1_to_NC;
wire[3:0] Tile_X1Y1_to_ND;
wire[3:0] Tile_X1Y1_to_NF;
wire[7:0] Tile_X1Y1_to_NG;
wire[7:0] Tile_X1Y1_to_NH;
wire[11:0] Tile_X1Y1_to_NI;
wire[3:0] Tile_X1Y1_to_SA;
wire[3:0] Tile_X1Y1_to_SB;
wire[3:0] Tile_X1Y1_to_SC;
wire[3:0] Tile_X1Y1_to_SD;
wire[3:0] Tile_X1Y1_to_SF;
wire[7:0] Tile_X1Y1_to_SG;
wire[7:0] Tile_X1Y1_to_SH;
wire[11:0] Tile_X1Y1_to_SI;
wire[3:0] Tile_X2Y1_to_EA;
wire[3:0] Tile_X2Y1_to_EB;
wire[3:0] Tile_X2Y1_to_EC;
wire[3:0] Tile_X2Y1_to_ED;
wire[3:0] Tile_X2Y1_to_EF;
wire[7:0] Tile_X2Y1_to_EG;
wire[7:0] Tile_X2Y1_to_EH;
wire[11:0] Tile_X2Y1_to_EI;
wire[3:0] Tile_X2Y1_to_WA;
wire[3:0] Tile_X2Y1_to_WB;
wire[3:0] Tile_X2Y1_to_WC;
wire[3:0] Tile_X2Y1_to_WD;
wire[3:0] Tile_X2Y1_to_WF;
wire[7:0] Tile_X2Y1_to_WG;
wire[7:0] Tile_X2Y1_to_WH;
wire[11:0] Tile_X2Y1_to_WI;
wire[3:0] Tile_X2Y1_to_NA;
wire[3:0] Tile_X2Y1_to_NB;
wire[3:0] Tile_X2Y1_to_NC;
wire[3:0] Tile_X2Y1_to_ND;
wire[3:0] Tile_X2Y1_to_NF;
wire[7:0] Tile_X2Y1_to_NG;
wire[7:0] Tile_X2Y1_to_NH;
wire[11:0] Tile_X2Y1_to_NI;
wire[3:0] Tile_X2Y1_to_SA;
wire[3:0] Tile_X2Y1_to_SB;
wire[3:0] Tile_X2Y1_to_SC;
wire[3:0] Tile_X2Y1_to_SD;
wire[3:0] Tile_X2Y1_to_SF;
wire[7:0] Tile_X2Y1_to_SG;
wire[7:0] Tile_X2Y1_to_SH;
wire[11:0] Tile_X2Y1_to_SI;
wire[3:0] Tile_X3Y1_to_EA;
wire[3:0] Tile_X3Y1_to_EB;
wire[3:0] Tile_X3Y1_to_EC;
wire[3:0] Tile_X3Y1_to_ED;
wire[3:0] Tile_X3Y1_to_EF;
wire[7:0] Tile_X3Y1_to_EG;
wire[7:0] Tile_X3Y1_to_EH;
wire[11:0] Tile_X3Y1_to_EI;
wire[3:0] Tile_X3Y1_to_WA;
wire[3:0] Tile_X3Y1_to_WB;
wire[3:0] Tile_X3Y1_to_WC;
wire[3:0] Tile_X3Y1_to_WD;
wire[3:0] Tile_X3Y1_to_WF;
wire[7:0] Tile_X3Y1_to_WG;
wire[7:0] Tile_X3Y1_to_WH;
wire[11:0] Tile_X3Y1_to_WI;
wire[3:0] Tile_X3Y1_to_NA;
wire[3:0] Tile_X3Y1_to_NB;
wire[3:0] Tile_X3Y1_to_NC;
wire[3:0] Tile_X3Y1_to_ND;
wire[3:0] Tile_X3Y1_to_NF;
wire[7:0] Tile_X3Y1_to_NG;
wire[7:0] Tile_X3Y1_to_NH;
wire[11:0] Tile_X3Y1_to_NI;
wire[3:0] Tile_X3Y1_to_SA;
wire[3:0] Tile_X3Y1_to_SB;
wire[3:0] Tile_X3Y1_to_SC;
wire[3:0] Tile_X3Y1_to_SD;
wire[3:0] Tile_X3Y1_to_SF;
wire[7:0] Tile_X3Y1_to_SG;
wire[7:0] Tile_X3Y1_to_SH;
wire[11:0] Tile_X3Y1_to_SI;
wire[3:0] Tile_X4Y1_to_EA;
wire[3:0] Tile_X4Y1_to_EB;
wire[3:0] Tile_X4Y1_to_EC;
wire[3:0] Tile_X4Y1_to_ED;
wire[3:0] Tile_X4Y1_to_EF;
wire[7:0] Tile_X4Y1_to_EG;
wire[7:0] Tile_X4Y1_to_EH;
wire[11:0] Tile_X4Y1_to_EI;
wire[3:0] Tile_X4Y1_to_WA;
wire[3:0] Tile_X4Y1_to_WB;
wire[3:0] Tile_X4Y1_to_WC;
wire[3:0] Tile_X4Y1_to_WD;
wire[3:0] Tile_X4Y1_to_WF;
wire[7:0] Tile_X4Y1_to_WG;
wire[7:0] Tile_X4Y1_to_WH;
wire[11:0] Tile_X4Y1_to_WI;
wire[3:0] Tile_X4Y1_to_NA;
wire[3:0] Tile_X4Y1_to_NB;
wire[3:0] Tile_X4Y1_to_NC;
wire[3:0] Tile_X4Y1_to_ND;
wire[3:0] Tile_X4Y1_to_NF;
wire[7:0] Tile_X4Y1_to_NG;
wire[7:0] Tile_X4Y1_to_NH;
wire[11:0] Tile_X4Y1_to_NI;
wire[3:0] Tile_X4Y1_to_SA;
wire[3:0] Tile_X4Y1_to_SB;
wire[3:0] Tile_X4Y1_to_SC;
wire[3:0] Tile_X4Y1_to_SD;
wire[3:0] Tile_X4Y1_to_SF;
wire[7:0] Tile_X4Y1_to_SG;
wire[7:0] Tile_X4Y1_to_SH;
wire[11:0] Tile_X4Y1_to_SI;
wire[3:0] Tile_X5Y1_to_EA;
wire[3:0] Tile_X5Y1_to_EB;
wire[3:0] Tile_X5Y1_to_EC;
wire[3:0] Tile_X5Y1_to_ED;
wire[3:0] Tile_X5Y1_to_EF;
wire[7:0] Tile_X5Y1_to_EG;
wire[7:0] Tile_X5Y1_to_EH;
wire[11:0] Tile_X5Y1_to_EI;
wire[3:0] Tile_X5Y1_to_WA;
wire[3:0] Tile_X5Y1_to_WB;
wire[3:0] Tile_X5Y1_to_WC;
wire[3:0] Tile_X5Y1_to_WD;
wire[3:0] Tile_X5Y1_to_WF;
wire[7:0] Tile_X5Y1_to_WG;
wire[7:0] Tile_X5Y1_to_WH;
wire[11:0] Tile_X5Y1_to_WI;
wire[3:0] Tile_X5Y1_to_NA;
wire[3:0] Tile_X5Y1_to_NB;
wire[3:0] Tile_X5Y1_to_NC;
wire[3:0] Tile_X5Y1_to_ND;
wire[3:0] Tile_X5Y1_to_NF;
wire[7:0] Tile_X5Y1_to_NG;
wire[7:0] Tile_X5Y1_to_NH;
wire[11:0] Tile_X5Y1_to_NI;
wire[3:0] Tile_X5Y1_to_SA;
wire[3:0] Tile_X5Y1_to_SB;
wire[3:0] Tile_X5Y1_to_SC;
wire[3:0] Tile_X5Y1_to_SD;
wire[3:0] Tile_X5Y1_to_SF;
wire[7:0] Tile_X5Y1_to_SG;
wire[7:0] Tile_X5Y1_to_SH;
wire[11:0] Tile_X5Y1_to_SI;
wire[3:0] Tile_X6Y1_to_EA;
wire[3:0] Tile_X6Y1_to_EB;
wire[3:0] Tile_X6Y1_to_EC;
wire[3:0] Tile_X6Y1_to_ED;
wire[3:0] Tile_X6Y1_to_EF;
wire[7:0] Tile_X6Y1_to_EG;
wire[7:0] Tile_X6Y1_to_EH;
wire[11:0] Tile_X6Y1_to_EI;
wire[3:0] Tile_X6Y1_to_WA;
wire[3:0] Tile_X6Y1_to_WB;
wire[3:0] Tile_X6Y1_to_WC;
wire[3:0] Tile_X6Y1_to_WD;
wire[3:0] Tile_X6Y1_to_WF;
wire[7:0] Tile_X6Y1_to_WG;
wire[7:0] Tile_X6Y1_to_WH;
wire[11:0] Tile_X6Y1_to_WI;
wire[3:0] Tile_X6Y1_to_NA;
wire[3:0] Tile_X6Y1_to_NB;
wire[3:0] Tile_X6Y1_to_NC;
wire[3:0] Tile_X6Y1_to_ND;
wire[3:0] Tile_X6Y1_to_NF;
wire[7:0] Tile_X6Y1_to_NG;
wire[7:0] Tile_X6Y1_to_NH;
wire[11:0] Tile_X6Y1_to_NI;
wire[3:0] Tile_X6Y1_to_SA;
wire[3:0] Tile_X6Y1_to_SB;
wire[3:0] Tile_X6Y1_to_SC;
wire[3:0] Tile_X6Y1_to_SD;
wire[3:0] Tile_X6Y1_to_SF;
wire[7:0] Tile_X6Y1_to_SG;
wire[7:0] Tile_X6Y1_to_SH;
wire[11:0] Tile_X6Y1_to_SI;
wire[3:0] Tile_X7Y1_to_EA;
wire[3:0] Tile_X7Y1_to_EB;
wire[3:0] Tile_X7Y1_to_EC;
wire[3:0] Tile_X7Y1_to_ED;
wire[3:0] Tile_X7Y1_to_EF;
wire[7:0] Tile_X7Y1_to_EG;
wire[7:0] Tile_X7Y1_to_EH;
wire[11:0] Tile_X7Y1_to_EI;
wire[3:0] Tile_X7Y1_to_WA;
wire[3:0] Tile_X7Y1_to_WB;
wire[3:0] Tile_X7Y1_to_WC;
wire[3:0] Tile_X7Y1_to_WD;
wire[3:0] Tile_X7Y1_to_WF;
wire[7:0] Tile_X7Y1_to_WG;
wire[7:0] Tile_X7Y1_to_WH;
wire[11:0] Tile_X7Y1_to_WI;
wire[3:0] Tile_X7Y1_to_NA;
wire[3:0] Tile_X7Y1_to_NB;
wire[3:0] Tile_X7Y1_to_NC;
wire[3:0] Tile_X7Y1_to_ND;
wire[3:0] Tile_X7Y1_to_NF;
wire[7:0] Tile_X7Y1_to_NG;
wire[7:0] Tile_X7Y1_to_NH;
wire[11:0] Tile_X7Y1_to_NI;
wire[3:0] Tile_X7Y1_to_SA;
wire[3:0] Tile_X7Y1_to_SB;
wire[3:0] Tile_X7Y1_to_SC;
wire[3:0] Tile_X7Y1_to_SD;
wire[3:0] Tile_X7Y1_to_SF;
wire[7:0] Tile_X7Y1_to_SG;
wire[7:0] Tile_X7Y1_to_SH;
wire[11:0] Tile_X7Y1_to_SI;
wire[3:0] Tile_X8Y1_to_WA;
wire[3:0] Tile_X8Y1_to_WB;
wire[3:0] Tile_X8Y1_to_WC;
wire[3:0] Tile_X8Y1_to_WD;
wire[3:0] Tile_X8Y1_to_WF;
wire[7:0] Tile_X8Y1_to_WG;
wire[7:0] Tile_X8Y1_to_WH;
wire[11:0] Tile_X8Y1_to_WI;
wire[3:0] Tile_X8Y1_to_NA;
wire[3:0] Tile_X8Y1_to_NB;
wire[3:0] Tile_X8Y1_to_NC;
wire[3:0] Tile_X8Y1_to_ND;
wire[3:0] Tile_X8Y1_to_NF;
wire[7:0] Tile_X8Y1_to_NG;
wire[7:0] Tile_X8Y1_to_NH;
wire[11:0] Tile_X8Y1_to_NI;
wire[3:0] Tile_X8Y1_to_SA;
wire[3:0] Tile_X8Y1_to_SB;
wire[3:0] Tile_X8Y1_to_SC;
wire[3:0] Tile_X8Y1_to_SD;
wire[3:0] Tile_X8Y1_to_SF;
wire[7:0] Tile_X8Y1_to_SG;
wire[7:0] Tile_X8Y1_to_SH;
wire[11:0] Tile_X8Y1_to_SI;
wire[1:0] Tile_X9Y1_to_EA_1s;
wire[1:0] Tile_X9Y1_to_EB_1s;
wire[1:0] Tile_X9Y1_to_EC_1s;
wire[1:0] Tile_X9Y1_to_ED_1s;
wire[1:0] Tile_X9Y1_to_EF_1s;
wire[1:0] Tile_X9Y1_to_EG_1s;
wire[1:0] Tile_X9Y1_to_EH_1s;
wire[1:0] Tile_X9Y1_to_EI_1s;
wire[1:0] Tile_X9Y1_to_WA_1s;
wire[1:0] Tile_X9Y1_to_WB_1s;
wire[1:0] Tile_X9Y1_to_WC_1s;
wire[1:0] Tile_X9Y1_to_WD_1s;
wire[1:0] Tile_X9Y1_to_WF_1s;
wire[1:0] Tile_X9Y1_to_WG_1s;
wire[1:0] Tile_X9Y1_to_WH_1s;
wire[1:0] Tile_X9Y1_to_WI_1s;
wire[1:0] Tile_X9Y1_to_NA_1s;
wire[1:0] Tile_X9Y1_to_NB_1s;
wire[1:0] Tile_X9Y1_to_NC_1s;
wire[1:0] Tile_X9Y1_to_ND_1s;
wire[1:0] Tile_X9Y1_to_NF_1s;
wire[1:0] Tile_X9Y1_to_NG_1s;
wire[1:0] Tile_X9Y1_to_NH_1s;
wire[1:0] Tile_X9Y1_to_NI_1s;
wire[1:0] Tile_X9Y1_to_SA_1s;
wire[1:0] Tile_X9Y1_to_SB_1s;
wire[1:0] Tile_X9Y1_to_SC_1s;
wire[1:0] Tile_X9Y1_to_SD_1s;
wire[1:0] Tile_X9Y1_to_SF_1s;
wire[1:0] Tile_X9Y1_to_SG_1s;
wire[1:0] Tile_X9Y1_to_SH_1s;
wire[1:0] Tile_X9Y1_to_SI_1s;
wire[1:0] Tile_X10Y1_to_WA_1s;
wire[1:0] Tile_X10Y1_to_WB_1s;
wire[1:0] Tile_X10Y1_to_WC_1s;
wire[1:0] Tile_X10Y1_to_WD_1s;
wire[1:0] Tile_X10Y1_to_WF_1s;
wire[1:0] Tile_X10Y1_to_WG_1s;
wire[1:0] Tile_X10Y1_to_WH_1s;
wire[1:0] Tile_X10Y1_to_WI_1s;
wire[3:0] Tile_X0Y2_to_EA;
wire[3:0] Tile_X0Y2_to_EB;
wire[3:0] Tile_X0Y2_to_EC;
wire[3:0] Tile_X0Y2_to_ED;
wire[3:0] Tile_X0Y2_to_EF;
wire[7:0] Tile_X0Y2_to_EG;
wire[7:0] Tile_X0Y2_to_EH;
wire[11:0] Tile_X0Y2_to_EI;
wire[3:0] Tile_X0Y2_to_NA;
wire[3:0] Tile_X0Y2_to_NB;
wire[3:0] Tile_X0Y2_to_NC;
wire[3:0] Tile_X0Y2_to_ND;
wire[3:0] Tile_X0Y2_to_NF;
wire[7:0] Tile_X0Y2_to_NG;
wire[7:0] Tile_X0Y2_to_NH;
wire[11:0] Tile_X0Y2_to_NI;
wire[3:0] Tile_X0Y2_to_SA;
wire[3:0] Tile_X0Y2_to_SB;
wire[3:0] Tile_X0Y2_to_SC;
wire[3:0] Tile_X0Y2_to_SD;
wire[3:0] Tile_X0Y2_to_SF;
wire[7:0] Tile_X0Y2_to_SG;
wire[7:0] Tile_X0Y2_to_SH;
wire[11:0] Tile_X0Y2_to_SI;
wire[3:0] Tile_X1Y2_to_EA;
wire[3:0] Tile_X1Y2_to_EB;
wire[3:0] Tile_X1Y2_to_EC;
wire[3:0] Tile_X1Y2_to_ED;
wire[3:0] Tile_X1Y2_to_EF;
wire[7:0] Tile_X1Y2_to_EG;
wire[7:0] Tile_X1Y2_to_EH;
wire[11:0] Tile_X1Y2_to_EI;
wire[3:0] Tile_X1Y2_to_WA;
wire[3:0] Tile_X1Y2_to_WB;
wire[3:0] Tile_X1Y2_to_WC;
wire[3:0] Tile_X1Y2_to_WD;
wire[3:0] Tile_X1Y2_to_WF;
wire[7:0] Tile_X1Y2_to_WG;
wire[7:0] Tile_X1Y2_to_WH;
wire[11:0] Tile_X1Y2_to_WI;
wire[3:0] Tile_X1Y2_to_NA;
wire[3:0] Tile_X1Y2_to_NB;
wire[3:0] Tile_X1Y2_to_NC;
wire[3:0] Tile_X1Y2_to_ND;
wire[3:0] Tile_X1Y2_to_NF;
wire[7:0] Tile_X1Y2_to_NG;
wire[7:0] Tile_X1Y2_to_NH;
wire[11:0] Tile_X1Y2_to_NI;
wire[3:0] Tile_X1Y2_to_SA;
wire[3:0] Tile_X1Y2_to_SB;
wire[3:0] Tile_X1Y2_to_SC;
wire[3:0] Tile_X1Y2_to_SD;
wire[3:0] Tile_X1Y2_to_SF;
wire[7:0] Tile_X1Y2_to_SG;
wire[7:0] Tile_X1Y2_to_SH;
wire[11:0] Tile_X1Y2_to_SI;
wire[3:0] Tile_X2Y2_to_EA;
wire[3:0] Tile_X2Y2_to_EB;
wire[3:0] Tile_X2Y2_to_EC;
wire[3:0] Tile_X2Y2_to_ED;
wire[3:0] Tile_X2Y2_to_EF;
wire[7:0] Tile_X2Y2_to_EG;
wire[7:0] Tile_X2Y2_to_EH;
wire[11:0] Tile_X2Y2_to_EI;
wire[3:0] Tile_X2Y2_to_WA;
wire[3:0] Tile_X2Y2_to_WB;
wire[3:0] Tile_X2Y2_to_WC;
wire[3:0] Tile_X2Y2_to_WD;
wire[3:0] Tile_X2Y2_to_WF;
wire[7:0] Tile_X2Y2_to_WG;
wire[7:0] Tile_X2Y2_to_WH;
wire[11:0] Tile_X2Y2_to_WI;
wire[3:0] Tile_X2Y2_to_NA;
wire[3:0] Tile_X2Y2_to_NB;
wire[3:0] Tile_X2Y2_to_NC;
wire[3:0] Tile_X2Y2_to_ND;
wire[3:0] Tile_X2Y2_to_NF;
wire[7:0] Tile_X2Y2_to_NG;
wire[7:0] Tile_X2Y2_to_NH;
wire[11:0] Tile_X2Y2_to_NI;
wire[3:0] Tile_X2Y2_to_SA;
wire[3:0] Tile_X2Y2_to_SB;
wire[3:0] Tile_X2Y2_to_SC;
wire[3:0] Tile_X2Y2_to_SD;
wire[3:0] Tile_X2Y2_to_SF;
wire[7:0] Tile_X2Y2_to_SG;
wire[7:0] Tile_X2Y2_to_SH;
wire[11:0] Tile_X2Y2_to_SI;
wire[3:0] Tile_X3Y2_to_EA;
wire[3:0] Tile_X3Y2_to_EB;
wire[3:0] Tile_X3Y2_to_EC;
wire[3:0] Tile_X3Y2_to_ED;
wire[3:0] Tile_X3Y2_to_EF;
wire[7:0] Tile_X3Y2_to_EG;
wire[7:0] Tile_X3Y2_to_EH;
wire[11:0] Tile_X3Y2_to_EI;
wire[3:0] Tile_X3Y2_to_WA;
wire[3:0] Tile_X3Y2_to_WB;
wire[3:0] Tile_X3Y2_to_WC;
wire[3:0] Tile_X3Y2_to_WD;
wire[3:0] Tile_X3Y2_to_WF;
wire[7:0] Tile_X3Y2_to_WG;
wire[7:0] Tile_X3Y2_to_WH;
wire[11:0] Tile_X3Y2_to_WI;
wire[3:0] Tile_X3Y2_to_NA;
wire[3:0] Tile_X3Y2_to_NB;
wire[3:0] Tile_X3Y2_to_NC;
wire[3:0] Tile_X3Y2_to_ND;
wire[3:0] Tile_X3Y2_to_NF;
wire[7:0] Tile_X3Y2_to_NG;
wire[7:0] Tile_X3Y2_to_NH;
wire[11:0] Tile_X3Y2_to_NI;
wire[3:0] Tile_X3Y2_to_SA;
wire[3:0] Tile_X3Y2_to_SB;
wire[3:0] Tile_X3Y2_to_SC;
wire[3:0] Tile_X3Y2_to_SD;
wire[3:0] Tile_X3Y2_to_SF;
wire[7:0] Tile_X3Y2_to_SG;
wire[7:0] Tile_X3Y2_to_SH;
wire[11:0] Tile_X3Y2_to_SI;
wire[3:0] Tile_X4Y2_to_EA;
wire[3:0] Tile_X4Y2_to_EB;
wire[3:0] Tile_X4Y2_to_EC;
wire[3:0] Tile_X4Y2_to_ED;
wire[3:0] Tile_X4Y2_to_EF;
wire[7:0] Tile_X4Y2_to_EG;
wire[7:0] Tile_X4Y2_to_EH;
wire[11:0] Tile_X4Y2_to_EI;
wire[3:0] Tile_X4Y2_to_WA;
wire[3:0] Tile_X4Y2_to_WB;
wire[3:0] Tile_X4Y2_to_WC;
wire[3:0] Tile_X4Y2_to_WD;
wire[3:0] Tile_X4Y2_to_WF;
wire[7:0] Tile_X4Y2_to_WG;
wire[7:0] Tile_X4Y2_to_WH;
wire[11:0] Tile_X4Y2_to_WI;
wire[3:0] Tile_X4Y2_to_NA;
wire[3:0] Tile_X4Y2_to_NB;
wire[3:0] Tile_X4Y2_to_NC;
wire[3:0] Tile_X4Y2_to_ND;
wire[3:0] Tile_X4Y2_to_NF;
wire[7:0] Tile_X4Y2_to_NG;
wire[7:0] Tile_X4Y2_to_NH;
wire[11:0] Tile_X4Y2_to_NI;
wire[3:0] Tile_X4Y2_to_SA;
wire[3:0] Tile_X4Y2_to_SB;
wire[3:0] Tile_X4Y2_to_SC;
wire[3:0] Tile_X4Y2_to_SD;
wire[3:0] Tile_X4Y2_to_SF;
wire[7:0] Tile_X4Y2_to_SG;
wire[7:0] Tile_X4Y2_to_SH;
wire[11:0] Tile_X4Y2_to_SI;
wire[3:0] Tile_X5Y2_to_EA;
wire[3:0] Tile_X5Y2_to_EB;
wire[3:0] Tile_X5Y2_to_EC;
wire[3:0] Tile_X5Y2_to_ED;
wire[3:0] Tile_X5Y2_to_EF;
wire[7:0] Tile_X5Y2_to_EG;
wire[7:0] Tile_X5Y2_to_EH;
wire[11:0] Tile_X5Y2_to_EI;
wire[3:0] Tile_X5Y2_to_WA;
wire[3:0] Tile_X5Y2_to_WB;
wire[3:0] Tile_X5Y2_to_WC;
wire[3:0] Tile_X5Y2_to_WD;
wire[3:0] Tile_X5Y2_to_WF;
wire[7:0] Tile_X5Y2_to_WG;
wire[7:0] Tile_X5Y2_to_WH;
wire[11:0] Tile_X5Y2_to_WI;
wire[3:0] Tile_X5Y2_to_NA;
wire[3:0] Tile_X5Y2_to_NB;
wire[3:0] Tile_X5Y2_to_NC;
wire[3:0] Tile_X5Y2_to_ND;
wire[3:0] Tile_X5Y2_to_NF;
wire[7:0] Tile_X5Y2_to_NG;
wire[7:0] Tile_X5Y2_to_NH;
wire[11:0] Tile_X5Y2_to_NI;
wire[3:0] Tile_X5Y2_to_SA;
wire[3:0] Tile_X5Y2_to_SB;
wire[3:0] Tile_X5Y2_to_SC;
wire[3:0] Tile_X5Y2_to_SD;
wire[3:0] Tile_X5Y2_to_SF;
wire[7:0] Tile_X5Y2_to_SG;
wire[7:0] Tile_X5Y2_to_SH;
wire[11:0] Tile_X5Y2_to_SI;
wire[3:0] Tile_X6Y2_to_EA;
wire[3:0] Tile_X6Y2_to_EB;
wire[3:0] Tile_X6Y2_to_EC;
wire[3:0] Tile_X6Y2_to_ED;
wire[3:0] Tile_X6Y2_to_EF;
wire[7:0] Tile_X6Y2_to_EG;
wire[7:0] Tile_X6Y2_to_EH;
wire[11:0] Tile_X6Y2_to_EI;
wire[3:0] Tile_X6Y2_to_WA;
wire[3:0] Tile_X6Y2_to_WB;
wire[3:0] Tile_X6Y2_to_WC;
wire[3:0] Tile_X6Y2_to_WD;
wire[3:0] Tile_X6Y2_to_WF;
wire[7:0] Tile_X6Y2_to_WG;
wire[7:0] Tile_X6Y2_to_WH;
wire[11:0] Tile_X6Y2_to_WI;
wire[3:0] Tile_X6Y2_to_NA;
wire[3:0] Tile_X6Y2_to_NB;
wire[3:0] Tile_X6Y2_to_NC;
wire[3:0] Tile_X6Y2_to_ND;
wire[3:0] Tile_X6Y2_to_NF;
wire[7:0] Tile_X6Y2_to_NG;
wire[7:0] Tile_X6Y2_to_NH;
wire[11:0] Tile_X6Y2_to_NI;
wire[3:0] Tile_X6Y2_to_SA;
wire[3:0] Tile_X6Y2_to_SB;
wire[3:0] Tile_X6Y2_to_SC;
wire[3:0] Tile_X6Y2_to_SD;
wire[3:0] Tile_X6Y2_to_SF;
wire[7:0] Tile_X6Y2_to_SG;
wire[7:0] Tile_X6Y2_to_SH;
wire[11:0] Tile_X6Y2_to_SI;
wire[3:0] Tile_X7Y2_to_EA;
wire[3:0] Tile_X7Y2_to_EB;
wire[3:0] Tile_X7Y2_to_EC;
wire[3:0] Tile_X7Y2_to_ED;
wire[3:0] Tile_X7Y2_to_EF;
wire[7:0] Tile_X7Y2_to_EG;
wire[7:0] Tile_X7Y2_to_EH;
wire[11:0] Tile_X7Y2_to_EI;
wire[3:0] Tile_X7Y2_to_WA;
wire[3:0] Tile_X7Y2_to_WB;
wire[3:0] Tile_X7Y2_to_WC;
wire[3:0] Tile_X7Y2_to_WD;
wire[3:0] Tile_X7Y2_to_WF;
wire[7:0] Tile_X7Y2_to_WG;
wire[7:0] Tile_X7Y2_to_WH;
wire[11:0] Tile_X7Y2_to_WI;
wire[3:0] Tile_X7Y2_to_NA;
wire[3:0] Tile_X7Y2_to_NB;
wire[3:0] Tile_X7Y2_to_NC;
wire[3:0] Tile_X7Y2_to_ND;
wire[3:0] Tile_X7Y2_to_NF;
wire[7:0] Tile_X7Y2_to_NG;
wire[7:0] Tile_X7Y2_to_NH;
wire[11:0] Tile_X7Y2_to_NI;
wire[3:0] Tile_X7Y2_to_SA;
wire[3:0] Tile_X7Y2_to_SB;
wire[3:0] Tile_X7Y2_to_SC;
wire[3:0] Tile_X7Y2_to_SD;
wire[3:0] Tile_X7Y2_to_SF;
wire[7:0] Tile_X7Y2_to_SG;
wire[7:0] Tile_X7Y2_to_SH;
wire[11:0] Tile_X7Y2_to_SI;
wire[3:0] Tile_X8Y2_to_WA;
wire[3:0] Tile_X8Y2_to_WB;
wire[3:0] Tile_X8Y2_to_WC;
wire[3:0] Tile_X8Y2_to_WD;
wire[3:0] Tile_X8Y2_to_WF;
wire[7:0] Tile_X8Y2_to_WG;
wire[7:0] Tile_X8Y2_to_WH;
wire[11:0] Tile_X8Y2_to_WI;
wire[3:0] Tile_X8Y2_to_NA;
wire[3:0] Tile_X8Y2_to_NB;
wire[3:0] Tile_X8Y2_to_NC;
wire[3:0] Tile_X8Y2_to_ND;
wire[3:0] Tile_X8Y2_to_NF;
wire[7:0] Tile_X8Y2_to_NG;
wire[7:0] Tile_X8Y2_to_NH;
wire[11:0] Tile_X8Y2_to_NI;
wire[3:0] Tile_X8Y2_to_SA;
wire[3:0] Tile_X8Y2_to_SB;
wire[3:0] Tile_X8Y2_to_SC;
wire[3:0] Tile_X8Y2_to_SD;
wire[3:0] Tile_X8Y2_to_SF;
wire[7:0] Tile_X8Y2_to_SG;
wire[7:0] Tile_X8Y2_to_SH;
wire[11:0] Tile_X8Y2_to_SI;
wire[1:0] Tile_X9Y2_to_EA_1s;
wire[1:0] Tile_X9Y2_to_EB_1s;
wire[1:0] Tile_X9Y2_to_EC_1s;
wire[1:0] Tile_X9Y2_to_ED_1s;
wire[1:0] Tile_X9Y2_to_EF_1s;
wire[1:0] Tile_X9Y2_to_EG_1s;
wire[1:0] Tile_X9Y2_to_EH_1s;
wire[1:0] Tile_X9Y2_to_EI_1s;
wire[1:0] Tile_X9Y2_to_WA_1s;
wire[1:0] Tile_X9Y2_to_WB_1s;
wire[1:0] Tile_X9Y2_to_WC_1s;
wire[1:0] Tile_X9Y2_to_WD_1s;
wire[1:0] Tile_X9Y2_to_WF_1s;
wire[1:0] Tile_X9Y2_to_WG_1s;
wire[1:0] Tile_X9Y2_to_WH_1s;
wire[1:0] Tile_X9Y2_to_WI_1s;
wire[1:0] Tile_X9Y2_to_NA_1s;
wire[1:0] Tile_X9Y2_to_NB_1s;
wire[1:0] Tile_X9Y2_to_NC_1s;
wire[1:0] Tile_X9Y2_to_ND_1s;
wire[1:0] Tile_X9Y2_to_NF_1s;
wire[1:0] Tile_X9Y2_to_NG_1s;
wire[1:0] Tile_X9Y2_to_NH_1s;
wire[1:0] Tile_X9Y2_to_NI_1s;
wire[1:0] Tile_X9Y2_to_SA_1s;
wire[1:0] Tile_X9Y2_to_SB_1s;
wire[1:0] Tile_X9Y2_to_SC_1s;
wire[1:0] Tile_X9Y2_to_SD_1s;
wire[1:0] Tile_X9Y2_to_SF_1s;
wire[1:0] Tile_X9Y2_to_SG_1s;
wire[1:0] Tile_X9Y2_to_SH_1s;
wire[1:0] Tile_X9Y2_to_SI_1s;
wire[1:0] Tile_X10Y2_to_WA_1s;
wire[1:0] Tile_X10Y2_to_WB_1s;
wire[1:0] Tile_X10Y2_to_WC_1s;
wire[1:0] Tile_X10Y2_to_WD_1s;
wire[1:0] Tile_X10Y2_to_WF_1s;
wire[1:0] Tile_X10Y2_to_WG_1s;
wire[1:0] Tile_X10Y2_to_WH_1s;
wire[1:0] Tile_X10Y2_to_WI_1s;
wire[3:0] Tile_X0Y3_to_EA;
wire[3:0] Tile_X0Y3_to_EB;
wire[3:0] Tile_X0Y3_to_EC;
wire[3:0] Tile_X0Y3_to_ED;
wire[3:0] Tile_X0Y3_to_EF;
wire[7:0] Tile_X0Y3_to_EG;
wire[7:0] Tile_X0Y3_to_EH;
wire[11:0] Tile_X0Y3_to_EI;
wire[3:0] Tile_X0Y3_to_NA;
wire[3:0] Tile_X0Y3_to_NB;
wire[3:0] Tile_X0Y3_to_NC;
wire[3:0] Tile_X0Y3_to_ND;
wire[3:0] Tile_X0Y3_to_NF;
wire[7:0] Tile_X0Y3_to_NG;
wire[7:0] Tile_X0Y3_to_NH;
wire[11:0] Tile_X0Y3_to_NI;
wire[3:0] Tile_X0Y3_to_SA;
wire[3:0] Tile_X0Y3_to_SB;
wire[3:0] Tile_X0Y3_to_SC;
wire[3:0] Tile_X0Y3_to_SD;
wire[3:0] Tile_X0Y3_to_SF;
wire[7:0] Tile_X0Y3_to_SG;
wire[7:0] Tile_X0Y3_to_SH;
wire[11:0] Tile_X0Y3_to_SI;
wire[3:0] Tile_X1Y3_to_EA;
wire[3:0] Tile_X1Y3_to_EB;
wire[3:0] Tile_X1Y3_to_EC;
wire[3:0] Tile_X1Y3_to_ED;
wire[3:0] Tile_X1Y3_to_EF;
wire[7:0] Tile_X1Y3_to_EG;
wire[7:0] Tile_X1Y3_to_EH;
wire[11:0] Tile_X1Y3_to_EI;
wire[3:0] Tile_X1Y3_to_WA;
wire[3:0] Tile_X1Y3_to_WB;
wire[3:0] Tile_X1Y3_to_WC;
wire[3:0] Tile_X1Y3_to_WD;
wire[3:0] Tile_X1Y3_to_WF;
wire[7:0] Tile_X1Y3_to_WG;
wire[7:0] Tile_X1Y3_to_WH;
wire[11:0] Tile_X1Y3_to_WI;
wire[3:0] Tile_X1Y3_to_NA;
wire[3:0] Tile_X1Y3_to_NB;
wire[3:0] Tile_X1Y3_to_NC;
wire[3:0] Tile_X1Y3_to_ND;
wire[3:0] Tile_X1Y3_to_NF;
wire[7:0] Tile_X1Y3_to_NG;
wire[7:0] Tile_X1Y3_to_NH;
wire[11:0] Tile_X1Y3_to_NI;
wire[3:0] Tile_X1Y3_to_SA;
wire[3:0] Tile_X1Y3_to_SB;
wire[3:0] Tile_X1Y3_to_SC;
wire[3:0] Tile_X1Y3_to_SD;
wire[3:0] Tile_X1Y3_to_SF;
wire[7:0] Tile_X1Y3_to_SG;
wire[7:0] Tile_X1Y3_to_SH;
wire[11:0] Tile_X1Y3_to_SI;
wire[3:0] Tile_X2Y3_to_EA;
wire[3:0] Tile_X2Y3_to_EB;
wire[3:0] Tile_X2Y3_to_EC;
wire[3:0] Tile_X2Y3_to_ED;
wire[3:0] Tile_X2Y3_to_EF;
wire[7:0] Tile_X2Y3_to_EG;
wire[7:0] Tile_X2Y3_to_EH;
wire[11:0] Tile_X2Y3_to_EI;
wire[3:0] Tile_X2Y3_to_WA;
wire[3:0] Tile_X2Y3_to_WB;
wire[3:0] Tile_X2Y3_to_WC;
wire[3:0] Tile_X2Y3_to_WD;
wire[3:0] Tile_X2Y3_to_WF;
wire[7:0] Tile_X2Y3_to_WG;
wire[7:0] Tile_X2Y3_to_WH;
wire[11:0] Tile_X2Y3_to_WI;
wire[3:0] Tile_X2Y3_to_NA;
wire[3:0] Tile_X2Y3_to_NB;
wire[3:0] Tile_X2Y3_to_NC;
wire[3:0] Tile_X2Y3_to_ND;
wire[3:0] Tile_X2Y3_to_NF;
wire[7:0] Tile_X2Y3_to_NG;
wire[7:0] Tile_X2Y3_to_NH;
wire[11:0] Tile_X2Y3_to_NI;
wire[3:0] Tile_X2Y3_to_SA;
wire[3:0] Tile_X2Y3_to_SB;
wire[3:0] Tile_X2Y3_to_SC;
wire[3:0] Tile_X2Y3_to_SD;
wire[3:0] Tile_X2Y3_to_SF;
wire[7:0] Tile_X2Y3_to_SG;
wire[7:0] Tile_X2Y3_to_SH;
wire[11:0] Tile_X2Y3_to_SI;
wire[3:0] Tile_X3Y3_to_EA;
wire[3:0] Tile_X3Y3_to_EB;
wire[3:0] Tile_X3Y3_to_EC;
wire[3:0] Tile_X3Y3_to_ED;
wire[3:0] Tile_X3Y3_to_EF;
wire[7:0] Tile_X3Y3_to_EG;
wire[7:0] Tile_X3Y3_to_EH;
wire[11:0] Tile_X3Y3_to_EI;
wire[3:0] Tile_X3Y3_to_WA;
wire[3:0] Tile_X3Y3_to_WB;
wire[3:0] Tile_X3Y3_to_WC;
wire[3:0] Tile_X3Y3_to_WD;
wire[3:0] Tile_X3Y3_to_WF;
wire[7:0] Tile_X3Y3_to_WG;
wire[7:0] Tile_X3Y3_to_WH;
wire[11:0] Tile_X3Y3_to_WI;
wire[3:0] Tile_X3Y3_to_NA;
wire[3:0] Tile_X3Y3_to_NB;
wire[3:0] Tile_X3Y3_to_NC;
wire[3:0] Tile_X3Y3_to_ND;
wire[3:0] Tile_X3Y3_to_NF;
wire[7:0] Tile_X3Y3_to_NG;
wire[7:0] Tile_X3Y3_to_NH;
wire[11:0] Tile_X3Y3_to_NI;
wire[3:0] Tile_X3Y3_to_SA;
wire[3:0] Tile_X3Y3_to_SB;
wire[3:0] Tile_X3Y3_to_SC;
wire[3:0] Tile_X3Y3_to_SD;
wire[3:0] Tile_X3Y3_to_SF;
wire[7:0] Tile_X3Y3_to_SG;
wire[7:0] Tile_X3Y3_to_SH;
wire[11:0] Tile_X3Y3_to_SI;
wire[3:0] Tile_X4Y3_to_EA;
wire[3:0] Tile_X4Y3_to_EB;
wire[3:0] Tile_X4Y3_to_EC;
wire[3:0] Tile_X4Y3_to_ED;
wire[3:0] Tile_X4Y3_to_EF;
wire[7:0] Tile_X4Y3_to_EG;
wire[7:0] Tile_X4Y3_to_EH;
wire[11:0] Tile_X4Y3_to_EI;
wire[3:0] Tile_X4Y3_to_WA;
wire[3:0] Tile_X4Y3_to_WB;
wire[3:0] Tile_X4Y3_to_WC;
wire[3:0] Tile_X4Y3_to_WD;
wire[3:0] Tile_X4Y3_to_WF;
wire[7:0] Tile_X4Y3_to_WG;
wire[7:0] Tile_X4Y3_to_WH;
wire[11:0] Tile_X4Y3_to_WI;
wire[3:0] Tile_X4Y3_to_NA;
wire[3:0] Tile_X4Y3_to_NB;
wire[3:0] Tile_X4Y3_to_NC;
wire[3:0] Tile_X4Y3_to_ND;
wire[3:0] Tile_X4Y3_to_NF;
wire[7:0] Tile_X4Y3_to_NG;
wire[7:0] Tile_X4Y3_to_NH;
wire[11:0] Tile_X4Y3_to_NI;
wire[3:0] Tile_X4Y3_to_SA;
wire[3:0] Tile_X4Y3_to_SB;
wire[3:0] Tile_X4Y3_to_SC;
wire[3:0] Tile_X4Y3_to_SD;
wire[3:0] Tile_X4Y3_to_SF;
wire[7:0] Tile_X4Y3_to_SG;
wire[7:0] Tile_X4Y3_to_SH;
wire[11:0] Tile_X4Y3_to_SI;
wire[3:0] Tile_X5Y3_to_EA;
wire[3:0] Tile_X5Y3_to_EB;
wire[3:0] Tile_X5Y3_to_EC;
wire[3:0] Tile_X5Y3_to_ED;
wire[3:0] Tile_X5Y3_to_EF;
wire[7:0] Tile_X5Y3_to_EG;
wire[7:0] Tile_X5Y3_to_EH;
wire[11:0] Tile_X5Y3_to_EI;
wire[3:0] Tile_X5Y3_to_WA;
wire[3:0] Tile_X5Y3_to_WB;
wire[3:0] Tile_X5Y3_to_WC;
wire[3:0] Tile_X5Y3_to_WD;
wire[3:0] Tile_X5Y3_to_WF;
wire[7:0] Tile_X5Y3_to_WG;
wire[7:0] Tile_X5Y3_to_WH;
wire[11:0] Tile_X5Y3_to_WI;
wire[3:0] Tile_X5Y3_to_NA;
wire[3:0] Tile_X5Y3_to_NB;
wire[3:0] Tile_X5Y3_to_NC;
wire[3:0] Tile_X5Y3_to_ND;
wire[3:0] Tile_X5Y3_to_NF;
wire[7:0] Tile_X5Y3_to_NG;
wire[7:0] Tile_X5Y3_to_NH;
wire[11:0] Tile_X5Y3_to_NI;
wire[3:0] Tile_X5Y3_to_SA;
wire[3:0] Tile_X5Y3_to_SB;
wire[3:0] Tile_X5Y3_to_SC;
wire[3:0] Tile_X5Y3_to_SD;
wire[3:0] Tile_X5Y3_to_SF;
wire[7:0] Tile_X5Y3_to_SG;
wire[7:0] Tile_X5Y3_to_SH;
wire[11:0] Tile_X5Y3_to_SI;
wire[3:0] Tile_X6Y3_to_EA;
wire[3:0] Tile_X6Y3_to_EB;
wire[3:0] Tile_X6Y3_to_EC;
wire[3:0] Tile_X6Y3_to_ED;
wire[3:0] Tile_X6Y3_to_EF;
wire[7:0] Tile_X6Y3_to_EG;
wire[7:0] Tile_X6Y3_to_EH;
wire[11:0] Tile_X6Y3_to_EI;
wire[3:0] Tile_X6Y3_to_WA;
wire[3:0] Tile_X6Y3_to_WB;
wire[3:0] Tile_X6Y3_to_WC;
wire[3:0] Tile_X6Y3_to_WD;
wire[3:0] Tile_X6Y3_to_WF;
wire[7:0] Tile_X6Y3_to_WG;
wire[7:0] Tile_X6Y3_to_WH;
wire[11:0] Tile_X6Y3_to_WI;
wire[3:0] Tile_X6Y3_to_NA;
wire[3:0] Tile_X6Y3_to_NB;
wire[3:0] Tile_X6Y3_to_NC;
wire[3:0] Tile_X6Y3_to_ND;
wire[3:0] Tile_X6Y3_to_NF;
wire[7:0] Tile_X6Y3_to_NG;
wire[7:0] Tile_X6Y3_to_NH;
wire[11:0] Tile_X6Y3_to_NI;
wire[3:0] Tile_X6Y3_to_SA;
wire[3:0] Tile_X6Y3_to_SB;
wire[3:0] Tile_X6Y3_to_SC;
wire[3:0] Tile_X6Y3_to_SD;
wire[3:0] Tile_X6Y3_to_SF;
wire[7:0] Tile_X6Y3_to_SG;
wire[7:0] Tile_X6Y3_to_SH;
wire[11:0] Tile_X6Y3_to_SI;
wire[3:0] Tile_X7Y3_to_EA;
wire[3:0] Tile_X7Y3_to_EB;
wire[3:0] Tile_X7Y3_to_EC;
wire[3:0] Tile_X7Y3_to_ED;
wire[3:0] Tile_X7Y3_to_EF;
wire[7:0] Tile_X7Y3_to_EG;
wire[7:0] Tile_X7Y3_to_EH;
wire[11:0] Tile_X7Y3_to_EI;
wire[3:0] Tile_X7Y3_to_WA;
wire[3:0] Tile_X7Y3_to_WB;
wire[3:0] Tile_X7Y3_to_WC;
wire[3:0] Tile_X7Y3_to_WD;
wire[3:0] Tile_X7Y3_to_WF;
wire[7:0] Tile_X7Y3_to_WG;
wire[7:0] Tile_X7Y3_to_WH;
wire[11:0] Tile_X7Y3_to_WI;
wire[3:0] Tile_X7Y3_to_NA;
wire[3:0] Tile_X7Y3_to_NB;
wire[3:0] Tile_X7Y3_to_NC;
wire[3:0] Tile_X7Y3_to_ND;
wire[3:0] Tile_X7Y3_to_NF;
wire[7:0] Tile_X7Y3_to_NG;
wire[7:0] Tile_X7Y3_to_NH;
wire[11:0] Tile_X7Y3_to_NI;
wire[3:0] Tile_X7Y3_to_SA;
wire[3:0] Tile_X7Y3_to_SB;
wire[3:0] Tile_X7Y3_to_SC;
wire[3:0] Tile_X7Y3_to_SD;
wire[3:0] Tile_X7Y3_to_SF;
wire[7:0] Tile_X7Y3_to_SG;
wire[7:0] Tile_X7Y3_to_SH;
wire[11:0] Tile_X7Y3_to_SI;
wire[3:0] Tile_X8Y3_to_WA;
wire[3:0] Tile_X8Y3_to_WB;
wire[3:0] Tile_X8Y3_to_WC;
wire[3:0] Tile_X8Y3_to_WD;
wire[3:0] Tile_X8Y3_to_WF;
wire[7:0] Tile_X8Y3_to_WG;
wire[7:0] Tile_X8Y3_to_WH;
wire[11:0] Tile_X8Y3_to_WI;
wire[3:0] Tile_X8Y3_to_NA;
wire[3:0] Tile_X8Y3_to_NB;
wire[3:0] Tile_X8Y3_to_NC;
wire[3:0] Tile_X8Y3_to_ND;
wire[3:0] Tile_X8Y3_to_NF;
wire[7:0] Tile_X8Y3_to_NG;
wire[7:0] Tile_X8Y3_to_NH;
wire[11:0] Tile_X8Y3_to_NI;
wire[3:0] Tile_X8Y3_to_SA;
wire[3:0] Tile_X8Y3_to_SB;
wire[3:0] Tile_X8Y3_to_SC;
wire[3:0] Tile_X8Y3_to_SD;
wire[3:0] Tile_X8Y3_to_SF;
wire[7:0] Tile_X8Y3_to_SG;
wire[7:0] Tile_X8Y3_to_SH;
wire[11:0] Tile_X8Y3_to_SI;
wire[1:0] Tile_X9Y3_to_EA_1s;
wire[1:0] Tile_X9Y3_to_EB_1s;
wire[1:0] Tile_X9Y3_to_EC_1s;
wire[1:0] Tile_X9Y3_to_ED_1s;
wire[1:0] Tile_X9Y3_to_EF_1s;
wire[1:0] Tile_X9Y3_to_EG_1s;
wire[1:0] Tile_X9Y3_to_EH_1s;
wire[1:0] Tile_X9Y3_to_EI_1s;
wire[1:0] Tile_X9Y3_to_WA_1s;
wire[1:0] Tile_X9Y3_to_WB_1s;
wire[1:0] Tile_X9Y3_to_WC_1s;
wire[1:0] Tile_X9Y3_to_WD_1s;
wire[1:0] Tile_X9Y3_to_WF_1s;
wire[1:0] Tile_X9Y3_to_WG_1s;
wire[1:0] Tile_X9Y3_to_WH_1s;
wire[1:0] Tile_X9Y3_to_WI_1s;
wire[1:0] Tile_X9Y3_to_NA_1s;
wire[1:0] Tile_X9Y3_to_NB_1s;
wire[1:0] Tile_X9Y3_to_NC_1s;
wire[1:0] Tile_X9Y3_to_ND_1s;
wire[1:0] Tile_X9Y3_to_NF_1s;
wire[1:0] Tile_X9Y3_to_NG_1s;
wire[1:0] Tile_X9Y3_to_NH_1s;
wire[1:0] Tile_X9Y3_to_NI_1s;
wire[1:0] Tile_X9Y3_to_SA_1s;
wire[1:0] Tile_X9Y3_to_SB_1s;
wire[1:0] Tile_X9Y3_to_SC_1s;
wire[1:0] Tile_X9Y3_to_SD_1s;
wire[1:0] Tile_X9Y3_to_SF_1s;
wire[1:0] Tile_X9Y3_to_SG_1s;
wire[1:0] Tile_X9Y3_to_SH_1s;
wire[1:0] Tile_X9Y3_to_SI_1s;
wire[1:0] Tile_X10Y3_to_WA_1s;
wire[1:0] Tile_X10Y3_to_WB_1s;
wire[1:0] Tile_X10Y3_to_WC_1s;
wire[1:0] Tile_X10Y3_to_WD_1s;
wire[1:0] Tile_X10Y3_to_WF_1s;
wire[1:0] Tile_X10Y3_to_WG_1s;
wire[1:0] Tile_X10Y3_to_WH_1s;
wire[1:0] Tile_X10Y3_to_WI_1s;
wire[3:0] Tile_X0Y4_to_EA;
wire[3:0] Tile_X0Y4_to_EB;
wire[3:0] Tile_X0Y4_to_EC;
wire[3:0] Tile_X0Y4_to_ED;
wire[3:0] Tile_X0Y4_to_EF;
wire[7:0] Tile_X0Y4_to_EG;
wire[7:0] Tile_X0Y4_to_EH;
wire[11:0] Tile_X0Y4_to_EI;
wire[3:0] Tile_X0Y4_to_NA;
wire[3:0] Tile_X0Y4_to_NB;
wire[3:0] Tile_X0Y4_to_NC;
wire[3:0] Tile_X0Y4_to_ND;
wire[3:0] Tile_X0Y4_to_NF;
wire[7:0] Tile_X0Y4_to_NG;
wire[7:0] Tile_X0Y4_to_NH;
wire[11:0] Tile_X0Y4_to_NI;
wire[3:0] Tile_X0Y4_to_SA;
wire[3:0] Tile_X0Y4_to_SB;
wire[3:0] Tile_X0Y4_to_SC;
wire[3:0] Tile_X0Y4_to_SD;
wire[3:0] Tile_X0Y4_to_SF;
wire[7:0] Tile_X0Y4_to_SG;
wire[7:0] Tile_X0Y4_to_SH;
wire[11:0] Tile_X0Y4_to_SI;
wire[3:0] Tile_X1Y4_to_EA;
wire[3:0] Tile_X1Y4_to_EB;
wire[3:0] Tile_X1Y4_to_EC;
wire[3:0] Tile_X1Y4_to_ED;
wire[3:0] Tile_X1Y4_to_EF;
wire[7:0] Tile_X1Y4_to_EG;
wire[7:0] Tile_X1Y4_to_EH;
wire[11:0] Tile_X1Y4_to_EI;
wire[3:0] Tile_X1Y4_to_WA;
wire[3:0] Tile_X1Y4_to_WB;
wire[3:0] Tile_X1Y4_to_WC;
wire[3:0] Tile_X1Y4_to_WD;
wire[3:0] Tile_X1Y4_to_WF;
wire[7:0] Tile_X1Y4_to_WG;
wire[7:0] Tile_X1Y4_to_WH;
wire[11:0] Tile_X1Y4_to_WI;
wire[3:0] Tile_X1Y4_to_NA;
wire[3:0] Tile_X1Y4_to_NB;
wire[3:0] Tile_X1Y4_to_NC;
wire[3:0] Tile_X1Y4_to_ND;
wire[3:0] Tile_X1Y4_to_NF;
wire[7:0] Tile_X1Y4_to_NG;
wire[7:0] Tile_X1Y4_to_NH;
wire[11:0] Tile_X1Y4_to_NI;
wire[3:0] Tile_X1Y4_to_SA;
wire[3:0] Tile_X1Y4_to_SB;
wire[3:0] Tile_X1Y4_to_SC;
wire[3:0] Tile_X1Y4_to_SD;
wire[3:0] Tile_X1Y4_to_SF;
wire[7:0] Tile_X1Y4_to_SG;
wire[7:0] Tile_X1Y4_to_SH;
wire[11:0] Tile_X1Y4_to_SI;
wire[3:0] Tile_X2Y4_to_EA;
wire[3:0] Tile_X2Y4_to_EB;
wire[3:0] Tile_X2Y4_to_EC;
wire[3:0] Tile_X2Y4_to_ED;
wire[3:0] Tile_X2Y4_to_EF;
wire[7:0] Tile_X2Y4_to_EG;
wire[7:0] Tile_X2Y4_to_EH;
wire[11:0] Tile_X2Y4_to_EI;
wire[3:0] Tile_X2Y4_to_WA;
wire[3:0] Tile_X2Y4_to_WB;
wire[3:0] Tile_X2Y4_to_WC;
wire[3:0] Tile_X2Y4_to_WD;
wire[3:0] Tile_X2Y4_to_WF;
wire[7:0] Tile_X2Y4_to_WG;
wire[7:0] Tile_X2Y4_to_WH;
wire[11:0] Tile_X2Y4_to_WI;
wire[3:0] Tile_X2Y4_to_NA;
wire[3:0] Tile_X2Y4_to_NB;
wire[3:0] Tile_X2Y4_to_NC;
wire[3:0] Tile_X2Y4_to_ND;
wire[3:0] Tile_X2Y4_to_NF;
wire[7:0] Tile_X2Y4_to_NG;
wire[7:0] Tile_X2Y4_to_NH;
wire[11:0] Tile_X2Y4_to_NI;
wire[3:0] Tile_X2Y4_to_SA;
wire[3:0] Tile_X2Y4_to_SB;
wire[3:0] Tile_X2Y4_to_SC;
wire[3:0] Tile_X2Y4_to_SD;
wire[3:0] Tile_X2Y4_to_SF;
wire[7:0] Tile_X2Y4_to_SG;
wire[7:0] Tile_X2Y4_to_SH;
wire[11:0] Tile_X2Y4_to_SI;
wire[3:0] Tile_X3Y4_to_EA;
wire[3:0] Tile_X3Y4_to_EB;
wire[3:0] Tile_X3Y4_to_EC;
wire[3:0] Tile_X3Y4_to_ED;
wire[3:0] Tile_X3Y4_to_EF;
wire[7:0] Tile_X3Y4_to_EG;
wire[7:0] Tile_X3Y4_to_EH;
wire[11:0] Tile_X3Y4_to_EI;
wire[3:0] Tile_X3Y4_to_WA;
wire[3:0] Tile_X3Y4_to_WB;
wire[3:0] Tile_X3Y4_to_WC;
wire[3:0] Tile_X3Y4_to_WD;
wire[3:0] Tile_X3Y4_to_WF;
wire[7:0] Tile_X3Y4_to_WG;
wire[7:0] Tile_X3Y4_to_WH;
wire[11:0] Tile_X3Y4_to_WI;
wire[3:0] Tile_X3Y4_to_NA;
wire[3:0] Tile_X3Y4_to_NB;
wire[3:0] Tile_X3Y4_to_NC;
wire[3:0] Tile_X3Y4_to_ND;
wire[3:0] Tile_X3Y4_to_NF;
wire[7:0] Tile_X3Y4_to_NG;
wire[7:0] Tile_X3Y4_to_NH;
wire[11:0] Tile_X3Y4_to_NI;
wire[3:0] Tile_X3Y4_to_SA;
wire[3:0] Tile_X3Y4_to_SB;
wire[3:0] Tile_X3Y4_to_SC;
wire[3:0] Tile_X3Y4_to_SD;
wire[3:0] Tile_X3Y4_to_SF;
wire[7:0] Tile_X3Y4_to_SG;
wire[7:0] Tile_X3Y4_to_SH;
wire[11:0] Tile_X3Y4_to_SI;
wire[3:0] Tile_X4Y4_to_EA;
wire[3:0] Tile_X4Y4_to_EB;
wire[3:0] Tile_X4Y4_to_EC;
wire[3:0] Tile_X4Y4_to_ED;
wire[3:0] Tile_X4Y4_to_EF;
wire[7:0] Tile_X4Y4_to_EG;
wire[7:0] Tile_X4Y4_to_EH;
wire[11:0] Tile_X4Y4_to_EI;
wire[3:0] Tile_X4Y4_to_WA;
wire[3:0] Tile_X4Y4_to_WB;
wire[3:0] Tile_X4Y4_to_WC;
wire[3:0] Tile_X4Y4_to_WD;
wire[3:0] Tile_X4Y4_to_WF;
wire[7:0] Tile_X4Y4_to_WG;
wire[7:0] Tile_X4Y4_to_WH;
wire[11:0] Tile_X4Y4_to_WI;
wire[3:0] Tile_X4Y4_to_NA;
wire[3:0] Tile_X4Y4_to_NB;
wire[3:0] Tile_X4Y4_to_NC;
wire[3:0] Tile_X4Y4_to_ND;
wire[3:0] Tile_X4Y4_to_NF;
wire[7:0] Tile_X4Y4_to_NG;
wire[7:0] Tile_X4Y4_to_NH;
wire[11:0] Tile_X4Y4_to_NI;
wire[3:0] Tile_X4Y4_to_SA;
wire[3:0] Tile_X4Y4_to_SB;
wire[3:0] Tile_X4Y4_to_SC;
wire[3:0] Tile_X4Y4_to_SD;
wire[3:0] Tile_X4Y4_to_SF;
wire[7:0] Tile_X4Y4_to_SG;
wire[7:0] Tile_X4Y4_to_SH;
wire[11:0] Tile_X4Y4_to_SI;
wire[3:0] Tile_X5Y4_to_EA;
wire[3:0] Tile_X5Y4_to_EB;
wire[3:0] Tile_X5Y4_to_EC;
wire[3:0] Tile_X5Y4_to_ED;
wire[3:0] Tile_X5Y4_to_EF;
wire[7:0] Tile_X5Y4_to_EG;
wire[7:0] Tile_X5Y4_to_EH;
wire[11:0] Tile_X5Y4_to_EI;
wire[3:0] Tile_X5Y4_to_WA;
wire[3:0] Tile_X5Y4_to_WB;
wire[3:0] Tile_X5Y4_to_WC;
wire[3:0] Tile_X5Y4_to_WD;
wire[3:0] Tile_X5Y4_to_WF;
wire[7:0] Tile_X5Y4_to_WG;
wire[7:0] Tile_X5Y4_to_WH;
wire[11:0] Tile_X5Y4_to_WI;
wire[3:0] Tile_X5Y4_to_NA;
wire[3:0] Tile_X5Y4_to_NB;
wire[3:0] Tile_X5Y4_to_NC;
wire[3:0] Tile_X5Y4_to_ND;
wire[3:0] Tile_X5Y4_to_NF;
wire[7:0] Tile_X5Y4_to_NG;
wire[7:0] Tile_X5Y4_to_NH;
wire[11:0] Tile_X5Y4_to_NI;
wire[3:0] Tile_X5Y4_to_SA;
wire[3:0] Tile_X5Y4_to_SB;
wire[3:0] Tile_X5Y4_to_SC;
wire[3:0] Tile_X5Y4_to_SD;
wire[3:0] Tile_X5Y4_to_SF;
wire[7:0] Tile_X5Y4_to_SG;
wire[7:0] Tile_X5Y4_to_SH;
wire[11:0] Tile_X5Y4_to_SI;
wire[3:0] Tile_X6Y4_to_EA;
wire[3:0] Tile_X6Y4_to_EB;
wire[3:0] Tile_X6Y4_to_EC;
wire[3:0] Tile_X6Y4_to_ED;
wire[3:0] Tile_X6Y4_to_EF;
wire[7:0] Tile_X6Y4_to_EG;
wire[7:0] Tile_X6Y4_to_EH;
wire[11:0] Tile_X6Y4_to_EI;
wire[3:0] Tile_X6Y4_to_WA;
wire[3:0] Tile_X6Y4_to_WB;
wire[3:0] Tile_X6Y4_to_WC;
wire[3:0] Tile_X6Y4_to_WD;
wire[3:0] Tile_X6Y4_to_WF;
wire[7:0] Tile_X6Y4_to_WG;
wire[7:0] Tile_X6Y4_to_WH;
wire[11:0] Tile_X6Y4_to_WI;
wire[3:0] Tile_X6Y4_to_NA;
wire[3:0] Tile_X6Y4_to_NB;
wire[3:0] Tile_X6Y4_to_NC;
wire[3:0] Tile_X6Y4_to_ND;
wire[3:0] Tile_X6Y4_to_NF;
wire[7:0] Tile_X6Y4_to_NG;
wire[7:0] Tile_X6Y4_to_NH;
wire[11:0] Tile_X6Y4_to_NI;
wire[3:0] Tile_X6Y4_to_SA;
wire[3:0] Tile_X6Y4_to_SB;
wire[3:0] Tile_X6Y4_to_SC;
wire[3:0] Tile_X6Y4_to_SD;
wire[3:0] Tile_X6Y4_to_SF;
wire[7:0] Tile_X6Y4_to_SG;
wire[7:0] Tile_X6Y4_to_SH;
wire[11:0] Tile_X6Y4_to_SI;
wire[3:0] Tile_X7Y4_to_EA;
wire[3:0] Tile_X7Y4_to_EB;
wire[3:0] Tile_X7Y4_to_EC;
wire[3:0] Tile_X7Y4_to_ED;
wire[3:0] Tile_X7Y4_to_EF;
wire[7:0] Tile_X7Y4_to_EG;
wire[7:0] Tile_X7Y4_to_EH;
wire[11:0] Tile_X7Y4_to_EI;
wire[3:0] Tile_X7Y4_to_WA;
wire[3:0] Tile_X7Y4_to_WB;
wire[3:0] Tile_X7Y4_to_WC;
wire[3:0] Tile_X7Y4_to_WD;
wire[3:0] Tile_X7Y4_to_WF;
wire[7:0] Tile_X7Y4_to_WG;
wire[7:0] Tile_X7Y4_to_WH;
wire[11:0] Tile_X7Y4_to_WI;
wire[3:0] Tile_X7Y4_to_NA;
wire[3:0] Tile_X7Y4_to_NB;
wire[3:0] Tile_X7Y4_to_NC;
wire[3:0] Tile_X7Y4_to_ND;
wire[3:0] Tile_X7Y4_to_NF;
wire[7:0] Tile_X7Y4_to_NG;
wire[7:0] Tile_X7Y4_to_NH;
wire[11:0] Tile_X7Y4_to_NI;
wire[3:0] Tile_X7Y4_to_SA;
wire[3:0] Tile_X7Y4_to_SB;
wire[3:0] Tile_X7Y4_to_SC;
wire[3:0] Tile_X7Y4_to_SD;
wire[3:0] Tile_X7Y4_to_SF;
wire[7:0] Tile_X7Y4_to_SG;
wire[7:0] Tile_X7Y4_to_SH;
wire[11:0] Tile_X7Y4_to_SI;
wire[3:0] Tile_X8Y4_to_WA;
wire[3:0] Tile_X8Y4_to_WB;
wire[3:0] Tile_X8Y4_to_WC;
wire[3:0] Tile_X8Y4_to_WD;
wire[3:0] Tile_X8Y4_to_WF;
wire[7:0] Tile_X8Y4_to_WG;
wire[7:0] Tile_X8Y4_to_WH;
wire[11:0] Tile_X8Y4_to_WI;
wire[3:0] Tile_X8Y4_to_NA;
wire[3:0] Tile_X8Y4_to_NB;
wire[3:0] Tile_X8Y4_to_NC;
wire[3:0] Tile_X8Y4_to_ND;
wire[3:0] Tile_X8Y4_to_NF;
wire[7:0] Tile_X8Y4_to_NG;
wire[7:0] Tile_X8Y4_to_NH;
wire[11:0] Tile_X8Y4_to_NI;
wire[3:0] Tile_X8Y4_to_SA;
wire[3:0] Tile_X8Y4_to_SB;
wire[3:0] Tile_X8Y4_to_SC;
wire[3:0] Tile_X8Y4_to_SD;
wire[3:0] Tile_X8Y4_to_SF;
wire[7:0] Tile_X8Y4_to_SG;
wire[7:0] Tile_X8Y4_to_SH;
wire[11:0] Tile_X8Y4_to_SI;
wire[1:0] Tile_X9Y4_to_EA_1s;
wire[1:0] Tile_X9Y4_to_EB_1s;
wire[1:0] Tile_X9Y4_to_EC_1s;
wire[1:0] Tile_X9Y4_to_ED_1s;
wire[1:0] Tile_X9Y4_to_EF_1s;
wire[1:0] Tile_X9Y4_to_EG_1s;
wire[1:0] Tile_X9Y4_to_EH_1s;
wire[1:0] Tile_X9Y4_to_EI_1s;
wire[1:0] Tile_X9Y4_to_WA_1s;
wire[1:0] Tile_X9Y4_to_WB_1s;
wire[1:0] Tile_X9Y4_to_WC_1s;
wire[1:0] Tile_X9Y4_to_WD_1s;
wire[1:0] Tile_X9Y4_to_WF_1s;
wire[1:0] Tile_X9Y4_to_WG_1s;
wire[1:0] Tile_X9Y4_to_WH_1s;
wire[1:0] Tile_X9Y4_to_WI_1s;
wire[1:0] Tile_X9Y4_to_NA_1s;
wire[1:0] Tile_X9Y4_to_NB_1s;
wire[1:0] Tile_X9Y4_to_NC_1s;
wire[1:0] Tile_X9Y4_to_ND_1s;
wire[1:0] Tile_X9Y4_to_NF_1s;
wire[1:0] Tile_X9Y4_to_NG_1s;
wire[1:0] Tile_X9Y4_to_NH_1s;
wire[1:0] Tile_X9Y4_to_NI_1s;
wire[1:0] Tile_X9Y4_to_SA_1s;
wire[1:0] Tile_X9Y4_to_SB_1s;
wire[1:0] Tile_X9Y4_to_SC_1s;
wire[1:0] Tile_X9Y4_to_SD_1s;
wire[1:0] Tile_X9Y4_to_SF_1s;
wire[1:0] Tile_X9Y4_to_SG_1s;
wire[1:0] Tile_X9Y4_to_SH_1s;
wire[1:0] Tile_X9Y4_to_SI_1s;
wire[1:0] Tile_X10Y4_to_WA_1s;
wire[1:0] Tile_X10Y4_to_WB_1s;
wire[1:0] Tile_X10Y4_to_WC_1s;
wire[1:0] Tile_X10Y4_to_WD_1s;
wire[1:0] Tile_X10Y4_to_WF_1s;
wire[1:0] Tile_X10Y4_to_WG_1s;
wire[1:0] Tile_X10Y4_to_WH_1s;
wire[1:0] Tile_X10Y4_to_WI_1s;
wire[3:0] Tile_X0Y5_to_EA;
wire[3:0] Tile_X0Y5_to_EB;
wire[3:0] Tile_X0Y5_to_EC;
wire[3:0] Tile_X0Y5_to_ED;
wire[3:0] Tile_X0Y5_to_EF;
wire[7:0] Tile_X0Y5_to_EG;
wire[7:0] Tile_X0Y5_to_EH;
wire[11:0] Tile_X0Y5_to_EI;
wire[3:0] Tile_X0Y5_to_NA;
wire[3:0] Tile_X0Y5_to_NB;
wire[3:0] Tile_X0Y5_to_NC;
wire[3:0] Tile_X0Y5_to_ND;
wire[3:0] Tile_X0Y5_to_NF;
wire[7:0] Tile_X0Y5_to_NG;
wire[7:0] Tile_X0Y5_to_NH;
wire[11:0] Tile_X0Y5_to_NI;
wire[3:0] Tile_X0Y5_to_SA;
wire[3:0] Tile_X0Y5_to_SB;
wire[3:0] Tile_X0Y5_to_SC;
wire[3:0] Tile_X0Y5_to_SD;
wire[3:0] Tile_X0Y5_to_SF;
wire[7:0] Tile_X0Y5_to_SG;
wire[7:0] Tile_X0Y5_to_SH;
wire[11:0] Tile_X0Y5_to_SI;
wire[3:0] Tile_X1Y5_to_EA;
wire[3:0] Tile_X1Y5_to_EB;
wire[3:0] Tile_X1Y5_to_EC;
wire[3:0] Tile_X1Y5_to_ED;
wire[3:0] Tile_X1Y5_to_EF;
wire[7:0] Tile_X1Y5_to_EG;
wire[7:0] Tile_X1Y5_to_EH;
wire[11:0] Tile_X1Y5_to_EI;
wire[3:0] Tile_X1Y5_to_WA;
wire[3:0] Tile_X1Y5_to_WB;
wire[3:0] Tile_X1Y5_to_WC;
wire[3:0] Tile_X1Y5_to_WD;
wire[3:0] Tile_X1Y5_to_WF;
wire[7:0] Tile_X1Y5_to_WG;
wire[7:0] Tile_X1Y5_to_WH;
wire[11:0] Tile_X1Y5_to_WI;
wire[3:0] Tile_X1Y5_to_NA;
wire[3:0] Tile_X1Y5_to_NB;
wire[3:0] Tile_X1Y5_to_NC;
wire[3:0] Tile_X1Y5_to_ND;
wire[3:0] Tile_X1Y5_to_NF;
wire[7:0] Tile_X1Y5_to_NG;
wire[7:0] Tile_X1Y5_to_NH;
wire[11:0] Tile_X1Y5_to_NI;
wire[3:0] Tile_X1Y5_to_SA;
wire[3:0] Tile_X1Y5_to_SB;
wire[3:0] Tile_X1Y5_to_SC;
wire[3:0] Tile_X1Y5_to_SD;
wire[3:0] Tile_X1Y5_to_SF;
wire[7:0] Tile_X1Y5_to_SG;
wire[7:0] Tile_X1Y5_to_SH;
wire[11:0] Tile_X1Y5_to_SI;
wire[3:0] Tile_X2Y5_to_EA;
wire[3:0] Tile_X2Y5_to_EB;
wire[3:0] Tile_X2Y5_to_EC;
wire[3:0] Tile_X2Y5_to_ED;
wire[3:0] Tile_X2Y5_to_EF;
wire[7:0] Tile_X2Y5_to_EG;
wire[7:0] Tile_X2Y5_to_EH;
wire[11:0] Tile_X2Y5_to_EI;
wire[3:0] Tile_X2Y5_to_WA;
wire[3:0] Tile_X2Y5_to_WB;
wire[3:0] Tile_X2Y5_to_WC;
wire[3:0] Tile_X2Y5_to_WD;
wire[3:0] Tile_X2Y5_to_WF;
wire[7:0] Tile_X2Y5_to_WG;
wire[7:0] Tile_X2Y5_to_WH;
wire[11:0] Tile_X2Y5_to_WI;
wire[3:0] Tile_X2Y5_to_NA;
wire[3:0] Tile_X2Y5_to_NB;
wire[3:0] Tile_X2Y5_to_NC;
wire[3:0] Tile_X2Y5_to_ND;
wire[3:0] Tile_X2Y5_to_NF;
wire[7:0] Tile_X2Y5_to_NG;
wire[7:0] Tile_X2Y5_to_NH;
wire[11:0] Tile_X2Y5_to_NI;
wire[3:0] Tile_X2Y5_to_SA;
wire[3:0] Tile_X2Y5_to_SB;
wire[3:0] Tile_X2Y5_to_SC;
wire[3:0] Tile_X2Y5_to_SD;
wire[3:0] Tile_X2Y5_to_SF;
wire[7:0] Tile_X2Y5_to_SG;
wire[7:0] Tile_X2Y5_to_SH;
wire[11:0] Tile_X2Y5_to_SI;
wire[3:0] Tile_X3Y5_to_EA;
wire[3:0] Tile_X3Y5_to_EB;
wire[3:0] Tile_X3Y5_to_EC;
wire[3:0] Tile_X3Y5_to_ED;
wire[3:0] Tile_X3Y5_to_EF;
wire[7:0] Tile_X3Y5_to_EG;
wire[7:0] Tile_X3Y5_to_EH;
wire[11:0] Tile_X3Y5_to_EI;
wire[3:0] Tile_X3Y5_to_WA;
wire[3:0] Tile_X3Y5_to_WB;
wire[3:0] Tile_X3Y5_to_WC;
wire[3:0] Tile_X3Y5_to_WD;
wire[3:0] Tile_X3Y5_to_WF;
wire[7:0] Tile_X3Y5_to_WG;
wire[7:0] Tile_X3Y5_to_WH;
wire[11:0] Tile_X3Y5_to_WI;
wire[3:0] Tile_X3Y5_to_NA;
wire[3:0] Tile_X3Y5_to_NB;
wire[3:0] Tile_X3Y5_to_NC;
wire[3:0] Tile_X3Y5_to_ND;
wire[3:0] Tile_X3Y5_to_NF;
wire[7:0] Tile_X3Y5_to_NG;
wire[7:0] Tile_X3Y5_to_NH;
wire[11:0] Tile_X3Y5_to_NI;
wire[3:0] Tile_X3Y5_to_SA;
wire[3:0] Tile_X3Y5_to_SB;
wire[3:0] Tile_X3Y5_to_SC;
wire[3:0] Tile_X3Y5_to_SD;
wire[3:0] Tile_X3Y5_to_SF;
wire[7:0] Tile_X3Y5_to_SG;
wire[7:0] Tile_X3Y5_to_SH;
wire[11:0] Tile_X3Y5_to_SI;
wire[3:0] Tile_X4Y5_to_EA;
wire[3:0] Tile_X4Y5_to_EB;
wire[3:0] Tile_X4Y5_to_EC;
wire[3:0] Tile_X4Y5_to_ED;
wire[3:0] Tile_X4Y5_to_EF;
wire[7:0] Tile_X4Y5_to_EG;
wire[7:0] Tile_X4Y5_to_EH;
wire[11:0] Tile_X4Y5_to_EI;
wire[3:0] Tile_X4Y5_to_WA;
wire[3:0] Tile_X4Y5_to_WB;
wire[3:0] Tile_X4Y5_to_WC;
wire[3:0] Tile_X4Y5_to_WD;
wire[3:0] Tile_X4Y5_to_WF;
wire[7:0] Tile_X4Y5_to_WG;
wire[7:0] Tile_X4Y5_to_WH;
wire[11:0] Tile_X4Y5_to_WI;
wire[3:0] Tile_X4Y5_to_NA;
wire[3:0] Tile_X4Y5_to_NB;
wire[3:0] Tile_X4Y5_to_NC;
wire[3:0] Tile_X4Y5_to_ND;
wire[3:0] Tile_X4Y5_to_NF;
wire[7:0] Tile_X4Y5_to_NG;
wire[7:0] Tile_X4Y5_to_NH;
wire[11:0] Tile_X4Y5_to_NI;
wire[3:0] Tile_X4Y5_to_SA;
wire[3:0] Tile_X4Y5_to_SB;
wire[3:0] Tile_X4Y5_to_SC;
wire[3:0] Tile_X4Y5_to_SD;
wire[3:0] Tile_X4Y5_to_SF;
wire[7:0] Tile_X4Y5_to_SG;
wire[7:0] Tile_X4Y5_to_SH;
wire[11:0] Tile_X4Y5_to_SI;
wire[3:0] Tile_X5Y5_to_EA;
wire[3:0] Tile_X5Y5_to_EB;
wire[3:0] Tile_X5Y5_to_EC;
wire[3:0] Tile_X5Y5_to_ED;
wire[3:0] Tile_X5Y5_to_EF;
wire[7:0] Tile_X5Y5_to_EG;
wire[7:0] Tile_X5Y5_to_EH;
wire[11:0] Tile_X5Y5_to_EI;
wire[3:0] Tile_X5Y5_to_WA;
wire[3:0] Tile_X5Y5_to_WB;
wire[3:0] Tile_X5Y5_to_WC;
wire[3:0] Tile_X5Y5_to_WD;
wire[3:0] Tile_X5Y5_to_WF;
wire[7:0] Tile_X5Y5_to_WG;
wire[7:0] Tile_X5Y5_to_WH;
wire[11:0] Tile_X5Y5_to_WI;
wire[3:0] Tile_X5Y5_to_NA;
wire[3:0] Tile_X5Y5_to_NB;
wire[3:0] Tile_X5Y5_to_NC;
wire[3:0] Tile_X5Y5_to_ND;
wire[3:0] Tile_X5Y5_to_NF;
wire[7:0] Tile_X5Y5_to_NG;
wire[7:0] Tile_X5Y5_to_NH;
wire[11:0] Tile_X5Y5_to_NI;
wire[3:0] Tile_X5Y5_to_SA;
wire[3:0] Tile_X5Y5_to_SB;
wire[3:0] Tile_X5Y5_to_SC;
wire[3:0] Tile_X5Y5_to_SD;
wire[3:0] Tile_X5Y5_to_SF;
wire[7:0] Tile_X5Y5_to_SG;
wire[7:0] Tile_X5Y5_to_SH;
wire[11:0] Tile_X5Y5_to_SI;
wire[3:0] Tile_X6Y5_to_EA;
wire[3:0] Tile_X6Y5_to_EB;
wire[3:0] Tile_X6Y5_to_EC;
wire[3:0] Tile_X6Y5_to_ED;
wire[3:0] Tile_X6Y5_to_EF;
wire[7:0] Tile_X6Y5_to_EG;
wire[7:0] Tile_X6Y5_to_EH;
wire[11:0] Tile_X6Y5_to_EI;
wire[3:0] Tile_X6Y5_to_WA;
wire[3:0] Tile_X6Y5_to_WB;
wire[3:0] Tile_X6Y5_to_WC;
wire[3:0] Tile_X6Y5_to_WD;
wire[3:0] Tile_X6Y5_to_WF;
wire[7:0] Tile_X6Y5_to_WG;
wire[7:0] Tile_X6Y5_to_WH;
wire[11:0] Tile_X6Y5_to_WI;
wire[3:0] Tile_X6Y5_to_NA;
wire[3:0] Tile_X6Y5_to_NB;
wire[3:0] Tile_X6Y5_to_NC;
wire[3:0] Tile_X6Y5_to_ND;
wire[3:0] Tile_X6Y5_to_NF;
wire[7:0] Tile_X6Y5_to_NG;
wire[7:0] Tile_X6Y5_to_NH;
wire[11:0] Tile_X6Y5_to_NI;
wire[3:0] Tile_X6Y5_to_SA;
wire[3:0] Tile_X6Y5_to_SB;
wire[3:0] Tile_X6Y5_to_SC;
wire[3:0] Tile_X6Y5_to_SD;
wire[3:0] Tile_X6Y5_to_SF;
wire[7:0] Tile_X6Y5_to_SG;
wire[7:0] Tile_X6Y5_to_SH;
wire[11:0] Tile_X6Y5_to_SI;
wire[3:0] Tile_X7Y5_to_EA;
wire[3:0] Tile_X7Y5_to_EB;
wire[3:0] Tile_X7Y5_to_EC;
wire[3:0] Tile_X7Y5_to_ED;
wire[3:0] Tile_X7Y5_to_EF;
wire[7:0] Tile_X7Y5_to_EG;
wire[7:0] Tile_X7Y5_to_EH;
wire[11:0] Tile_X7Y5_to_EI;
wire[3:0] Tile_X7Y5_to_WA;
wire[3:0] Tile_X7Y5_to_WB;
wire[3:0] Tile_X7Y5_to_WC;
wire[3:0] Tile_X7Y5_to_WD;
wire[3:0] Tile_X7Y5_to_WF;
wire[7:0] Tile_X7Y5_to_WG;
wire[7:0] Tile_X7Y5_to_WH;
wire[11:0] Tile_X7Y5_to_WI;
wire[3:0] Tile_X7Y5_to_NA;
wire[3:0] Tile_X7Y5_to_NB;
wire[3:0] Tile_X7Y5_to_NC;
wire[3:0] Tile_X7Y5_to_ND;
wire[3:0] Tile_X7Y5_to_NF;
wire[7:0] Tile_X7Y5_to_NG;
wire[7:0] Tile_X7Y5_to_NH;
wire[11:0] Tile_X7Y5_to_NI;
wire[3:0] Tile_X7Y5_to_SA;
wire[3:0] Tile_X7Y5_to_SB;
wire[3:0] Tile_X7Y5_to_SC;
wire[3:0] Tile_X7Y5_to_SD;
wire[3:0] Tile_X7Y5_to_SF;
wire[7:0] Tile_X7Y5_to_SG;
wire[7:0] Tile_X7Y5_to_SH;
wire[11:0] Tile_X7Y5_to_SI;
wire[3:0] Tile_X8Y5_to_WA;
wire[3:0] Tile_X8Y5_to_WB;
wire[3:0] Tile_X8Y5_to_WC;
wire[3:0] Tile_X8Y5_to_WD;
wire[3:0] Tile_X8Y5_to_WF;
wire[7:0] Tile_X8Y5_to_WG;
wire[7:0] Tile_X8Y5_to_WH;
wire[11:0] Tile_X8Y5_to_WI;
wire[3:0] Tile_X8Y5_to_NA;
wire[3:0] Tile_X8Y5_to_NB;
wire[3:0] Tile_X8Y5_to_NC;
wire[3:0] Tile_X8Y5_to_ND;
wire[3:0] Tile_X8Y5_to_NF;
wire[7:0] Tile_X8Y5_to_NG;
wire[7:0] Tile_X8Y5_to_NH;
wire[11:0] Tile_X8Y5_to_NI;
wire[3:0] Tile_X8Y5_to_SA;
wire[3:0] Tile_X8Y5_to_SB;
wire[3:0] Tile_X8Y5_to_SC;
wire[3:0] Tile_X8Y5_to_SD;
wire[3:0] Tile_X8Y5_to_SF;
wire[7:0] Tile_X8Y5_to_SG;
wire[7:0] Tile_X8Y5_to_SH;
wire[11:0] Tile_X8Y5_to_SI;
wire[1:0] Tile_X9Y5_to_EA_1s;
wire[1:0] Tile_X9Y5_to_EB_1s;
wire[1:0] Tile_X9Y5_to_EC_1s;
wire[1:0] Tile_X9Y5_to_ED_1s;
wire[1:0] Tile_X9Y5_to_EF_1s;
wire[1:0] Tile_X9Y5_to_EG_1s;
wire[1:0] Tile_X9Y5_to_EH_1s;
wire[1:0] Tile_X9Y5_to_EI_1s;
wire[1:0] Tile_X9Y5_to_WA_1s;
wire[1:0] Tile_X9Y5_to_WB_1s;
wire[1:0] Tile_X9Y5_to_WC_1s;
wire[1:0] Tile_X9Y5_to_WD_1s;
wire[1:0] Tile_X9Y5_to_WF_1s;
wire[1:0] Tile_X9Y5_to_WG_1s;
wire[1:0] Tile_X9Y5_to_WH_1s;
wire[1:0] Tile_X9Y5_to_WI_1s;
wire[1:0] Tile_X9Y5_to_NA_1s;
wire[1:0] Tile_X9Y5_to_NB_1s;
wire[1:0] Tile_X9Y5_to_NC_1s;
wire[1:0] Tile_X9Y5_to_ND_1s;
wire[1:0] Tile_X9Y5_to_NF_1s;
wire[1:0] Tile_X9Y5_to_NG_1s;
wire[1:0] Tile_X9Y5_to_NH_1s;
wire[1:0] Tile_X9Y5_to_NI_1s;
wire[1:0] Tile_X9Y5_to_SA_1s;
wire[1:0] Tile_X9Y5_to_SB_1s;
wire[1:0] Tile_X9Y5_to_SC_1s;
wire[1:0] Tile_X9Y5_to_SD_1s;
wire[1:0] Tile_X9Y5_to_SF_1s;
wire[1:0] Tile_X9Y5_to_SG_1s;
wire[1:0] Tile_X9Y5_to_SH_1s;
wire[1:0] Tile_X9Y5_to_SI_1s;
wire[1:0] Tile_X10Y5_to_WA_1s;
wire[1:0] Tile_X10Y5_to_WB_1s;
wire[1:0] Tile_X10Y5_to_WC_1s;
wire[1:0] Tile_X10Y5_to_WD_1s;
wire[1:0] Tile_X10Y5_to_WF_1s;
wire[1:0] Tile_X10Y5_to_WG_1s;
wire[1:0] Tile_X10Y5_to_WH_1s;
wire[1:0] Tile_X10Y5_to_WI_1s;
wire[3:0] Tile_X0Y6_to_EA;
wire[3:0] Tile_X0Y6_to_EB;
wire[3:0] Tile_X0Y6_to_EC;
wire[3:0] Tile_X0Y6_to_ED;
wire[3:0] Tile_X0Y6_to_EF;
wire[7:0] Tile_X0Y6_to_EG;
wire[7:0] Tile_X0Y6_to_EH;
wire[11:0] Tile_X0Y6_to_EI;
wire[3:0] Tile_X0Y6_to_NA;
wire[3:0] Tile_X0Y6_to_NB;
wire[3:0] Tile_X0Y6_to_NC;
wire[3:0] Tile_X0Y6_to_ND;
wire[3:0] Tile_X0Y6_to_NF;
wire[7:0] Tile_X0Y6_to_NG;
wire[7:0] Tile_X0Y6_to_NH;
wire[11:0] Tile_X0Y6_to_NI;
wire[3:0] Tile_X0Y6_to_SA;
wire[3:0] Tile_X0Y6_to_SB;
wire[3:0] Tile_X0Y6_to_SC;
wire[3:0] Tile_X0Y6_to_SD;
wire[3:0] Tile_X0Y6_to_SF;
wire[7:0] Tile_X0Y6_to_SG;
wire[7:0] Tile_X0Y6_to_SH;
wire[11:0] Tile_X0Y6_to_SI;
wire[3:0] Tile_X1Y6_to_EA;
wire[3:0] Tile_X1Y6_to_EB;
wire[3:0] Tile_X1Y6_to_EC;
wire[3:0] Tile_X1Y6_to_ED;
wire[3:0] Tile_X1Y6_to_EF;
wire[7:0] Tile_X1Y6_to_EG;
wire[7:0] Tile_X1Y6_to_EH;
wire[11:0] Tile_X1Y6_to_EI;
wire[3:0] Tile_X1Y6_to_WA;
wire[3:0] Tile_X1Y6_to_WB;
wire[3:0] Tile_X1Y6_to_WC;
wire[3:0] Tile_X1Y6_to_WD;
wire[3:0] Tile_X1Y6_to_WF;
wire[7:0] Tile_X1Y6_to_WG;
wire[7:0] Tile_X1Y6_to_WH;
wire[11:0] Tile_X1Y6_to_WI;
wire[3:0] Tile_X1Y6_to_NA;
wire[3:0] Tile_X1Y6_to_NB;
wire[3:0] Tile_X1Y6_to_NC;
wire[3:0] Tile_X1Y6_to_ND;
wire[3:0] Tile_X1Y6_to_NF;
wire[7:0] Tile_X1Y6_to_NG;
wire[7:0] Tile_X1Y6_to_NH;
wire[11:0] Tile_X1Y6_to_NI;
wire[3:0] Tile_X1Y6_to_SA;
wire[3:0] Tile_X1Y6_to_SB;
wire[3:0] Tile_X1Y6_to_SC;
wire[3:0] Tile_X1Y6_to_SD;
wire[3:0] Tile_X1Y6_to_SF;
wire[7:0] Tile_X1Y6_to_SG;
wire[7:0] Tile_X1Y6_to_SH;
wire[11:0] Tile_X1Y6_to_SI;
wire[3:0] Tile_X2Y6_to_EA;
wire[3:0] Tile_X2Y6_to_EB;
wire[3:0] Tile_X2Y6_to_EC;
wire[3:0] Tile_X2Y6_to_ED;
wire[3:0] Tile_X2Y6_to_EF;
wire[7:0] Tile_X2Y6_to_EG;
wire[7:0] Tile_X2Y6_to_EH;
wire[11:0] Tile_X2Y6_to_EI;
wire[3:0] Tile_X2Y6_to_WA;
wire[3:0] Tile_X2Y6_to_WB;
wire[3:0] Tile_X2Y6_to_WC;
wire[3:0] Tile_X2Y6_to_WD;
wire[3:0] Tile_X2Y6_to_WF;
wire[7:0] Tile_X2Y6_to_WG;
wire[7:0] Tile_X2Y6_to_WH;
wire[11:0] Tile_X2Y6_to_WI;
wire[3:0] Tile_X2Y6_to_NA;
wire[3:0] Tile_X2Y6_to_NB;
wire[3:0] Tile_X2Y6_to_NC;
wire[3:0] Tile_X2Y6_to_ND;
wire[3:0] Tile_X2Y6_to_NF;
wire[7:0] Tile_X2Y6_to_NG;
wire[7:0] Tile_X2Y6_to_NH;
wire[11:0] Tile_X2Y6_to_NI;
wire[3:0] Tile_X2Y6_to_SA;
wire[3:0] Tile_X2Y6_to_SB;
wire[3:0] Tile_X2Y6_to_SC;
wire[3:0] Tile_X2Y6_to_SD;
wire[3:0] Tile_X2Y6_to_SF;
wire[7:0] Tile_X2Y6_to_SG;
wire[7:0] Tile_X2Y6_to_SH;
wire[11:0] Tile_X2Y6_to_SI;
wire[3:0] Tile_X3Y6_to_EA;
wire[3:0] Tile_X3Y6_to_EB;
wire[3:0] Tile_X3Y6_to_EC;
wire[3:0] Tile_X3Y6_to_ED;
wire[3:0] Tile_X3Y6_to_EF;
wire[7:0] Tile_X3Y6_to_EG;
wire[7:0] Tile_X3Y6_to_EH;
wire[11:0] Tile_X3Y6_to_EI;
wire[3:0] Tile_X3Y6_to_WA;
wire[3:0] Tile_X3Y6_to_WB;
wire[3:0] Tile_X3Y6_to_WC;
wire[3:0] Tile_X3Y6_to_WD;
wire[3:0] Tile_X3Y6_to_WF;
wire[7:0] Tile_X3Y6_to_WG;
wire[7:0] Tile_X3Y6_to_WH;
wire[11:0] Tile_X3Y6_to_WI;
wire[3:0] Tile_X3Y6_to_NA;
wire[3:0] Tile_X3Y6_to_NB;
wire[3:0] Tile_X3Y6_to_NC;
wire[3:0] Tile_X3Y6_to_ND;
wire[3:0] Tile_X3Y6_to_NF;
wire[7:0] Tile_X3Y6_to_NG;
wire[7:0] Tile_X3Y6_to_NH;
wire[11:0] Tile_X3Y6_to_NI;
wire[3:0] Tile_X3Y6_to_SA;
wire[3:0] Tile_X3Y6_to_SB;
wire[3:0] Tile_X3Y6_to_SC;
wire[3:0] Tile_X3Y6_to_SD;
wire[3:0] Tile_X3Y6_to_SF;
wire[7:0] Tile_X3Y6_to_SG;
wire[7:0] Tile_X3Y6_to_SH;
wire[11:0] Tile_X3Y6_to_SI;
wire[3:0] Tile_X4Y6_to_EA;
wire[3:0] Tile_X4Y6_to_EB;
wire[3:0] Tile_X4Y6_to_EC;
wire[3:0] Tile_X4Y6_to_ED;
wire[3:0] Tile_X4Y6_to_EF;
wire[7:0] Tile_X4Y6_to_EG;
wire[7:0] Tile_X4Y6_to_EH;
wire[11:0] Tile_X4Y6_to_EI;
wire[3:0] Tile_X4Y6_to_WA;
wire[3:0] Tile_X4Y6_to_WB;
wire[3:0] Tile_X4Y6_to_WC;
wire[3:0] Tile_X4Y6_to_WD;
wire[3:0] Tile_X4Y6_to_WF;
wire[7:0] Tile_X4Y6_to_WG;
wire[7:0] Tile_X4Y6_to_WH;
wire[11:0] Tile_X4Y6_to_WI;
wire[3:0] Tile_X4Y6_to_NA;
wire[3:0] Tile_X4Y6_to_NB;
wire[3:0] Tile_X4Y6_to_NC;
wire[3:0] Tile_X4Y6_to_ND;
wire[3:0] Tile_X4Y6_to_NF;
wire[7:0] Tile_X4Y6_to_NG;
wire[7:0] Tile_X4Y6_to_NH;
wire[11:0] Tile_X4Y6_to_NI;
wire[3:0] Tile_X4Y6_to_SA;
wire[3:0] Tile_X4Y6_to_SB;
wire[3:0] Tile_X4Y6_to_SC;
wire[3:0] Tile_X4Y6_to_SD;
wire[3:0] Tile_X4Y6_to_SF;
wire[7:0] Tile_X4Y6_to_SG;
wire[7:0] Tile_X4Y6_to_SH;
wire[11:0] Tile_X4Y6_to_SI;
wire[3:0] Tile_X5Y6_to_EA;
wire[3:0] Tile_X5Y6_to_EB;
wire[3:0] Tile_X5Y6_to_EC;
wire[3:0] Tile_X5Y6_to_ED;
wire[3:0] Tile_X5Y6_to_EF;
wire[7:0] Tile_X5Y6_to_EG;
wire[7:0] Tile_X5Y6_to_EH;
wire[11:0] Tile_X5Y6_to_EI;
wire[3:0] Tile_X5Y6_to_WA;
wire[3:0] Tile_X5Y6_to_WB;
wire[3:0] Tile_X5Y6_to_WC;
wire[3:0] Tile_X5Y6_to_WD;
wire[3:0] Tile_X5Y6_to_WF;
wire[7:0] Tile_X5Y6_to_WG;
wire[7:0] Tile_X5Y6_to_WH;
wire[11:0] Tile_X5Y6_to_WI;
wire[3:0] Tile_X5Y6_to_NA;
wire[3:0] Tile_X5Y6_to_NB;
wire[3:0] Tile_X5Y6_to_NC;
wire[3:0] Tile_X5Y6_to_ND;
wire[3:0] Tile_X5Y6_to_NF;
wire[7:0] Tile_X5Y6_to_NG;
wire[7:0] Tile_X5Y6_to_NH;
wire[11:0] Tile_X5Y6_to_NI;
wire[3:0] Tile_X5Y6_to_SA;
wire[3:0] Tile_X5Y6_to_SB;
wire[3:0] Tile_X5Y6_to_SC;
wire[3:0] Tile_X5Y6_to_SD;
wire[3:0] Tile_X5Y6_to_SF;
wire[7:0] Tile_X5Y6_to_SG;
wire[7:0] Tile_X5Y6_to_SH;
wire[11:0] Tile_X5Y6_to_SI;
wire[3:0] Tile_X6Y6_to_EA;
wire[3:0] Tile_X6Y6_to_EB;
wire[3:0] Tile_X6Y6_to_EC;
wire[3:0] Tile_X6Y6_to_ED;
wire[3:0] Tile_X6Y6_to_EF;
wire[7:0] Tile_X6Y6_to_EG;
wire[7:0] Tile_X6Y6_to_EH;
wire[11:0] Tile_X6Y6_to_EI;
wire[3:0] Tile_X6Y6_to_WA;
wire[3:0] Tile_X6Y6_to_WB;
wire[3:0] Tile_X6Y6_to_WC;
wire[3:0] Tile_X6Y6_to_WD;
wire[3:0] Tile_X6Y6_to_WF;
wire[7:0] Tile_X6Y6_to_WG;
wire[7:0] Tile_X6Y6_to_WH;
wire[11:0] Tile_X6Y6_to_WI;
wire[3:0] Tile_X6Y6_to_NA;
wire[3:0] Tile_X6Y6_to_NB;
wire[3:0] Tile_X6Y6_to_NC;
wire[3:0] Tile_X6Y6_to_ND;
wire[3:0] Tile_X6Y6_to_NF;
wire[7:0] Tile_X6Y6_to_NG;
wire[7:0] Tile_X6Y6_to_NH;
wire[11:0] Tile_X6Y6_to_NI;
wire[3:0] Tile_X6Y6_to_SA;
wire[3:0] Tile_X6Y6_to_SB;
wire[3:0] Tile_X6Y6_to_SC;
wire[3:0] Tile_X6Y6_to_SD;
wire[3:0] Tile_X6Y6_to_SF;
wire[7:0] Tile_X6Y6_to_SG;
wire[7:0] Tile_X6Y6_to_SH;
wire[11:0] Tile_X6Y6_to_SI;
wire[3:0] Tile_X7Y6_to_EA;
wire[3:0] Tile_X7Y6_to_EB;
wire[3:0] Tile_X7Y6_to_EC;
wire[3:0] Tile_X7Y6_to_ED;
wire[3:0] Tile_X7Y6_to_EF;
wire[7:0] Tile_X7Y6_to_EG;
wire[7:0] Tile_X7Y6_to_EH;
wire[11:0] Tile_X7Y6_to_EI;
wire[3:0] Tile_X7Y6_to_WA;
wire[3:0] Tile_X7Y6_to_WB;
wire[3:0] Tile_X7Y6_to_WC;
wire[3:0] Tile_X7Y6_to_WD;
wire[3:0] Tile_X7Y6_to_WF;
wire[7:0] Tile_X7Y6_to_WG;
wire[7:0] Tile_X7Y6_to_WH;
wire[11:0] Tile_X7Y6_to_WI;
wire[3:0] Tile_X7Y6_to_NA;
wire[3:0] Tile_X7Y6_to_NB;
wire[3:0] Tile_X7Y6_to_NC;
wire[3:0] Tile_X7Y6_to_ND;
wire[3:0] Tile_X7Y6_to_NF;
wire[7:0] Tile_X7Y6_to_NG;
wire[7:0] Tile_X7Y6_to_NH;
wire[11:0] Tile_X7Y6_to_NI;
wire[3:0] Tile_X7Y6_to_SA;
wire[3:0] Tile_X7Y6_to_SB;
wire[3:0] Tile_X7Y6_to_SC;
wire[3:0] Tile_X7Y6_to_SD;
wire[3:0] Tile_X7Y6_to_SF;
wire[7:0] Tile_X7Y6_to_SG;
wire[7:0] Tile_X7Y6_to_SH;
wire[11:0] Tile_X7Y6_to_SI;
wire[3:0] Tile_X8Y6_to_WA;
wire[3:0] Tile_X8Y6_to_WB;
wire[3:0] Tile_X8Y6_to_WC;
wire[3:0] Tile_X8Y6_to_WD;
wire[3:0] Tile_X8Y6_to_WF;
wire[7:0] Tile_X8Y6_to_WG;
wire[7:0] Tile_X8Y6_to_WH;
wire[11:0] Tile_X8Y6_to_WI;
wire[3:0] Tile_X8Y6_to_NA;
wire[3:0] Tile_X8Y6_to_NB;
wire[3:0] Tile_X8Y6_to_NC;
wire[3:0] Tile_X8Y6_to_ND;
wire[3:0] Tile_X8Y6_to_NF;
wire[7:0] Tile_X8Y6_to_NG;
wire[7:0] Tile_X8Y6_to_NH;
wire[11:0] Tile_X8Y6_to_NI;
wire[3:0] Tile_X8Y6_to_SA;
wire[3:0] Tile_X8Y6_to_SB;
wire[3:0] Tile_X8Y6_to_SC;
wire[3:0] Tile_X8Y6_to_SD;
wire[3:0] Tile_X8Y6_to_SF;
wire[7:0] Tile_X8Y6_to_SG;
wire[7:0] Tile_X8Y6_to_SH;
wire[11:0] Tile_X8Y6_to_SI;
wire[1:0] Tile_X9Y6_to_EA_1s;
wire[1:0] Tile_X9Y6_to_EB_1s;
wire[1:0] Tile_X9Y6_to_EC_1s;
wire[1:0] Tile_X9Y6_to_ED_1s;
wire[1:0] Tile_X9Y6_to_EF_1s;
wire[1:0] Tile_X9Y6_to_EG_1s;
wire[1:0] Tile_X9Y6_to_EH_1s;
wire[1:0] Tile_X9Y6_to_EI_1s;
wire[1:0] Tile_X9Y6_to_WA_1s;
wire[1:0] Tile_X9Y6_to_WB_1s;
wire[1:0] Tile_X9Y6_to_WC_1s;
wire[1:0] Tile_X9Y6_to_WD_1s;
wire[1:0] Tile_X9Y6_to_WF_1s;
wire[1:0] Tile_X9Y6_to_WG_1s;
wire[1:0] Tile_X9Y6_to_WH_1s;
wire[1:0] Tile_X9Y6_to_WI_1s;
wire[1:0] Tile_X9Y6_to_NA_1s;
wire[1:0] Tile_X9Y6_to_NB_1s;
wire[1:0] Tile_X9Y6_to_NC_1s;
wire[1:0] Tile_X9Y6_to_ND_1s;
wire[1:0] Tile_X9Y6_to_NF_1s;
wire[1:0] Tile_X9Y6_to_NG_1s;
wire[1:0] Tile_X9Y6_to_NH_1s;
wire[1:0] Tile_X9Y6_to_NI_1s;
wire[1:0] Tile_X9Y6_to_SA_1s;
wire[1:0] Tile_X9Y6_to_SB_1s;
wire[1:0] Tile_X9Y6_to_SC_1s;
wire[1:0] Tile_X9Y6_to_SD_1s;
wire[1:0] Tile_X9Y6_to_SF_1s;
wire[1:0] Tile_X9Y6_to_SG_1s;
wire[1:0] Tile_X9Y6_to_SH_1s;
wire[1:0] Tile_X9Y6_to_SI_1s;
wire[1:0] Tile_X10Y6_to_WA_1s;
wire[1:0] Tile_X10Y6_to_WB_1s;
wire[1:0] Tile_X10Y6_to_WC_1s;
wire[1:0] Tile_X10Y6_to_WD_1s;
wire[1:0] Tile_X10Y6_to_WF_1s;
wire[1:0] Tile_X10Y6_to_WG_1s;
wire[1:0] Tile_X10Y6_to_WH_1s;
wire[1:0] Tile_X10Y6_to_WI_1s;
wire[3:0] Tile_X0Y7_to_EA;
wire[3:0] Tile_X0Y7_to_EB;
wire[3:0] Tile_X0Y7_to_EC;
wire[3:0] Tile_X0Y7_to_ED;
wire[3:0] Tile_X0Y7_to_EF;
wire[7:0] Tile_X0Y7_to_EG;
wire[7:0] Tile_X0Y7_to_EH;
wire[11:0] Tile_X0Y7_to_EI;
wire[3:0] Tile_X0Y7_to_NA;
wire[3:0] Tile_X0Y7_to_NB;
wire[3:0] Tile_X0Y7_to_NC;
wire[3:0] Tile_X0Y7_to_ND;
wire[3:0] Tile_X0Y7_to_NF;
wire[7:0] Tile_X0Y7_to_NG;
wire[7:0] Tile_X0Y7_to_NH;
wire[11:0] Tile_X0Y7_to_NI;
wire[3:0] Tile_X0Y7_to_SA;
wire[3:0] Tile_X0Y7_to_SB;
wire[3:0] Tile_X0Y7_to_SC;
wire[3:0] Tile_X0Y7_to_SD;
wire[3:0] Tile_X0Y7_to_SF;
wire[7:0] Tile_X0Y7_to_SG;
wire[7:0] Tile_X0Y7_to_SH;
wire[11:0] Tile_X0Y7_to_SI;
wire[3:0] Tile_X1Y7_to_EA;
wire[3:0] Tile_X1Y7_to_EB;
wire[3:0] Tile_X1Y7_to_EC;
wire[3:0] Tile_X1Y7_to_ED;
wire[3:0] Tile_X1Y7_to_EF;
wire[7:0] Tile_X1Y7_to_EG;
wire[7:0] Tile_X1Y7_to_EH;
wire[11:0] Tile_X1Y7_to_EI;
wire[3:0] Tile_X1Y7_to_WA;
wire[3:0] Tile_X1Y7_to_WB;
wire[3:0] Tile_X1Y7_to_WC;
wire[3:0] Tile_X1Y7_to_WD;
wire[3:0] Tile_X1Y7_to_WF;
wire[7:0] Tile_X1Y7_to_WG;
wire[7:0] Tile_X1Y7_to_WH;
wire[11:0] Tile_X1Y7_to_WI;
wire[3:0] Tile_X1Y7_to_NA;
wire[3:0] Tile_X1Y7_to_NB;
wire[3:0] Tile_X1Y7_to_NC;
wire[3:0] Tile_X1Y7_to_ND;
wire[3:0] Tile_X1Y7_to_NF;
wire[7:0] Tile_X1Y7_to_NG;
wire[7:0] Tile_X1Y7_to_NH;
wire[11:0] Tile_X1Y7_to_NI;
wire[3:0] Tile_X1Y7_to_SA;
wire[3:0] Tile_X1Y7_to_SB;
wire[3:0] Tile_X1Y7_to_SC;
wire[3:0] Tile_X1Y7_to_SD;
wire[3:0] Tile_X1Y7_to_SF;
wire[7:0] Tile_X1Y7_to_SG;
wire[7:0] Tile_X1Y7_to_SH;
wire[11:0] Tile_X1Y7_to_SI;
wire[3:0] Tile_X2Y7_to_EA;
wire[3:0] Tile_X2Y7_to_EB;
wire[3:0] Tile_X2Y7_to_EC;
wire[3:0] Tile_X2Y7_to_ED;
wire[3:0] Tile_X2Y7_to_EF;
wire[7:0] Tile_X2Y7_to_EG;
wire[7:0] Tile_X2Y7_to_EH;
wire[11:0] Tile_X2Y7_to_EI;
wire[3:0] Tile_X2Y7_to_WA;
wire[3:0] Tile_X2Y7_to_WB;
wire[3:0] Tile_X2Y7_to_WC;
wire[3:0] Tile_X2Y7_to_WD;
wire[3:0] Tile_X2Y7_to_WF;
wire[7:0] Tile_X2Y7_to_WG;
wire[7:0] Tile_X2Y7_to_WH;
wire[11:0] Tile_X2Y7_to_WI;
wire[3:0] Tile_X2Y7_to_NA;
wire[3:0] Tile_X2Y7_to_NB;
wire[3:0] Tile_X2Y7_to_NC;
wire[3:0] Tile_X2Y7_to_ND;
wire[3:0] Tile_X2Y7_to_NF;
wire[7:0] Tile_X2Y7_to_NG;
wire[7:0] Tile_X2Y7_to_NH;
wire[11:0] Tile_X2Y7_to_NI;
wire[3:0] Tile_X2Y7_to_SA;
wire[3:0] Tile_X2Y7_to_SB;
wire[3:0] Tile_X2Y7_to_SC;
wire[3:0] Tile_X2Y7_to_SD;
wire[3:0] Tile_X2Y7_to_SF;
wire[7:0] Tile_X2Y7_to_SG;
wire[7:0] Tile_X2Y7_to_SH;
wire[11:0] Tile_X2Y7_to_SI;
wire[3:0] Tile_X3Y7_to_EA;
wire[3:0] Tile_X3Y7_to_EB;
wire[3:0] Tile_X3Y7_to_EC;
wire[3:0] Tile_X3Y7_to_ED;
wire[3:0] Tile_X3Y7_to_EF;
wire[7:0] Tile_X3Y7_to_EG;
wire[7:0] Tile_X3Y7_to_EH;
wire[11:0] Tile_X3Y7_to_EI;
wire[3:0] Tile_X3Y7_to_WA;
wire[3:0] Tile_X3Y7_to_WB;
wire[3:0] Tile_X3Y7_to_WC;
wire[3:0] Tile_X3Y7_to_WD;
wire[3:0] Tile_X3Y7_to_WF;
wire[7:0] Tile_X3Y7_to_WG;
wire[7:0] Tile_X3Y7_to_WH;
wire[11:0] Tile_X3Y7_to_WI;
wire[3:0] Tile_X3Y7_to_NA;
wire[3:0] Tile_X3Y7_to_NB;
wire[3:0] Tile_X3Y7_to_NC;
wire[3:0] Tile_X3Y7_to_ND;
wire[3:0] Tile_X3Y7_to_NF;
wire[7:0] Tile_X3Y7_to_NG;
wire[7:0] Tile_X3Y7_to_NH;
wire[11:0] Tile_X3Y7_to_NI;
wire[3:0] Tile_X3Y7_to_SA;
wire[3:0] Tile_X3Y7_to_SB;
wire[3:0] Tile_X3Y7_to_SC;
wire[3:0] Tile_X3Y7_to_SD;
wire[3:0] Tile_X3Y7_to_SF;
wire[7:0] Tile_X3Y7_to_SG;
wire[7:0] Tile_X3Y7_to_SH;
wire[11:0] Tile_X3Y7_to_SI;
wire[3:0] Tile_X4Y7_to_EA;
wire[3:0] Tile_X4Y7_to_EB;
wire[3:0] Tile_X4Y7_to_EC;
wire[3:0] Tile_X4Y7_to_ED;
wire[3:0] Tile_X4Y7_to_EF;
wire[7:0] Tile_X4Y7_to_EG;
wire[7:0] Tile_X4Y7_to_EH;
wire[11:0] Tile_X4Y7_to_EI;
wire[3:0] Tile_X4Y7_to_WA;
wire[3:0] Tile_X4Y7_to_WB;
wire[3:0] Tile_X4Y7_to_WC;
wire[3:0] Tile_X4Y7_to_WD;
wire[3:0] Tile_X4Y7_to_WF;
wire[7:0] Tile_X4Y7_to_WG;
wire[7:0] Tile_X4Y7_to_WH;
wire[11:0] Tile_X4Y7_to_WI;
wire[3:0] Tile_X4Y7_to_NA;
wire[3:0] Tile_X4Y7_to_NB;
wire[3:0] Tile_X4Y7_to_NC;
wire[3:0] Tile_X4Y7_to_ND;
wire[3:0] Tile_X4Y7_to_NF;
wire[7:0] Tile_X4Y7_to_NG;
wire[7:0] Tile_X4Y7_to_NH;
wire[11:0] Tile_X4Y7_to_NI;
wire[3:0] Tile_X4Y7_to_SA;
wire[3:0] Tile_X4Y7_to_SB;
wire[3:0] Tile_X4Y7_to_SC;
wire[3:0] Tile_X4Y7_to_SD;
wire[3:0] Tile_X4Y7_to_SF;
wire[7:0] Tile_X4Y7_to_SG;
wire[7:0] Tile_X4Y7_to_SH;
wire[11:0] Tile_X4Y7_to_SI;
wire[3:0] Tile_X5Y7_to_EA;
wire[3:0] Tile_X5Y7_to_EB;
wire[3:0] Tile_X5Y7_to_EC;
wire[3:0] Tile_X5Y7_to_ED;
wire[3:0] Tile_X5Y7_to_EF;
wire[7:0] Tile_X5Y7_to_EG;
wire[7:0] Tile_X5Y7_to_EH;
wire[11:0] Tile_X5Y7_to_EI;
wire[3:0] Tile_X5Y7_to_WA;
wire[3:0] Tile_X5Y7_to_WB;
wire[3:0] Tile_X5Y7_to_WC;
wire[3:0] Tile_X5Y7_to_WD;
wire[3:0] Tile_X5Y7_to_WF;
wire[7:0] Tile_X5Y7_to_WG;
wire[7:0] Tile_X5Y7_to_WH;
wire[11:0] Tile_X5Y7_to_WI;
wire[3:0] Tile_X5Y7_to_NA;
wire[3:0] Tile_X5Y7_to_NB;
wire[3:0] Tile_X5Y7_to_NC;
wire[3:0] Tile_X5Y7_to_ND;
wire[3:0] Tile_X5Y7_to_NF;
wire[7:0] Tile_X5Y7_to_NG;
wire[7:0] Tile_X5Y7_to_NH;
wire[11:0] Tile_X5Y7_to_NI;
wire[3:0] Tile_X5Y7_to_SA;
wire[3:0] Tile_X5Y7_to_SB;
wire[3:0] Tile_X5Y7_to_SC;
wire[3:0] Tile_X5Y7_to_SD;
wire[3:0] Tile_X5Y7_to_SF;
wire[7:0] Tile_X5Y7_to_SG;
wire[7:0] Tile_X5Y7_to_SH;
wire[11:0] Tile_X5Y7_to_SI;
wire[3:0] Tile_X6Y7_to_EA;
wire[3:0] Tile_X6Y7_to_EB;
wire[3:0] Tile_X6Y7_to_EC;
wire[3:0] Tile_X6Y7_to_ED;
wire[3:0] Tile_X6Y7_to_EF;
wire[7:0] Tile_X6Y7_to_EG;
wire[7:0] Tile_X6Y7_to_EH;
wire[11:0] Tile_X6Y7_to_EI;
wire[3:0] Tile_X6Y7_to_WA;
wire[3:0] Tile_X6Y7_to_WB;
wire[3:0] Tile_X6Y7_to_WC;
wire[3:0] Tile_X6Y7_to_WD;
wire[3:0] Tile_X6Y7_to_WF;
wire[7:0] Tile_X6Y7_to_WG;
wire[7:0] Tile_X6Y7_to_WH;
wire[11:0] Tile_X6Y7_to_WI;
wire[3:0] Tile_X6Y7_to_NA;
wire[3:0] Tile_X6Y7_to_NB;
wire[3:0] Tile_X6Y7_to_NC;
wire[3:0] Tile_X6Y7_to_ND;
wire[3:0] Tile_X6Y7_to_NF;
wire[7:0] Tile_X6Y7_to_NG;
wire[7:0] Tile_X6Y7_to_NH;
wire[11:0] Tile_X6Y7_to_NI;
wire[3:0] Tile_X6Y7_to_SA;
wire[3:0] Tile_X6Y7_to_SB;
wire[3:0] Tile_X6Y7_to_SC;
wire[3:0] Tile_X6Y7_to_SD;
wire[3:0] Tile_X6Y7_to_SF;
wire[7:0] Tile_X6Y7_to_SG;
wire[7:0] Tile_X6Y7_to_SH;
wire[11:0] Tile_X6Y7_to_SI;
wire[3:0] Tile_X7Y7_to_EA;
wire[3:0] Tile_X7Y7_to_EB;
wire[3:0] Tile_X7Y7_to_EC;
wire[3:0] Tile_X7Y7_to_ED;
wire[3:0] Tile_X7Y7_to_EF;
wire[7:0] Tile_X7Y7_to_EG;
wire[7:0] Tile_X7Y7_to_EH;
wire[11:0] Tile_X7Y7_to_EI;
wire[3:0] Tile_X7Y7_to_WA;
wire[3:0] Tile_X7Y7_to_WB;
wire[3:0] Tile_X7Y7_to_WC;
wire[3:0] Tile_X7Y7_to_WD;
wire[3:0] Tile_X7Y7_to_WF;
wire[7:0] Tile_X7Y7_to_WG;
wire[7:0] Tile_X7Y7_to_WH;
wire[11:0] Tile_X7Y7_to_WI;
wire[3:0] Tile_X7Y7_to_NA;
wire[3:0] Tile_X7Y7_to_NB;
wire[3:0] Tile_X7Y7_to_NC;
wire[3:0] Tile_X7Y7_to_ND;
wire[3:0] Tile_X7Y7_to_NF;
wire[7:0] Tile_X7Y7_to_NG;
wire[7:0] Tile_X7Y7_to_NH;
wire[11:0] Tile_X7Y7_to_NI;
wire[3:0] Tile_X7Y7_to_SA;
wire[3:0] Tile_X7Y7_to_SB;
wire[3:0] Tile_X7Y7_to_SC;
wire[3:0] Tile_X7Y7_to_SD;
wire[3:0] Tile_X7Y7_to_SF;
wire[7:0] Tile_X7Y7_to_SG;
wire[7:0] Tile_X7Y7_to_SH;
wire[11:0] Tile_X7Y7_to_SI;
wire[3:0] Tile_X8Y7_to_WA;
wire[3:0] Tile_X8Y7_to_WB;
wire[3:0] Tile_X8Y7_to_WC;
wire[3:0] Tile_X8Y7_to_WD;
wire[3:0] Tile_X8Y7_to_WF;
wire[7:0] Tile_X8Y7_to_WG;
wire[7:0] Tile_X8Y7_to_WH;
wire[11:0] Tile_X8Y7_to_WI;
wire[3:0] Tile_X8Y7_to_NA;
wire[3:0] Tile_X8Y7_to_NB;
wire[3:0] Tile_X8Y7_to_NC;
wire[3:0] Tile_X8Y7_to_ND;
wire[3:0] Tile_X8Y7_to_NF;
wire[7:0] Tile_X8Y7_to_NG;
wire[7:0] Tile_X8Y7_to_NH;
wire[11:0] Tile_X8Y7_to_NI;
wire[3:0] Tile_X8Y7_to_SA;
wire[3:0] Tile_X8Y7_to_SB;
wire[3:0] Tile_X8Y7_to_SC;
wire[3:0] Tile_X8Y7_to_SD;
wire[3:0] Tile_X8Y7_to_SF;
wire[7:0] Tile_X8Y7_to_SG;
wire[7:0] Tile_X8Y7_to_SH;
wire[11:0] Tile_X8Y7_to_SI;
wire[1:0] Tile_X9Y7_to_EA_1s;
wire[1:0] Tile_X9Y7_to_EB_1s;
wire[1:0] Tile_X9Y7_to_EC_1s;
wire[1:0] Tile_X9Y7_to_ED_1s;
wire[1:0] Tile_X9Y7_to_EF_1s;
wire[1:0] Tile_X9Y7_to_EG_1s;
wire[1:0] Tile_X9Y7_to_EH_1s;
wire[1:0] Tile_X9Y7_to_EI_1s;
wire[1:0] Tile_X9Y7_to_WA_1s;
wire[1:0] Tile_X9Y7_to_WB_1s;
wire[1:0] Tile_X9Y7_to_WC_1s;
wire[1:0] Tile_X9Y7_to_WD_1s;
wire[1:0] Tile_X9Y7_to_WF_1s;
wire[1:0] Tile_X9Y7_to_WG_1s;
wire[1:0] Tile_X9Y7_to_WH_1s;
wire[1:0] Tile_X9Y7_to_WI_1s;
wire[1:0] Tile_X9Y7_to_NA_1s;
wire[1:0] Tile_X9Y7_to_NB_1s;
wire[1:0] Tile_X9Y7_to_NC_1s;
wire[1:0] Tile_X9Y7_to_ND_1s;
wire[1:0] Tile_X9Y7_to_NF_1s;
wire[1:0] Tile_X9Y7_to_NG_1s;
wire[1:0] Tile_X9Y7_to_NH_1s;
wire[1:0] Tile_X9Y7_to_NI_1s;
wire[1:0] Tile_X9Y7_to_SA_1s;
wire[1:0] Tile_X9Y7_to_SB_1s;
wire[1:0] Tile_X9Y7_to_SC_1s;
wire[1:0] Tile_X9Y7_to_SD_1s;
wire[1:0] Tile_X9Y7_to_SF_1s;
wire[1:0] Tile_X9Y7_to_SG_1s;
wire[1:0] Tile_X9Y7_to_SH_1s;
wire[1:0] Tile_X9Y7_to_SI_1s;
wire[1:0] Tile_X10Y7_to_WA_1s;
wire[1:0] Tile_X10Y7_to_WB_1s;
wire[1:0] Tile_X10Y7_to_WC_1s;
wire[1:0] Tile_X10Y7_to_WD_1s;
wire[1:0] Tile_X10Y7_to_WF_1s;
wire[1:0] Tile_X10Y7_to_WG_1s;
wire[1:0] Tile_X10Y7_to_WH_1s;
wire[1:0] Tile_X10Y7_to_WI_1s;
wire[3:0] Tile_X0Y8_to_EA;
wire[3:0] Tile_X0Y8_to_EB;
wire[3:0] Tile_X0Y8_to_EC;
wire[3:0] Tile_X0Y8_to_ED;
wire[3:0] Tile_X0Y8_to_EF;
wire[7:0] Tile_X0Y8_to_EG;
wire[7:0] Tile_X0Y8_to_EH;
wire[11:0] Tile_X0Y8_to_EI;
wire[3:0] Tile_X0Y8_to_NA;
wire[3:0] Tile_X0Y8_to_NB;
wire[3:0] Tile_X0Y8_to_NC;
wire[3:0] Tile_X0Y8_to_ND;
wire[3:0] Tile_X0Y8_to_NF;
wire[7:0] Tile_X0Y8_to_NG;
wire[7:0] Tile_X0Y8_to_NH;
wire[11:0] Tile_X0Y8_to_NI;
wire[3:0] Tile_X0Y8_to_SA;
wire[3:0] Tile_X0Y8_to_SB;
wire[3:0] Tile_X0Y8_to_SC;
wire[3:0] Tile_X0Y8_to_SD;
wire[3:0] Tile_X0Y8_to_SF;
wire[7:0] Tile_X0Y8_to_SG;
wire[7:0] Tile_X0Y8_to_SH;
wire[11:0] Tile_X0Y8_to_SI;
wire[3:0] Tile_X1Y8_to_EA;
wire[3:0] Tile_X1Y8_to_EB;
wire[3:0] Tile_X1Y8_to_EC;
wire[3:0] Tile_X1Y8_to_ED;
wire[3:0] Tile_X1Y8_to_EF;
wire[7:0] Tile_X1Y8_to_EG;
wire[7:0] Tile_X1Y8_to_EH;
wire[11:0] Tile_X1Y8_to_EI;
wire[3:0] Tile_X1Y8_to_WA;
wire[3:0] Tile_X1Y8_to_WB;
wire[3:0] Tile_X1Y8_to_WC;
wire[3:0] Tile_X1Y8_to_WD;
wire[3:0] Tile_X1Y8_to_WF;
wire[7:0] Tile_X1Y8_to_WG;
wire[7:0] Tile_X1Y8_to_WH;
wire[11:0] Tile_X1Y8_to_WI;
wire[3:0] Tile_X1Y8_to_NA;
wire[3:0] Tile_X1Y8_to_NB;
wire[3:0] Tile_X1Y8_to_NC;
wire[3:0] Tile_X1Y8_to_ND;
wire[3:0] Tile_X1Y8_to_NF;
wire[7:0] Tile_X1Y8_to_NG;
wire[7:0] Tile_X1Y8_to_NH;
wire[11:0] Tile_X1Y8_to_NI;
wire[3:0] Tile_X1Y8_to_SA;
wire[3:0] Tile_X1Y8_to_SB;
wire[3:0] Tile_X1Y8_to_SC;
wire[3:0] Tile_X1Y8_to_SD;
wire[3:0] Tile_X1Y8_to_SF;
wire[7:0] Tile_X1Y8_to_SG;
wire[7:0] Tile_X1Y8_to_SH;
wire[11:0] Tile_X1Y8_to_SI;
wire[3:0] Tile_X2Y8_to_EA;
wire[3:0] Tile_X2Y8_to_EB;
wire[3:0] Tile_X2Y8_to_EC;
wire[3:0] Tile_X2Y8_to_ED;
wire[3:0] Tile_X2Y8_to_EF;
wire[7:0] Tile_X2Y8_to_EG;
wire[7:0] Tile_X2Y8_to_EH;
wire[11:0] Tile_X2Y8_to_EI;
wire[3:0] Tile_X2Y8_to_WA;
wire[3:0] Tile_X2Y8_to_WB;
wire[3:0] Tile_X2Y8_to_WC;
wire[3:0] Tile_X2Y8_to_WD;
wire[3:0] Tile_X2Y8_to_WF;
wire[7:0] Tile_X2Y8_to_WG;
wire[7:0] Tile_X2Y8_to_WH;
wire[11:0] Tile_X2Y8_to_WI;
wire[3:0] Tile_X2Y8_to_NA;
wire[3:0] Tile_X2Y8_to_NB;
wire[3:0] Tile_X2Y8_to_NC;
wire[3:0] Tile_X2Y8_to_ND;
wire[3:0] Tile_X2Y8_to_NF;
wire[7:0] Tile_X2Y8_to_NG;
wire[7:0] Tile_X2Y8_to_NH;
wire[11:0] Tile_X2Y8_to_NI;
wire[3:0] Tile_X2Y8_to_SA;
wire[3:0] Tile_X2Y8_to_SB;
wire[3:0] Tile_X2Y8_to_SC;
wire[3:0] Tile_X2Y8_to_SD;
wire[3:0] Tile_X2Y8_to_SF;
wire[7:0] Tile_X2Y8_to_SG;
wire[7:0] Tile_X2Y8_to_SH;
wire[11:0] Tile_X2Y8_to_SI;
wire[3:0] Tile_X3Y8_to_EA;
wire[3:0] Tile_X3Y8_to_EB;
wire[3:0] Tile_X3Y8_to_EC;
wire[3:0] Tile_X3Y8_to_ED;
wire[3:0] Tile_X3Y8_to_EF;
wire[7:0] Tile_X3Y8_to_EG;
wire[7:0] Tile_X3Y8_to_EH;
wire[11:0] Tile_X3Y8_to_EI;
wire[3:0] Tile_X3Y8_to_WA;
wire[3:0] Tile_X3Y8_to_WB;
wire[3:0] Tile_X3Y8_to_WC;
wire[3:0] Tile_X3Y8_to_WD;
wire[3:0] Tile_X3Y8_to_WF;
wire[7:0] Tile_X3Y8_to_WG;
wire[7:0] Tile_X3Y8_to_WH;
wire[11:0] Tile_X3Y8_to_WI;
wire[3:0] Tile_X3Y8_to_NA;
wire[3:0] Tile_X3Y8_to_NB;
wire[3:0] Tile_X3Y8_to_NC;
wire[3:0] Tile_X3Y8_to_ND;
wire[3:0] Tile_X3Y8_to_NF;
wire[7:0] Tile_X3Y8_to_NG;
wire[7:0] Tile_X3Y8_to_NH;
wire[11:0] Tile_X3Y8_to_NI;
wire[3:0] Tile_X3Y8_to_SA;
wire[3:0] Tile_X3Y8_to_SB;
wire[3:0] Tile_X3Y8_to_SC;
wire[3:0] Tile_X3Y8_to_SD;
wire[3:0] Tile_X3Y8_to_SF;
wire[7:0] Tile_X3Y8_to_SG;
wire[7:0] Tile_X3Y8_to_SH;
wire[11:0] Tile_X3Y8_to_SI;
wire[3:0] Tile_X4Y8_to_EA;
wire[3:0] Tile_X4Y8_to_EB;
wire[3:0] Tile_X4Y8_to_EC;
wire[3:0] Tile_X4Y8_to_ED;
wire[3:0] Tile_X4Y8_to_EF;
wire[7:0] Tile_X4Y8_to_EG;
wire[7:0] Tile_X4Y8_to_EH;
wire[11:0] Tile_X4Y8_to_EI;
wire[3:0] Tile_X4Y8_to_WA;
wire[3:0] Tile_X4Y8_to_WB;
wire[3:0] Tile_X4Y8_to_WC;
wire[3:0] Tile_X4Y8_to_WD;
wire[3:0] Tile_X4Y8_to_WF;
wire[7:0] Tile_X4Y8_to_WG;
wire[7:0] Tile_X4Y8_to_WH;
wire[11:0] Tile_X4Y8_to_WI;
wire[3:0] Tile_X4Y8_to_NA;
wire[3:0] Tile_X4Y8_to_NB;
wire[3:0] Tile_X4Y8_to_NC;
wire[3:0] Tile_X4Y8_to_ND;
wire[3:0] Tile_X4Y8_to_NF;
wire[7:0] Tile_X4Y8_to_NG;
wire[7:0] Tile_X4Y8_to_NH;
wire[11:0] Tile_X4Y8_to_NI;
wire[3:0] Tile_X4Y8_to_SA;
wire[3:0] Tile_X4Y8_to_SB;
wire[3:0] Tile_X4Y8_to_SC;
wire[3:0] Tile_X4Y8_to_SD;
wire[3:0] Tile_X4Y8_to_SF;
wire[7:0] Tile_X4Y8_to_SG;
wire[7:0] Tile_X4Y8_to_SH;
wire[11:0] Tile_X4Y8_to_SI;
wire[3:0] Tile_X5Y8_to_EA;
wire[3:0] Tile_X5Y8_to_EB;
wire[3:0] Tile_X5Y8_to_EC;
wire[3:0] Tile_X5Y8_to_ED;
wire[3:0] Tile_X5Y8_to_EF;
wire[7:0] Tile_X5Y8_to_EG;
wire[7:0] Tile_X5Y8_to_EH;
wire[11:0] Tile_X5Y8_to_EI;
wire[3:0] Tile_X5Y8_to_WA;
wire[3:0] Tile_X5Y8_to_WB;
wire[3:0] Tile_X5Y8_to_WC;
wire[3:0] Tile_X5Y8_to_WD;
wire[3:0] Tile_X5Y8_to_WF;
wire[7:0] Tile_X5Y8_to_WG;
wire[7:0] Tile_X5Y8_to_WH;
wire[11:0] Tile_X5Y8_to_WI;
wire[3:0] Tile_X5Y8_to_NA;
wire[3:0] Tile_X5Y8_to_NB;
wire[3:0] Tile_X5Y8_to_NC;
wire[3:0] Tile_X5Y8_to_ND;
wire[3:0] Tile_X5Y8_to_NF;
wire[7:0] Tile_X5Y8_to_NG;
wire[7:0] Tile_X5Y8_to_NH;
wire[11:0] Tile_X5Y8_to_NI;
wire[3:0] Tile_X5Y8_to_SA;
wire[3:0] Tile_X5Y8_to_SB;
wire[3:0] Tile_X5Y8_to_SC;
wire[3:0] Tile_X5Y8_to_SD;
wire[3:0] Tile_X5Y8_to_SF;
wire[7:0] Tile_X5Y8_to_SG;
wire[7:0] Tile_X5Y8_to_SH;
wire[11:0] Tile_X5Y8_to_SI;
wire[3:0] Tile_X6Y8_to_EA;
wire[3:0] Tile_X6Y8_to_EB;
wire[3:0] Tile_X6Y8_to_EC;
wire[3:0] Tile_X6Y8_to_ED;
wire[3:0] Tile_X6Y8_to_EF;
wire[7:0] Tile_X6Y8_to_EG;
wire[7:0] Tile_X6Y8_to_EH;
wire[11:0] Tile_X6Y8_to_EI;
wire[3:0] Tile_X6Y8_to_WA;
wire[3:0] Tile_X6Y8_to_WB;
wire[3:0] Tile_X6Y8_to_WC;
wire[3:0] Tile_X6Y8_to_WD;
wire[3:0] Tile_X6Y8_to_WF;
wire[7:0] Tile_X6Y8_to_WG;
wire[7:0] Tile_X6Y8_to_WH;
wire[11:0] Tile_X6Y8_to_WI;
wire[3:0] Tile_X6Y8_to_NA;
wire[3:0] Tile_X6Y8_to_NB;
wire[3:0] Tile_X6Y8_to_NC;
wire[3:0] Tile_X6Y8_to_ND;
wire[3:0] Tile_X6Y8_to_NF;
wire[7:0] Tile_X6Y8_to_NG;
wire[7:0] Tile_X6Y8_to_NH;
wire[11:0] Tile_X6Y8_to_NI;
wire[3:0] Tile_X6Y8_to_SA;
wire[3:0] Tile_X6Y8_to_SB;
wire[3:0] Tile_X6Y8_to_SC;
wire[3:0] Tile_X6Y8_to_SD;
wire[3:0] Tile_X6Y8_to_SF;
wire[7:0] Tile_X6Y8_to_SG;
wire[7:0] Tile_X6Y8_to_SH;
wire[11:0] Tile_X6Y8_to_SI;
wire[3:0] Tile_X7Y8_to_EA;
wire[3:0] Tile_X7Y8_to_EB;
wire[3:0] Tile_X7Y8_to_EC;
wire[3:0] Tile_X7Y8_to_ED;
wire[3:0] Tile_X7Y8_to_EF;
wire[7:0] Tile_X7Y8_to_EG;
wire[7:0] Tile_X7Y8_to_EH;
wire[11:0] Tile_X7Y8_to_EI;
wire[3:0] Tile_X7Y8_to_WA;
wire[3:0] Tile_X7Y8_to_WB;
wire[3:0] Tile_X7Y8_to_WC;
wire[3:0] Tile_X7Y8_to_WD;
wire[3:0] Tile_X7Y8_to_WF;
wire[7:0] Tile_X7Y8_to_WG;
wire[7:0] Tile_X7Y8_to_WH;
wire[11:0] Tile_X7Y8_to_WI;
wire[3:0] Tile_X7Y8_to_NA;
wire[3:0] Tile_X7Y8_to_NB;
wire[3:0] Tile_X7Y8_to_NC;
wire[3:0] Tile_X7Y8_to_ND;
wire[3:0] Tile_X7Y8_to_NF;
wire[7:0] Tile_X7Y8_to_NG;
wire[7:0] Tile_X7Y8_to_NH;
wire[11:0] Tile_X7Y8_to_NI;
wire[3:0] Tile_X7Y8_to_SA;
wire[3:0] Tile_X7Y8_to_SB;
wire[3:0] Tile_X7Y8_to_SC;
wire[3:0] Tile_X7Y8_to_SD;
wire[3:0] Tile_X7Y8_to_SF;
wire[7:0] Tile_X7Y8_to_SG;
wire[7:0] Tile_X7Y8_to_SH;
wire[11:0] Tile_X7Y8_to_SI;
wire[3:0] Tile_X8Y8_to_WA;
wire[3:0] Tile_X8Y8_to_WB;
wire[3:0] Tile_X8Y8_to_WC;
wire[3:0] Tile_X8Y8_to_WD;
wire[3:0] Tile_X8Y8_to_WF;
wire[7:0] Tile_X8Y8_to_WG;
wire[7:0] Tile_X8Y8_to_WH;
wire[11:0] Tile_X8Y8_to_WI;
wire[3:0] Tile_X8Y8_to_NA;
wire[3:0] Tile_X8Y8_to_NB;
wire[3:0] Tile_X8Y8_to_NC;
wire[3:0] Tile_X8Y8_to_ND;
wire[3:0] Tile_X8Y8_to_NF;
wire[7:0] Tile_X8Y8_to_NG;
wire[7:0] Tile_X8Y8_to_NH;
wire[11:0] Tile_X8Y8_to_NI;
wire[3:0] Tile_X8Y8_to_SA;
wire[3:0] Tile_X8Y8_to_SB;
wire[3:0] Tile_X8Y8_to_SC;
wire[3:0] Tile_X8Y8_to_SD;
wire[3:0] Tile_X8Y8_to_SF;
wire[7:0] Tile_X8Y8_to_SG;
wire[7:0] Tile_X8Y8_to_SH;
wire[11:0] Tile_X8Y8_to_SI;
wire[1:0] Tile_X9Y8_to_EA_1s;
wire[1:0] Tile_X9Y8_to_EB_1s;
wire[1:0] Tile_X9Y8_to_EC_1s;
wire[1:0] Tile_X9Y8_to_ED_1s;
wire[1:0] Tile_X9Y8_to_EF_1s;
wire[1:0] Tile_X9Y8_to_EG_1s;
wire[1:0] Tile_X9Y8_to_EH_1s;
wire[1:0] Tile_X9Y8_to_EI_1s;
wire[1:0] Tile_X9Y8_to_WA_1s;
wire[1:0] Tile_X9Y8_to_WB_1s;
wire[1:0] Tile_X9Y8_to_WC_1s;
wire[1:0] Tile_X9Y8_to_WD_1s;
wire[1:0] Tile_X9Y8_to_WF_1s;
wire[1:0] Tile_X9Y8_to_WG_1s;
wire[1:0] Tile_X9Y8_to_WH_1s;
wire[1:0] Tile_X9Y8_to_WI_1s;
wire[1:0] Tile_X9Y8_to_NA_1s;
wire[1:0] Tile_X9Y8_to_NB_1s;
wire[1:0] Tile_X9Y8_to_NC_1s;
wire[1:0] Tile_X9Y8_to_ND_1s;
wire[1:0] Tile_X9Y8_to_NF_1s;
wire[1:0] Tile_X9Y8_to_NG_1s;
wire[1:0] Tile_X9Y8_to_NH_1s;
wire[1:0] Tile_X9Y8_to_NI_1s;
wire[1:0] Tile_X9Y8_to_SA_1s;
wire[1:0] Tile_X9Y8_to_SB_1s;
wire[1:0] Tile_X9Y8_to_SC_1s;
wire[1:0] Tile_X9Y8_to_SD_1s;
wire[1:0] Tile_X9Y8_to_SF_1s;
wire[1:0] Tile_X9Y8_to_SG_1s;
wire[1:0] Tile_X9Y8_to_SH_1s;
wire[1:0] Tile_X9Y8_to_SI_1s;
wire[1:0] Tile_X10Y8_to_WA_1s;
wire[1:0] Tile_X10Y8_to_WB_1s;
wire[1:0] Tile_X10Y8_to_WC_1s;
wire[1:0] Tile_X10Y8_to_WD_1s;
wire[1:0] Tile_X10Y8_to_WF_1s;
wire[1:0] Tile_X10Y8_to_WG_1s;
wire[1:0] Tile_X10Y8_to_WH_1s;
wire[1:0] Tile_X10Y8_to_WI_1s;
wire[3:0] Tile_X0Y9_to_EA;
wire[3:0] Tile_X0Y9_to_EB;
wire[3:0] Tile_X0Y9_to_EC;
wire[3:0] Tile_X0Y9_to_ED;
wire[3:0] Tile_X0Y9_to_EF;
wire[7:0] Tile_X0Y9_to_EG;
wire[7:0] Tile_X0Y9_to_EH;
wire[11:0] Tile_X0Y9_to_EI;
wire[3:0] Tile_X0Y9_to_NA;
wire[3:0] Tile_X0Y9_to_NB;
wire[3:0] Tile_X0Y9_to_NC;
wire[3:0] Tile_X0Y9_to_ND;
wire[3:0] Tile_X0Y9_to_NF;
wire[7:0] Tile_X0Y9_to_NG;
wire[7:0] Tile_X0Y9_to_NH;
wire[11:0] Tile_X0Y9_to_NI;
wire[3:0] Tile_X0Y9_to_SA;
wire[3:0] Tile_X0Y9_to_SB;
wire[3:0] Tile_X0Y9_to_SC;
wire[3:0] Tile_X0Y9_to_SD;
wire[3:0] Tile_X0Y9_to_SF;
wire[7:0] Tile_X0Y9_to_SG;
wire[7:0] Tile_X0Y9_to_SH;
wire[11:0] Tile_X0Y9_to_SI;
wire[3:0] Tile_X1Y9_to_EA;
wire[3:0] Tile_X1Y9_to_EB;
wire[3:0] Tile_X1Y9_to_EC;
wire[3:0] Tile_X1Y9_to_ED;
wire[3:0] Tile_X1Y9_to_EF;
wire[7:0] Tile_X1Y9_to_EG;
wire[7:0] Tile_X1Y9_to_EH;
wire[11:0] Tile_X1Y9_to_EI;
wire[3:0] Tile_X1Y9_to_WA;
wire[3:0] Tile_X1Y9_to_WB;
wire[3:0] Tile_X1Y9_to_WC;
wire[3:0] Tile_X1Y9_to_WD;
wire[3:0] Tile_X1Y9_to_WF;
wire[7:0] Tile_X1Y9_to_WG;
wire[7:0] Tile_X1Y9_to_WH;
wire[11:0] Tile_X1Y9_to_WI;
wire[3:0] Tile_X1Y9_to_NA;
wire[3:0] Tile_X1Y9_to_NB;
wire[3:0] Tile_X1Y9_to_NC;
wire[3:0] Tile_X1Y9_to_ND;
wire[3:0] Tile_X1Y9_to_NF;
wire[7:0] Tile_X1Y9_to_NG;
wire[7:0] Tile_X1Y9_to_NH;
wire[11:0] Tile_X1Y9_to_NI;
wire[3:0] Tile_X1Y9_to_SA;
wire[3:0] Tile_X1Y9_to_SB;
wire[3:0] Tile_X1Y9_to_SC;
wire[3:0] Tile_X1Y9_to_SD;
wire[3:0] Tile_X1Y9_to_SF;
wire[7:0] Tile_X1Y9_to_SG;
wire[7:0] Tile_X1Y9_to_SH;
wire[11:0] Tile_X1Y9_to_SI;
wire[3:0] Tile_X2Y9_to_EA;
wire[3:0] Tile_X2Y9_to_EB;
wire[3:0] Tile_X2Y9_to_EC;
wire[3:0] Tile_X2Y9_to_ED;
wire[3:0] Tile_X2Y9_to_EF;
wire[7:0] Tile_X2Y9_to_EG;
wire[7:0] Tile_X2Y9_to_EH;
wire[11:0] Tile_X2Y9_to_EI;
wire[3:0] Tile_X2Y9_to_WA;
wire[3:0] Tile_X2Y9_to_WB;
wire[3:0] Tile_X2Y9_to_WC;
wire[3:0] Tile_X2Y9_to_WD;
wire[3:0] Tile_X2Y9_to_WF;
wire[7:0] Tile_X2Y9_to_WG;
wire[7:0] Tile_X2Y9_to_WH;
wire[11:0] Tile_X2Y9_to_WI;
wire[3:0] Tile_X2Y9_to_NA;
wire[3:0] Tile_X2Y9_to_NB;
wire[3:0] Tile_X2Y9_to_NC;
wire[3:0] Tile_X2Y9_to_ND;
wire[3:0] Tile_X2Y9_to_NF;
wire[7:0] Tile_X2Y9_to_NG;
wire[7:0] Tile_X2Y9_to_NH;
wire[11:0] Tile_X2Y9_to_NI;
wire[3:0] Tile_X2Y9_to_SA;
wire[3:0] Tile_X2Y9_to_SB;
wire[3:0] Tile_X2Y9_to_SC;
wire[3:0] Tile_X2Y9_to_SD;
wire[3:0] Tile_X2Y9_to_SF;
wire[7:0] Tile_X2Y9_to_SG;
wire[7:0] Tile_X2Y9_to_SH;
wire[11:0] Tile_X2Y9_to_SI;
wire[3:0] Tile_X3Y9_to_EA;
wire[3:0] Tile_X3Y9_to_EB;
wire[3:0] Tile_X3Y9_to_EC;
wire[3:0] Tile_X3Y9_to_ED;
wire[3:0] Tile_X3Y9_to_EF;
wire[7:0] Tile_X3Y9_to_EG;
wire[7:0] Tile_X3Y9_to_EH;
wire[11:0] Tile_X3Y9_to_EI;
wire[3:0] Tile_X3Y9_to_WA;
wire[3:0] Tile_X3Y9_to_WB;
wire[3:0] Tile_X3Y9_to_WC;
wire[3:0] Tile_X3Y9_to_WD;
wire[3:0] Tile_X3Y9_to_WF;
wire[7:0] Tile_X3Y9_to_WG;
wire[7:0] Tile_X3Y9_to_WH;
wire[11:0] Tile_X3Y9_to_WI;
wire[3:0] Tile_X3Y9_to_NA;
wire[3:0] Tile_X3Y9_to_NB;
wire[3:0] Tile_X3Y9_to_NC;
wire[3:0] Tile_X3Y9_to_ND;
wire[3:0] Tile_X3Y9_to_NF;
wire[7:0] Tile_X3Y9_to_NG;
wire[7:0] Tile_X3Y9_to_NH;
wire[11:0] Tile_X3Y9_to_NI;
wire[3:0] Tile_X3Y9_to_SA;
wire[3:0] Tile_X3Y9_to_SB;
wire[3:0] Tile_X3Y9_to_SC;
wire[3:0] Tile_X3Y9_to_SD;
wire[3:0] Tile_X3Y9_to_SF;
wire[7:0] Tile_X3Y9_to_SG;
wire[7:0] Tile_X3Y9_to_SH;
wire[11:0] Tile_X3Y9_to_SI;
wire[3:0] Tile_X4Y9_to_EA;
wire[3:0] Tile_X4Y9_to_EB;
wire[3:0] Tile_X4Y9_to_EC;
wire[3:0] Tile_X4Y9_to_ED;
wire[3:0] Tile_X4Y9_to_EF;
wire[7:0] Tile_X4Y9_to_EG;
wire[7:0] Tile_X4Y9_to_EH;
wire[11:0] Tile_X4Y9_to_EI;
wire[3:0] Tile_X4Y9_to_WA;
wire[3:0] Tile_X4Y9_to_WB;
wire[3:0] Tile_X4Y9_to_WC;
wire[3:0] Tile_X4Y9_to_WD;
wire[3:0] Tile_X4Y9_to_WF;
wire[7:0] Tile_X4Y9_to_WG;
wire[7:0] Tile_X4Y9_to_WH;
wire[11:0] Tile_X4Y9_to_WI;
wire[3:0] Tile_X4Y9_to_NA;
wire[3:0] Tile_X4Y9_to_NB;
wire[3:0] Tile_X4Y9_to_NC;
wire[3:0] Tile_X4Y9_to_ND;
wire[3:0] Tile_X4Y9_to_NF;
wire[7:0] Tile_X4Y9_to_NG;
wire[7:0] Tile_X4Y9_to_NH;
wire[11:0] Tile_X4Y9_to_NI;
wire[3:0] Tile_X4Y9_to_SA;
wire[3:0] Tile_X4Y9_to_SB;
wire[3:0] Tile_X4Y9_to_SC;
wire[3:0] Tile_X4Y9_to_SD;
wire[3:0] Tile_X4Y9_to_SF;
wire[7:0] Tile_X4Y9_to_SG;
wire[7:0] Tile_X4Y9_to_SH;
wire[11:0] Tile_X4Y9_to_SI;
wire[3:0] Tile_X5Y9_to_EA;
wire[3:0] Tile_X5Y9_to_EB;
wire[3:0] Tile_X5Y9_to_EC;
wire[3:0] Tile_X5Y9_to_ED;
wire[3:0] Tile_X5Y9_to_EF;
wire[7:0] Tile_X5Y9_to_EG;
wire[7:0] Tile_X5Y9_to_EH;
wire[11:0] Tile_X5Y9_to_EI;
wire[3:0] Tile_X5Y9_to_WA;
wire[3:0] Tile_X5Y9_to_WB;
wire[3:0] Tile_X5Y9_to_WC;
wire[3:0] Tile_X5Y9_to_WD;
wire[3:0] Tile_X5Y9_to_WF;
wire[7:0] Tile_X5Y9_to_WG;
wire[7:0] Tile_X5Y9_to_WH;
wire[11:0] Tile_X5Y9_to_WI;
wire[3:0] Tile_X5Y9_to_NA;
wire[3:0] Tile_X5Y9_to_NB;
wire[3:0] Tile_X5Y9_to_NC;
wire[3:0] Tile_X5Y9_to_ND;
wire[3:0] Tile_X5Y9_to_NF;
wire[7:0] Tile_X5Y9_to_NG;
wire[7:0] Tile_X5Y9_to_NH;
wire[11:0] Tile_X5Y9_to_NI;
wire[3:0] Tile_X5Y9_to_SA;
wire[3:0] Tile_X5Y9_to_SB;
wire[3:0] Tile_X5Y9_to_SC;
wire[3:0] Tile_X5Y9_to_SD;
wire[3:0] Tile_X5Y9_to_SF;
wire[7:0] Tile_X5Y9_to_SG;
wire[7:0] Tile_X5Y9_to_SH;
wire[11:0] Tile_X5Y9_to_SI;
wire[3:0] Tile_X6Y9_to_EA;
wire[3:0] Tile_X6Y9_to_EB;
wire[3:0] Tile_X6Y9_to_EC;
wire[3:0] Tile_X6Y9_to_ED;
wire[3:0] Tile_X6Y9_to_EF;
wire[7:0] Tile_X6Y9_to_EG;
wire[7:0] Tile_X6Y9_to_EH;
wire[11:0] Tile_X6Y9_to_EI;
wire[3:0] Tile_X6Y9_to_WA;
wire[3:0] Tile_X6Y9_to_WB;
wire[3:0] Tile_X6Y9_to_WC;
wire[3:0] Tile_X6Y9_to_WD;
wire[3:0] Tile_X6Y9_to_WF;
wire[7:0] Tile_X6Y9_to_WG;
wire[7:0] Tile_X6Y9_to_WH;
wire[11:0] Tile_X6Y9_to_WI;
wire[3:0] Tile_X6Y9_to_NA;
wire[3:0] Tile_X6Y9_to_NB;
wire[3:0] Tile_X6Y9_to_NC;
wire[3:0] Tile_X6Y9_to_ND;
wire[3:0] Tile_X6Y9_to_NF;
wire[7:0] Tile_X6Y9_to_NG;
wire[7:0] Tile_X6Y9_to_NH;
wire[11:0] Tile_X6Y9_to_NI;
wire[3:0] Tile_X6Y9_to_SA;
wire[3:0] Tile_X6Y9_to_SB;
wire[3:0] Tile_X6Y9_to_SC;
wire[3:0] Tile_X6Y9_to_SD;
wire[3:0] Tile_X6Y9_to_SF;
wire[7:0] Tile_X6Y9_to_SG;
wire[7:0] Tile_X6Y9_to_SH;
wire[11:0] Tile_X6Y9_to_SI;
wire[3:0] Tile_X7Y9_to_EA;
wire[3:0] Tile_X7Y9_to_EB;
wire[3:0] Tile_X7Y9_to_EC;
wire[3:0] Tile_X7Y9_to_ED;
wire[3:0] Tile_X7Y9_to_EF;
wire[7:0] Tile_X7Y9_to_EG;
wire[7:0] Tile_X7Y9_to_EH;
wire[11:0] Tile_X7Y9_to_EI;
wire[3:0] Tile_X7Y9_to_WA;
wire[3:0] Tile_X7Y9_to_WB;
wire[3:0] Tile_X7Y9_to_WC;
wire[3:0] Tile_X7Y9_to_WD;
wire[3:0] Tile_X7Y9_to_WF;
wire[7:0] Tile_X7Y9_to_WG;
wire[7:0] Tile_X7Y9_to_WH;
wire[11:0] Tile_X7Y9_to_WI;
wire[3:0] Tile_X7Y9_to_NA;
wire[3:0] Tile_X7Y9_to_NB;
wire[3:0] Tile_X7Y9_to_NC;
wire[3:0] Tile_X7Y9_to_ND;
wire[3:0] Tile_X7Y9_to_NF;
wire[7:0] Tile_X7Y9_to_NG;
wire[7:0] Tile_X7Y9_to_NH;
wire[11:0] Tile_X7Y9_to_NI;
wire[3:0] Tile_X7Y9_to_SA;
wire[3:0] Tile_X7Y9_to_SB;
wire[3:0] Tile_X7Y9_to_SC;
wire[3:0] Tile_X7Y9_to_SD;
wire[3:0] Tile_X7Y9_to_SF;
wire[7:0] Tile_X7Y9_to_SG;
wire[7:0] Tile_X7Y9_to_SH;
wire[11:0] Tile_X7Y9_to_SI;
wire[3:0] Tile_X8Y9_to_WA;
wire[3:0] Tile_X8Y9_to_WB;
wire[3:0] Tile_X8Y9_to_WC;
wire[3:0] Tile_X8Y9_to_WD;
wire[3:0] Tile_X8Y9_to_WF;
wire[7:0] Tile_X8Y9_to_WG;
wire[7:0] Tile_X8Y9_to_WH;
wire[11:0] Tile_X8Y9_to_WI;
wire[3:0] Tile_X8Y9_to_NA;
wire[3:0] Tile_X8Y9_to_NB;
wire[3:0] Tile_X8Y9_to_NC;
wire[3:0] Tile_X8Y9_to_ND;
wire[3:0] Tile_X8Y9_to_NF;
wire[7:0] Tile_X8Y9_to_NG;
wire[7:0] Tile_X8Y9_to_NH;
wire[11:0] Tile_X8Y9_to_NI;
wire[3:0] Tile_X8Y9_to_SA;
wire[3:0] Tile_X8Y9_to_SB;
wire[3:0] Tile_X8Y9_to_SC;
wire[3:0] Tile_X8Y9_to_SD;
wire[3:0] Tile_X8Y9_to_SF;
wire[7:0] Tile_X8Y9_to_SG;
wire[7:0] Tile_X8Y9_to_SH;
wire[11:0] Tile_X8Y9_to_SI;
wire[1:0] Tile_X9Y9_to_EA_1s;
wire[1:0] Tile_X9Y9_to_EB_1s;
wire[1:0] Tile_X9Y9_to_EC_1s;
wire[1:0] Tile_X9Y9_to_ED_1s;
wire[1:0] Tile_X9Y9_to_EF_1s;
wire[1:0] Tile_X9Y9_to_EG_1s;
wire[1:0] Tile_X9Y9_to_EH_1s;
wire[1:0] Tile_X9Y9_to_EI_1s;
wire[1:0] Tile_X9Y9_to_WA_1s;
wire[1:0] Tile_X9Y9_to_WB_1s;
wire[1:0] Tile_X9Y9_to_WC_1s;
wire[1:0] Tile_X9Y9_to_WD_1s;
wire[1:0] Tile_X9Y9_to_WF_1s;
wire[1:0] Tile_X9Y9_to_WG_1s;
wire[1:0] Tile_X9Y9_to_WH_1s;
wire[1:0] Tile_X9Y9_to_WI_1s;
wire[1:0] Tile_X9Y9_to_NA_1s;
wire[1:0] Tile_X9Y9_to_NB_1s;
wire[1:0] Tile_X9Y9_to_NC_1s;
wire[1:0] Tile_X9Y9_to_ND_1s;
wire[1:0] Tile_X9Y9_to_NF_1s;
wire[1:0] Tile_X9Y9_to_NG_1s;
wire[1:0] Tile_X9Y9_to_NH_1s;
wire[1:0] Tile_X9Y9_to_NI_1s;
wire[1:0] Tile_X9Y9_to_SA_1s;
wire[1:0] Tile_X9Y9_to_SB_1s;
wire[1:0] Tile_X9Y9_to_SC_1s;
wire[1:0] Tile_X9Y9_to_SD_1s;
wire[1:0] Tile_X9Y9_to_SF_1s;
wire[1:0] Tile_X9Y9_to_SG_1s;
wire[1:0] Tile_X9Y9_to_SH_1s;
wire[1:0] Tile_X9Y9_to_SI_1s;
wire[1:0] Tile_X10Y9_to_WA_1s;
wire[1:0] Tile_X10Y9_to_WB_1s;
wire[1:0] Tile_X10Y9_to_WC_1s;
wire[1:0] Tile_X10Y9_to_WD_1s;
wire[1:0] Tile_X10Y9_to_WF_1s;
wire[1:0] Tile_X10Y9_to_WG_1s;
wire[1:0] Tile_X10Y9_to_WH_1s;
wire[1:0] Tile_X10Y9_to_WI_1s;
wire[3:0] Tile_X0Y10_to_EA;
wire[3:0] Tile_X0Y10_to_EB;
wire[3:0] Tile_X0Y10_to_EC;
wire[3:0] Tile_X0Y10_to_ED;
wire[3:0] Tile_X0Y10_to_EF;
wire[7:0] Tile_X0Y10_to_EG;
wire[7:0] Tile_X0Y10_to_EH;
wire[11:0] Tile_X0Y10_to_EI;
wire[3:0] Tile_X0Y10_to_NA;
wire[3:0] Tile_X0Y10_to_NB;
wire[3:0] Tile_X0Y10_to_NC;
wire[3:0] Tile_X0Y10_to_ND;
wire[3:0] Tile_X0Y10_to_NF;
wire[7:0] Tile_X0Y10_to_NG;
wire[7:0] Tile_X0Y10_to_NH;
wire[11:0] Tile_X0Y10_to_NI;
wire[3:0] Tile_X0Y10_to_SA;
wire[3:0] Tile_X0Y10_to_SB;
wire[3:0] Tile_X0Y10_to_SC;
wire[3:0] Tile_X0Y10_to_SD;
wire[3:0] Tile_X0Y10_to_SF;
wire[7:0] Tile_X0Y10_to_SG;
wire[7:0] Tile_X0Y10_to_SH;
wire[11:0] Tile_X0Y10_to_SI;
wire[3:0] Tile_X1Y10_to_EA;
wire[3:0] Tile_X1Y10_to_EB;
wire[3:0] Tile_X1Y10_to_EC;
wire[3:0] Tile_X1Y10_to_ED;
wire[3:0] Tile_X1Y10_to_EF;
wire[7:0] Tile_X1Y10_to_EG;
wire[7:0] Tile_X1Y10_to_EH;
wire[11:0] Tile_X1Y10_to_EI;
wire[3:0] Tile_X1Y10_to_WA;
wire[3:0] Tile_X1Y10_to_WB;
wire[3:0] Tile_X1Y10_to_WC;
wire[3:0] Tile_X1Y10_to_WD;
wire[3:0] Tile_X1Y10_to_WF;
wire[7:0] Tile_X1Y10_to_WG;
wire[7:0] Tile_X1Y10_to_WH;
wire[11:0] Tile_X1Y10_to_WI;
wire[3:0] Tile_X1Y10_to_NA;
wire[3:0] Tile_X1Y10_to_NB;
wire[3:0] Tile_X1Y10_to_NC;
wire[3:0] Tile_X1Y10_to_ND;
wire[3:0] Tile_X1Y10_to_NF;
wire[7:0] Tile_X1Y10_to_NG;
wire[7:0] Tile_X1Y10_to_NH;
wire[11:0] Tile_X1Y10_to_NI;
wire[3:0] Tile_X1Y10_to_SA;
wire[3:0] Tile_X1Y10_to_SB;
wire[3:0] Tile_X1Y10_to_SC;
wire[3:0] Tile_X1Y10_to_SD;
wire[3:0] Tile_X1Y10_to_SF;
wire[7:0] Tile_X1Y10_to_SG;
wire[7:0] Tile_X1Y10_to_SH;
wire[11:0] Tile_X1Y10_to_SI;
wire[3:0] Tile_X2Y10_to_EA;
wire[3:0] Tile_X2Y10_to_EB;
wire[3:0] Tile_X2Y10_to_EC;
wire[3:0] Tile_X2Y10_to_ED;
wire[3:0] Tile_X2Y10_to_EF;
wire[7:0] Tile_X2Y10_to_EG;
wire[7:0] Tile_X2Y10_to_EH;
wire[11:0] Tile_X2Y10_to_EI;
wire[3:0] Tile_X2Y10_to_WA;
wire[3:0] Tile_X2Y10_to_WB;
wire[3:0] Tile_X2Y10_to_WC;
wire[3:0] Tile_X2Y10_to_WD;
wire[3:0] Tile_X2Y10_to_WF;
wire[7:0] Tile_X2Y10_to_WG;
wire[7:0] Tile_X2Y10_to_WH;
wire[11:0] Tile_X2Y10_to_WI;
wire[3:0] Tile_X2Y10_to_NA;
wire[3:0] Tile_X2Y10_to_NB;
wire[3:0] Tile_X2Y10_to_NC;
wire[3:0] Tile_X2Y10_to_ND;
wire[3:0] Tile_X2Y10_to_NF;
wire[7:0] Tile_X2Y10_to_NG;
wire[7:0] Tile_X2Y10_to_NH;
wire[11:0] Tile_X2Y10_to_NI;
wire[3:0] Tile_X2Y10_to_SA;
wire[3:0] Tile_X2Y10_to_SB;
wire[3:0] Tile_X2Y10_to_SC;
wire[3:0] Tile_X2Y10_to_SD;
wire[3:0] Tile_X2Y10_to_SF;
wire[7:0] Tile_X2Y10_to_SG;
wire[7:0] Tile_X2Y10_to_SH;
wire[11:0] Tile_X2Y10_to_SI;
wire[3:0] Tile_X3Y10_to_EA;
wire[3:0] Tile_X3Y10_to_EB;
wire[3:0] Tile_X3Y10_to_EC;
wire[3:0] Tile_X3Y10_to_ED;
wire[3:0] Tile_X3Y10_to_EF;
wire[7:0] Tile_X3Y10_to_EG;
wire[7:0] Tile_X3Y10_to_EH;
wire[11:0] Tile_X3Y10_to_EI;
wire[3:0] Tile_X3Y10_to_WA;
wire[3:0] Tile_X3Y10_to_WB;
wire[3:0] Tile_X3Y10_to_WC;
wire[3:0] Tile_X3Y10_to_WD;
wire[3:0] Tile_X3Y10_to_WF;
wire[7:0] Tile_X3Y10_to_WG;
wire[7:0] Tile_X3Y10_to_WH;
wire[11:0] Tile_X3Y10_to_WI;
wire[3:0] Tile_X3Y10_to_NA;
wire[3:0] Tile_X3Y10_to_NB;
wire[3:0] Tile_X3Y10_to_NC;
wire[3:0] Tile_X3Y10_to_ND;
wire[3:0] Tile_X3Y10_to_NF;
wire[7:0] Tile_X3Y10_to_NG;
wire[7:0] Tile_X3Y10_to_NH;
wire[11:0] Tile_X3Y10_to_NI;
wire[3:0] Tile_X3Y10_to_SA;
wire[3:0] Tile_X3Y10_to_SB;
wire[3:0] Tile_X3Y10_to_SC;
wire[3:0] Tile_X3Y10_to_SD;
wire[3:0] Tile_X3Y10_to_SF;
wire[7:0] Tile_X3Y10_to_SG;
wire[7:0] Tile_X3Y10_to_SH;
wire[11:0] Tile_X3Y10_to_SI;
wire[3:0] Tile_X4Y10_to_EA;
wire[3:0] Tile_X4Y10_to_EB;
wire[3:0] Tile_X4Y10_to_EC;
wire[3:0] Tile_X4Y10_to_ED;
wire[3:0] Tile_X4Y10_to_EF;
wire[7:0] Tile_X4Y10_to_EG;
wire[7:0] Tile_X4Y10_to_EH;
wire[11:0] Tile_X4Y10_to_EI;
wire[3:0] Tile_X4Y10_to_WA;
wire[3:0] Tile_X4Y10_to_WB;
wire[3:0] Tile_X4Y10_to_WC;
wire[3:0] Tile_X4Y10_to_WD;
wire[3:0] Tile_X4Y10_to_WF;
wire[7:0] Tile_X4Y10_to_WG;
wire[7:0] Tile_X4Y10_to_WH;
wire[11:0] Tile_X4Y10_to_WI;
wire[3:0] Tile_X4Y10_to_NA;
wire[3:0] Tile_X4Y10_to_NB;
wire[3:0] Tile_X4Y10_to_NC;
wire[3:0] Tile_X4Y10_to_ND;
wire[3:0] Tile_X4Y10_to_NF;
wire[7:0] Tile_X4Y10_to_NG;
wire[7:0] Tile_X4Y10_to_NH;
wire[11:0] Tile_X4Y10_to_NI;
wire[3:0] Tile_X4Y10_to_SA;
wire[3:0] Tile_X4Y10_to_SB;
wire[3:0] Tile_X4Y10_to_SC;
wire[3:0] Tile_X4Y10_to_SD;
wire[3:0] Tile_X4Y10_to_SF;
wire[7:0] Tile_X4Y10_to_SG;
wire[7:0] Tile_X4Y10_to_SH;
wire[11:0] Tile_X4Y10_to_SI;
wire[3:0] Tile_X5Y10_to_EA;
wire[3:0] Tile_X5Y10_to_EB;
wire[3:0] Tile_X5Y10_to_EC;
wire[3:0] Tile_X5Y10_to_ED;
wire[3:0] Tile_X5Y10_to_EF;
wire[7:0] Tile_X5Y10_to_EG;
wire[7:0] Tile_X5Y10_to_EH;
wire[11:0] Tile_X5Y10_to_EI;
wire[3:0] Tile_X5Y10_to_WA;
wire[3:0] Tile_X5Y10_to_WB;
wire[3:0] Tile_X5Y10_to_WC;
wire[3:0] Tile_X5Y10_to_WD;
wire[3:0] Tile_X5Y10_to_WF;
wire[7:0] Tile_X5Y10_to_WG;
wire[7:0] Tile_X5Y10_to_WH;
wire[11:0] Tile_X5Y10_to_WI;
wire[3:0] Tile_X5Y10_to_NA;
wire[3:0] Tile_X5Y10_to_NB;
wire[3:0] Tile_X5Y10_to_NC;
wire[3:0] Tile_X5Y10_to_ND;
wire[3:0] Tile_X5Y10_to_NF;
wire[7:0] Tile_X5Y10_to_NG;
wire[7:0] Tile_X5Y10_to_NH;
wire[11:0] Tile_X5Y10_to_NI;
wire[3:0] Tile_X5Y10_to_SA;
wire[3:0] Tile_X5Y10_to_SB;
wire[3:0] Tile_X5Y10_to_SC;
wire[3:0] Tile_X5Y10_to_SD;
wire[3:0] Tile_X5Y10_to_SF;
wire[7:0] Tile_X5Y10_to_SG;
wire[7:0] Tile_X5Y10_to_SH;
wire[11:0] Tile_X5Y10_to_SI;
wire[3:0] Tile_X6Y10_to_EA;
wire[3:0] Tile_X6Y10_to_EB;
wire[3:0] Tile_X6Y10_to_EC;
wire[3:0] Tile_X6Y10_to_ED;
wire[3:0] Tile_X6Y10_to_EF;
wire[7:0] Tile_X6Y10_to_EG;
wire[7:0] Tile_X6Y10_to_EH;
wire[11:0] Tile_X6Y10_to_EI;
wire[3:0] Tile_X6Y10_to_WA;
wire[3:0] Tile_X6Y10_to_WB;
wire[3:0] Tile_X6Y10_to_WC;
wire[3:0] Tile_X6Y10_to_WD;
wire[3:0] Tile_X6Y10_to_WF;
wire[7:0] Tile_X6Y10_to_WG;
wire[7:0] Tile_X6Y10_to_WH;
wire[11:0] Tile_X6Y10_to_WI;
wire[3:0] Tile_X6Y10_to_NA;
wire[3:0] Tile_X6Y10_to_NB;
wire[3:0] Tile_X6Y10_to_NC;
wire[3:0] Tile_X6Y10_to_ND;
wire[3:0] Tile_X6Y10_to_NF;
wire[7:0] Tile_X6Y10_to_NG;
wire[7:0] Tile_X6Y10_to_NH;
wire[11:0] Tile_X6Y10_to_NI;
wire[3:0] Tile_X6Y10_to_SA;
wire[3:0] Tile_X6Y10_to_SB;
wire[3:0] Tile_X6Y10_to_SC;
wire[3:0] Tile_X6Y10_to_SD;
wire[3:0] Tile_X6Y10_to_SF;
wire[7:0] Tile_X6Y10_to_SG;
wire[7:0] Tile_X6Y10_to_SH;
wire[11:0] Tile_X6Y10_to_SI;
wire[3:0] Tile_X7Y10_to_EA;
wire[3:0] Tile_X7Y10_to_EB;
wire[3:0] Tile_X7Y10_to_EC;
wire[3:0] Tile_X7Y10_to_ED;
wire[3:0] Tile_X7Y10_to_EF;
wire[7:0] Tile_X7Y10_to_EG;
wire[7:0] Tile_X7Y10_to_EH;
wire[11:0] Tile_X7Y10_to_EI;
wire[3:0] Tile_X7Y10_to_WA;
wire[3:0] Tile_X7Y10_to_WB;
wire[3:0] Tile_X7Y10_to_WC;
wire[3:0] Tile_X7Y10_to_WD;
wire[3:0] Tile_X7Y10_to_WF;
wire[7:0] Tile_X7Y10_to_WG;
wire[7:0] Tile_X7Y10_to_WH;
wire[11:0] Tile_X7Y10_to_WI;
wire[3:0] Tile_X7Y10_to_NA;
wire[3:0] Tile_X7Y10_to_NB;
wire[3:0] Tile_X7Y10_to_NC;
wire[3:0] Tile_X7Y10_to_ND;
wire[3:0] Tile_X7Y10_to_NF;
wire[7:0] Tile_X7Y10_to_NG;
wire[7:0] Tile_X7Y10_to_NH;
wire[11:0] Tile_X7Y10_to_NI;
wire[3:0] Tile_X7Y10_to_SA;
wire[3:0] Tile_X7Y10_to_SB;
wire[3:0] Tile_X7Y10_to_SC;
wire[3:0] Tile_X7Y10_to_SD;
wire[3:0] Tile_X7Y10_to_SF;
wire[7:0] Tile_X7Y10_to_SG;
wire[7:0] Tile_X7Y10_to_SH;
wire[11:0] Tile_X7Y10_to_SI;
wire[3:0] Tile_X8Y10_to_WA;
wire[3:0] Tile_X8Y10_to_WB;
wire[3:0] Tile_X8Y10_to_WC;
wire[3:0] Tile_X8Y10_to_WD;
wire[3:0] Tile_X8Y10_to_WF;
wire[7:0] Tile_X8Y10_to_WG;
wire[7:0] Tile_X8Y10_to_WH;
wire[11:0] Tile_X8Y10_to_WI;
wire[3:0] Tile_X8Y10_to_NA;
wire[3:0] Tile_X8Y10_to_NB;
wire[3:0] Tile_X8Y10_to_NC;
wire[3:0] Tile_X8Y10_to_ND;
wire[3:0] Tile_X8Y10_to_NF;
wire[7:0] Tile_X8Y10_to_NG;
wire[7:0] Tile_X8Y10_to_NH;
wire[11:0] Tile_X8Y10_to_NI;
wire[3:0] Tile_X8Y10_to_SA;
wire[3:0] Tile_X8Y10_to_SB;
wire[3:0] Tile_X8Y10_to_SC;
wire[3:0] Tile_X8Y10_to_SD;
wire[3:0] Tile_X8Y10_to_SF;
wire[7:0] Tile_X8Y10_to_SG;
wire[7:0] Tile_X8Y10_to_SH;
wire[11:0] Tile_X8Y10_to_SI;
wire[1:0] Tile_X9Y10_to_EA_1s;
wire[1:0] Tile_X9Y10_to_EB_1s;
wire[1:0] Tile_X9Y10_to_EC_1s;
wire[1:0] Tile_X9Y10_to_ED_1s;
wire[1:0] Tile_X9Y10_to_EF_1s;
wire[1:0] Tile_X9Y10_to_EG_1s;
wire[1:0] Tile_X9Y10_to_EH_1s;
wire[1:0] Tile_X9Y10_to_EI_1s;
wire[1:0] Tile_X9Y10_to_WA_1s;
wire[1:0] Tile_X9Y10_to_WB_1s;
wire[1:0] Tile_X9Y10_to_WC_1s;
wire[1:0] Tile_X9Y10_to_WD_1s;
wire[1:0] Tile_X9Y10_to_WF_1s;
wire[1:0] Tile_X9Y10_to_WG_1s;
wire[1:0] Tile_X9Y10_to_WH_1s;
wire[1:0] Tile_X9Y10_to_WI_1s;
wire[1:0] Tile_X9Y10_to_NA_1s;
wire[1:0] Tile_X9Y10_to_NB_1s;
wire[1:0] Tile_X9Y10_to_NC_1s;
wire[1:0] Tile_X9Y10_to_ND_1s;
wire[1:0] Tile_X9Y10_to_NF_1s;
wire[1:0] Tile_X9Y10_to_NG_1s;
wire[1:0] Tile_X9Y10_to_NH_1s;
wire[1:0] Tile_X9Y10_to_NI_1s;
wire[1:0] Tile_X9Y10_to_SA_1s;
wire[1:0] Tile_X9Y10_to_SB_1s;
wire[1:0] Tile_X9Y10_to_SC_1s;
wire[1:0] Tile_X9Y10_to_SD_1s;
wire[1:0] Tile_X9Y10_to_SF_1s;
wire[1:0] Tile_X9Y10_to_SG_1s;
wire[1:0] Tile_X9Y10_to_SH_1s;
wire[1:0] Tile_X9Y10_to_SI_1s;
wire[1:0] Tile_X10Y10_to_WA_1s;
wire[1:0] Tile_X10Y10_to_WB_1s;
wire[1:0] Tile_X10Y10_to_WC_1s;
wire[1:0] Tile_X10Y10_to_WD_1s;
wire[1:0] Tile_X10Y10_to_WF_1s;
wire[1:0] Tile_X10Y10_to_WG_1s;
wire[1:0] Tile_X10Y10_to_WH_1s;
wire[1:0] Tile_X10Y10_to_WI_1s;
wire[3:0] Tile_X0Y11_to_EA;
wire[3:0] Tile_X0Y11_to_EB;
wire[3:0] Tile_X0Y11_to_EC;
wire[3:0] Tile_X0Y11_to_ED;
wire[3:0] Tile_X0Y11_to_EF;
wire[7:0] Tile_X0Y11_to_EG;
wire[7:0] Tile_X0Y11_to_EH;
wire[11:0] Tile_X0Y11_to_EI;
wire[3:0] Tile_X0Y11_to_NA;
wire[3:0] Tile_X0Y11_to_NB;
wire[3:0] Tile_X0Y11_to_NC;
wire[3:0] Tile_X0Y11_to_ND;
wire[3:0] Tile_X0Y11_to_NF;
wire[7:0] Tile_X0Y11_to_NG;
wire[7:0] Tile_X0Y11_to_NH;
wire[11:0] Tile_X0Y11_to_NI;
wire[3:0] Tile_X0Y11_to_SA;
wire[3:0] Tile_X0Y11_to_SB;
wire[3:0] Tile_X0Y11_to_SC;
wire[3:0] Tile_X0Y11_to_SD;
wire[3:0] Tile_X0Y11_to_SF;
wire[7:0] Tile_X0Y11_to_SG;
wire[7:0] Tile_X0Y11_to_SH;
wire[11:0] Tile_X0Y11_to_SI;
wire[3:0] Tile_X1Y11_to_EA;
wire[3:0] Tile_X1Y11_to_EB;
wire[3:0] Tile_X1Y11_to_EC;
wire[3:0] Tile_X1Y11_to_ED;
wire[3:0] Tile_X1Y11_to_EF;
wire[7:0] Tile_X1Y11_to_EG;
wire[7:0] Tile_X1Y11_to_EH;
wire[11:0] Tile_X1Y11_to_EI;
wire[3:0] Tile_X1Y11_to_WA;
wire[3:0] Tile_X1Y11_to_WB;
wire[3:0] Tile_X1Y11_to_WC;
wire[3:0] Tile_X1Y11_to_WD;
wire[3:0] Tile_X1Y11_to_WF;
wire[7:0] Tile_X1Y11_to_WG;
wire[7:0] Tile_X1Y11_to_WH;
wire[11:0] Tile_X1Y11_to_WI;
wire[3:0] Tile_X1Y11_to_NA;
wire[3:0] Tile_X1Y11_to_NB;
wire[3:0] Tile_X1Y11_to_NC;
wire[3:0] Tile_X1Y11_to_ND;
wire[3:0] Tile_X1Y11_to_NF;
wire[7:0] Tile_X1Y11_to_NG;
wire[7:0] Tile_X1Y11_to_NH;
wire[11:0] Tile_X1Y11_to_NI;
wire[3:0] Tile_X1Y11_to_SA;
wire[3:0] Tile_X1Y11_to_SB;
wire[3:0] Tile_X1Y11_to_SC;
wire[3:0] Tile_X1Y11_to_SD;
wire[3:0] Tile_X1Y11_to_SF;
wire[7:0] Tile_X1Y11_to_SG;
wire[7:0] Tile_X1Y11_to_SH;
wire[11:0] Tile_X1Y11_to_SI;
wire[3:0] Tile_X2Y11_to_EA;
wire[3:0] Tile_X2Y11_to_EB;
wire[3:0] Tile_X2Y11_to_EC;
wire[3:0] Tile_X2Y11_to_ED;
wire[3:0] Tile_X2Y11_to_EF;
wire[7:0] Tile_X2Y11_to_EG;
wire[7:0] Tile_X2Y11_to_EH;
wire[11:0] Tile_X2Y11_to_EI;
wire[3:0] Tile_X2Y11_to_WA;
wire[3:0] Tile_X2Y11_to_WB;
wire[3:0] Tile_X2Y11_to_WC;
wire[3:0] Tile_X2Y11_to_WD;
wire[3:0] Tile_X2Y11_to_WF;
wire[7:0] Tile_X2Y11_to_WG;
wire[7:0] Tile_X2Y11_to_WH;
wire[11:0] Tile_X2Y11_to_WI;
wire[3:0] Tile_X2Y11_to_NA;
wire[3:0] Tile_X2Y11_to_NB;
wire[3:0] Tile_X2Y11_to_NC;
wire[3:0] Tile_X2Y11_to_ND;
wire[3:0] Tile_X2Y11_to_NF;
wire[7:0] Tile_X2Y11_to_NG;
wire[7:0] Tile_X2Y11_to_NH;
wire[11:0] Tile_X2Y11_to_NI;
wire[3:0] Tile_X2Y11_to_SA;
wire[3:0] Tile_X2Y11_to_SB;
wire[3:0] Tile_X2Y11_to_SC;
wire[3:0] Tile_X2Y11_to_SD;
wire[3:0] Tile_X2Y11_to_SF;
wire[7:0] Tile_X2Y11_to_SG;
wire[7:0] Tile_X2Y11_to_SH;
wire[11:0] Tile_X2Y11_to_SI;
wire[3:0] Tile_X3Y11_to_EA;
wire[3:0] Tile_X3Y11_to_EB;
wire[3:0] Tile_X3Y11_to_EC;
wire[3:0] Tile_X3Y11_to_ED;
wire[3:0] Tile_X3Y11_to_EF;
wire[7:0] Tile_X3Y11_to_EG;
wire[7:0] Tile_X3Y11_to_EH;
wire[11:0] Tile_X3Y11_to_EI;
wire[3:0] Tile_X3Y11_to_WA;
wire[3:0] Tile_X3Y11_to_WB;
wire[3:0] Tile_X3Y11_to_WC;
wire[3:0] Tile_X3Y11_to_WD;
wire[3:0] Tile_X3Y11_to_WF;
wire[7:0] Tile_X3Y11_to_WG;
wire[7:0] Tile_X3Y11_to_WH;
wire[11:0] Tile_X3Y11_to_WI;
wire[3:0] Tile_X3Y11_to_NA;
wire[3:0] Tile_X3Y11_to_NB;
wire[3:0] Tile_X3Y11_to_NC;
wire[3:0] Tile_X3Y11_to_ND;
wire[3:0] Tile_X3Y11_to_NF;
wire[7:0] Tile_X3Y11_to_NG;
wire[7:0] Tile_X3Y11_to_NH;
wire[11:0] Tile_X3Y11_to_NI;
wire[3:0] Tile_X3Y11_to_SA;
wire[3:0] Tile_X3Y11_to_SB;
wire[3:0] Tile_X3Y11_to_SC;
wire[3:0] Tile_X3Y11_to_SD;
wire[3:0] Tile_X3Y11_to_SF;
wire[7:0] Tile_X3Y11_to_SG;
wire[7:0] Tile_X3Y11_to_SH;
wire[11:0] Tile_X3Y11_to_SI;
wire[3:0] Tile_X4Y11_to_EA;
wire[3:0] Tile_X4Y11_to_EB;
wire[3:0] Tile_X4Y11_to_EC;
wire[3:0] Tile_X4Y11_to_ED;
wire[3:0] Tile_X4Y11_to_EF;
wire[7:0] Tile_X4Y11_to_EG;
wire[7:0] Tile_X4Y11_to_EH;
wire[11:0] Tile_X4Y11_to_EI;
wire[3:0] Tile_X4Y11_to_WA;
wire[3:0] Tile_X4Y11_to_WB;
wire[3:0] Tile_X4Y11_to_WC;
wire[3:0] Tile_X4Y11_to_WD;
wire[3:0] Tile_X4Y11_to_WF;
wire[7:0] Tile_X4Y11_to_WG;
wire[7:0] Tile_X4Y11_to_WH;
wire[11:0] Tile_X4Y11_to_WI;
wire[3:0] Tile_X4Y11_to_NA;
wire[3:0] Tile_X4Y11_to_NB;
wire[3:0] Tile_X4Y11_to_NC;
wire[3:0] Tile_X4Y11_to_ND;
wire[3:0] Tile_X4Y11_to_NF;
wire[7:0] Tile_X4Y11_to_NG;
wire[7:0] Tile_X4Y11_to_NH;
wire[11:0] Tile_X4Y11_to_NI;
wire[3:0] Tile_X4Y11_to_SA;
wire[3:0] Tile_X4Y11_to_SB;
wire[3:0] Tile_X4Y11_to_SC;
wire[3:0] Tile_X4Y11_to_SD;
wire[3:0] Tile_X4Y11_to_SF;
wire[7:0] Tile_X4Y11_to_SG;
wire[7:0] Tile_X4Y11_to_SH;
wire[11:0] Tile_X4Y11_to_SI;
wire[3:0] Tile_X5Y11_to_EA;
wire[3:0] Tile_X5Y11_to_EB;
wire[3:0] Tile_X5Y11_to_EC;
wire[3:0] Tile_X5Y11_to_ED;
wire[3:0] Tile_X5Y11_to_EF;
wire[7:0] Tile_X5Y11_to_EG;
wire[7:0] Tile_X5Y11_to_EH;
wire[11:0] Tile_X5Y11_to_EI;
wire[3:0] Tile_X5Y11_to_WA;
wire[3:0] Tile_X5Y11_to_WB;
wire[3:0] Tile_X5Y11_to_WC;
wire[3:0] Tile_X5Y11_to_WD;
wire[3:0] Tile_X5Y11_to_WF;
wire[7:0] Tile_X5Y11_to_WG;
wire[7:0] Tile_X5Y11_to_WH;
wire[11:0] Tile_X5Y11_to_WI;
wire[3:0] Tile_X5Y11_to_NA;
wire[3:0] Tile_X5Y11_to_NB;
wire[3:0] Tile_X5Y11_to_NC;
wire[3:0] Tile_X5Y11_to_ND;
wire[3:0] Tile_X5Y11_to_NF;
wire[7:0] Tile_X5Y11_to_NG;
wire[7:0] Tile_X5Y11_to_NH;
wire[11:0] Tile_X5Y11_to_NI;
wire[3:0] Tile_X5Y11_to_SA;
wire[3:0] Tile_X5Y11_to_SB;
wire[3:0] Tile_X5Y11_to_SC;
wire[3:0] Tile_X5Y11_to_SD;
wire[3:0] Tile_X5Y11_to_SF;
wire[7:0] Tile_X5Y11_to_SG;
wire[7:0] Tile_X5Y11_to_SH;
wire[11:0] Tile_X5Y11_to_SI;
wire[3:0] Tile_X6Y11_to_EA;
wire[3:0] Tile_X6Y11_to_EB;
wire[3:0] Tile_X6Y11_to_EC;
wire[3:0] Tile_X6Y11_to_ED;
wire[3:0] Tile_X6Y11_to_EF;
wire[7:0] Tile_X6Y11_to_EG;
wire[7:0] Tile_X6Y11_to_EH;
wire[11:0] Tile_X6Y11_to_EI;
wire[3:0] Tile_X6Y11_to_WA;
wire[3:0] Tile_X6Y11_to_WB;
wire[3:0] Tile_X6Y11_to_WC;
wire[3:0] Tile_X6Y11_to_WD;
wire[3:0] Tile_X6Y11_to_WF;
wire[7:0] Tile_X6Y11_to_WG;
wire[7:0] Tile_X6Y11_to_WH;
wire[11:0] Tile_X6Y11_to_WI;
wire[3:0] Tile_X6Y11_to_NA;
wire[3:0] Tile_X6Y11_to_NB;
wire[3:0] Tile_X6Y11_to_NC;
wire[3:0] Tile_X6Y11_to_ND;
wire[3:0] Tile_X6Y11_to_NF;
wire[7:0] Tile_X6Y11_to_NG;
wire[7:0] Tile_X6Y11_to_NH;
wire[11:0] Tile_X6Y11_to_NI;
wire[3:0] Tile_X6Y11_to_SA;
wire[3:0] Tile_X6Y11_to_SB;
wire[3:0] Tile_X6Y11_to_SC;
wire[3:0] Tile_X6Y11_to_SD;
wire[3:0] Tile_X6Y11_to_SF;
wire[7:0] Tile_X6Y11_to_SG;
wire[7:0] Tile_X6Y11_to_SH;
wire[11:0] Tile_X6Y11_to_SI;
wire[3:0] Tile_X7Y11_to_EA;
wire[3:0] Tile_X7Y11_to_EB;
wire[3:0] Tile_X7Y11_to_EC;
wire[3:0] Tile_X7Y11_to_ED;
wire[3:0] Tile_X7Y11_to_EF;
wire[7:0] Tile_X7Y11_to_EG;
wire[7:0] Tile_X7Y11_to_EH;
wire[11:0] Tile_X7Y11_to_EI;
wire[3:0] Tile_X7Y11_to_WA;
wire[3:0] Tile_X7Y11_to_WB;
wire[3:0] Tile_X7Y11_to_WC;
wire[3:0] Tile_X7Y11_to_WD;
wire[3:0] Tile_X7Y11_to_WF;
wire[7:0] Tile_X7Y11_to_WG;
wire[7:0] Tile_X7Y11_to_WH;
wire[11:0] Tile_X7Y11_to_WI;
wire[3:0] Tile_X7Y11_to_NA;
wire[3:0] Tile_X7Y11_to_NB;
wire[3:0] Tile_X7Y11_to_NC;
wire[3:0] Tile_X7Y11_to_ND;
wire[3:0] Tile_X7Y11_to_NF;
wire[7:0] Tile_X7Y11_to_NG;
wire[7:0] Tile_X7Y11_to_NH;
wire[11:0] Tile_X7Y11_to_NI;
wire[3:0] Tile_X7Y11_to_SA;
wire[3:0] Tile_X7Y11_to_SB;
wire[3:0] Tile_X7Y11_to_SC;
wire[3:0] Tile_X7Y11_to_SD;
wire[3:0] Tile_X7Y11_to_SF;
wire[7:0] Tile_X7Y11_to_SG;
wire[7:0] Tile_X7Y11_to_SH;
wire[11:0] Tile_X7Y11_to_SI;
wire[3:0] Tile_X8Y11_to_WA;
wire[3:0] Tile_X8Y11_to_WB;
wire[3:0] Tile_X8Y11_to_WC;
wire[3:0] Tile_X8Y11_to_WD;
wire[3:0] Tile_X8Y11_to_WF;
wire[7:0] Tile_X8Y11_to_WG;
wire[7:0] Tile_X8Y11_to_WH;
wire[11:0] Tile_X8Y11_to_WI;
wire[3:0] Tile_X8Y11_to_NA;
wire[3:0] Tile_X8Y11_to_NB;
wire[3:0] Tile_X8Y11_to_NC;
wire[3:0] Tile_X8Y11_to_ND;
wire[3:0] Tile_X8Y11_to_NF;
wire[7:0] Tile_X8Y11_to_NG;
wire[7:0] Tile_X8Y11_to_NH;
wire[11:0] Tile_X8Y11_to_NI;
wire[3:0] Tile_X8Y11_to_SA;
wire[3:0] Tile_X8Y11_to_SB;
wire[3:0] Tile_X8Y11_to_SC;
wire[3:0] Tile_X8Y11_to_SD;
wire[3:0] Tile_X8Y11_to_SF;
wire[7:0] Tile_X8Y11_to_SG;
wire[7:0] Tile_X8Y11_to_SH;
wire[11:0] Tile_X8Y11_to_SI;
wire[1:0] Tile_X9Y11_to_EA_1s;
wire[1:0] Tile_X9Y11_to_EB_1s;
wire[1:0] Tile_X9Y11_to_EC_1s;
wire[1:0] Tile_X9Y11_to_ED_1s;
wire[1:0] Tile_X9Y11_to_EF_1s;
wire[1:0] Tile_X9Y11_to_EG_1s;
wire[1:0] Tile_X9Y11_to_EH_1s;
wire[1:0] Tile_X9Y11_to_EI_1s;
wire[1:0] Tile_X9Y11_to_WA_1s;
wire[1:0] Tile_X9Y11_to_WB_1s;
wire[1:0] Tile_X9Y11_to_WC_1s;
wire[1:0] Tile_X9Y11_to_WD_1s;
wire[1:0] Tile_X9Y11_to_WF_1s;
wire[1:0] Tile_X9Y11_to_WG_1s;
wire[1:0] Tile_X9Y11_to_WH_1s;
wire[1:0] Tile_X9Y11_to_WI_1s;
wire[1:0] Tile_X9Y11_to_NA_1s;
wire[1:0] Tile_X9Y11_to_NB_1s;
wire[1:0] Tile_X9Y11_to_NC_1s;
wire[1:0] Tile_X9Y11_to_ND_1s;
wire[1:0] Tile_X9Y11_to_NF_1s;
wire[1:0] Tile_X9Y11_to_NG_1s;
wire[1:0] Tile_X9Y11_to_NH_1s;
wire[1:0] Tile_X9Y11_to_NI_1s;
wire[1:0] Tile_X9Y11_to_SA_1s;
wire[1:0] Tile_X9Y11_to_SB_1s;
wire[1:0] Tile_X9Y11_to_SC_1s;
wire[1:0] Tile_X9Y11_to_SD_1s;
wire[1:0] Tile_X9Y11_to_SF_1s;
wire[1:0] Tile_X9Y11_to_SG_1s;
wire[1:0] Tile_X9Y11_to_SH_1s;
wire[1:0] Tile_X9Y11_to_SI_1s;
wire[1:0] Tile_X10Y11_to_WA_1s;
wire[1:0] Tile_X10Y11_to_WB_1s;
wire[1:0] Tile_X10Y11_to_WC_1s;
wire[1:0] Tile_X10Y11_to_WD_1s;
wire[1:0] Tile_X10Y11_to_WF_1s;
wire[1:0] Tile_X10Y11_to_WG_1s;
wire[1:0] Tile_X10Y11_to_WH_1s;
wire[1:0] Tile_X10Y11_to_WI_1s;
wire[3:0] Tile_X0Y12_to_EA;
wire[3:0] Tile_X0Y12_to_EB;
wire[3:0] Tile_X0Y12_to_EC;
wire[3:0] Tile_X0Y12_to_ED;
wire[3:0] Tile_X0Y12_to_EF;
wire[7:0] Tile_X0Y12_to_EG;
wire[7:0] Tile_X0Y12_to_EH;
wire[11:0] Tile_X0Y12_to_EI;
wire[3:0] Tile_X0Y12_to_NA;
wire[3:0] Tile_X0Y12_to_NB;
wire[3:0] Tile_X0Y12_to_NC;
wire[3:0] Tile_X0Y12_to_ND;
wire[3:0] Tile_X0Y12_to_NF;
wire[7:0] Tile_X0Y12_to_NG;
wire[7:0] Tile_X0Y12_to_NH;
wire[11:0] Tile_X0Y12_to_NI;
wire[3:0] Tile_X0Y12_to_SA;
wire[3:0] Tile_X0Y12_to_SB;
wire[3:0] Tile_X0Y12_to_SC;
wire[3:0] Tile_X0Y12_to_SD;
wire[3:0] Tile_X0Y12_to_SF;
wire[7:0] Tile_X0Y12_to_SG;
wire[7:0] Tile_X0Y12_to_SH;
wire[11:0] Tile_X0Y12_to_SI;
wire[3:0] Tile_X1Y12_to_EA;
wire[3:0] Tile_X1Y12_to_EB;
wire[3:0] Tile_X1Y12_to_EC;
wire[3:0] Tile_X1Y12_to_ED;
wire[3:0] Tile_X1Y12_to_EF;
wire[7:0] Tile_X1Y12_to_EG;
wire[7:0] Tile_X1Y12_to_EH;
wire[11:0] Tile_X1Y12_to_EI;
wire[3:0] Tile_X1Y12_to_WA;
wire[3:0] Tile_X1Y12_to_WB;
wire[3:0] Tile_X1Y12_to_WC;
wire[3:0] Tile_X1Y12_to_WD;
wire[3:0] Tile_X1Y12_to_WF;
wire[7:0] Tile_X1Y12_to_WG;
wire[7:0] Tile_X1Y12_to_WH;
wire[11:0] Tile_X1Y12_to_WI;
wire[3:0] Tile_X1Y12_to_NA;
wire[3:0] Tile_X1Y12_to_NB;
wire[3:0] Tile_X1Y12_to_NC;
wire[3:0] Tile_X1Y12_to_ND;
wire[3:0] Tile_X1Y12_to_NF;
wire[7:0] Tile_X1Y12_to_NG;
wire[7:0] Tile_X1Y12_to_NH;
wire[11:0] Tile_X1Y12_to_NI;
wire[3:0] Tile_X1Y12_to_SA;
wire[3:0] Tile_X1Y12_to_SB;
wire[3:0] Tile_X1Y12_to_SC;
wire[3:0] Tile_X1Y12_to_SD;
wire[3:0] Tile_X1Y12_to_SF;
wire[7:0] Tile_X1Y12_to_SG;
wire[7:0] Tile_X1Y12_to_SH;
wire[11:0] Tile_X1Y12_to_SI;
wire[3:0] Tile_X2Y12_to_EA;
wire[3:0] Tile_X2Y12_to_EB;
wire[3:0] Tile_X2Y12_to_EC;
wire[3:0] Tile_X2Y12_to_ED;
wire[3:0] Tile_X2Y12_to_EF;
wire[7:0] Tile_X2Y12_to_EG;
wire[7:0] Tile_X2Y12_to_EH;
wire[11:0] Tile_X2Y12_to_EI;
wire[3:0] Tile_X2Y12_to_WA;
wire[3:0] Tile_X2Y12_to_WB;
wire[3:0] Tile_X2Y12_to_WC;
wire[3:0] Tile_X2Y12_to_WD;
wire[3:0] Tile_X2Y12_to_WF;
wire[7:0] Tile_X2Y12_to_WG;
wire[7:0] Tile_X2Y12_to_WH;
wire[11:0] Tile_X2Y12_to_WI;
wire[3:0] Tile_X2Y12_to_NA;
wire[3:0] Tile_X2Y12_to_NB;
wire[3:0] Tile_X2Y12_to_NC;
wire[3:0] Tile_X2Y12_to_ND;
wire[3:0] Tile_X2Y12_to_NF;
wire[7:0] Tile_X2Y12_to_NG;
wire[7:0] Tile_X2Y12_to_NH;
wire[11:0] Tile_X2Y12_to_NI;
wire[3:0] Tile_X2Y12_to_SA;
wire[3:0] Tile_X2Y12_to_SB;
wire[3:0] Tile_X2Y12_to_SC;
wire[3:0] Tile_X2Y12_to_SD;
wire[3:0] Tile_X2Y12_to_SF;
wire[7:0] Tile_X2Y12_to_SG;
wire[7:0] Tile_X2Y12_to_SH;
wire[11:0] Tile_X2Y12_to_SI;
wire[3:0] Tile_X3Y12_to_EA;
wire[3:0] Tile_X3Y12_to_EB;
wire[3:0] Tile_X3Y12_to_EC;
wire[3:0] Tile_X3Y12_to_ED;
wire[3:0] Tile_X3Y12_to_EF;
wire[7:0] Tile_X3Y12_to_EG;
wire[7:0] Tile_X3Y12_to_EH;
wire[11:0] Tile_X3Y12_to_EI;
wire[3:0] Tile_X3Y12_to_WA;
wire[3:0] Tile_X3Y12_to_WB;
wire[3:0] Tile_X3Y12_to_WC;
wire[3:0] Tile_X3Y12_to_WD;
wire[3:0] Tile_X3Y12_to_WF;
wire[7:0] Tile_X3Y12_to_WG;
wire[7:0] Tile_X3Y12_to_WH;
wire[11:0] Tile_X3Y12_to_WI;
wire[3:0] Tile_X3Y12_to_NA;
wire[3:0] Tile_X3Y12_to_NB;
wire[3:0] Tile_X3Y12_to_NC;
wire[3:0] Tile_X3Y12_to_ND;
wire[3:0] Tile_X3Y12_to_NF;
wire[7:0] Tile_X3Y12_to_NG;
wire[7:0] Tile_X3Y12_to_NH;
wire[11:0] Tile_X3Y12_to_NI;
wire[3:0] Tile_X3Y12_to_SA;
wire[3:0] Tile_X3Y12_to_SB;
wire[3:0] Tile_X3Y12_to_SC;
wire[3:0] Tile_X3Y12_to_SD;
wire[3:0] Tile_X3Y12_to_SF;
wire[7:0] Tile_X3Y12_to_SG;
wire[7:0] Tile_X3Y12_to_SH;
wire[11:0] Tile_X3Y12_to_SI;
wire[3:0] Tile_X4Y12_to_EA;
wire[3:0] Tile_X4Y12_to_EB;
wire[3:0] Tile_X4Y12_to_EC;
wire[3:0] Tile_X4Y12_to_ED;
wire[3:0] Tile_X4Y12_to_EF;
wire[7:0] Tile_X4Y12_to_EG;
wire[7:0] Tile_X4Y12_to_EH;
wire[11:0] Tile_X4Y12_to_EI;
wire[3:0] Tile_X4Y12_to_WA;
wire[3:0] Tile_X4Y12_to_WB;
wire[3:0] Tile_X4Y12_to_WC;
wire[3:0] Tile_X4Y12_to_WD;
wire[3:0] Tile_X4Y12_to_WF;
wire[7:0] Tile_X4Y12_to_WG;
wire[7:0] Tile_X4Y12_to_WH;
wire[11:0] Tile_X4Y12_to_WI;
wire[3:0] Tile_X4Y12_to_NA;
wire[3:0] Tile_X4Y12_to_NB;
wire[3:0] Tile_X4Y12_to_NC;
wire[3:0] Tile_X4Y12_to_ND;
wire[3:0] Tile_X4Y12_to_NF;
wire[7:0] Tile_X4Y12_to_NG;
wire[7:0] Tile_X4Y12_to_NH;
wire[11:0] Tile_X4Y12_to_NI;
wire[3:0] Tile_X4Y12_to_SA;
wire[3:0] Tile_X4Y12_to_SB;
wire[3:0] Tile_X4Y12_to_SC;
wire[3:0] Tile_X4Y12_to_SD;
wire[3:0] Tile_X4Y12_to_SF;
wire[7:0] Tile_X4Y12_to_SG;
wire[7:0] Tile_X4Y12_to_SH;
wire[11:0] Tile_X4Y12_to_SI;
wire[3:0] Tile_X5Y12_to_EA;
wire[3:0] Tile_X5Y12_to_EB;
wire[3:0] Tile_X5Y12_to_EC;
wire[3:0] Tile_X5Y12_to_ED;
wire[3:0] Tile_X5Y12_to_EF;
wire[7:0] Tile_X5Y12_to_EG;
wire[7:0] Tile_X5Y12_to_EH;
wire[11:0] Tile_X5Y12_to_EI;
wire[3:0] Tile_X5Y12_to_WA;
wire[3:0] Tile_X5Y12_to_WB;
wire[3:0] Tile_X5Y12_to_WC;
wire[3:0] Tile_X5Y12_to_WD;
wire[3:0] Tile_X5Y12_to_WF;
wire[7:0] Tile_X5Y12_to_WG;
wire[7:0] Tile_X5Y12_to_WH;
wire[11:0] Tile_X5Y12_to_WI;
wire[3:0] Tile_X5Y12_to_NA;
wire[3:0] Tile_X5Y12_to_NB;
wire[3:0] Tile_X5Y12_to_NC;
wire[3:0] Tile_X5Y12_to_ND;
wire[3:0] Tile_X5Y12_to_NF;
wire[7:0] Tile_X5Y12_to_NG;
wire[7:0] Tile_X5Y12_to_NH;
wire[11:0] Tile_X5Y12_to_NI;
wire[3:0] Tile_X5Y12_to_SA;
wire[3:0] Tile_X5Y12_to_SB;
wire[3:0] Tile_X5Y12_to_SC;
wire[3:0] Tile_X5Y12_to_SD;
wire[3:0] Tile_X5Y12_to_SF;
wire[7:0] Tile_X5Y12_to_SG;
wire[7:0] Tile_X5Y12_to_SH;
wire[11:0] Tile_X5Y12_to_SI;
wire[3:0] Tile_X6Y12_to_EA;
wire[3:0] Tile_X6Y12_to_EB;
wire[3:0] Tile_X6Y12_to_EC;
wire[3:0] Tile_X6Y12_to_ED;
wire[3:0] Tile_X6Y12_to_EF;
wire[7:0] Tile_X6Y12_to_EG;
wire[7:0] Tile_X6Y12_to_EH;
wire[11:0] Tile_X6Y12_to_EI;
wire[3:0] Tile_X6Y12_to_WA;
wire[3:0] Tile_X6Y12_to_WB;
wire[3:0] Tile_X6Y12_to_WC;
wire[3:0] Tile_X6Y12_to_WD;
wire[3:0] Tile_X6Y12_to_WF;
wire[7:0] Tile_X6Y12_to_WG;
wire[7:0] Tile_X6Y12_to_WH;
wire[11:0] Tile_X6Y12_to_WI;
wire[3:0] Tile_X6Y12_to_NA;
wire[3:0] Tile_X6Y12_to_NB;
wire[3:0] Tile_X6Y12_to_NC;
wire[3:0] Tile_X6Y12_to_ND;
wire[3:0] Tile_X6Y12_to_NF;
wire[7:0] Tile_X6Y12_to_NG;
wire[7:0] Tile_X6Y12_to_NH;
wire[11:0] Tile_X6Y12_to_NI;
wire[3:0] Tile_X6Y12_to_SA;
wire[3:0] Tile_X6Y12_to_SB;
wire[3:0] Tile_X6Y12_to_SC;
wire[3:0] Tile_X6Y12_to_SD;
wire[3:0] Tile_X6Y12_to_SF;
wire[7:0] Tile_X6Y12_to_SG;
wire[7:0] Tile_X6Y12_to_SH;
wire[11:0] Tile_X6Y12_to_SI;
wire[3:0] Tile_X7Y12_to_EA;
wire[3:0] Tile_X7Y12_to_EB;
wire[3:0] Tile_X7Y12_to_EC;
wire[3:0] Tile_X7Y12_to_ED;
wire[3:0] Tile_X7Y12_to_EF;
wire[7:0] Tile_X7Y12_to_EG;
wire[7:0] Tile_X7Y12_to_EH;
wire[11:0] Tile_X7Y12_to_EI;
wire[3:0] Tile_X7Y12_to_WA;
wire[3:0] Tile_X7Y12_to_WB;
wire[3:0] Tile_X7Y12_to_WC;
wire[3:0] Tile_X7Y12_to_WD;
wire[3:0] Tile_X7Y12_to_WF;
wire[7:0] Tile_X7Y12_to_WG;
wire[7:0] Tile_X7Y12_to_WH;
wire[11:0] Tile_X7Y12_to_WI;
wire[3:0] Tile_X7Y12_to_NA;
wire[3:0] Tile_X7Y12_to_NB;
wire[3:0] Tile_X7Y12_to_NC;
wire[3:0] Tile_X7Y12_to_ND;
wire[3:0] Tile_X7Y12_to_NF;
wire[7:0] Tile_X7Y12_to_NG;
wire[7:0] Tile_X7Y12_to_NH;
wire[11:0] Tile_X7Y12_to_NI;
wire[3:0] Tile_X7Y12_to_SA;
wire[3:0] Tile_X7Y12_to_SB;
wire[3:0] Tile_X7Y12_to_SC;
wire[3:0] Tile_X7Y12_to_SD;
wire[3:0] Tile_X7Y12_to_SF;
wire[7:0] Tile_X7Y12_to_SG;
wire[7:0] Tile_X7Y12_to_SH;
wire[11:0] Tile_X7Y12_to_SI;
wire[3:0] Tile_X8Y12_to_WA;
wire[3:0] Tile_X8Y12_to_WB;
wire[3:0] Tile_X8Y12_to_WC;
wire[3:0] Tile_X8Y12_to_WD;
wire[3:0] Tile_X8Y12_to_WF;
wire[7:0] Tile_X8Y12_to_WG;
wire[7:0] Tile_X8Y12_to_WH;
wire[11:0] Tile_X8Y12_to_WI;
wire[3:0] Tile_X8Y12_to_NA;
wire[3:0] Tile_X8Y12_to_NB;
wire[3:0] Tile_X8Y12_to_NC;
wire[3:0] Tile_X8Y12_to_ND;
wire[3:0] Tile_X8Y12_to_NF;
wire[7:0] Tile_X8Y12_to_NG;
wire[7:0] Tile_X8Y12_to_NH;
wire[11:0] Tile_X8Y12_to_NI;
wire[3:0] Tile_X8Y12_to_SA;
wire[3:0] Tile_X8Y12_to_SB;
wire[3:0] Tile_X8Y12_to_SC;
wire[3:0] Tile_X8Y12_to_SD;
wire[3:0] Tile_X8Y12_to_SF;
wire[7:0] Tile_X8Y12_to_SG;
wire[7:0] Tile_X8Y12_to_SH;
wire[11:0] Tile_X8Y12_to_SI;
wire[1:0] Tile_X9Y12_to_EA_1s;
wire[1:0] Tile_X9Y12_to_EB_1s;
wire[1:0] Tile_X9Y12_to_EC_1s;
wire[1:0] Tile_X9Y12_to_ED_1s;
wire[1:0] Tile_X9Y12_to_EF_1s;
wire[1:0] Tile_X9Y12_to_EG_1s;
wire[1:0] Tile_X9Y12_to_EH_1s;
wire[1:0] Tile_X9Y12_to_EI_1s;
wire[1:0] Tile_X9Y12_to_WA_1s;
wire[1:0] Tile_X9Y12_to_WB_1s;
wire[1:0] Tile_X9Y12_to_WC_1s;
wire[1:0] Tile_X9Y12_to_WD_1s;
wire[1:0] Tile_X9Y12_to_WF_1s;
wire[1:0] Tile_X9Y12_to_WG_1s;
wire[1:0] Tile_X9Y12_to_WH_1s;
wire[1:0] Tile_X9Y12_to_WI_1s;
wire[1:0] Tile_X9Y12_to_NA_1s;
wire[1:0] Tile_X9Y12_to_NB_1s;
wire[1:0] Tile_X9Y12_to_NC_1s;
wire[1:0] Tile_X9Y12_to_ND_1s;
wire[1:0] Tile_X9Y12_to_NF_1s;
wire[1:0] Tile_X9Y12_to_NG_1s;
wire[1:0] Tile_X9Y12_to_NH_1s;
wire[1:0] Tile_X9Y12_to_NI_1s;
wire[1:0] Tile_X9Y12_to_SA_1s;
wire[1:0] Tile_X9Y12_to_SB_1s;
wire[1:0] Tile_X9Y12_to_SC_1s;
wire[1:0] Tile_X9Y12_to_SD_1s;
wire[1:0] Tile_X9Y12_to_SF_1s;
wire[1:0] Tile_X9Y12_to_SG_1s;
wire[1:0] Tile_X9Y12_to_SH_1s;
wire[1:0] Tile_X9Y12_to_SI_1s;
wire[1:0] Tile_X10Y12_to_WA_1s;
wire[1:0] Tile_X10Y12_to_WB_1s;
wire[1:0] Tile_X10Y12_to_WC_1s;
wire[1:0] Tile_X10Y12_to_WD_1s;
wire[1:0] Tile_X10Y12_to_WF_1s;
wire[1:0] Tile_X10Y12_to_WG_1s;
wire[1:0] Tile_X10Y12_to_WH_1s;
wire[1:0] Tile_X10Y12_to_WI_1s;
wire[3:0] Tile_X0Y13_to_EA;
wire[3:0] Tile_X0Y13_to_EB;
wire[3:0] Tile_X0Y13_to_EC;
wire[3:0] Tile_X0Y13_to_ED;
wire[3:0] Tile_X0Y13_to_EF;
wire[7:0] Tile_X0Y13_to_EG;
wire[7:0] Tile_X0Y13_to_EH;
wire[11:0] Tile_X0Y13_to_EI;
wire[3:0] Tile_X0Y13_to_NA;
wire[3:0] Tile_X0Y13_to_NB;
wire[3:0] Tile_X0Y13_to_NC;
wire[3:0] Tile_X0Y13_to_ND;
wire[3:0] Tile_X0Y13_to_NF;
wire[7:0] Tile_X0Y13_to_NG;
wire[7:0] Tile_X0Y13_to_NH;
wire[11:0] Tile_X0Y13_to_NI;
wire[3:0] Tile_X0Y13_to_SA;
wire[3:0] Tile_X0Y13_to_SB;
wire[3:0] Tile_X0Y13_to_SC;
wire[3:0] Tile_X0Y13_to_SD;
wire[3:0] Tile_X0Y13_to_SF;
wire[7:0] Tile_X0Y13_to_SG;
wire[7:0] Tile_X0Y13_to_SH;
wire[11:0] Tile_X0Y13_to_SI;
wire[3:0] Tile_X1Y13_to_EA;
wire[3:0] Tile_X1Y13_to_EB;
wire[3:0] Tile_X1Y13_to_EC;
wire[3:0] Tile_X1Y13_to_ED;
wire[3:0] Tile_X1Y13_to_EF;
wire[7:0] Tile_X1Y13_to_EG;
wire[7:0] Tile_X1Y13_to_EH;
wire[11:0] Tile_X1Y13_to_EI;
wire[3:0] Tile_X1Y13_to_WA;
wire[3:0] Tile_X1Y13_to_WB;
wire[3:0] Tile_X1Y13_to_WC;
wire[3:0] Tile_X1Y13_to_WD;
wire[3:0] Tile_X1Y13_to_WF;
wire[7:0] Tile_X1Y13_to_WG;
wire[7:0] Tile_X1Y13_to_WH;
wire[11:0] Tile_X1Y13_to_WI;
wire[3:0] Tile_X1Y13_to_NA;
wire[3:0] Tile_X1Y13_to_NB;
wire[3:0] Tile_X1Y13_to_NC;
wire[3:0] Tile_X1Y13_to_ND;
wire[3:0] Tile_X1Y13_to_NF;
wire[7:0] Tile_X1Y13_to_NG;
wire[7:0] Tile_X1Y13_to_NH;
wire[11:0] Tile_X1Y13_to_NI;
wire[3:0] Tile_X1Y13_to_SA;
wire[3:0] Tile_X1Y13_to_SB;
wire[3:0] Tile_X1Y13_to_SC;
wire[3:0] Tile_X1Y13_to_SD;
wire[3:0] Tile_X1Y13_to_SF;
wire[7:0] Tile_X1Y13_to_SG;
wire[7:0] Tile_X1Y13_to_SH;
wire[11:0] Tile_X1Y13_to_SI;
wire[3:0] Tile_X2Y13_to_EA;
wire[3:0] Tile_X2Y13_to_EB;
wire[3:0] Tile_X2Y13_to_EC;
wire[3:0] Tile_X2Y13_to_ED;
wire[3:0] Tile_X2Y13_to_EF;
wire[7:0] Tile_X2Y13_to_EG;
wire[7:0] Tile_X2Y13_to_EH;
wire[11:0] Tile_X2Y13_to_EI;
wire[3:0] Tile_X2Y13_to_WA;
wire[3:0] Tile_X2Y13_to_WB;
wire[3:0] Tile_X2Y13_to_WC;
wire[3:0] Tile_X2Y13_to_WD;
wire[3:0] Tile_X2Y13_to_WF;
wire[7:0] Tile_X2Y13_to_WG;
wire[7:0] Tile_X2Y13_to_WH;
wire[11:0] Tile_X2Y13_to_WI;
wire[3:0] Tile_X2Y13_to_NA;
wire[3:0] Tile_X2Y13_to_NB;
wire[3:0] Tile_X2Y13_to_NC;
wire[3:0] Tile_X2Y13_to_ND;
wire[3:0] Tile_X2Y13_to_NF;
wire[7:0] Tile_X2Y13_to_NG;
wire[7:0] Tile_X2Y13_to_NH;
wire[11:0] Tile_X2Y13_to_NI;
wire[3:0] Tile_X2Y13_to_SA;
wire[3:0] Tile_X2Y13_to_SB;
wire[3:0] Tile_X2Y13_to_SC;
wire[3:0] Tile_X2Y13_to_SD;
wire[3:0] Tile_X2Y13_to_SF;
wire[7:0] Tile_X2Y13_to_SG;
wire[7:0] Tile_X2Y13_to_SH;
wire[11:0] Tile_X2Y13_to_SI;
wire[3:0] Tile_X3Y13_to_EA;
wire[3:0] Tile_X3Y13_to_EB;
wire[3:0] Tile_X3Y13_to_EC;
wire[3:0] Tile_X3Y13_to_ED;
wire[3:0] Tile_X3Y13_to_EF;
wire[7:0] Tile_X3Y13_to_EG;
wire[7:0] Tile_X3Y13_to_EH;
wire[11:0] Tile_X3Y13_to_EI;
wire[3:0] Tile_X3Y13_to_WA;
wire[3:0] Tile_X3Y13_to_WB;
wire[3:0] Tile_X3Y13_to_WC;
wire[3:0] Tile_X3Y13_to_WD;
wire[3:0] Tile_X3Y13_to_WF;
wire[7:0] Tile_X3Y13_to_WG;
wire[7:0] Tile_X3Y13_to_WH;
wire[11:0] Tile_X3Y13_to_WI;
wire[3:0] Tile_X3Y13_to_NA;
wire[3:0] Tile_X3Y13_to_NB;
wire[3:0] Tile_X3Y13_to_NC;
wire[3:0] Tile_X3Y13_to_ND;
wire[3:0] Tile_X3Y13_to_NF;
wire[7:0] Tile_X3Y13_to_NG;
wire[7:0] Tile_X3Y13_to_NH;
wire[11:0] Tile_X3Y13_to_NI;
wire[3:0] Tile_X3Y13_to_SA;
wire[3:0] Tile_X3Y13_to_SB;
wire[3:0] Tile_X3Y13_to_SC;
wire[3:0] Tile_X3Y13_to_SD;
wire[3:0] Tile_X3Y13_to_SF;
wire[7:0] Tile_X3Y13_to_SG;
wire[7:0] Tile_X3Y13_to_SH;
wire[11:0] Tile_X3Y13_to_SI;
wire[3:0] Tile_X4Y13_to_EA;
wire[3:0] Tile_X4Y13_to_EB;
wire[3:0] Tile_X4Y13_to_EC;
wire[3:0] Tile_X4Y13_to_ED;
wire[3:0] Tile_X4Y13_to_EF;
wire[7:0] Tile_X4Y13_to_EG;
wire[7:0] Tile_X4Y13_to_EH;
wire[11:0] Tile_X4Y13_to_EI;
wire[3:0] Tile_X4Y13_to_WA;
wire[3:0] Tile_X4Y13_to_WB;
wire[3:0] Tile_X4Y13_to_WC;
wire[3:0] Tile_X4Y13_to_WD;
wire[3:0] Tile_X4Y13_to_WF;
wire[7:0] Tile_X4Y13_to_WG;
wire[7:0] Tile_X4Y13_to_WH;
wire[11:0] Tile_X4Y13_to_WI;
wire[3:0] Tile_X4Y13_to_NA;
wire[3:0] Tile_X4Y13_to_NB;
wire[3:0] Tile_X4Y13_to_NC;
wire[3:0] Tile_X4Y13_to_ND;
wire[3:0] Tile_X4Y13_to_NF;
wire[7:0] Tile_X4Y13_to_NG;
wire[7:0] Tile_X4Y13_to_NH;
wire[11:0] Tile_X4Y13_to_NI;
wire[3:0] Tile_X4Y13_to_SA;
wire[3:0] Tile_X4Y13_to_SB;
wire[3:0] Tile_X4Y13_to_SC;
wire[3:0] Tile_X4Y13_to_SD;
wire[3:0] Tile_X4Y13_to_SF;
wire[7:0] Tile_X4Y13_to_SG;
wire[7:0] Tile_X4Y13_to_SH;
wire[11:0] Tile_X4Y13_to_SI;
wire[3:0] Tile_X5Y13_to_EA;
wire[3:0] Tile_X5Y13_to_EB;
wire[3:0] Tile_X5Y13_to_EC;
wire[3:0] Tile_X5Y13_to_ED;
wire[3:0] Tile_X5Y13_to_EF;
wire[7:0] Tile_X5Y13_to_EG;
wire[7:0] Tile_X5Y13_to_EH;
wire[11:0] Tile_X5Y13_to_EI;
wire[3:0] Tile_X5Y13_to_WA;
wire[3:0] Tile_X5Y13_to_WB;
wire[3:0] Tile_X5Y13_to_WC;
wire[3:0] Tile_X5Y13_to_WD;
wire[3:0] Tile_X5Y13_to_WF;
wire[7:0] Tile_X5Y13_to_WG;
wire[7:0] Tile_X5Y13_to_WH;
wire[11:0] Tile_X5Y13_to_WI;
wire[3:0] Tile_X5Y13_to_NA;
wire[3:0] Tile_X5Y13_to_NB;
wire[3:0] Tile_X5Y13_to_NC;
wire[3:0] Tile_X5Y13_to_ND;
wire[3:0] Tile_X5Y13_to_NF;
wire[7:0] Tile_X5Y13_to_NG;
wire[7:0] Tile_X5Y13_to_NH;
wire[11:0] Tile_X5Y13_to_NI;
wire[3:0] Tile_X5Y13_to_SA;
wire[3:0] Tile_X5Y13_to_SB;
wire[3:0] Tile_X5Y13_to_SC;
wire[3:0] Tile_X5Y13_to_SD;
wire[3:0] Tile_X5Y13_to_SF;
wire[7:0] Tile_X5Y13_to_SG;
wire[7:0] Tile_X5Y13_to_SH;
wire[11:0] Tile_X5Y13_to_SI;
wire[3:0] Tile_X6Y13_to_EA;
wire[3:0] Tile_X6Y13_to_EB;
wire[3:0] Tile_X6Y13_to_EC;
wire[3:0] Tile_X6Y13_to_ED;
wire[3:0] Tile_X6Y13_to_EF;
wire[7:0] Tile_X6Y13_to_EG;
wire[7:0] Tile_X6Y13_to_EH;
wire[11:0] Tile_X6Y13_to_EI;
wire[3:0] Tile_X6Y13_to_WA;
wire[3:0] Tile_X6Y13_to_WB;
wire[3:0] Tile_X6Y13_to_WC;
wire[3:0] Tile_X6Y13_to_WD;
wire[3:0] Tile_X6Y13_to_WF;
wire[7:0] Tile_X6Y13_to_WG;
wire[7:0] Tile_X6Y13_to_WH;
wire[11:0] Tile_X6Y13_to_WI;
wire[3:0] Tile_X6Y13_to_NA;
wire[3:0] Tile_X6Y13_to_NB;
wire[3:0] Tile_X6Y13_to_NC;
wire[3:0] Tile_X6Y13_to_ND;
wire[3:0] Tile_X6Y13_to_NF;
wire[7:0] Tile_X6Y13_to_NG;
wire[7:0] Tile_X6Y13_to_NH;
wire[11:0] Tile_X6Y13_to_NI;
wire[3:0] Tile_X6Y13_to_SA;
wire[3:0] Tile_X6Y13_to_SB;
wire[3:0] Tile_X6Y13_to_SC;
wire[3:0] Tile_X6Y13_to_SD;
wire[3:0] Tile_X6Y13_to_SF;
wire[7:0] Tile_X6Y13_to_SG;
wire[7:0] Tile_X6Y13_to_SH;
wire[11:0] Tile_X6Y13_to_SI;
wire[3:0] Tile_X7Y13_to_EA;
wire[3:0] Tile_X7Y13_to_EB;
wire[3:0] Tile_X7Y13_to_EC;
wire[3:0] Tile_X7Y13_to_ED;
wire[3:0] Tile_X7Y13_to_EF;
wire[7:0] Tile_X7Y13_to_EG;
wire[7:0] Tile_X7Y13_to_EH;
wire[11:0] Tile_X7Y13_to_EI;
wire[3:0] Tile_X7Y13_to_WA;
wire[3:0] Tile_X7Y13_to_WB;
wire[3:0] Tile_X7Y13_to_WC;
wire[3:0] Tile_X7Y13_to_WD;
wire[3:0] Tile_X7Y13_to_WF;
wire[7:0] Tile_X7Y13_to_WG;
wire[7:0] Tile_X7Y13_to_WH;
wire[11:0] Tile_X7Y13_to_WI;
wire[3:0] Tile_X7Y13_to_NA;
wire[3:0] Tile_X7Y13_to_NB;
wire[3:0] Tile_X7Y13_to_NC;
wire[3:0] Tile_X7Y13_to_ND;
wire[3:0] Tile_X7Y13_to_NF;
wire[7:0] Tile_X7Y13_to_NG;
wire[7:0] Tile_X7Y13_to_NH;
wire[11:0] Tile_X7Y13_to_NI;
wire[3:0] Tile_X7Y13_to_SA;
wire[3:0] Tile_X7Y13_to_SB;
wire[3:0] Tile_X7Y13_to_SC;
wire[3:0] Tile_X7Y13_to_SD;
wire[3:0] Tile_X7Y13_to_SF;
wire[7:0] Tile_X7Y13_to_SG;
wire[7:0] Tile_X7Y13_to_SH;
wire[11:0] Tile_X7Y13_to_SI;
wire[3:0] Tile_X8Y13_to_WA;
wire[3:0] Tile_X8Y13_to_WB;
wire[3:0] Tile_X8Y13_to_WC;
wire[3:0] Tile_X8Y13_to_WD;
wire[3:0] Tile_X8Y13_to_WF;
wire[7:0] Tile_X8Y13_to_WG;
wire[7:0] Tile_X8Y13_to_WH;
wire[11:0] Tile_X8Y13_to_WI;
wire[3:0] Tile_X8Y13_to_NA;
wire[3:0] Tile_X8Y13_to_NB;
wire[3:0] Tile_X8Y13_to_NC;
wire[3:0] Tile_X8Y13_to_ND;
wire[3:0] Tile_X8Y13_to_NF;
wire[7:0] Tile_X8Y13_to_NG;
wire[7:0] Tile_X8Y13_to_NH;
wire[11:0] Tile_X8Y13_to_NI;
wire[3:0] Tile_X8Y13_to_SA;
wire[3:0] Tile_X8Y13_to_SB;
wire[3:0] Tile_X8Y13_to_SC;
wire[3:0] Tile_X8Y13_to_SD;
wire[3:0] Tile_X8Y13_to_SF;
wire[7:0] Tile_X8Y13_to_SG;
wire[7:0] Tile_X8Y13_to_SH;
wire[11:0] Tile_X8Y13_to_SI;
wire[1:0] Tile_X9Y13_to_EA_1s;
wire[1:0] Tile_X9Y13_to_EB_1s;
wire[1:0] Tile_X9Y13_to_EC_1s;
wire[1:0] Tile_X9Y13_to_ED_1s;
wire[1:0] Tile_X9Y13_to_EF_1s;
wire[1:0] Tile_X9Y13_to_EG_1s;
wire[1:0] Tile_X9Y13_to_EH_1s;
wire[1:0] Tile_X9Y13_to_EI_1s;
wire[1:0] Tile_X9Y13_to_WA_1s;
wire[1:0] Tile_X9Y13_to_WB_1s;
wire[1:0] Tile_X9Y13_to_WC_1s;
wire[1:0] Tile_X9Y13_to_WD_1s;
wire[1:0] Tile_X9Y13_to_WF_1s;
wire[1:0] Tile_X9Y13_to_WG_1s;
wire[1:0] Tile_X9Y13_to_WH_1s;
wire[1:0] Tile_X9Y13_to_WI_1s;
wire[1:0] Tile_X9Y13_to_NA_1s;
wire[1:0] Tile_X9Y13_to_NB_1s;
wire[1:0] Tile_X9Y13_to_NC_1s;
wire[1:0] Tile_X9Y13_to_ND_1s;
wire[1:0] Tile_X9Y13_to_NF_1s;
wire[1:0] Tile_X9Y13_to_NG_1s;
wire[1:0] Tile_X9Y13_to_NH_1s;
wire[1:0] Tile_X9Y13_to_NI_1s;
wire[1:0] Tile_X9Y13_to_SA_1s;
wire[1:0] Tile_X9Y13_to_SB_1s;
wire[1:0] Tile_X9Y13_to_SC_1s;
wire[1:0] Tile_X9Y13_to_SD_1s;
wire[1:0] Tile_X9Y13_to_SF_1s;
wire[1:0] Tile_X9Y13_to_SG_1s;
wire[1:0] Tile_X9Y13_to_SH_1s;
wire[1:0] Tile_X9Y13_to_SI_1s;
wire[1:0] Tile_X10Y13_to_WA_1s;
wire[1:0] Tile_X10Y13_to_WB_1s;
wire[1:0] Tile_X10Y13_to_WC_1s;
wire[1:0] Tile_X10Y13_to_WD_1s;
wire[1:0] Tile_X10Y13_to_WF_1s;
wire[1:0] Tile_X10Y13_to_WG_1s;
wire[1:0] Tile_X10Y13_to_WH_1s;
wire[1:0] Tile_X10Y13_to_WI_1s;
wire[3:0] Tile_X0Y14_to_EA;
wire[3:0] Tile_X0Y14_to_EB;
wire[3:0] Tile_X0Y14_to_EC;
wire[3:0] Tile_X0Y14_to_ED;
wire[3:0] Tile_X0Y14_to_EF;
wire[7:0] Tile_X0Y14_to_EG;
wire[7:0] Tile_X0Y14_to_EH;
wire[11:0] Tile_X0Y14_to_EI;
wire[3:0] Tile_X0Y14_to_NA;
wire[3:0] Tile_X0Y14_to_NB;
wire[3:0] Tile_X0Y14_to_NC;
wire[3:0] Tile_X0Y14_to_ND;
wire[3:0] Tile_X0Y14_to_NF;
wire[7:0] Tile_X0Y14_to_NG;
wire[7:0] Tile_X0Y14_to_NH;
wire[11:0] Tile_X0Y14_to_NI;
wire[3:0] Tile_X0Y14_to_SA;
wire[3:0] Tile_X0Y14_to_SB;
wire[3:0] Tile_X0Y14_to_SC;
wire[3:0] Tile_X0Y14_to_SD;
wire[3:0] Tile_X0Y14_to_SF;
wire[7:0] Tile_X0Y14_to_SG;
wire[7:0] Tile_X0Y14_to_SH;
wire[11:0] Tile_X0Y14_to_SI;
wire[3:0] Tile_X1Y14_to_EA;
wire[3:0] Tile_X1Y14_to_EB;
wire[3:0] Tile_X1Y14_to_EC;
wire[3:0] Tile_X1Y14_to_ED;
wire[3:0] Tile_X1Y14_to_EF;
wire[7:0] Tile_X1Y14_to_EG;
wire[7:0] Tile_X1Y14_to_EH;
wire[11:0] Tile_X1Y14_to_EI;
wire[3:0] Tile_X1Y14_to_WA;
wire[3:0] Tile_X1Y14_to_WB;
wire[3:0] Tile_X1Y14_to_WC;
wire[3:0] Tile_X1Y14_to_WD;
wire[3:0] Tile_X1Y14_to_WF;
wire[7:0] Tile_X1Y14_to_WG;
wire[7:0] Tile_X1Y14_to_WH;
wire[11:0] Tile_X1Y14_to_WI;
wire[3:0] Tile_X1Y14_to_NA;
wire[3:0] Tile_X1Y14_to_NB;
wire[3:0] Tile_X1Y14_to_NC;
wire[3:0] Tile_X1Y14_to_ND;
wire[3:0] Tile_X1Y14_to_NF;
wire[7:0] Tile_X1Y14_to_NG;
wire[7:0] Tile_X1Y14_to_NH;
wire[11:0] Tile_X1Y14_to_NI;
wire[3:0] Tile_X1Y14_to_SA;
wire[3:0] Tile_X1Y14_to_SB;
wire[3:0] Tile_X1Y14_to_SC;
wire[3:0] Tile_X1Y14_to_SD;
wire[3:0] Tile_X1Y14_to_SF;
wire[7:0] Tile_X1Y14_to_SG;
wire[7:0] Tile_X1Y14_to_SH;
wire[11:0] Tile_X1Y14_to_SI;
wire[3:0] Tile_X2Y14_to_EA;
wire[3:0] Tile_X2Y14_to_EB;
wire[3:0] Tile_X2Y14_to_EC;
wire[3:0] Tile_X2Y14_to_ED;
wire[3:0] Tile_X2Y14_to_EF;
wire[7:0] Tile_X2Y14_to_EG;
wire[7:0] Tile_X2Y14_to_EH;
wire[11:0] Tile_X2Y14_to_EI;
wire[3:0] Tile_X2Y14_to_WA;
wire[3:0] Tile_X2Y14_to_WB;
wire[3:0] Tile_X2Y14_to_WC;
wire[3:0] Tile_X2Y14_to_WD;
wire[3:0] Tile_X2Y14_to_WF;
wire[7:0] Tile_X2Y14_to_WG;
wire[7:0] Tile_X2Y14_to_WH;
wire[11:0] Tile_X2Y14_to_WI;
wire[3:0] Tile_X2Y14_to_NA;
wire[3:0] Tile_X2Y14_to_NB;
wire[3:0] Tile_X2Y14_to_NC;
wire[3:0] Tile_X2Y14_to_ND;
wire[3:0] Tile_X2Y14_to_NF;
wire[7:0] Tile_X2Y14_to_NG;
wire[7:0] Tile_X2Y14_to_NH;
wire[11:0] Tile_X2Y14_to_NI;
wire[3:0] Tile_X2Y14_to_SA;
wire[3:0] Tile_X2Y14_to_SB;
wire[3:0] Tile_X2Y14_to_SC;
wire[3:0] Tile_X2Y14_to_SD;
wire[3:0] Tile_X2Y14_to_SF;
wire[7:0] Tile_X2Y14_to_SG;
wire[7:0] Tile_X2Y14_to_SH;
wire[11:0] Tile_X2Y14_to_SI;
wire[3:0] Tile_X3Y14_to_EA;
wire[3:0] Tile_X3Y14_to_EB;
wire[3:0] Tile_X3Y14_to_EC;
wire[3:0] Tile_X3Y14_to_ED;
wire[3:0] Tile_X3Y14_to_EF;
wire[7:0] Tile_X3Y14_to_EG;
wire[7:0] Tile_X3Y14_to_EH;
wire[11:0] Tile_X3Y14_to_EI;
wire[3:0] Tile_X3Y14_to_WA;
wire[3:0] Tile_X3Y14_to_WB;
wire[3:0] Tile_X3Y14_to_WC;
wire[3:0] Tile_X3Y14_to_WD;
wire[3:0] Tile_X3Y14_to_WF;
wire[7:0] Tile_X3Y14_to_WG;
wire[7:0] Tile_X3Y14_to_WH;
wire[11:0] Tile_X3Y14_to_WI;
wire[3:0] Tile_X3Y14_to_NA;
wire[3:0] Tile_X3Y14_to_NB;
wire[3:0] Tile_X3Y14_to_NC;
wire[3:0] Tile_X3Y14_to_ND;
wire[3:0] Tile_X3Y14_to_NF;
wire[7:0] Tile_X3Y14_to_NG;
wire[7:0] Tile_X3Y14_to_NH;
wire[11:0] Tile_X3Y14_to_NI;
wire[3:0] Tile_X3Y14_to_SA;
wire[3:0] Tile_X3Y14_to_SB;
wire[3:0] Tile_X3Y14_to_SC;
wire[3:0] Tile_X3Y14_to_SD;
wire[3:0] Tile_X3Y14_to_SF;
wire[7:0] Tile_X3Y14_to_SG;
wire[7:0] Tile_X3Y14_to_SH;
wire[11:0] Tile_X3Y14_to_SI;
wire[3:0] Tile_X4Y14_to_EA;
wire[3:0] Tile_X4Y14_to_EB;
wire[3:0] Tile_X4Y14_to_EC;
wire[3:0] Tile_X4Y14_to_ED;
wire[3:0] Tile_X4Y14_to_EF;
wire[7:0] Tile_X4Y14_to_EG;
wire[7:0] Tile_X4Y14_to_EH;
wire[11:0] Tile_X4Y14_to_EI;
wire[3:0] Tile_X4Y14_to_WA;
wire[3:0] Tile_X4Y14_to_WB;
wire[3:0] Tile_X4Y14_to_WC;
wire[3:0] Tile_X4Y14_to_WD;
wire[3:0] Tile_X4Y14_to_WF;
wire[7:0] Tile_X4Y14_to_WG;
wire[7:0] Tile_X4Y14_to_WH;
wire[11:0] Tile_X4Y14_to_WI;
wire[3:0] Tile_X4Y14_to_NA;
wire[3:0] Tile_X4Y14_to_NB;
wire[3:0] Tile_X4Y14_to_NC;
wire[3:0] Tile_X4Y14_to_ND;
wire[3:0] Tile_X4Y14_to_NF;
wire[7:0] Tile_X4Y14_to_NG;
wire[7:0] Tile_X4Y14_to_NH;
wire[11:0] Tile_X4Y14_to_NI;
wire[3:0] Tile_X4Y14_to_SA;
wire[3:0] Tile_X4Y14_to_SB;
wire[3:0] Tile_X4Y14_to_SC;
wire[3:0] Tile_X4Y14_to_SD;
wire[3:0] Tile_X4Y14_to_SF;
wire[7:0] Tile_X4Y14_to_SG;
wire[7:0] Tile_X4Y14_to_SH;
wire[11:0] Tile_X4Y14_to_SI;
wire[3:0] Tile_X5Y14_to_EA;
wire[3:0] Tile_X5Y14_to_EB;
wire[3:0] Tile_X5Y14_to_EC;
wire[3:0] Tile_X5Y14_to_ED;
wire[3:0] Tile_X5Y14_to_EF;
wire[7:0] Tile_X5Y14_to_EG;
wire[7:0] Tile_X5Y14_to_EH;
wire[11:0] Tile_X5Y14_to_EI;
wire[3:0] Tile_X5Y14_to_WA;
wire[3:0] Tile_X5Y14_to_WB;
wire[3:0] Tile_X5Y14_to_WC;
wire[3:0] Tile_X5Y14_to_WD;
wire[3:0] Tile_X5Y14_to_WF;
wire[7:0] Tile_X5Y14_to_WG;
wire[7:0] Tile_X5Y14_to_WH;
wire[11:0] Tile_X5Y14_to_WI;
wire[3:0] Tile_X5Y14_to_NA;
wire[3:0] Tile_X5Y14_to_NB;
wire[3:0] Tile_X5Y14_to_NC;
wire[3:0] Tile_X5Y14_to_ND;
wire[3:0] Tile_X5Y14_to_NF;
wire[7:0] Tile_X5Y14_to_NG;
wire[7:0] Tile_X5Y14_to_NH;
wire[11:0] Tile_X5Y14_to_NI;
wire[3:0] Tile_X5Y14_to_SA;
wire[3:0] Tile_X5Y14_to_SB;
wire[3:0] Tile_X5Y14_to_SC;
wire[3:0] Tile_X5Y14_to_SD;
wire[3:0] Tile_X5Y14_to_SF;
wire[7:0] Tile_X5Y14_to_SG;
wire[7:0] Tile_X5Y14_to_SH;
wire[11:0] Tile_X5Y14_to_SI;
wire[3:0] Tile_X6Y14_to_EA;
wire[3:0] Tile_X6Y14_to_EB;
wire[3:0] Tile_X6Y14_to_EC;
wire[3:0] Tile_X6Y14_to_ED;
wire[3:0] Tile_X6Y14_to_EF;
wire[7:0] Tile_X6Y14_to_EG;
wire[7:0] Tile_X6Y14_to_EH;
wire[11:0] Tile_X6Y14_to_EI;
wire[3:0] Tile_X6Y14_to_WA;
wire[3:0] Tile_X6Y14_to_WB;
wire[3:0] Tile_X6Y14_to_WC;
wire[3:0] Tile_X6Y14_to_WD;
wire[3:0] Tile_X6Y14_to_WF;
wire[7:0] Tile_X6Y14_to_WG;
wire[7:0] Tile_X6Y14_to_WH;
wire[11:0] Tile_X6Y14_to_WI;
wire[3:0] Tile_X6Y14_to_NA;
wire[3:0] Tile_X6Y14_to_NB;
wire[3:0] Tile_X6Y14_to_NC;
wire[3:0] Tile_X6Y14_to_ND;
wire[3:0] Tile_X6Y14_to_NF;
wire[7:0] Tile_X6Y14_to_NG;
wire[7:0] Tile_X6Y14_to_NH;
wire[11:0] Tile_X6Y14_to_NI;
wire[3:0] Tile_X6Y14_to_SA;
wire[3:0] Tile_X6Y14_to_SB;
wire[3:0] Tile_X6Y14_to_SC;
wire[3:0] Tile_X6Y14_to_SD;
wire[3:0] Tile_X6Y14_to_SF;
wire[7:0] Tile_X6Y14_to_SG;
wire[7:0] Tile_X6Y14_to_SH;
wire[11:0] Tile_X6Y14_to_SI;
wire[3:0] Tile_X7Y14_to_EA;
wire[3:0] Tile_X7Y14_to_EB;
wire[3:0] Tile_X7Y14_to_EC;
wire[3:0] Tile_X7Y14_to_ED;
wire[3:0] Tile_X7Y14_to_EF;
wire[7:0] Tile_X7Y14_to_EG;
wire[7:0] Tile_X7Y14_to_EH;
wire[11:0] Tile_X7Y14_to_EI;
wire[3:0] Tile_X7Y14_to_WA;
wire[3:0] Tile_X7Y14_to_WB;
wire[3:0] Tile_X7Y14_to_WC;
wire[3:0] Tile_X7Y14_to_WD;
wire[3:0] Tile_X7Y14_to_WF;
wire[7:0] Tile_X7Y14_to_WG;
wire[7:0] Tile_X7Y14_to_WH;
wire[11:0] Tile_X7Y14_to_WI;
wire[3:0] Tile_X7Y14_to_NA;
wire[3:0] Tile_X7Y14_to_NB;
wire[3:0] Tile_X7Y14_to_NC;
wire[3:0] Tile_X7Y14_to_ND;
wire[3:0] Tile_X7Y14_to_NF;
wire[7:0] Tile_X7Y14_to_NG;
wire[7:0] Tile_X7Y14_to_NH;
wire[11:0] Tile_X7Y14_to_NI;
wire[3:0] Tile_X7Y14_to_SA;
wire[3:0] Tile_X7Y14_to_SB;
wire[3:0] Tile_X7Y14_to_SC;
wire[3:0] Tile_X7Y14_to_SD;
wire[3:0] Tile_X7Y14_to_SF;
wire[7:0] Tile_X7Y14_to_SG;
wire[7:0] Tile_X7Y14_to_SH;
wire[11:0] Tile_X7Y14_to_SI;
wire[3:0] Tile_X8Y14_to_WA;
wire[3:0] Tile_X8Y14_to_WB;
wire[3:0] Tile_X8Y14_to_WC;
wire[3:0] Tile_X8Y14_to_WD;
wire[3:0] Tile_X8Y14_to_WF;
wire[7:0] Tile_X8Y14_to_WG;
wire[7:0] Tile_X8Y14_to_WH;
wire[11:0] Tile_X8Y14_to_WI;
wire[3:0] Tile_X8Y14_to_NA;
wire[3:0] Tile_X8Y14_to_NB;
wire[3:0] Tile_X8Y14_to_NC;
wire[3:0] Tile_X8Y14_to_ND;
wire[3:0] Tile_X8Y14_to_NF;
wire[7:0] Tile_X8Y14_to_NG;
wire[7:0] Tile_X8Y14_to_NH;
wire[11:0] Tile_X8Y14_to_NI;
wire[3:0] Tile_X8Y14_to_SA;
wire[3:0] Tile_X8Y14_to_SB;
wire[3:0] Tile_X8Y14_to_SC;
wire[3:0] Tile_X8Y14_to_SD;
wire[3:0] Tile_X8Y14_to_SF;
wire[7:0] Tile_X8Y14_to_SG;
wire[7:0] Tile_X8Y14_to_SH;
wire[11:0] Tile_X8Y14_to_SI;
wire[1:0] Tile_X9Y14_to_EA_1s;
wire[1:0] Tile_X9Y14_to_EB_1s;
wire[1:0] Tile_X9Y14_to_EC_1s;
wire[1:0] Tile_X9Y14_to_ED_1s;
wire[1:0] Tile_X9Y14_to_EF_1s;
wire[1:0] Tile_X9Y14_to_EG_1s;
wire[1:0] Tile_X9Y14_to_EH_1s;
wire[1:0] Tile_X9Y14_to_EI_1s;
wire[1:0] Tile_X9Y14_to_WA_1s;
wire[1:0] Tile_X9Y14_to_WB_1s;
wire[1:0] Tile_X9Y14_to_WC_1s;
wire[1:0] Tile_X9Y14_to_WD_1s;
wire[1:0] Tile_X9Y14_to_WF_1s;
wire[1:0] Tile_X9Y14_to_WG_1s;
wire[1:0] Tile_X9Y14_to_WH_1s;
wire[1:0] Tile_X9Y14_to_WI_1s;
wire[1:0] Tile_X9Y14_to_NA_1s;
wire[1:0] Tile_X9Y14_to_NB_1s;
wire[1:0] Tile_X9Y14_to_NC_1s;
wire[1:0] Tile_X9Y14_to_ND_1s;
wire[1:0] Tile_X9Y14_to_NF_1s;
wire[1:0] Tile_X9Y14_to_NG_1s;
wire[1:0] Tile_X9Y14_to_NH_1s;
wire[1:0] Tile_X9Y14_to_NI_1s;
wire[1:0] Tile_X9Y14_to_SA_1s;
wire[1:0] Tile_X9Y14_to_SB_1s;
wire[1:0] Tile_X9Y14_to_SC_1s;
wire[1:0] Tile_X9Y14_to_SD_1s;
wire[1:0] Tile_X9Y14_to_SF_1s;
wire[1:0] Tile_X9Y14_to_SG_1s;
wire[1:0] Tile_X9Y14_to_SH_1s;
wire[1:0] Tile_X9Y14_to_SI_1s;
wire[1:0] Tile_X10Y14_to_WA_1s;
wire[1:0] Tile_X10Y14_to_WB_1s;
wire[1:0] Tile_X10Y14_to_WC_1s;
wire[1:0] Tile_X10Y14_to_WD_1s;
wire[1:0] Tile_X10Y14_to_WF_1s;
wire[1:0] Tile_X10Y14_to_WG_1s;
wire[1:0] Tile_X10Y14_to_WH_1s;
wire[1:0] Tile_X10Y14_to_WI_1s;
wire[3:0] Tile_X0Y15_to_EA;
wire[3:0] Tile_X0Y15_to_EB;
wire[3:0] Tile_X0Y15_to_EC;
wire[3:0] Tile_X0Y15_to_ED;
wire[3:0] Tile_X0Y15_to_EF;
wire[7:0] Tile_X0Y15_to_EG;
wire[7:0] Tile_X0Y15_to_EH;
wire[11:0] Tile_X0Y15_to_EI;
wire[3:0] Tile_X0Y15_to_NA;
wire[3:0] Tile_X0Y15_to_NB;
wire[3:0] Tile_X0Y15_to_NC;
wire[3:0] Tile_X0Y15_to_ND;
wire[3:0] Tile_X0Y15_to_NF;
wire[7:0] Tile_X0Y15_to_NG;
wire[7:0] Tile_X0Y15_to_NH;
wire[11:0] Tile_X0Y15_to_NI;
wire[3:0] Tile_X0Y15_to_SA;
wire[3:0] Tile_X0Y15_to_SB;
wire[3:0] Tile_X0Y15_to_SC;
wire[3:0] Tile_X0Y15_to_SD;
wire[3:0] Tile_X0Y15_to_SF;
wire[7:0] Tile_X0Y15_to_SG;
wire[7:0] Tile_X0Y15_to_SH;
wire[11:0] Tile_X0Y15_to_SI;
wire[3:0] Tile_X1Y15_to_EA;
wire[3:0] Tile_X1Y15_to_EB;
wire[3:0] Tile_X1Y15_to_EC;
wire[3:0] Tile_X1Y15_to_ED;
wire[3:0] Tile_X1Y15_to_EF;
wire[7:0] Tile_X1Y15_to_EG;
wire[7:0] Tile_X1Y15_to_EH;
wire[11:0] Tile_X1Y15_to_EI;
wire[3:0] Tile_X1Y15_to_WA;
wire[3:0] Tile_X1Y15_to_WB;
wire[3:0] Tile_X1Y15_to_WC;
wire[3:0] Tile_X1Y15_to_WD;
wire[3:0] Tile_X1Y15_to_WF;
wire[7:0] Tile_X1Y15_to_WG;
wire[7:0] Tile_X1Y15_to_WH;
wire[11:0] Tile_X1Y15_to_WI;
wire[3:0] Tile_X1Y15_to_NA;
wire[3:0] Tile_X1Y15_to_NB;
wire[3:0] Tile_X1Y15_to_NC;
wire[3:0] Tile_X1Y15_to_ND;
wire[3:0] Tile_X1Y15_to_NF;
wire[7:0] Tile_X1Y15_to_NG;
wire[7:0] Tile_X1Y15_to_NH;
wire[11:0] Tile_X1Y15_to_NI;
wire[3:0] Tile_X1Y15_to_SA;
wire[3:0] Tile_X1Y15_to_SB;
wire[3:0] Tile_X1Y15_to_SC;
wire[3:0] Tile_X1Y15_to_SD;
wire[3:0] Tile_X1Y15_to_SF;
wire[7:0] Tile_X1Y15_to_SG;
wire[7:0] Tile_X1Y15_to_SH;
wire[11:0] Tile_X1Y15_to_SI;
wire[3:0] Tile_X2Y15_to_EA;
wire[3:0] Tile_X2Y15_to_EB;
wire[3:0] Tile_X2Y15_to_EC;
wire[3:0] Tile_X2Y15_to_ED;
wire[3:0] Tile_X2Y15_to_EF;
wire[7:0] Tile_X2Y15_to_EG;
wire[7:0] Tile_X2Y15_to_EH;
wire[11:0] Tile_X2Y15_to_EI;
wire[3:0] Tile_X2Y15_to_WA;
wire[3:0] Tile_X2Y15_to_WB;
wire[3:0] Tile_X2Y15_to_WC;
wire[3:0] Tile_X2Y15_to_WD;
wire[3:0] Tile_X2Y15_to_WF;
wire[7:0] Tile_X2Y15_to_WG;
wire[7:0] Tile_X2Y15_to_WH;
wire[11:0] Tile_X2Y15_to_WI;
wire[3:0] Tile_X2Y15_to_NA;
wire[3:0] Tile_X2Y15_to_NB;
wire[3:0] Tile_X2Y15_to_NC;
wire[3:0] Tile_X2Y15_to_ND;
wire[3:0] Tile_X2Y15_to_NF;
wire[7:0] Tile_X2Y15_to_NG;
wire[7:0] Tile_X2Y15_to_NH;
wire[11:0] Tile_X2Y15_to_NI;
wire[3:0] Tile_X2Y15_to_SA;
wire[3:0] Tile_X2Y15_to_SB;
wire[3:0] Tile_X2Y15_to_SC;
wire[3:0] Tile_X2Y15_to_SD;
wire[3:0] Tile_X2Y15_to_SF;
wire[7:0] Tile_X2Y15_to_SG;
wire[7:0] Tile_X2Y15_to_SH;
wire[11:0] Tile_X2Y15_to_SI;
wire[3:0] Tile_X3Y15_to_EA;
wire[3:0] Tile_X3Y15_to_EB;
wire[3:0] Tile_X3Y15_to_EC;
wire[3:0] Tile_X3Y15_to_ED;
wire[3:0] Tile_X3Y15_to_EF;
wire[7:0] Tile_X3Y15_to_EG;
wire[7:0] Tile_X3Y15_to_EH;
wire[11:0] Tile_X3Y15_to_EI;
wire[3:0] Tile_X3Y15_to_WA;
wire[3:0] Tile_X3Y15_to_WB;
wire[3:0] Tile_X3Y15_to_WC;
wire[3:0] Tile_X3Y15_to_WD;
wire[3:0] Tile_X3Y15_to_WF;
wire[7:0] Tile_X3Y15_to_WG;
wire[7:0] Tile_X3Y15_to_WH;
wire[11:0] Tile_X3Y15_to_WI;
wire[3:0] Tile_X3Y15_to_NA;
wire[3:0] Tile_X3Y15_to_NB;
wire[3:0] Tile_X3Y15_to_NC;
wire[3:0] Tile_X3Y15_to_ND;
wire[3:0] Tile_X3Y15_to_NF;
wire[7:0] Tile_X3Y15_to_NG;
wire[7:0] Tile_X3Y15_to_NH;
wire[11:0] Tile_X3Y15_to_NI;
wire[3:0] Tile_X3Y15_to_SA;
wire[3:0] Tile_X3Y15_to_SB;
wire[3:0] Tile_X3Y15_to_SC;
wire[3:0] Tile_X3Y15_to_SD;
wire[3:0] Tile_X3Y15_to_SF;
wire[7:0] Tile_X3Y15_to_SG;
wire[7:0] Tile_X3Y15_to_SH;
wire[11:0] Tile_X3Y15_to_SI;
wire[3:0] Tile_X4Y15_to_EA;
wire[3:0] Tile_X4Y15_to_EB;
wire[3:0] Tile_X4Y15_to_EC;
wire[3:0] Tile_X4Y15_to_ED;
wire[3:0] Tile_X4Y15_to_EF;
wire[7:0] Tile_X4Y15_to_EG;
wire[7:0] Tile_X4Y15_to_EH;
wire[11:0] Tile_X4Y15_to_EI;
wire[3:0] Tile_X4Y15_to_WA;
wire[3:0] Tile_X4Y15_to_WB;
wire[3:0] Tile_X4Y15_to_WC;
wire[3:0] Tile_X4Y15_to_WD;
wire[3:0] Tile_X4Y15_to_WF;
wire[7:0] Tile_X4Y15_to_WG;
wire[7:0] Tile_X4Y15_to_WH;
wire[11:0] Tile_X4Y15_to_WI;
wire[3:0] Tile_X4Y15_to_NA;
wire[3:0] Tile_X4Y15_to_NB;
wire[3:0] Tile_X4Y15_to_NC;
wire[3:0] Tile_X4Y15_to_ND;
wire[3:0] Tile_X4Y15_to_NF;
wire[7:0] Tile_X4Y15_to_NG;
wire[7:0] Tile_X4Y15_to_NH;
wire[11:0] Tile_X4Y15_to_NI;
wire[3:0] Tile_X4Y15_to_SA;
wire[3:0] Tile_X4Y15_to_SB;
wire[3:0] Tile_X4Y15_to_SC;
wire[3:0] Tile_X4Y15_to_SD;
wire[3:0] Tile_X4Y15_to_SF;
wire[7:0] Tile_X4Y15_to_SG;
wire[7:0] Tile_X4Y15_to_SH;
wire[11:0] Tile_X4Y15_to_SI;
wire[3:0] Tile_X5Y15_to_EA;
wire[3:0] Tile_X5Y15_to_EB;
wire[3:0] Tile_X5Y15_to_EC;
wire[3:0] Tile_X5Y15_to_ED;
wire[3:0] Tile_X5Y15_to_EF;
wire[7:0] Tile_X5Y15_to_EG;
wire[7:0] Tile_X5Y15_to_EH;
wire[11:0] Tile_X5Y15_to_EI;
wire[3:0] Tile_X5Y15_to_WA;
wire[3:0] Tile_X5Y15_to_WB;
wire[3:0] Tile_X5Y15_to_WC;
wire[3:0] Tile_X5Y15_to_WD;
wire[3:0] Tile_X5Y15_to_WF;
wire[7:0] Tile_X5Y15_to_WG;
wire[7:0] Tile_X5Y15_to_WH;
wire[11:0] Tile_X5Y15_to_WI;
wire[3:0] Tile_X5Y15_to_NA;
wire[3:0] Tile_X5Y15_to_NB;
wire[3:0] Tile_X5Y15_to_NC;
wire[3:0] Tile_X5Y15_to_ND;
wire[3:0] Tile_X5Y15_to_NF;
wire[7:0] Tile_X5Y15_to_NG;
wire[7:0] Tile_X5Y15_to_NH;
wire[11:0] Tile_X5Y15_to_NI;
wire[3:0] Tile_X5Y15_to_SA;
wire[3:0] Tile_X5Y15_to_SB;
wire[3:0] Tile_X5Y15_to_SC;
wire[3:0] Tile_X5Y15_to_SD;
wire[3:0] Tile_X5Y15_to_SF;
wire[7:0] Tile_X5Y15_to_SG;
wire[7:0] Tile_X5Y15_to_SH;
wire[11:0] Tile_X5Y15_to_SI;
wire[3:0] Tile_X6Y15_to_EA;
wire[3:0] Tile_X6Y15_to_EB;
wire[3:0] Tile_X6Y15_to_EC;
wire[3:0] Tile_X6Y15_to_ED;
wire[3:0] Tile_X6Y15_to_EF;
wire[7:0] Tile_X6Y15_to_EG;
wire[7:0] Tile_X6Y15_to_EH;
wire[11:0] Tile_X6Y15_to_EI;
wire[3:0] Tile_X6Y15_to_WA;
wire[3:0] Tile_X6Y15_to_WB;
wire[3:0] Tile_X6Y15_to_WC;
wire[3:0] Tile_X6Y15_to_WD;
wire[3:0] Tile_X6Y15_to_WF;
wire[7:0] Tile_X6Y15_to_WG;
wire[7:0] Tile_X6Y15_to_WH;
wire[11:0] Tile_X6Y15_to_WI;
wire[3:0] Tile_X6Y15_to_NA;
wire[3:0] Tile_X6Y15_to_NB;
wire[3:0] Tile_X6Y15_to_NC;
wire[3:0] Tile_X6Y15_to_ND;
wire[3:0] Tile_X6Y15_to_NF;
wire[7:0] Tile_X6Y15_to_NG;
wire[7:0] Tile_X6Y15_to_NH;
wire[11:0] Tile_X6Y15_to_NI;
wire[3:0] Tile_X6Y15_to_SA;
wire[3:0] Tile_X6Y15_to_SB;
wire[3:0] Tile_X6Y15_to_SC;
wire[3:0] Tile_X6Y15_to_SD;
wire[3:0] Tile_X6Y15_to_SF;
wire[7:0] Tile_X6Y15_to_SG;
wire[7:0] Tile_X6Y15_to_SH;
wire[11:0] Tile_X6Y15_to_SI;
wire[3:0] Tile_X7Y15_to_EA;
wire[3:0] Tile_X7Y15_to_EB;
wire[3:0] Tile_X7Y15_to_EC;
wire[3:0] Tile_X7Y15_to_ED;
wire[3:0] Tile_X7Y15_to_EF;
wire[7:0] Tile_X7Y15_to_EG;
wire[7:0] Tile_X7Y15_to_EH;
wire[11:0] Tile_X7Y15_to_EI;
wire[3:0] Tile_X7Y15_to_WA;
wire[3:0] Tile_X7Y15_to_WB;
wire[3:0] Tile_X7Y15_to_WC;
wire[3:0] Tile_X7Y15_to_WD;
wire[3:0] Tile_X7Y15_to_WF;
wire[7:0] Tile_X7Y15_to_WG;
wire[7:0] Tile_X7Y15_to_WH;
wire[11:0] Tile_X7Y15_to_WI;
wire[3:0] Tile_X7Y15_to_NA;
wire[3:0] Tile_X7Y15_to_NB;
wire[3:0] Tile_X7Y15_to_NC;
wire[3:0] Tile_X7Y15_to_ND;
wire[3:0] Tile_X7Y15_to_NF;
wire[7:0] Tile_X7Y15_to_NG;
wire[7:0] Tile_X7Y15_to_NH;
wire[11:0] Tile_X7Y15_to_NI;
wire[3:0] Tile_X7Y15_to_SA;
wire[3:0] Tile_X7Y15_to_SB;
wire[3:0] Tile_X7Y15_to_SC;
wire[3:0] Tile_X7Y15_to_SD;
wire[3:0] Tile_X7Y15_to_SF;
wire[7:0] Tile_X7Y15_to_SG;
wire[7:0] Tile_X7Y15_to_SH;
wire[11:0] Tile_X7Y15_to_SI;
wire[3:0] Tile_X8Y15_to_WA;
wire[3:0] Tile_X8Y15_to_WB;
wire[3:0] Tile_X8Y15_to_WC;
wire[3:0] Tile_X8Y15_to_WD;
wire[3:0] Tile_X8Y15_to_WF;
wire[7:0] Tile_X8Y15_to_WG;
wire[7:0] Tile_X8Y15_to_WH;
wire[11:0] Tile_X8Y15_to_WI;
wire[3:0] Tile_X8Y15_to_NA;
wire[3:0] Tile_X8Y15_to_NB;
wire[3:0] Tile_X8Y15_to_NC;
wire[3:0] Tile_X8Y15_to_ND;
wire[3:0] Tile_X8Y15_to_NF;
wire[7:0] Tile_X8Y15_to_NG;
wire[7:0] Tile_X8Y15_to_NH;
wire[11:0] Tile_X8Y15_to_NI;
wire[3:0] Tile_X8Y15_to_SA;
wire[3:0] Tile_X8Y15_to_SB;
wire[3:0] Tile_X8Y15_to_SC;
wire[3:0] Tile_X8Y15_to_SD;
wire[3:0] Tile_X8Y15_to_SF;
wire[7:0] Tile_X8Y15_to_SG;
wire[7:0] Tile_X8Y15_to_SH;
wire[11:0] Tile_X8Y15_to_SI;
wire[1:0] Tile_X9Y15_to_EA_1s;
wire[1:0] Tile_X9Y15_to_EB_1s;
wire[1:0] Tile_X9Y15_to_EC_1s;
wire[1:0] Tile_X9Y15_to_ED_1s;
wire[1:0] Tile_X9Y15_to_EF_1s;
wire[1:0] Tile_X9Y15_to_EG_1s;
wire[1:0] Tile_X9Y15_to_EH_1s;
wire[1:0] Tile_X9Y15_to_EI_1s;
wire[1:0] Tile_X9Y15_to_WA_1s;
wire[1:0] Tile_X9Y15_to_WB_1s;
wire[1:0] Tile_X9Y15_to_WC_1s;
wire[1:0] Tile_X9Y15_to_WD_1s;
wire[1:0] Tile_X9Y15_to_WF_1s;
wire[1:0] Tile_X9Y15_to_WG_1s;
wire[1:0] Tile_X9Y15_to_WH_1s;
wire[1:0] Tile_X9Y15_to_WI_1s;
wire[1:0] Tile_X9Y15_to_NA_1s;
wire[1:0] Tile_X9Y15_to_NB_1s;
wire[1:0] Tile_X9Y15_to_NC_1s;
wire[1:0] Tile_X9Y15_to_ND_1s;
wire[1:0] Tile_X9Y15_to_NF_1s;
wire[1:0] Tile_X9Y15_to_NG_1s;
wire[1:0] Tile_X9Y15_to_NH_1s;
wire[1:0] Tile_X9Y15_to_NI_1s;
wire[1:0] Tile_X9Y15_to_SA_1s;
wire[1:0] Tile_X9Y15_to_SB_1s;
wire[1:0] Tile_X9Y15_to_SC_1s;
wire[1:0] Tile_X9Y15_to_SD_1s;
wire[1:0] Tile_X9Y15_to_SF_1s;
wire[1:0] Tile_X9Y15_to_SG_1s;
wire[1:0] Tile_X9Y15_to_SH_1s;
wire[1:0] Tile_X9Y15_to_SI_1s;
wire[1:0] Tile_X10Y15_to_WA_1s;
wire[1:0] Tile_X10Y15_to_WB_1s;
wire[1:0] Tile_X10Y15_to_WC_1s;
wire[1:0] Tile_X10Y15_to_WD_1s;
wire[1:0] Tile_X10Y15_to_WF_1s;
wire[1:0] Tile_X10Y15_to_WG_1s;
wire[1:0] Tile_X10Y15_to_WH_1s;
wire[1:0] Tile_X10Y15_to_WI_1s;
wire[3:0] Tile_X0Y16_to_EA;
wire[3:0] Tile_X0Y16_to_EB;
wire[3:0] Tile_X0Y16_to_EC;
wire[3:0] Tile_X0Y16_to_ED;
wire[3:0] Tile_X0Y16_to_EF;
wire[7:0] Tile_X0Y16_to_EG;
wire[7:0] Tile_X0Y16_to_EH;
wire[11:0] Tile_X0Y16_to_EI;
wire[3:0] Tile_X0Y16_to_NA;
wire[3:0] Tile_X0Y16_to_NB;
wire[3:0] Tile_X0Y16_to_NC;
wire[3:0] Tile_X0Y16_to_ND;
wire[3:0] Tile_X0Y16_to_NF;
wire[7:0] Tile_X0Y16_to_NG;
wire[7:0] Tile_X0Y16_to_NH;
wire[11:0] Tile_X0Y16_to_NI;
wire[3:0] Tile_X0Y16_to_SA;
wire[3:0] Tile_X0Y16_to_SB;
wire[3:0] Tile_X0Y16_to_SC;
wire[3:0] Tile_X0Y16_to_SD;
wire[3:0] Tile_X0Y16_to_SF;
wire[7:0] Tile_X0Y16_to_SG;
wire[7:0] Tile_X0Y16_to_SH;
wire[11:0] Tile_X0Y16_to_SI;
wire[3:0] Tile_X1Y16_to_EA;
wire[3:0] Tile_X1Y16_to_EB;
wire[3:0] Tile_X1Y16_to_EC;
wire[3:0] Tile_X1Y16_to_ED;
wire[3:0] Tile_X1Y16_to_EF;
wire[7:0] Tile_X1Y16_to_EG;
wire[7:0] Tile_X1Y16_to_EH;
wire[11:0] Tile_X1Y16_to_EI;
wire[3:0] Tile_X1Y16_to_WA;
wire[3:0] Tile_X1Y16_to_WB;
wire[3:0] Tile_X1Y16_to_WC;
wire[3:0] Tile_X1Y16_to_WD;
wire[3:0] Tile_X1Y16_to_WF;
wire[7:0] Tile_X1Y16_to_WG;
wire[7:0] Tile_X1Y16_to_WH;
wire[11:0] Tile_X1Y16_to_WI;
wire[3:0] Tile_X1Y16_to_NA;
wire[3:0] Tile_X1Y16_to_NB;
wire[3:0] Tile_X1Y16_to_NC;
wire[3:0] Tile_X1Y16_to_ND;
wire[3:0] Tile_X1Y16_to_NF;
wire[7:0] Tile_X1Y16_to_NG;
wire[7:0] Tile_X1Y16_to_NH;
wire[11:0] Tile_X1Y16_to_NI;
wire[3:0] Tile_X1Y16_to_SA;
wire[3:0] Tile_X1Y16_to_SB;
wire[3:0] Tile_X1Y16_to_SC;
wire[3:0] Tile_X1Y16_to_SD;
wire[3:0] Tile_X1Y16_to_SF;
wire[7:0] Tile_X1Y16_to_SG;
wire[7:0] Tile_X1Y16_to_SH;
wire[11:0] Tile_X1Y16_to_SI;
wire[3:0] Tile_X2Y16_to_EA;
wire[3:0] Tile_X2Y16_to_EB;
wire[3:0] Tile_X2Y16_to_EC;
wire[3:0] Tile_X2Y16_to_ED;
wire[3:0] Tile_X2Y16_to_EF;
wire[7:0] Tile_X2Y16_to_EG;
wire[7:0] Tile_X2Y16_to_EH;
wire[11:0] Tile_X2Y16_to_EI;
wire[3:0] Tile_X2Y16_to_WA;
wire[3:0] Tile_X2Y16_to_WB;
wire[3:0] Tile_X2Y16_to_WC;
wire[3:0] Tile_X2Y16_to_WD;
wire[3:0] Tile_X2Y16_to_WF;
wire[7:0] Tile_X2Y16_to_WG;
wire[7:0] Tile_X2Y16_to_WH;
wire[11:0] Tile_X2Y16_to_WI;
wire[3:0] Tile_X2Y16_to_NA;
wire[3:0] Tile_X2Y16_to_NB;
wire[3:0] Tile_X2Y16_to_NC;
wire[3:0] Tile_X2Y16_to_ND;
wire[3:0] Tile_X2Y16_to_NF;
wire[7:0] Tile_X2Y16_to_NG;
wire[7:0] Tile_X2Y16_to_NH;
wire[11:0] Tile_X2Y16_to_NI;
wire[3:0] Tile_X2Y16_to_SA;
wire[3:0] Tile_X2Y16_to_SB;
wire[3:0] Tile_X2Y16_to_SC;
wire[3:0] Tile_X2Y16_to_SD;
wire[3:0] Tile_X2Y16_to_SF;
wire[7:0] Tile_X2Y16_to_SG;
wire[7:0] Tile_X2Y16_to_SH;
wire[11:0] Tile_X2Y16_to_SI;
wire[3:0] Tile_X3Y16_to_EA;
wire[3:0] Tile_X3Y16_to_EB;
wire[3:0] Tile_X3Y16_to_EC;
wire[3:0] Tile_X3Y16_to_ED;
wire[3:0] Tile_X3Y16_to_EF;
wire[7:0] Tile_X3Y16_to_EG;
wire[7:0] Tile_X3Y16_to_EH;
wire[11:0] Tile_X3Y16_to_EI;
wire[3:0] Tile_X3Y16_to_WA;
wire[3:0] Tile_X3Y16_to_WB;
wire[3:0] Tile_X3Y16_to_WC;
wire[3:0] Tile_X3Y16_to_WD;
wire[3:0] Tile_X3Y16_to_WF;
wire[7:0] Tile_X3Y16_to_WG;
wire[7:0] Tile_X3Y16_to_WH;
wire[11:0] Tile_X3Y16_to_WI;
wire[3:0] Tile_X3Y16_to_NA;
wire[3:0] Tile_X3Y16_to_NB;
wire[3:0] Tile_X3Y16_to_NC;
wire[3:0] Tile_X3Y16_to_ND;
wire[3:0] Tile_X3Y16_to_NF;
wire[7:0] Tile_X3Y16_to_NG;
wire[7:0] Tile_X3Y16_to_NH;
wire[11:0] Tile_X3Y16_to_NI;
wire[3:0] Tile_X3Y16_to_SA;
wire[3:0] Tile_X3Y16_to_SB;
wire[3:0] Tile_X3Y16_to_SC;
wire[3:0] Tile_X3Y16_to_SD;
wire[3:0] Tile_X3Y16_to_SF;
wire[7:0] Tile_X3Y16_to_SG;
wire[7:0] Tile_X3Y16_to_SH;
wire[11:0] Tile_X3Y16_to_SI;
wire[3:0] Tile_X4Y16_to_EA;
wire[3:0] Tile_X4Y16_to_EB;
wire[3:0] Tile_X4Y16_to_EC;
wire[3:0] Tile_X4Y16_to_ED;
wire[3:0] Tile_X4Y16_to_EF;
wire[7:0] Tile_X4Y16_to_EG;
wire[7:0] Tile_X4Y16_to_EH;
wire[11:0] Tile_X4Y16_to_EI;
wire[3:0] Tile_X4Y16_to_WA;
wire[3:0] Tile_X4Y16_to_WB;
wire[3:0] Tile_X4Y16_to_WC;
wire[3:0] Tile_X4Y16_to_WD;
wire[3:0] Tile_X4Y16_to_WF;
wire[7:0] Tile_X4Y16_to_WG;
wire[7:0] Tile_X4Y16_to_WH;
wire[11:0] Tile_X4Y16_to_WI;
wire[3:0] Tile_X4Y16_to_NA;
wire[3:0] Tile_X4Y16_to_NB;
wire[3:0] Tile_X4Y16_to_NC;
wire[3:0] Tile_X4Y16_to_ND;
wire[3:0] Tile_X4Y16_to_NF;
wire[7:0] Tile_X4Y16_to_NG;
wire[7:0] Tile_X4Y16_to_NH;
wire[11:0] Tile_X4Y16_to_NI;
wire[3:0] Tile_X4Y16_to_SA;
wire[3:0] Tile_X4Y16_to_SB;
wire[3:0] Tile_X4Y16_to_SC;
wire[3:0] Tile_X4Y16_to_SD;
wire[3:0] Tile_X4Y16_to_SF;
wire[7:0] Tile_X4Y16_to_SG;
wire[7:0] Tile_X4Y16_to_SH;
wire[11:0] Tile_X4Y16_to_SI;
wire[3:0] Tile_X5Y16_to_EA;
wire[3:0] Tile_X5Y16_to_EB;
wire[3:0] Tile_X5Y16_to_EC;
wire[3:0] Tile_X5Y16_to_ED;
wire[3:0] Tile_X5Y16_to_EF;
wire[7:0] Tile_X5Y16_to_EG;
wire[7:0] Tile_X5Y16_to_EH;
wire[11:0] Tile_X5Y16_to_EI;
wire[3:0] Tile_X5Y16_to_WA;
wire[3:0] Tile_X5Y16_to_WB;
wire[3:0] Tile_X5Y16_to_WC;
wire[3:0] Tile_X5Y16_to_WD;
wire[3:0] Tile_X5Y16_to_WF;
wire[7:0] Tile_X5Y16_to_WG;
wire[7:0] Tile_X5Y16_to_WH;
wire[11:0] Tile_X5Y16_to_WI;
wire[3:0] Tile_X5Y16_to_NA;
wire[3:0] Tile_X5Y16_to_NB;
wire[3:0] Tile_X5Y16_to_NC;
wire[3:0] Tile_X5Y16_to_ND;
wire[3:0] Tile_X5Y16_to_NF;
wire[7:0] Tile_X5Y16_to_NG;
wire[7:0] Tile_X5Y16_to_NH;
wire[11:0] Tile_X5Y16_to_NI;
wire[3:0] Tile_X5Y16_to_SA;
wire[3:0] Tile_X5Y16_to_SB;
wire[3:0] Tile_X5Y16_to_SC;
wire[3:0] Tile_X5Y16_to_SD;
wire[3:0] Tile_X5Y16_to_SF;
wire[7:0] Tile_X5Y16_to_SG;
wire[7:0] Tile_X5Y16_to_SH;
wire[11:0] Tile_X5Y16_to_SI;
wire[3:0] Tile_X6Y16_to_EA;
wire[3:0] Tile_X6Y16_to_EB;
wire[3:0] Tile_X6Y16_to_EC;
wire[3:0] Tile_X6Y16_to_ED;
wire[3:0] Tile_X6Y16_to_EF;
wire[7:0] Tile_X6Y16_to_EG;
wire[7:0] Tile_X6Y16_to_EH;
wire[11:0] Tile_X6Y16_to_EI;
wire[3:0] Tile_X6Y16_to_WA;
wire[3:0] Tile_X6Y16_to_WB;
wire[3:0] Tile_X6Y16_to_WC;
wire[3:0] Tile_X6Y16_to_WD;
wire[3:0] Tile_X6Y16_to_WF;
wire[7:0] Tile_X6Y16_to_WG;
wire[7:0] Tile_X6Y16_to_WH;
wire[11:0] Tile_X6Y16_to_WI;
wire[3:0] Tile_X6Y16_to_NA;
wire[3:0] Tile_X6Y16_to_NB;
wire[3:0] Tile_X6Y16_to_NC;
wire[3:0] Tile_X6Y16_to_ND;
wire[3:0] Tile_X6Y16_to_NF;
wire[7:0] Tile_X6Y16_to_NG;
wire[7:0] Tile_X6Y16_to_NH;
wire[11:0] Tile_X6Y16_to_NI;
wire[3:0] Tile_X6Y16_to_SA;
wire[3:0] Tile_X6Y16_to_SB;
wire[3:0] Tile_X6Y16_to_SC;
wire[3:0] Tile_X6Y16_to_SD;
wire[3:0] Tile_X6Y16_to_SF;
wire[7:0] Tile_X6Y16_to_SG;
wire[7:0] Tile_X6Y16_to_SH;
wire[11:0] Tile_X6Y16_to_SI;
wire[3:0] Tile_X7Y16_to_EA;
wire[3:0] Tile_X7Y16_to_EB;
wire[3:0] Tile_X7Y16_to_EC;
wire[3:0] Tile_X7Y16_to_ED;
wire[3:0] Tile_X7Y16_to_EF;
wire[7:0] Tile_X7Y16_to_EG;
wire[7:0] Tile_X7Y16_to_EH;
wire[11:0] Tile_X7Y16_to_EI;
wire[3:0] Tile_X7Y16_to_WA;
wire[3:0] Tile_X7Y16_to_WB;
wire[3:0] Tile_X7Y16_to_WC;
wire[3:0] Tile_X7Y16_to_WD;
wire[3:0] Tile_X7Y16_to_WF;
wire[7:0] Tile_X7Y16_to_WG;
wire[7:0] Tile_X7Y16_to_WH;
wire[11:0] Tile_X7Y16_to_WI;
wire[3:0] Tile_X7Y16_to_NA;
wire[3:0] Tile_X7Y16_to_NB;
wire[3:0] Tile_X7Y16_to_NC;
wire[3:0] Tile_X7Y16_to_ND;
wire[3:0] Tile_X7Y16_to_NF;
wire[7:0] Tile_X7Y16_to_NG;
wire[7:0] Tile_X7Y16_to_NH;
wire[11:0] Tile_X7Y16_to_NI;
wire[3:0] Tile_X7Y16_to_SA;
wire[3:0] Tile_X7Y16_to_SB;
wire[3:0] Tile_X7Y16_to_SC;
wire[3:0] Tile_X7Y16_to_SD;
wire[3:0] Tile_X7Y16_to_SF;
wire[7:0] Tile_X7Y16_to_SG;
wire[7:0] Tile_X7Y16_to_SH;
wire[11:0] Tile_X7Y16_to_SI;
wire[3:0] Tile_X8Y16_to_WA;
wire[3:0] Tile_X8Y16_to_WB;
wire[3:0] Tile_X8Y16_to_WC;
wire[3:0] Tile_X8Y16_to_WD;
wire[3:0] Tile_X8Y16_to_WF;
wire[7:0] Tile_X8Y16_to_WG;
wire[7:0] Tile_X8Y16_to_WH;
wire[11:0] Tile_X8Y16_to_WI;
wire[3:0] Tile_X8Y16_to_NA;
wire[3:0] Tile_X8Y16_to_NB;
wire[3:0] Tile_X8Y16_to_NC;
wire[3:0] Tile_X8Y16_to_ND;
wire[3:0] Tile_X8Y16_to_NF;
wire[7:0] Tile_X8Y16_to_NG;
wire[7:0] Tile_X8Y16_to_NH;
wire[11:0] Tile_X8Y16_to_NI;
wire[3:0] Tile_X8Y16_to_SA;
wire[3:0] Tile_X8Y16_to_SB;
wire[3:0] Tile_X8Y16_to_SC;
wire[3:0] Tile_X8Y16_to_SD;
wire[3:0] Tile_X8Y16_to_SF;
wire[7:0] Tile_X8Y16_to_SG;
wire[7:0] Tile_X8Y16_to_SH;
wire[11:0] Tile_X8Y16_to_SI;
wire[1:0] Tile_X9Y16_to_EA_1s;
wire[1:0] Tile_X9Y16_to_EB_1s;
wire[1:0] Tile_X9Y16_to_EC_1s;
wire[1:0] Tile_X9Y16_to_ED_1s;
wire[1:0] Tile_X9Y16_to_EF_1s;
wire[1:0] Tile_X9Y16_to_EG_1s;
wire[1:0] Tile_X9Y16_to_EH_1s;
wire[1:0] Tile_X9Y16_to_EI_1s;
wire[1:0] Tile_X9Y16_to_WA_1s;
wire[1:0] Tile_X9Y16_to_WB_1s;
wire[1:0] Tile_X9Y16_to_WC_1s;
wire[1:0] Tile_X9Y16_to_WD_1s;
wire[1:0] Tile_X9Y16_to_WF_1s;
wire[1:0] Tile_X9Y16_to_WG_1s;
wire[1:0] Tile_X9Y16_to_WH_1s;
wire[1:0] Tile_X9Y16_to_WI_1s;
wire[1:0] Tile_X9Y16_to_NA_1s;
wire[1:0] Tile_X9Y16_to_NB_1s;
wire[1:0] Tile_X9Y16_to_NC_1s;
wire[1:0] Tile_X9Y16_to_ND_1s;
wire[1:0] Tile_X9Y16_to_NF_1s;
wire[1:0] Tile_X9Y16_to_NG_1s;
wire[1:0] Tile_X9Y16_to_NH_1s;
wire[1:0] Tile_X9Y16_to_NI_1s;
wire[1:0] Tile_X9Y16_to_SA_1s;
wire[1:0] Tile_X9Y16_to_SB_1s;
wire[1:0] Tile_X9Y16_to_SC_1s;
wire[1:0] Tile_X9Y16_to_SD_1s;
wire[1:0] Tile_X9Y16_to_SF_1s;
wire[1:0] Tile_X9Y16_to_SG_1s;
wire[1:0] Tile_X9Y16_to_SH_1s;
wire[1:0] Tile_X9Y16_to_SI_1s;
wire[1:0] Tile_X10Y16_to_WA_1s;
wire[1:0] Tile_X10Y16_to_WB_1s;
wire[1:0] Tile_X10Y16_to_WC_1s;
wire[1:0] Tile_X10Y16_to_WD_1s;
wire[1:0] Tile_X10Y16_to_WF_1s;
wire[1:0] Tile_X10Y16_to_WG_1s;
wire[1:0] Tile_X10Y16_to_WH_1s;
wire[1:0] Tile_X10Y16_to_WI_1s;
wire[3:0] Tile_X0Y17_to_EA;
wire[3:0] Tile_X0Y17_to_EB;
wire[3:0] Tile_X0Y17_to_EC;
wire[3:0] Tile_X0Y17_to_ED;
wire[3:0] Tile_X0Y17_to_EF;
wire[7:0] Tile_X0Y17_to_EG;
wire[7:0] Tile_X0Y17_to_EH;
wire[11:0] Tile_X0Y17_to_EI;
wire[3:0] Tile_X0Y17_to_NA;
wire[3:0] Tile_X0Y17_to_NB;
wire[3:0] Tile_X0Y17_to_NC;
wire[3:0] Tile_X0Y17_to_ND;
wire[3:0] Tile_X0Y17_to_NF;
wire[7:0] Tile_X0Y17_to_NG;
wire[7:0] Tile_X0Y17_to_NH;
wire[11:0] Tile_X0Y17_to_NI;
wire[3:0] Tile_X0Y17_to_SA;
wire[3:0] Tile_X0Y17_to_SB;
wire[3:0] Tile_X0Y17_to_SC;
wire[3:0] Tile_X0Y17_to_SD;
wire[3:0] Tile_X0Y17_to_SF;
wire[7:0] Tile_X0Y17_to_SG;
wire[7:0] Tile_X0Y17_to_SH;
wire[11:0] Tile_X0Y17_to_SI;
wire[3:0] Tile_X1Y17_to_EA;
wire[3:0] Tile_X1Y17_to_EB;
wire[3:0] Tile_X1Y17_to_EC;
wire[3:0] Tile_X1Y17_to_ED;
wire[3:0] Tile_X1Y17_to_EF;
wire[7:0] Tile_X1Y17_to_EG;
wire[7:0] Tile_X1Y17_to_EH;
wire[11:0] Tile_X1Y17_to_EI;
wire[3:0] Tile_X1Y17_to_WA;
wire[3:0] Tile_X1Y17_to_WB;
wire[3:0] Tile_X1Y17_to_WC;
wire[3:0] Tile_X1Y17_to_WD;
wire[3:0] Tile_X1Y17_to_WF;
wire[7:0] Tile_X1Y17_to_WG;
wire[7:0] Tile_X1Y17_to_WH;
wire[11:0] Tile_X1Y17_to_WI;
wire[3:0] Tile_X1Y17_to_NA;
wire[3:0] Tile_X1Y17_to_NB;
wire[3:0] Tile_X1Y17_to_NC;
wire[3:0] Tile_X1Y17_to_ND;
wire[3:0] Tile_X1Y17_to_NF;
wire[7:0] Tile_X1Y17_to_NG;
wire[7:0] Tile_X1Y17_to_NH;
wire[11:0] Tile_X1Y17_to_NI;
wire[3:0] Tile_X1Y17_to_SA;
wire[3:0] Tile_X1Y17_to_SB;
wire[3:0] Tile_X1Y17_to_SC;
wire[3:0] Tile_X1Y17_to_SD;
wire[3:0] Tile_X1Y17_to_SF;
wire[7:0] Tile_X1Y17_to_SG;
wire[7:0] Tile_X1Y17_to_SH;
wire[11:0] Tile_X1Y17_to_SI;
wire[3:0] Tile_X2Y17_to_EA;
wire[3:0] Tile_X2Y17_to_EB;
wire[3:0] Tile_X2Y17_to_EC;
wire[3:0] Tile_X2Y17_to_ED;
wire[3:0] Tile_X2Y17_to_EF;
wire[7:0] Tile_X2Y17_to_EG;
wire[7:0] Tile_X2Y17_to_EH;
wire[11:0] Tile_X2Y17_to_EI;
wire[3:0] Tile_X2Y17_to_WA;
wire[3:0] Tile_X2Y17_to_WB;
wire[3:0] Tile_X2Y17_to_WC;
wire[3:0] Tile_X2Y17_to_WD;
wire[3:0] Tile_X2Y17_to_WF;
wire[7:0] Tile_X2Y17_to_WG;
wire[7:0] Tile_X2Y17_to_WH;
wire[11:0] Tile_X2Y17_to_WI;
wire[3:0] Tile_X2Y17_to_NA;
wire[3:0] Tile_X2Y17_to_NB;
wire[3:0] Tile_X2Y17_to_NC;
wire[3:0] Tile_X2Y17_to_ND;
wire[3:0] Tile_X2Y17_to_NF;
wire[7:0] Tile_X2Y17_to_NG;
wire[7:0] Tile_X2Y17_to_NH;
wire[11:0] Tile_X2Y17_to_NI;
wire[3:0] Tile_X2Y17_to_SA;
wire[3:0] Tile_X2Y17_to_SB;
wire[3:0] Tile_X2Y17_to_SC;
wire[3:0] Tile_X2Y17_to_SD;
wire[3:0] Tile_X2Y17_to_SF;
wire[7:0] Tile_X2Y17_to_SG;
wire[7:0] Tile_X2Y17_to_SH;
wire[11:0] Tile_X2Y17_to_SI;
wire[3:0] Tile_X3Y17_to_EA;
wire[3:0] Tile_X3Y17_to_EB;
wire[3:0] Tile_X3Y17_to_EC;
wire[3:0] Tile_X3Y17_to_ED;
wire[3:0] Tile_X3Y17_to_EF;
wire[7:0] Tile_X3Y17_to_EG;
wire[7:0] Tile_X3Y17_to_EH;
wire[11:0] Tile_X3Y17_to_EI;
wire[3:0] Tile_X3Y17_to_WA;
wire[3:0] Tile_X3Y17_to_WB;
wire[3:0] Tile_X3Y17_to_WC;
wire[3:0] Tile_X3Y17_to_WD;
wire[3:0] Tile_X3Y17_to_WF;
wire[7:0] Tile_X3Y17_to_WG;
wire[7:0] Tile_X3Y17_to_WH;
wire[11:0] Tile_X3Y17_to_WI;
wire[3:0] Tile_X3Y17_to_NA;
wire[3:0] Tile_X3Y17_to_NB;
wire[3:0] Tile_X3Y17_to_NC;
wire[3:0] Tile_X3Y17_to_ND;
wire[3:0] Tile_X3Y17_to_NF;
wire[7:0] Tile_X3Y17_to_NG;
wire[7:0] Tile_X3Y17_to_NH;
wire[11:0] Tile_X3Y17_to_NI;
wire[3:0] Tile_X3Y17_to_SA;
wire[3:0] Tile_X3Y17_to_SB;
wire[3:0] Tile_X3Y17_to_SC;
wire[3:0] Tile_X3Y17_to_SD;
wire[3:0] Tile_X3Y17_to_SF;
wire[7:0] Tile_X3Y17_to_SG;
wire[7:0] Tile_X3Y17_to_SH;
wire[11:0] Tile_X3Y17_to_SI;
wire[3:0] Tile_X4Y17_to_EA;
wire[3:0] Tile_X4Y17_to_EB;
wire[3:0] Tile_X4Y17_to_EC;
wire[3:0] Tile_X4Y17_to_ED;
wire[3:0] Tile_X4Y17_to_EF;
wire[7:0] Tile_X4Y17_to_EG;
wire[7:0] Tile_X4Y17_to_EH;
wire[11:0] Tile_X4Y17_to_EI;
wire[3:0] Tile_X4Y17_to_WA;
wire[3:0] Tile_X4Y17_to_WB;
wire[3:0] Tile_X4Y17_to_WC;
wire[3:0] Tile_X4Y17_to_WD;
wire[3:0] Tile_X4Y17_to_WF;
wire[7:0] Tile_X4Y17_to_WG;
wire[7:0] Tile_X4Y17_to_WH;
wire[11:0] Tile_X4Y17_to_WI;
wire[3:0] Tile_X4Y17_to_NA;
wire[3:0] Tile_X4Y17_to_NB;
wire[3:0] Tile_X4Y17_to_NC;
wire[3:0] Tile_X4Y17_to_ND;
wire[3:0] Tile_X4Y17_to_NF;
wire[7:0] Tile_X4Y17_to_NG;
wire[7:0] Tile_X4Y17_to_NH;
wire[11:0] Tile_X4Y17_to_NI;
wire[3:0] Tile_X4Y17_to_SA;
wire[3:0] Tile_X4Y17_to_SB;
wire[3:0] Tile_X4Y17_to_SC;
wire[3:0] Tile_X4Y17_to_SD;
wire[3:0] Tile_X4Y17_to_SF;
wire[7:0] Tile_X4Y17_to_SG;
wire[7:0] Tile_X4Y17_to_SH;
wire[11:0] Tile_X4Y17_to_SI;
wire[3:0] Tile_X5Y17_to_EA;
wire[3:0] Tile_X5Y17_to_EB;
wire[3:0] Tile_X5Y17_to_EC;
wire[3:0] Tile_X5Y17_to_ED;
wire[3:0] Tile_X5Y17_to_EF;
wire[7:0] Tile_X5Y17_to_EG;
wire[7:0] Tile_X5Y17_to_EH;
wire[11:0] Tile_X5Y17_to_EI;
wire[3:0] Tile_X5Y17_to_WA;
wire[3:0] Tile_X5Y17_to_WB;
wire[3:0] Tile_X5Y17_to_WC;
wire[3:0] Tile_X5Y17_to_WD;
wire[3:0] Tile_X5Y17_to_WF;
wire[7:0] Tile_X5Y17_to_WG;
wire[7:0] Tile_X5Y17_to_WH;
wire[11:0] Tile_X5Y17_to_WI;
wire[3:0] Tile_X5Y17_to_NA;
wire[3:0] Tile_X5Y17_to_NB;
wire[3:0] Tile_X5Y17_to_NC;
wire[3:0] Tile_X5Y17_to_ND;
wire[3:0] Tile_X5Y17_to_NF;
wire[7:0] Tile_X5Y17_to_NG;
wire[7:0] Tile_X5Y17_to_NH;
wire[11:0] Tile_X5Y17_to_NI;
wire[3:0] Tile_X5Y17_to_SA;
wire[3:0] Tile_X5Y17_to_SB;
wire[3:0] Tile_X5Y17_to_SC;
wire[3:0] Tile_X5Y17_to_SD;
wire[3:0] Tile_X5Y17_to_SF;
wire[7:0] Tile_X5Y17_to_SG;
wire[7:0] Tile_X5Y17_to_SH;
wire[11:0] Tile_X5Y17_to_SI;
wire[3:0] Tile_X6Y17_to_EA;
wire[3:0] Tile_X6Y17_to_EB;
wire[3:0] Tile_X6Y17_to_EC;
wire[3:0] Tile_X6Y17_to_ED;
wire[3:0] Tile_X6Y17_to_EF;
wire[7:0] Tile_X6Y17_to_EG;
wire[7:0] Tile_X6Y17_to_EH;
wire[11:0] Tile_X6Y17_to_EI;
wire[3:0] Tile_X6Y17_to_WA;
wire[3:0] Tile_X6Y17_to_WB;
wire[3:0] Tile_X6Y17_to_WC;
wire[3:0] Tile_X6Y17_to_WD;
wire[3:0] Tile_X6Y17_to_WF;
wire[7:0] Tile_X6Y17_to_WG;
wire[7:0] Tile_X6Y17_to_WH;
wire[11:0] Tile_X6Y17_to_WI;
wire[3:0] Tile_X6Y17_to_NA;
wire[3:0] Tile_X6Y17_to_NB;
wire[3:0] Tile_X6Y17_to_NC;
wire[3:0] Tile_X6Y17_to_ND;
wire[3:0] Tile_X6Y17_to_NF;
wire[7:0] Tile_X6Y17_to_NG;
wire[7:0] Tile_X6Y17_to_NH;
wire[11:0] Tile_X6Y17_to_NI;
wire[3:0] Tile_X6Y17_to_SA;
wire[3:0] Tile_X6Y17_to_SB;
wire[3:0] Tile_X6Y17_to_SC;
wire[3:0] Tile_X6Y17_to_SD;
wire[3:0] Tile_X6Y17_to_SF;
wire[7:0] Tile_X6Y17_to_SG;
wire[7:0] Tile_X6Y17_to_SH;
wire[11:0] Tile_X6Y17_to_SI;
wire[3:0] Tile_X7Y17_to_EA;
wire[3:0] Tile_X7Y17_to_EB;
wire[3:0] Tile_X7Y17_to_EC;
wire[3:0] Tile_X7Y17_to_ED;
wire[3:0] Tile_X7Y17_to_EF;
wire[7:0] Tile_X7Y17_to_EG;
wire[7:0] Tile_X7Y17_to_EH;
wire[11:0] Tile_X7Y17_to_EI;
wire[3:0] Tile_X7Y17_to_WA;
wire[3:0] Tile_X7Y17_to_WB;
wire[3:0] Tile_X7Y17_to_WC;
wire[3:0] Tile_X7Y17_to_WD;
wire[3:0] Tile_X7Y17_to_WF;
wire[7:0] Tile_X7Y17_to_WG;
wire[7:0] Tile_X7Y17_to_WH;
wire[11:0] Tile_X7Y17_to_WI;
wire[3:0] Tile_X7Y17_to_NA;
wire[3:0] Tile_X7Y17_to_NB;
wire[3:0] Tile_X7Y17_to_NC;
wire[3:0] Tile_X7Y17_to_ND;
wire[3:0] Tile_X7Y17_to_NF;
wire[7:0] Tile_X7Y17_to_NG;
wire[7:0] Tile_X7Y17_to_NH;
wire[11:0] Tile_X7Y17_to_NI;
wire[3:0] Tile_X7Y17_to_SA;
wire[3:0] Tile_X7Y17_to_SB;
wire[3:0] Tile_X7Y17_to_SC;
wire[3:0] Tile_X7Y17_to_SD;
wire[3:0] Tile_X7Y17_to_SF;
wire[7:0] Tile_X7Y17_to_SG;
wire[7:0] Tile_X7Y17_to_SH;
wire[11:0] Tile_X7Y17_to_SI;
wire[3:0] Tile_X8Y17_to_WA;
wire[3:0] Tile_X8Y17_to_WB;
wire[3:0] Tile_X8Y17_to_WC;
wire[3:0] Tile_X8Y17_to_WD;
wire[3:0] Tile_X8Y17_to_WF;
wire[7:0] Tile_X8Y17_to_WG;
wire[7:0] Tile_X8Y17_to_WH;
wire[11:0] Tile_X8Y17_to_WI;
wire[3:0] Tile_X8Y17_to_NA;
wire[3:0] Tile_X8Y17_to_NB;
wire[3:0] Tile_X8Y17_to_NC;
wire[3:0] Tile_X8Y17_to_ND;
wire[3:0] Tile_X8Y17_to_NF;
wire[7:0] Tile_X8Y17_to_NG;
wire[7:0] Tile_X8Y17_to_NH;
wire[11:0] Tile_X8Y17_to_NI;
wire[3:0] Tile_X8Y17_to_SA;
wire[3:0] Tile_X8Y17_to_SB;
wire[3:0] Tile_X8Y17_to_SC;
wire[3:0] Tile_X8Y17_to_SD;
wire[3:0] Tile_X8Y17_to_SF;
wire[7:0] Tile_X8Y17_to_SG;
wire[7:0] Tile_X8Y17_to_SH;
wire[11:0] Tile_X8Y17_to_SI;
wire[1:0] Tile_X9Y17_to_EA_1s;
wire[1:0] Tile_X9Y17_to_EB_1s;
wire[1:0] Tile_X9Y17_to_EC_1s;
wire[1:0] Tile_X9Y17_to_ED_1s;
wire[1:0] Tile_X9Y17_to_EF_1s;
wire[1:0] Tile_X9Y17_to_EG_1s;
wire[1:0] Tile_X9Y17_to_EH_1s;
wire[1:0] Tile_X9Y17_to_EI_1s;
wire[1:0] Tile_X9Y17_to_WA_1s;
wire[1:0] Tile_X9Y17_to_WB_1s;
wire[1:0] Tile_X9Y17_to_WC_1s;
wire[1:0] Tile_X9Y17_to_WD_1s;
wire[1:0] Tile_X9Y17_to_WF_1s;
wire[1:0] Tile_X9Y17_to_WG_1s;
wire[1:0] Tile_X9Y17_to_WH_1s;
wire[1:0] Tile_X9Y17_to_WI_1s;
wire[1:0] Tile_X9Y17_to_NA_1s;
wire[1:0] Tile_X9Y17_to_NB_1s;
wire[1:0] Tile_X9Y17_to_NC_1s;
wire[1:0] Tile_X9Y17_to_ND_1s;
wire[1:0] Tile_X9Y17_to_NF_1s;
wire[1:0] Tile_X9Y17_to_NG_1s;
wire[1:0] Tile_X9Y17_to_NH_1s;
wire[1:0] Tile_X9Y17_to_NI_1s;
wire[1:0] Tile_X9Y17_to_SA_1s;
wire[1:0] Tile_X9Y17_to_SB_1s;
wire[1:0] Tile_X9Y17_to_SC_1s;
wire[1:0] Tile_X9Y17_to_SD_1s;
wire[1:0] Tile_X9Y17_to_SF_1s;
wire[1:0] Tile_X9Y17_to_SG_1s;
wire[1:0] Tile_X9Y17_to_SH_1s;
wire[1:0] Tile_X9Y17_to_SI_1s;
wire[1:0] Tile_X10Y17_to_WA_1s;
wire[1:0] Tile_X10Y17_to_WB_1s;
wire[1:0] Tile_X10Y17_to_WC_1s;
wire[1:0] Tile_X10Y17_to_WD_1s;
wire[1:0] Tile_X10Y17_to_WF_1s;
wire[1:0] Tile_X10Y17_to_WG_1s;
wire[1:0] Tile_X10Y17_to_WH_1s;
wire[1:0] Tile_X10Y17_to_WI_1s;
wire[3:0] Tile_X0Y18_to_EA;
wire[3:0] Tile_X0Y18_to_EB;
wire[3:0] Tile_X0Y18_to_EC;
wire[3:0] Tile_X0Y18_to_ED;
wire[3:0] Tile_X0Y18_to_EF;
wire[7:0] Tile_X0Y18_to_EG;
wire[7:0] Tile_X0Y18_to_EH;
wire[11:0] Tile_X0Y18_to_EI;
wire[3:0] Tile_X0Y18_to_NA;
wire[3:0] Tile_X0Y18_to_NB;
wire[3:0] Tile_X0Y18_to_NC;
wire[3:0] Tile_X0Y18_to_ND;
wire[3:0] Tile_X0Y18_to_NF;
wire[7:0] Tile_X0Y18_to_NG;
wire[7:0] Tile_X0Y18_to_NH;
wire[11:0] Tile_X0Y18_to_NI;
wire[3:0] Tile_X0Y18_to_SA;
wire[3:0] Tile_X0Y18_to_SB;
wire[3:0] Tile_X0Y18_to_SC;
wire[3:0] Tile_X0Y18_to_SD;
wire[3:0] Tile_X0Y18_to_SF;
wire[7:0] Tile_X0Y18_to_SG;
wire[7:0] Tile_X0Y18_to_SH;
wire[11:0] Tile_X0Y18_to_SI;
wire[3:0] Tile_X1Y18_to_EA;
wire[3:0] Tile_X1Y18_to_EB;
wire[3:0] Tile_X1Y18_to_EC;
wire[3:0] Tile_X1Y18_to_ED;
wire[3:0] Tile_X1Y18_to_EF;
wire[7:0] Tile_X1Y18_to_EG;
wire[7:0] Tile_X1Y18_to_EH;
wire[11:0] Tile_X1Y18_to_EI;
wire[3:0] Tile_X1Y18_to_WA;
wire[3:0] Tile_X1Y18_to_WB;
wire[3:0] Tile_X1Y18_to_WC;
wire[3:0] Tile_X1Y18_to_WD;
wire[3:0] Tile_X1Y18_to_WF;
wire[7:0] Tile_X1Y18_to_WG;
wire[7:0] Tile_X1Y18_to_WH;
wire[11:0] Tile_X1Y18_to_WI;
wire[3:0] Tile_X1Y18_to_NA;
wire[3:0] Tile_X1Y18_to_NB;
wire[3:0] Tile_X1Y18_to_NC;
wire[3:0] Tile_X1Y18_to_ND;
wire[3:0] Tile_X1Y18_to_NF;
wire[7:0] Tile_X1Y18_to_NG;
wire[7:0] Tile_X1Y18_to_NH;
wire[11:0] Tile_X1Y18_to_NI;
wire[3:0] Tile_X1Y18_to_SA;
wire[3:0] Tile_X1Y18_to_SB;
wire[3:0] Tile_X1Y18_to_SC;
wire[3:0] Tile_X1Y18_to_SD;
wire[3:0] Tile_X1Y18_to_SF;
wire[7:0] Tile_X1Y18_to_SG;
wire[7:0] Tile_X1Y18_to_SH;
wire[11:0] Tile_X1Y18_to_SI;
wire[3:0] Tile_X2Y18_to_EA;
wire[3:0] Tile_X2Y18_to_EB;
wire[3:0] Tile_X2Y18_to_EC;
wire[3:0] Tile_X2Y18_to_ED;
wire[3:0] Tile_X2Y18_to_EF;
wire[7:0] Tile_X2Y18_to_EG;
wire[7:0] Tile_X2Y18_to_EH;
wire[11:0] Tile_X2Y18_to_EI;
wire[3:0] Tile_X2Y18_to_WA;
wire[3:0] Tile_X2Y18_to_WB;
wire[3:0] Tile_X2Y18_to_WC;
wire[3:0] Tile_X2Y18_to_WD;
wire[3:0] Tile_X2Y18_to_WF;
wire[7:0] Tile_X2Y18_to_WG;
wire[7:0] Tile_X2Y18_to_WH;
wire[11:0] Tile_X2Y18_to_WI;
wire[3:0] Tile_X2Y18_to_NA;
wire[3:0] Tile_X2Y18_to_NB;
wire[3:0] Tile_X2Y18_to_NC;
wire[3:0] Tile_X2Y18_to_ND;
wire[3:0] Tile_X2Y18_to_NF;
wire[7:0] Tile_X2Y18_to_NG;
wire[7:0] Tile_X2Y18_to_NH;
wire[11:0] Tile_X2Y18_to_NI;
wire[3:0] Tile_X2Y18_to_SA;
wire[3:0] Tile_X2Y18_to_SB;
wire[3:0] Tile_X2Y18_to_SC;
wire[3:0] Tile_X2Y18_to_SD;
wire[3:0] Tile_X2Y18_to_SF;
wire[7:0] Tile_X2Y18_to_SG;
wire[7:0] Tile_X2Y18_to_SH;
wire[11:0] Tile_X2Y18_to_SI;
wire[3:0] Tile_X3Y18_to_EA;
wire[3:0] Tile_X3Y18_to_EB;
wire[3:0] Tile_X3Y18_to_EC;
wire[3:0] Tile_X3Y18_to_ED;
wire[3:0] Tile_X3Y18_to_EF;
wire[7:0] Tile_X3Y18_to_EG;
wire[7:0] Tile_X3Y18_to_EH;
wire[11:0] Tile_X3Y18_to_EI;
wire[3:0] Tile_X3Y18_to_WA;
wire[3:0] Tile_X3Y18_to_WB;
wire[3:0] Tile_X3Y18_to_WC;
wire[3:0] Tile_X3Y18_to_WD;
wire[3:0] Tile_X3Y18_to_WF;
wire[7:0] Tile_X3Y18_to_WG;
wire[7:0] Tile_X3Y18_to_WH;
wire[11:0] Tile_X3Y18_to_WI;
wire[3:0] Tile_X3Y18_to_NA;
wire[3:0] Tile_X3Y18_to_NB;
wire[3:0] Tile_X3Y18_to_NC;
wire[3:0] Tile_X3Y18_to_ND;
wire[3:0] Tile_X3Y18_to_NF;
wire[7:0] Tile_X3Y18_to_NG;
wire[7:0] Tile_X3Y18_to_NH;
wire[11:0] Tile_X3Y18_to_NI;
wire[3:0] Tile_X3Y18_to_SA;
wire[3:0] Tile_X3Y18_to_SB;
wire[3:0] Tile_X3Y18_to_SC;
wire[3:0] Tile_X3Y18_to_SD;
wire[3:0] Tile_X3Y18_to_SF;
wire[7:0] Tile_X3Y18_to_SG;
wire[7:0] Tile_X3Y18_to_SH;
wire[11:0] Tile_X3Y18_to_SI;
wire[3:0] Tile_X4Y18_to_EA;
wire[3:0] Tile_X4Y18_to_EB;
wire[3:0] Tile_X4Y18_to_EC;
wire[3:0] Tile_X4Y18_to_ED;
wire[3:0] Tile_X4Y18_to_EF;
wire[7:0] Tile_X4Y18_to_EG;
wire[7:0] Tile_X4Y18_to_EH;
wire[11:0] Tile_X4Y18_to_EI;
wire[3:0] Tile_X4Y18_to_WA;
wire[3:0] Tile_X4Y18_to_WB;
wire[3:0] Tile_X4Y18_to_WC;
wire[3:0] Tile_X4Y18_to_WD;
wire[3:0] Tile_X4Y18_to_WF;
wire[7:0] Tile_X4Y18_to_WG;
wire[7:0] Tile_X4Y18_to_WH;
wire[11:0] Tile_X4Y18_to_WI;
wire[3:0] Tile_X4Y18_to_NA;
wire[3:0] Tile_X4Y18_to_NB;
wire[3:0] Tile_X4Y18_to_NC;
wire[3:0] Tile_X4Y18_to_ND;
wire[3:0] Tile_X4Y18_to_NF;
wire[7:0] Tile_X4Y18_to_NG;
wire[7:0] Tile_X4Y18_to_NH;
wire[11:0] Tile_X4Y18_to_NI;
wire[3:0] Tile_X4Y18_to_SA;
wire[3:0] Tile_X4Y18_to_SB;
wire[3:0] Tile_X4Y18_to_SC;
wire[3:0] Tile_X4Y18_to_SD;
wire[3:0] Tile_X4Y18_to_SF;
wire[7:0] Tile_X4Y18_to_SG;
wire[7:0] Tile_X4Y18_to_SH;
wire[11:0] Tile_X4Y18_to_SI;
wire[3:0] Tile_X5Y18_to_EA;
wire[3:0] Tile_X5Y18_to_EB;
wire[3:0] Tile_X5Y18_to_EC;
wire[3:0] Tile_X5Y18_to_ED;
wire[3:0] Tile_X5Y18_to_EF;
wire[7:0] Tile_X5Y18_to_EG;
wire[7:0] Tile_X5Y18_to_EH;
wire[11:0] Tile_X5Y18_to_EI;
wire[3:0] Tile_X5Y18_to_WA;
wire[3:0] Tile_X5Y18_to_WB;
wire[3:0] Tile_X5Y18_to_WC;
wire[3:0] Tile_X5Y18_to_WD;
wire[3:0] Tile_X5Y18_to_WF;
wire[7:0] Tile_X5Y18_to_WG;
wire[7:0] Tile_X5Y18_to_WH;
wire[11:0] Tile_X5Y18_to_WI;
wire[3:0] Tile_X5Y18_to_NA;
wire[3:0] Tile_X5Y18_to_NB;
wire[3:0] Tile_X5Y18_to_NC;
wire[3:0] Tile_X5Y18_to_ND;
wire[3:0] Tile_X5Y18_to_NF;
wire[7:0] Tile_X5Y18_to_NG;
wire[7:0] Tile_X5Y18_to_NH;
wire[11:0] Tile_X5Y18_to_NI;
wire[3:0] Tile_X5Y18_to_SA;
wire[3:0] Tile_X5Y18_to_SB;
wire[3:0] Tile_X5Y18_to_SC;
wire[3:0] Tile_X5Y18_to_SD;
wire[3:0] Tile_X5Y18_to_SF;
wire[7:0] Tile_X5Y18_to_SG;
wire[7:0] Tile_X5Y18_to_SH;
wire[11:0] Tile_X5Y18_to_SI;
wire[3:0] Tile_X6Y18_to_EA;
wire[3:0] Tile_X6Y18_to_EB;
wire[3:0] Tile_X6Y18_to_EC;
wire[3:0] Tile_X6Y18_to_ED;
wire[3:0] Tile_X6Y18_to_EF;
wire[7:0] Tile_X6Y18_to_EG;
wire[7:0] Tile_X6Y18_to_EH;
wire[11:0] Tile_X6Y18_to_EI;
wire[3:0] Tile_X6Y18_to_WA;
wire[3:0] Tile_X6Y18_to_WB;
wire[3:0] Tile_X6Y18_to_WC;
wire[3:0] Tile_X6Y18_to_WD;
wire[3:0] Tile_X6Y18_to_WF;
wire[7:0] Tile_X6Y18_to_WG;
wire[7:0] Tile_X6Y18_to_WH;
wire[11:0] Tile_X6Y18_to_WI;
wire[3:0] Tile_X6Y18_to_NA;
wire[3:0] Tile_X6Y18_to_NB;
wire[3:0] Tile_X6Y18_to_NC;
wire[3:0] Tile_X6Y18_to_ND;
wire[3:0] Tile_X6Y18_to_NF;
wire[7:0] Tile_X6Y18_to_NG;
wire[7:0] Tile_X6Y18_to_NH;
wire[11:0] Tile_X6Y18_to_NI;
wire[3:0] Tile_X6Y18_to_SA;
wire[3:0] Tile_X6Y18_to_SB;
wire[3:0] Tile_X6Y18_to_SC;
wire[3:0] Tile_X6Y18_to_SD;
wire[3:0] Tile_X6Y18_to_SF;
wire[7:0] Tile_X6Y18_to_SG;
wire[7:0] Tile_X6Y18_to_SH;
wire[11:0] Tile_X6Y18_to_SI;
wire[3:0] Tile_X7Y18_to_EA;
wire[3:0] Tile_X7Y18_to_EB;
wire[3:0] Tile_X7Y18_to_EC;
wire[3:0] Tile_X7Y18_to_ED;
wire[3:0] Tile_X7Y18_to_EF;
wire[7:0] Tile_X7Y18_to_EG;
wire[7:0] Tile_X7Y18_to_EH;
wire[11:0] Tile_X7Y18_to_EI;
wire[3:0] Tile_X7Y18_to_WA;
wire[3:0] Tile_X7Y18_to_WB;
wire[3:0] Tile_X7Y18_to_WC;
wire[3:0] Tile_X7Y18_to_WD;
wire[3:0] Tile_X7Y18_to_WF;
wire[7:0] Tile_X7Y18_to_WG;
wire[7:0] Tile_X7Y18_to_WH;
wire[11:0] Tile_X7Y18_to_WI;
wire[3:0] Tile_X7Y18_to_NA;
wire[3:0] Tile_X7Y18_to_NB;
wire[3:0] Tile_X7Y18_to_NC;
wire[3:0] Tile_X7Y18_to_ND;
wire[3:0] Tile_X7Y18_to_NF;
wire[7:0] Tile_X7Y18_to_NG;
wire[7:0] Tile_X7Y18_to_NH;
wire[11:0] Tile_X7Y18_to_NI;
wire[3:0] Tile_X7Y18_to_SA;
wire[3:0] Tile_X7Y18_to_SB;
wire[3:0] Tile_X7Y18_to_SC;
wire[3:0] Tile_X7Y18_to_SD;
wire[3:0] Tile_X7Y18_to_SF;
wire[7:0] Tile_X7Y18_to_SG;
wire[7:0] Tile_X7Y18_to_SH;
wire[11:0] Tile_X7Y18_to_SI;
wire[3:0] Tile_X8Y18_to_WA;
wire[3:0] Tile_X8Y18_to_WB;
wire[3:0] Tile_X8Y18_to_WC;
wire[3:0] Tile_X8Y18_to_WD;
wire[3:0] Tile_X8Y18_to_WF;
wire[7:0] Tile_X8Y18_to_WG;
wire[7:0] Tile_X8Y18_to_WH;
wire[11:0] Tile_X8Y18_to_WI;
wire[3:0] Tile_X8Y18_to_NA;
wire[3:0] Tile_X8Y18_to_NB;
wire[3:0] Tile_X8Y18_to_NC;
wire[3:0] Tile_X8Y18_to_ND;
wire[3:0] Tile_X8Y18_to_NF;
wire[7:0] Tile_X8Y18_to_NG;
wire[7:0] Tile_X8Y18_to_NH;
wire[11:0] Tile_X8Y18_to_NI;
wire[3:0] Tile_X8Y18_to_SA;
wire[3:0] Tile_X8Y18_to_SB;
wire[3:0] Tile_X8Y18_to_SC;
wire[3:0] Tile_X8Y18_to_SD;
wire[3:0] Tile_X8Y18_to_SF;
wire[7:0] Tile_X8Y18_to_SG;
wire[7:0] Tile_X8Y18_to_SH;
wire[11:0] Tile_X8Y18_to_SI;
wire[1:0] Tile_X9Y18_to_EA_1s;
wire[1:0] Tile_X9Y18_to_EB_1s;
wire[1:0] Tile_X9Y18_to_EC_1s;
wire[1:0] Tile_X9Y18_to_ED_1s;
wire[1:0] Tile_X9Y18_to_EF_1s;
wire[1:0] Tile_X9Y18_to_EG_1s;
wire[1:0] Tile_X9Y18_to_EH_1s;
wire[1:0] Tile_X9Y18_to_EI_1s;
wire[1:0] Tile_X9Y18_to_WA_1s;
wire[1:0] Tile_X9Y18_to_WB_1s;
wire[1:0] Tile_X9Y18_to_WC_1s;
wire[1:0] Tile_X9Y18_to_WD_1s;
wire[1:0] Tile_X9Y18_to_WF_1s;
wire[1:0] Tile_X9Y18_to_WG_1s;
wire[1:0] Tile_X9Y18_to_WH_1s;
wire[1:0] Tile_X9Y18_to_WI_1s;
wire[1:0] Tile_X9Y18_to_NA_1s;
wire[1:0] Tile_X9Y18_to_NB_1s;
wire[1:0] Tile_X9Y18_to_NC_1s;
wire[1:0] Tile_X9Y18_to_ND_1s;
wire[1:0] Tile_X9Y18_to_NF_1s;
wire[1:0] Tile_X9Y18_to_NG_1s;
wire[1:0] Tile_X9Y18_to_NH_1s;
wire[1:0] Tile_X9Y18_to_NI_1s;
wire[1:0] Tile_X9Y18_to_SA_1s;
wire[1:0] Tile_X9Y18_to_SB_1s;
wire[1:0] Tile_X9Y18_to_SC_1s;
wire[1:0] Tile_X9Y18_to_SD_1s;
wire[1:0] Tile_X9Y18_to_SF_1s;
wire[1:0] Tile_X9Y18_to_SG_1s;
wire[1:0] Tile_X9Y18_to_SH_1s;
wire[1:0] Tile_X9Y18_to_SI_1s;
wire[1:0] Tile_X10Y18_to_WA_1s;
wire[1:0] Tile_X10Y18_to_WB_1s;
wire[1:0] Tile_X10Y18_to_WC_1s;
wire[1:0] Tile_X10Y18_to_WD_1s;
wire[1:0] Tile_X10Y18_to_WF_1s;
wire[1:0] Tile_X10Y18_to_WG_1s;
wire[1:0] Tile_X10Y18_to_WH_1s;
wire[1:0] Tile_X10Y18_to_WI_1s;
wire[3:0] Tile_X0Y19_to_EA;
wire[3:0] Tile_X0Y19_to_EB;
wire[3:0] Tile_X0Y19_to_EC;
wire[3:0] Tile_X0Y19_to_ED;
wire[3:0] Tile_X0Y19_to_EF;
wire[7:0] Tile_X0Y19_to_EG;
wire[7:0] Tile_X0Y19_to_EH;
wire[11:0] Tile_X0Y19_to_EI;
wire[3:0] Tile_X0Y19_to_NA;
wire[3:0] Tile_X0Y19_to_NB;
wire[3:0] Tile_X0Y19_to_NC;
wire[3:0] Tile_X0Y19_to_ND;
wire[3:0] Tile_X0Y19_to_NF;
wire[7:0] Tile_X0Y19_to_NG;
wire[7:0] Tile_X0Y19_to_NH;
wire[11:0] Tile_X0Y19_to_NI;
wire[3:0] Tile_X0Y19_to_SA;
wire[3:0] Tile_X0Y19_to_SB;
wire[3:0] Tile_X0Y19_to_SC;
wire[3:0] Tile_X0Y19_to_SD;
wire[3:0] Tile_X0Y19_to_SF;
wire[7:0] Tile_X0Y19_to_SG;
wire[7:0] Tile_X0Y19_to_SH;
wire[11:0] Tile_X0Y19_to_SI;
wire[3:0] Tile_X1Y19_to_EA;
wire[3:0] Tile_X1Y19_to_EB;
wire[3:0] Tile_X1Y19_to_EC;
wire[3:0] Tile_X1Y19_to_ED;
wire[3:0] Tile_X1Y19_to_EF;
wire[7:0] Tile_X1Y19_to_EG;
wire[7:0] Tile_X1Y19_to_EH;
wire[11:0] Tile_X1Y19_to_EI;
wire[3:0] Tile_X1Y19_to_WA;
wire[3:0] Tile_X1Y19_to_WB;
wire[3:0] Tile_X1Y19_to_WC;
wire[3:0] Tile_X1Y19_to_WD;
wire[3:0] Tile_X1Y19_to_WF;
wire[7:0] Tile_X1Y19_to_WG;
wire[7:0] Tile_X1Y19_to_WH;
wire[11:0] Tile_X1Y19_to_WI;
wire[3:0] Tile_X1Y19_to_NA;
wire[3:0] Tile_X1Y19_to_NB;
wire[3:0] Tile_X1Y19_to_NC;
wire[3:0] Tile_X1Y19_to_ND;
wire[3:0] Tile_X1Y19_to_NF;
wire[7:0] Tile_X1Y19_to_NG;
wire[7:0] Tile_X1Y19_to_NH;
wire[11:0] Tile_X1Y19_to_NI;
wire[3:0] Tile_X1Y19_to_SA;
wire[3:0] Tile_X1Y19_to_SB;
wire[3:0] Tile_X1Y19_to_SC;
wire[3:0] Tile_X1Y19_to_SD;
wire[3:0] Tile_X1Y19_to_SF;
wire[7:0] Tile_X1Y19_to_SG;
wire[7:0] Tile_X1Y19_to_SH;
wire[11:0] Tile_X1Y19_to_SI;
wire[3:0] Tile_X2Y19_to_EA;
wire[3:0] Tile_X2Y19_to_EB;
wire[3:0] Tile_X2Y19_to_EC;
wire[3:0] Tile_X2Y19_to_ED;
wire[3:0] Tile_X2Y19_to_EF;
wire[7:0] Tile_X2Y19_to_EG;
wire[7:0] Tile_X2Y19_to_EH;
wire[11:0] Tile_X2Y19_to_EI;
wire[3:0] Tile_X2Y19_to_WA;
wire[3:0] Tile_X2Y19_to_WB;
wire[3:0] Tile_X2Y19_to_WC;
wire[3:0] Tile_X2Y19_to_WD;
wire[3:0] Tile_X2Y19_to_WF;
wire[7:0] Tile_X2Y19_to_WG;
wire[7:0] Tile_X2Y19_to_WH;
wire[11:0] Tile_X2Y19_to_WI;
wire[3:0] Tile_X2Y19_to_NA;
wire[3:0] Tile_X2Y19_to_NB;
wire[3:0] Tile_X2Y19_to_NC;
wire[3:0] Tile_X2Y19_to_ND;
wire[3:0] Tile_X2Y19_to_NF;
wire[7:0] Tile_X2Y19_to_NG;
wire[7:0] Tile_X2Y19_to_NH;
wire[11:0] Tile_X2Y19_to_NI;
wire[3:0] Tile_X2Y19_to_SA;
wire[3:0] Tile_X2Y19_to_SB;
wire[3:0] Tile_X2Y19_to_SC;
wire[3:0] Tile_X2Y19_to_SD;
wire[3:0] Tile_X2Y19_to_SF;
wire[7:0] Tile_X2Y19_to_SG;
wire[7:0] Tile_X2Y19_to_SH;
wire[11:0] Tile_X2Y19_to_SI;
wire[3:0] Tile_X3Y19_to_EA;
wire[3:0] Tile_X3Y19_to_EB;
wire[3:0] Tile_X3Y19_to_EC;
wire[3:0] Tile_X3Y19_to_ED;
wire[3:0] Tile_X3Y19_to_EF;
wire[7:0] Tile_X3Y19_to_EG;
wire[7:0] Tile_X3Y19_to_EH;
wire[11:0] Tile_X3Y19_to_EI;
wire[3:0] Tile_X3Y19_to_WA;
wire[3:0] Tile_X3Y19_to_WB;
wire[3:0] Tile_X3Y19_to_WC;
wire[3:0] Tile_X3Y19_to_WD;
wire[3:0] Tile_X3Y19_to_WF;
wire[7:0] Tile_X3Y19_to_WG;
wire[7:0] Tile_X3Y19_to_WH;
wire[11:0] Tile_X3Y19_to_WI;
wire[3:0] Tile_X3Y19_to_NA;
wire[3:0] Tile_X3Y19_to_NB;
wire[3:0] Tile_X3Y19_to_NC;
wire[3:0] Tile_X3Y19_to_ND;
wire[3:0] Tile_X3Y19_to_NF;
wire[7:0] Tile_X3Y19_to_NG;
wire[7:0] Tile_X3Y19_to_NH;
wire[11:0] Tile_X3Y19_to_NI;
wire[3:0] Tile_X3Y19_to_SA;
wire[3:0] Tile_X3Y19_to_SB;
wire[3:0] Tile_X3Y19_to_SC;
wire[3:0] Tile_X3Y19_to_SD;
wire[3:0] Tile_X3Y19_to_SF;
wire[7:0] Tile_X3Y19_to_SG;
wire[7:0] Tile_X3Y19_to_SH;
wire[11:0] Tile_X3Y19_to_SI;
wire[3:0] Tile_X4Y19_to_EA;
wire[3:0] Tile_X4Y19_to_EB;
wire[3:0] Tile_X4Y19_to_EC;
wire[3:0] Tile_X4Y19_to_ED;
wire[3:0] Tile_X4Y19_to_EF;
wire[7:0] Tile_X4Y19_to_EG;
wire[7:0] Tile_X4Y19_to_EH;
wire[11:0] Tile_X4Y19_to_EI;
wire[3:0] Tile_X4Y19_to_WA;
wire[3:0] Tile_X4Y19_to_WB;
wire[3:0] Tile_X4Y19_to_WC;
wire[3:0] Tile_X4Y19_to_WD;
wire[3:0] Tile_X4Y19_to_WF;
wire[7:0] Tile_X4Y19_to_WG;
wire[7:0] Tile_X4Y19_to_WH;
wire[11:0] Tile_X4Y19_to_WI;
wire[3:0] Tile_X4Y19_to_NA;
wire[3:0] Tile_X4Y19_to_NB;
wire[3:0] Tile_X4Y19_to_NC;
wire[3:0] Tile_X4Y19_to_ND;
wire[3:0] Tile_X4Y19_to_NF;
wire[7:0] Tile_X4Y19_to_NG;
wire[7:0] Tile_X4Y19_to_NH;
wire[11:0] Tile_X4Y19_to_NI;
wire[3:0] Tile_X4Y19_to_SA;
wire[3:0] Tile_X4Y19_to_SB;
wire[3:0] Tile_X4Y19_to_SC;
wire[3:0] Tile_X4Y19_to_SD;
wire[3:0] Tile_X4Y19_to_SF;
wire[7:0] Tile_X4Y19_to_SG;
wire[7:0] Tile_X4Y19_to_SH;
wire[11:0] Tile_X4Y19_to_SI;
wire[3:0] Tile_X5Y19_to_EA;
wire[3:0] Tile_X5Y19_to_EB;
wire[3:0] Tile_X5Y19_to_EC;
wire[3:0] Tile_X5Y19_to_ED;
wire[3:0] Tile_X5Y19_to_EF;
wire[7:0] Tile_X5Y19_to_EG;
wire[7:0] Tile_X5Y19_to_EH;
wire[11:0] Tile_X5Y19_to_EI;
wire[3:0] Tile_X5Y19_to_WA;
wire[3:0] Tile_X5Y19_to_WB;
wire[3:0] Tile_X5Y19_to_WC;
wire[3:0] Tile_X5Y19_to_WD;
wire[3:0] Tile_X5Y19_to_WF;
wire[7:0] Tile_X5Y19_to_WG;
wire[7:0] Tile_X5Y19_to_WH;
wire[11:0] Tile_X5Y19_to_WI;
wire[3:0] Tile_X5Y19_to_NA;
wire[3:0] Tile_X5Y19_to_NB;
wire[3:0] Tile_X5Y19_to_NC;
wire[3:0] Tile_X5Y19_to_ND;
wire[3:0] Tile_X5Y19_to_NF;
wire[7:0] Tile_X5Y19_to_NG;
wire[7:0] Tile_X5Y19_to_NH;
wire[11:0] Tile_X5Y19_to_NI;
wire[3:0] Tile_X5Y19_to_SA;
wire[3:0] Tile_X5Y19_to_SB;
wire[3:0] Tile_X5Y19_to_SC;
wire[3:0] Tile_X5Y19_to_SD;
wire[3:0] Tile_X5Y19_to_SF;
wire[7:0] Tile_X5Y19_to_SG;
wire[7:0] Tile_X5Y19_to_SH;
wire[11:0] Tile_X5Y19_to_SI;
wire[3:0] Tile_X6Y19_to_EA;
wire[3:0] Tile_X6Y19_to_EB;
wire[3:0] Tile_X6Y19_to_EC;
wire[3:0] Tile_X6Y19_to_ED;
wire[3:0] Tile_X6Y19_to_EF;
wire[7:0] Tile_X6Y19_to_EG;
wire[7:0] Tile_X6Y19_to_EH;
wire[11:0] Tile_X6Y19_to_EI;
wire[3:0] Tile_X6Y19_to_WA;
wire[3:0] Tile_X6Y19_to_WB;
wire[3:0] Tile_X6Y19_to_WC;
wire[3:0] Tile_X6Y19_to_WD;
wire[3:0] Tile_X6Y19_to_WF;
wire[7:0] Tile_X6Y19_to_WG;
wire[7:0] Tile_X6Y19_to_WH;
wire[11:0] Tile_X6Y19_to_WI;
wire[3:0] Tile_X6Y19_to_NA;
wire[3:0] Tile_X6Y19_to_NB;
wire[3:0] Tile_X6Y19_to_NC;
wire[3:0] Tile_X6Y19_to_ND;
wire[3:0] Tile_X6Y19_to_NF;
wire[7:0] Tile_X6Y19_to_NG;
wire[7:0] Tile_X6Y19_to_NH;
wire[11:0] Tile_X6Y19_to_NI;
wire[3:0] Tile_X6Y19_to_SA;
wire[3:0] Tile_X6Y19_to_SB;
wire[3:0] Tile_X6Y19_to_SC;
wire[3:0] Tile_X6Y19_to_SD;
wire[3:0] Tile_X6Y19_to_SF;
wire[7:0] Tile_X6Y19_to_SG;
wire[7:0] Tile_X6Y19_to_SH;
wire[11:0] Tile_X6Y19_to_SI;
wire[3:0] Tile_X7Y19_to_EA;
wire[3:0] Tile_X7Y19_to_EB;
wire[3:0] Tile_X7Y19_to_EC;
wire[3:0] Tile_X7Y19_to_ED;
wire[3:0] Tile_X7Y19_to_EF;
wire[7:0] Tile_X7Y19_to_EG;
wire[7:0] Tile_X7Y19_to_EH;
wire[11:0] Tile_X7Y19_to_EI;
wire[3:0] Tile_X7Y19_to_WA;
wire[3:0] Tile_X7Y19_to_WB;
wire[3:0] Tile_X7Y19_to_WC;
wire[3:0] Tile_X7Y19_to_WD;
wire[3:0] Tile_X7Y19_to_WF;
wire[7:0] Tile_X7Y19_to_WG;
wire[7:0] Tile_X7Y19_to_WH;
wire[11:0] Tile_X7Y19_to_WI;
wire[3:0] Tile_X7Y19_to_NA;
wire[3:0] Tile_X7Y19_to_NB;
wire[3:0] Tile_X7Y19_to_NC;
wire[3:0] Tile_X7Y19_to_ND;
wire[3:0] Tile_X7Y19_to_NF;
wire[7:0] Tile_X7Y19_to_NG;
wire[7:0] Tile_X7Y19_to_NH;
wire[11:0] Tile_X7Y19_to_NI;
wire[3:0] Tile_X7Y19_to_SA;
wire[3:0] Tile_X7Y19_to_SB;
wire[3:0] Tile_X7Y19_to_SC;
wire[3:0] Tile_X7Y19_to_SD;
wire[3:0] Tile_X7Y19_to_SF;
wire[7:0] Tile_X7Y19_to_SG;
wire[7:0] Tile_X7Y19_to_SH;
wire[11:0] Tile_X7Y19_to_SI;
wire[3:0] Tile_X8Y19_to_WA;
wire[3:0] Tile_X8Y19_to_WB;
wire[3:0] Tile_X8Y19_to_WC;
wire[3:0] Tile_X8Y19_to_WD;
wire[3:0] Tile_X8Y19_to_WF;
wire[7:0] Tile_X8Y19_to_WG;
wire[7:0] Tile_X8Y19_to_WH;
wire[11:0] Tile_X8Y19_to_WI;
wire[3:0] Tile_X8Y19_to_NA;
wire[3:0] Tile_X8Y19_to_NB;
wire[3:0] Tile_X8Y19_to_NC;
wire[3:0] Tile_X8Y19_to_ND;
wire[3:0] Tile_X8Y19_to_NF;
wire[7:0] Tile_X8Y19_to_NG;
wire[7:0] Tile_X8Y19_to_NH;
wire[11:0] Tile_X8Y19_to_NI;
wire[3:0] Tile_X8Y19_to_SA;
wire[3:0] Tile_X8Y19_to_SB;
wire[3:0] Tile_X8Y19_to_SC;
wire[3:0] Tile_X8Y19_to_SD;
wire[3:0] Tile_X8Y19_to_SF;
wire[7:0] Tile_X8Y19_to_SG;
wire[7:0] Tile_X8Y19_to_SH;
wire[11:0] Tile_X8Y19_to_SI;
wire[1:0] Tile_X9Y19_to_EA_1s;
wire[1:0] Tile_X9Y19_to_EB_1s;
wire[1:0] Tile_X9Y19_to_EC_1s;
wire[1:0] Tile_X9Y19_to_ED_1s;
wire[1:0] Tile_X9Y19_to_EF_1s;
wire[1:0] Tile_X9Y19_to_EG_1s;
wire[1:0] Tile_X9Y19_to_EH_1s;
wire[1:0] Tile_X9Y19_to_EI_1s;
wire[1:0] Tile_X9Y19_to_WA_1s;
wire[1:0] Tile_X9Y19_to_WB_1s;
wire[1:0] Tile_X9Y19_to_WC_1s;
wire[1:0] Tile_X9Y19_to_WD_1s;
wire[1:0] Tile_X9Y19_to_WF_1s;
wire[1:0] Tile_X9Y19_to_WG_1s;
wire[1:0] Tile_X9Y19_to_WH_1s;
wire[1:0] Tile_X9Y19_to_WI_1s;
wire[1:0] Tile_X9Y19_to_NA_1s;
wire[1:0] Tile_X9Y19_to_NB_1s;
wire[1:0] Tile_X9Y19_to_NC_1s;
wire[1:0] Tile_X9Y19_to_ND_1s;
wire[1:0] Tile_X9Y19_to_NF_1s;
wire[1:0] Tile_X9Y19_to_NG_1s;
wire[1:0] Tile_X9Y19_to_NH_1s;
wire[1:0] Tile_X9Y19_to_NI_1s;
wire[1:0] Tile_X9Y19_to_SA_1s;
wire[1:0] Tile_X9Y19_to_SB_1s;
wire[1:0] Tile_X9Y19_to_SC_1s;
wire[1:0] Tile_X9Y19_to_SD_1s;
wire[1:0] Tile_X9Y19_to_SF_1s;
wire[1:0] Tile_X9Y19_to_SG_1s;
wire[1:0] Tile_X9Y19_to_SH_1s;
wire[1:0] Tile_X9Y19_to_SI_1s;
wire[1:0] Tile_X10Y19_to_WA_1s;
wire[1:0] Tile_X10Y19_to_WB_1s;
wire[1:0] Tile_X10Y19_to_WC_1s;
wire[1:0] Tile_X10Y19_to_WD_1s;
wire[1:0] Tile_X10Y19_to_WF_1s;
wire[1:0] Tile_X10Y19_to_WG_1s;
wire[1:0] Tile_X10Y19_to_WH_1s;
wire[1:0] Tile_X10Y19_to_WI_1s;
wire[3:0] Tile_X0Y20_to_EA;
wire[3:0] Tile_X0Y20_to_EB;
wire[3:0] Tile_X0Y20_to_EC;
wire[3:0] Tile_X0Y20_to_ED;
wire[3:0] Tile_X0Y20_to_EF;
wire[7:0] Tile_X0Y20_to_EG;
wire[7:0] Tile_X0Y20_to_EH;
wire[11:0] Tile_X0Y20_to_EI;
wire[3:0] Tile_X0Y20_to_NA;
wire[3:0] Tile_X0Y20_to_NB;
wire[3:0] Tile_X0Y20_to_NC;
wire[3:0] Tile_X0Y20_to_ND;
wire[3:0] Tile_X0Y20_to_NF;
wire[7:0] Tile_X0Y20_to_NG;
wire[7:0] Tile_X0Y20_to_NH;
wire[11:0] Tile_X0Y20_to_NI;
wire[3:0] Tile_X0Y20_to_SA;
wire[3:0] Tile_X0Y20_to_SB;
wire[3:0] Tile_X0Y20_to_SC;
wire[3:0] Tile_X0Y20_to_SD;
wire[3:0] Tile_X0Y20_to_SF;
wire[7:0] Tile_X0Y20_to_SG;
wire[7:0] Tile_X0Y20_to_SH;
wire[11:0] Tile_X0Y20_to_SI;
wire[3:0] Tile_X1Y20_to_EA;
wire[3:0] Tile_X1Y20_to_EB;
wire[3:0] Tile_X1Y20_to_EC;
wire[3:0] Tile_X1Y20_to_ED;
wire[3:0] Tile_X1Y20_to_EF;
wire[7:0] Tile_X1Y20_to_EG;
wire[7:0] Tile_X1Y20_to_EH;
wire[11:0] Tile_X1Y20_to_EI;
wire[3:0] Tile_X1Y20_to_WA;
wire[3:0] Tile_X1Y20_to_WB;
wire[3:0] Tile_X1Y20_to_WC;
wire[3:0] Tile_X1Y20_to_WD;
wire[3:0] Tile_X1Y20_to_WF;
wire[7:0] Tile_X1Y20_to_WG;
wire[7:0] Tile_X1Y20_to_WH;
wire[11:0] Tile_X1Y20_to_WI;
wire[3:0] Tile_X1Y20_to_NA;
wire[3:0] Tile_X1Y20_to_NB;
wire[3:0] Tile_X1Y20_to_NC;
wire[3:0] Tile_X1Y20_to_ND;
wire[3:0] Tile_X1Y20_to_NF;
wire[7:0] Tile_X1Y20_to_NG;
wire[7:0] Tile_X1Y20_to_NH;
wire[11:0] Tile_X1Y20_to_NI;
wire[3:0] Tile_X1Y20_to_SA;
wire[3:0] Tile_X1Y20_to_SB;
wire[3:0] Tile_X1Y20_to_SC;
wire[3:0] Tile_X1Y20_to_SD;
wire[3:0] Tile_X1Y20_to_SF;
wire[7:0] Tile_X1Y20_to_SG;
wire[7:0] Tile_X1Y20_to_SH;
wire[11:0] Tile_X1Y20_to_SI;
wire[3:0] Tile_X2Y20_to_EA;
wire[3:0] Tile_X2Y20_to_EB;
wire[3:0] Tile_X2Y20_to_EC;
wire[3:0] Tile_X2Y20_to_ED;
wire[3:0] Tile_X2Y20_to_EF;
wire[7:0] Tile_X2Y20_to_EG;
wire[7:0] Tile_X2Y20_to_EH;
wire[11:0] Tile_X2Y20_to_EI;
wire[3:0] Tile_X2Y20_to_WA;
wire[3:0] Tile_X2Y20_to_WB;
wire[3:0] Tile_X2Y20_to_WC;
wire[3:0] Tile_X2Y20_to_WD;
wire[3:0] Tile_X2Y20_to_WF;
wire[7:0] Tile_X2Y20_to_WG;
wire[7:0] Tile_X2Y20_to_WH;
wire[11:0] Tile_X2Y20_to_WI;
wire[3:0] Tile_X2Y20_to_NA;
wire[3:0] Tile_X2Y20_to_NB;
wire[3:0] Tile_X2Y20_to_NC;
wire[3:0] Tile_X2Y20_to_ND;
wire[3:0] Tile_X2Y20_to_NF;
wire[7:0] Tile_X2Y20_to_NG;
wire[7:0] Tile_X2Y20_to_NH;
wire[11:0] Tile_X2Y20_to_NI;
wire[3:0] Tile_X2Y20_to_SA;
wire[3:0] Tile_X2Y20_to_SB;
wire[3:0] Tile_X2Y20_to_SC;
wire[3:0] Tile_X2Y20_to_SD;
wire[3:0] Tile_X2Y20_to_SF;
wire[7:0] Tile_X2Y20_to_SG;
wire[7:0] Tile_X2Y20_to_SH;
wire[11:0] Tile_X2Y20_to_SI;
wire[3:0] Tile_X3Y20_to_EA;
wire[3:0] Tile_X3Y20_to_EB;
wire[3:0] Tile_X3Y20_to_EC;
wire[3:0] Tile_X3Y20_to_ED;
wire[3:0] Tile_X3Y20_to_EF;
wire[7:0] Tile_X3Y20_to_EG;
wire[7:0] Tile_X3Y20_to_EH;
wire[11:0] Tile_X3Y20_to_EI;
wire[3:0] Tile_X3Y20_to_WA;
wire[3:0] Tile_X3Y20_to_WB;
wire[3:0] Tile_X3Y20_to_WC;
wire[3:0] Tile_X3Y20_to_WD;
wire[3:0] Tile_X3Y20_to_WF;
wire[7:0] Tile_X3Y20_to_WG;
wire[7:0] Tile_X3Y20_to_WH;
wire[11:0] Tile_X3Y20_to_WI;
wire[3:0] Tile_X3Y20_to_NA;
wire[3:0] Tile_X3Y20_to_NB;
wire[3:0] Tile_X3Y20_to_NC;
wire[3:0] Tile_X3Y20_to_ND;
wire[3:0] Tile_X3Y20_to_NF;
wire[7:0] Tile_X3Y20_to_NG;
wire[7:0] Tile_X3Y20_to_NH;
wire[11:0] Tile_X3Y20_to_NI;
wire[3:0] Tile_X3Y20_to_SA;
wire[3:0] Tile_X3Y20_to_SB;
wire[3:0] Tile_X3Y20_to_SC;
wire[3:0] Tile_X3Y20_to_SD;
wire[3:0] Tile_X3Y20_to_SF;
wire[7:0] Tile_X3Y20_to_SG;
wire[7:0] Tile_X3Y20_to_SH;
wire[11:0] Tile_X3Y20_to_SI;
wire[3:0] Tile_X4Y20_to_EA;
wire[3:0] Tile_X4Y20_to_EB;
wire[3:0] Tile_X4Y20_to_EC;
wire[3:0] Tile_X4Y20_to_ED;
wire[3:0] Tile_X4Y20_to_EF;
wire[7:0] Tile_X4Y20_to_EG;
wire[7:0] Tile_X4Y20_to_EH;
wire[11:0] Tile_X4Y20_to_EI;
wire[3:0] Tile_X4Y20_to_WA;
wire[3:0] Tile_X4Y20_to_WB;
wire[3:0] Tile_X4Y20_to_WC;
wire[3:0] Tile_X4Y20_to_WD;
wire[3:0] Tile_X4Y20_to_WF;
wire[7:0] Tile_X4Y20_to_WG;
wire[7:0] Tile_X4Y20_to_WH;
wire[11:0] Tile_X4Y20_to_WI;
wire[3:0] Tile_X4Y20_to_NA;
wire[3:0] Tile_X4Y20_to_NB;
wire[3:0] Tile_X4Y20_to_NC;
wire[3:0] Tile_X4Y20_to_ND;
wire[3:0] Tile_X4Y20_to_NF;
wire[7:0] Tile_X4Y20_to_NG;
wire[7:0] Tile_X4Y20_to_NH;
wire[11:0] Tile_X4Y20_to_NI;
wire[3:0] Tile_X4Y20_to_SA;
wire[3:0] Tile_X4Y20_to_SB;
wire[3:0] Tile_X4Y20_to_SC;
wire[3:0] Tile_X4Y20_to_SD;
wire[3:0] Tile_X4Y20_to_SF;
wire[7:0] Tile_X4Y20_to_SG;
wire[7:0] Tile_X4Y20_to_SH;
wire[11:0] Tile_X4Y20_to_SI;
wire[3:0] Tile_X5Y20_to_EA;
wire[3:0] Tile_X5Y20_to_EB;
wire[3:0] Tile_X5Y20_to_EC;
wire[3:0] Tile_X5Y20_to_ED;
wire[3:0] Tile_X5Y20_to_EF;
wire[7:0] Tile_X5Y20_to_EG;
wire[7:0] Tile_X5Y20_to_EH;
wire[11:0] Tile_X5Y20_to_EI;
wire[3:0] Tile_X5Y20_to_WA;
wire[3:0] Tile_X5Y20_to_WB;
wire[3:0] Tile_X5Y20_to_WC;
wire[3:0] Tile_X5Y20_to_WD;
wire[3:0] Tile_X5Y20_to_WF;
wire[7:0] Tile_X5Y20_to_WG;
wire[7:0] Tile_X5Y20_to_WH;
wire[11:0] Tile_X5Y20_to_WI;
wire[3:0] Tile_X5Y20_to_NA;
wire[3:0] Tile_X5Y20_to_NB;
wire[3:0] Tile_X5Y20_to_NC;
wire[3:0] Tile_X5Y20_to_ND;
wire[3:0] Tile_X5Y20_to_NF;
wire[7:0] Tile_X5Y20_to_NG;
wire[7:0] Tile_X5Y20_to_NH;
wire[11:0] Tile_X5Y20_to_NI;
wire[3:0] Tile_X5Y20_to_SA;
wire[3:0] Tile_X5Y20_to_SB;
wire[3:0] Tile_X5Y20_to_SC;
wire[3:0] Tile_X5Y20_to_SD;
wire[3:0] Tile_X5Y20_to_SF;
wire[7:0] Tile_X5Y20_to_SG;
wire[7:0] Tile_X5Y20_to_SH;
wire[11:0] Tile_X5Y20_to_SI;
wire[3:0] Tile_X6Y20_to_EA;
wire[3:0] Tile_X6Y20_to_EB;
wire[3:0] Tile_X6Y20_to_EC;
wire[3:0] Tile_X6Y20_to_ED;
wire[3:0] Tile_X6Y20_to_EF;
wire[7:0] Tile_X6Y20_to_EG;
wire[7:0] Tile_X6Y20_to_EH;
wire[11:0] Tile_X6Y20_to_EI;
wire[3:0] Tile_X6Y20_to_WA;
wire[3:0] Tile_X6Y20_to_WB;
wire[3:0] Tile_X6Y20_to_WC;
wire[3:0] Tile_X6Y20_to_WD;
wire[3:0] Tile_X6Y20_to_WF;
wire[7:0] Tile_X6Y20_to_WG;
wire[7:0] Tile_X6Y20_to_WH;
wire[11:0] Tile_X6Y20_to_WI;
wire[3:0] Tile_X6Y20_to_NA;
wire[3:0] Tile_X6Y20_to_NB;
wire[3:0] Tile_X6Y20_to_NC;
wire[3:0] Tile_X6Y20_to_ND;
wire[3:0] Tile_X6Y20_to_NF;
wire[7:0] Tile_X6Y20_to_NG;
wire[7:0] Tile_X6Y20_to_NH;
wire[11:0] Tile_X6Y20_to_NI;
wire[3:0] Tile_X6Y20_to_SA;
wire[3:0] Tile_X6Y20_to_SB;
wire[3:0] Tile_X6Y20_to_SC;
wire[3:0] Tile_X6Y20_to_SD;
wire[3:0] Tile_X6Y20_to_SF;
wire[7:0] Tile_X6Y20_to_SG;
wire[7:0] Tile_X6Y20_to_SH;
wire[11:0] Tile_X6Y20_to_SI;
wire[3:0] Tile_X7Y20_to_EA;
wire[3:0] Tile_X7Y20_to_EB;
wire[3:0] Tile_X7Y20_to_EC;
wire[3:0] Tile_X7Y20_to_ED;
wire[3:0] Tile_X7Y20_to_EF;
wire[7:0] Tile_X7Y20_to_EG;
wire[7:0] Tile_X7Y20_to_EH;
wire[11:0] Tile_X7Y20_to_EI;
wire[3:0] Tile_X7Y20_to_WA;
wire[3:0] Tile_X7Y20_to_WB;
wire[3:0] Tile_X7Y20_to_WC;
wire[3:0] Tile_X7Y20_to_WD;
wire[3:0] Tile_X7Y20_to_WF;
wire[7:0] Tile_X7Y20_to_WG;
wire[7:0] Tile_X7Y20_to_WH;
wire[11:0] Tile_X7Y20_to_WI;
wire[3:0] Tile_X7Y20_to_NA;
wire[3:0] Tile_X7Y20_to_NB;
wire[3:0] Tile_X7Y20_to_NC;
wire[3:0] Tile_X7Y20_to_ND;
wire[3:0] Tile_X7Y20_to_NF;
wire[7:0] Tile_X7Y20_to_NG;
wire[7:0] Tile_X7Y20_to_NH;
wire[11:0] Tile_X7Y20_to_NI;
wire[3:0] Tile_X7Y20_to_SA;
wire[3:0] Tile_X7Y20_to_SB;
wire[3:0] Tile_X7Y20_to_SC;
wire[3:0] Tile_X7Y20_to_SD;
wire[3:0] Tile_X7Y20_to_SF;
wire[7:0] Tile_X7Y20_to_SG;
wire[7:0] Tile_X7Y20_to_SH;
wire[11:0] Tile_X7Y20_to_SI;
wire[3:0] Tile_X8Y20_to_WA;
wire[3:0] Tile_X8Y20_to_WB;
wire[3:0] Tile_X8Y20_to_WC;
wire[3:0] Tile_X8Y20_to_WD;
wire[3:0] Tile_X8Y20_to_WF;
wire[7:0] Tile_X8Y20_to_WG;
wire[7:0] Tile_X8Y20_to_WH;
wire[11:0] Tile_X8Y20_to_WI;
wire[3:0] Tile_X8Y20_to_NA;
wire[3:0] Tile_X8Y20_to_NB;
wire[3:0] Tile_X8Y20_to_NC;
wire[3:0] Tile_X8Y20_to_ND;
wire[3:0] Tile_X8Y20_to_NF;
wire[7:0] Tile_X8Y20_to_NG;
wire[7:0] Tile_X8Y20_to_NH;
wire[11:0] Tile_X8Y20_to_NI;
wire[3:0] Tile_X8Y20_to_SA;
wire[3:0] Tile_X8Y20_to_SB;
wire[3:0] Tile_X8Y20_to_SC;
wire[3:0] Tile_X8Y20_to_SD;
wire[3:0] Tile_X8Y20_to_SF;
wire[7:0] Tile_X8Y20_to_SG;
wire[7:0] Tile_X8Y20_to_SH;
wire[11:0] Tile_X8Y20_to_SI;
wire[1:0] Tile_X9Y20_to_EA_1s;
wire[1:0] Tile_X9Y20_to_EB_1s;
wire[1:0] Tile_X9Y20_to_EC_1s;
wire[1:0] Tile_X9Y20_to_ED_1s;
wire[1:0] Tile_X9Y20_to_EF_1s;
wire[1:0] Tile_X9Y20_to_EG_1s;
wire[1:0] Tile_X9Y20_to_EH_1s;
wire[1:0] Tile_X9Y20_to_EI_1s;
wire[1:0] Tile_X9Y20_to_WA_1s;
wire[1:0] Tile_X9Y20_to_WB_1s;
wire[1:0] Tile_X9Y20_to_WC_1s;
wire[1:0] Tile_X9Y20_to_WD_1s;
wire[1:0] Tile_X9Y20_to_WF_1s;
wire[1:0] Tile_X9Y20_to_WG_1s;
wire[1:0] Tile_X9Y20_to_WH_1s;
wire[1:0] Tile_X9Y20_to_WI_1s;
wire[1:0] Tile_X9Y20_to_NA_1s;
wire[1:0] Tile_X9Y20_to_NB_1s;
wire[1:0] Tile_X9Y20_to_NC_1s;
wire[1:0] Tile_X9Y20_to_ND_1s;
wire[1:0] Tile_X9Y20_to_NF_1s;
wire[1:0] Tile_X9Y20_to_NG_1s;
wire[1:0] Tile_X9Y20_to_NH_1s;
wire[1:0] Tile_X9Y20_to_NI_1s;
wire[1:0] Tile_X9Y20_to_SA_1s;
wire[1:0] Tile_X9Y20_to_SB_1s;
wire[1:0] Tile_X9Y20_to_SC_1s;
wire[1:0] Tile_X9Y20_to_SD_1s;
wire[1:0] Tile_X9Y20_to_SF_1s;
wire[1:0] Tile_X9Y20_to_SG_1s;
wire[1:0] Tile_X9Y20_to_SH_1s;
wire[1:0] Tile_X9Y20_to_SI_1s;
wire[1:0] Tile_X10Y20_to_WA_1s;
wire[1:0] Tile_X10Y20_to_WB_1s;
wire[1:0] Tile_X10Y20_to_WC_1s;
wire[1:0] Tile_X10Y20_to_WD_1s;
wire[1:0] Tile_X10Y20_to_WF_1s;
wire[1:0] Tile_X10Y20_to_WG_1s;
wire[1:0] Tile_X10Y20_to_WH_1s;
wire[1:0] Tile_X10Y20_to_WI_1s;
wire[3:0] Tile_X0Y21_to_EA;
wire[3:0] Tile_X0Y21_to_EB;
wire[3:0] Tile_X0Y21_to_EC;
wire[3:0] Tile_X0Y21_to_ED;
wire[3:0] Tile_X0Y21_to_EF;
wire[7:0] Tile_X0Y21_to_EG;
wire[7:0] Tile_X0Y21_to_EH;
wire[11:0] Tile_X0Y21_to_EI;
wire[3:0] Tile_X0Y21_to_NA;
wire[3:0] Tile_X0Y21_to_NB;
wire[3:0] Tile_X0Y21_to_NC;
wire[3:0] Tile_X0Y21_to_ND;
wire[3:0] Tile_X0Y21_to_NF;
wire[7:0] Tile_X0Y21_to_NG;
wire[7:0] Tile_X0Y21_to_NH;
wire[11:0] Tile_X0Y21_to_NI;
wire[3:0] Tile_X0Y21_to_SA;
wire[3:0] Tile_X0Y21_to_SB;
wire[3:0] Tile_X0Y21_to_SC;
wire[3:0] Tile_X0Y21_to_SD;
wire[3:0] Tile_X0Y21_to_SF;
wire[7:0] Tile_X0Y21_to_SG;
wire[7:0] Tile_X0Y21_to_SH;
wire[11:0] Tile_X0Y21_to_SI;
wire[3:0] Tile_X1Y21_to_EA;
wire[3:0] Tile_X1Y21_to_EB;
wire[3:0] Tile_X1Y21_to_EC;
wire[3:0] Tile_X1Y21_to_ED;
wire[3:0] Tile_X1Y21_to_EF;
wire[7:0] Tile_X1Y21_to_EG;
wire[7:0] Tile_X1Y21_to_EH;
wire[11:0] Tile_X1Y21_to_EI;
wire[3:0] Tile_X1Y21_to_WA;
wire[3:0] Tile_X1Y21_to_WB;
wire[3:0] Tile_X1Y21_to_WC;
wire[3:0] Tile_X1Y21_to_WD;
wire[3:0] Tile_X1Y21_to_WF;
wire[7:0] Tile_X1Y21_to_WG;
wire[7:0] Tile_X1Y21_to_WH;
wire[11:0] Tile_X1Y21_to_WI;
wire[3:0] Tile_X1Y21_to_NA;
wire[3:0] Tile_X1Y21_to_NB;
wire[3:0] Tile_X1Y21_to_NC;
wire[3:0] Tile_X1Y21_to_ND;
wire[3:0] Tile_X1Y21_to_NF;
wire[7:0] Tile_X1Y21_to_NG;
wire[7:0] Tile_X1Y21_to_NH;
wire[11:0] Tile_X1Y21_to_NI;
wire[3:0] Tile_X1Y21_to_SA;
wire[3:0] Tile_X1Y21_to_SB;
wire[3:0] Tile_X1Y21_to_SC;
wire[3:0] Tile_X1Y21_to_SD;
wire[3:0] Tile_X1Y21_to_SF;
wire[7:0] Tile_X1Y21_to_SG;
wire[7:0] Tile_X1Y21_to_SH;
wire[11:0] Tile_X1Y21_to_SI;
wire[3:0] Tile_X2Y21_to_EA;
wire[3:0] Tile_X2Y21_to_EB;
wire[3:0] Tile_X2Y21_to_EC;
wire[3:0] Tile_X2Y21_to_ED;
wire[3:0] Tile_X2Y21_to_EF;
wire[7:0] Tile_X2Y21_to_EG;
wire[7:0] Tile_X2Y21_to_EH;
wire[11:0] Tile_X2Y21_to_EI;
wire[3:0] Tile_X2Y21_to_WA;
wire[3:0] Tile_X2Y21_to_WB;
wire[3:0] Tile_X2Y21_to_WC;
wire[3:0] Tile_X2Y21_to_WD;
wire[3:0] Tile_X2Y21_to_WF;
wire[7:0] Tile_X2Y21_to_WG;
wire[7:0] Tile_X2Y21_to_WH;
wire[11:0] Tile_X2Y21_to_WI;
wire[3:0] Tile_X2Y21_to_NA;
wire[3:0] Tile_X2Y21_to_NB;
wire[3:0] Tile_X2Y21_to_NC;
wire[3:0] Tile_X2Y21_to_ND;
wire[3:0] Tile_X2Y21_to_NF;
wire[7:0] Tile_X2Y21_to_NG;
wire[7:0] Tile_X2Y21_to_NH;
wire[11:0] Tile_X2Y21_to_NI;
wire[3:0] Tile_X2Y21_to_SA;
wire[3:0] Tile_X2Y21_to_SB;
wire[3:0] Tile_X2Y21_to_SC;
wire[3:0] Tile_X2Y21_to_SD;
wire[3:0] Tile_X2Y21_to_SF;
wire[7:0] Tile_X2Y21_to_SG;
wire[7:0] Tile_X2Y21_to_SH;
wire[11:0] Tile_X2Y21_to_SI;
wire[3:0] Tile_X3Y21_to_EA;
wire[3:0] Tile_X3Y21_to_EB;
wire[3:0] Tile_X3Y21_to_EC;
wire[3:0] Tile_X3Y21_to_ED;
wire[3:0] Tile_X3Y21_to_EF;
wire[7:0] Tile_X3Y21_to_EG;
wire[7:0] Tile_X3Y21_to_EH;
wire[11:0] Tile_X3Y21_to_EI;
wire[3:0] Tile_X3Y21_to_WA;
wire[3:0] Tile_X3Y21_to_WB;
wire[3:0] Tile_X3Y21_to_WC;
wire[3:0] Tile_X3Y21_to_WD;
wire[3:0] Tile_X3Y21_to_WF;
wire[7:0] Tile_X3Y21_to_WG;
wire[7:0] Tile_X3Y21_to_WH;
wire[11:0] Tile_X3Y21_to_WI;
wire[3:0] Tile_X3Y21_to_NA;
wire[3:0] Tile_X3Y21_to_NB;
wire[3:0] Tile_X3Y21_to_NC;
wire[3:0] Tile_X3Y21_to_ND;
wire[3:0] Tile_X3Y21_to_NF;
wire[7:0] Tile_X3Y21_to_NG;
wire[7:0] Tile_X3Y21_to_NH;
wire[11:0] Tile_X3Y21_to_NI;
wire[3:0] Tile_X3Y21_to_SA;
wire[3:0] Tile_X3Y21_to_SB;
wire[3:0] Tile_X3Y21_to_SC;
wire[3:0] Tile_X3Y21_to_SD;
wire[3:0] Tile_X3Y21_to_SF;
wire[7:0] Tile_X3Y21_to_SG;
wire[7:0] Tile_X3Y21_to_SH;
wire[11:0] Tile_X3Y21_to_SI;
wire[3:0] Tile_X4Y21_to_EA;
wire[3:0] Tile_X4Y21_to_EB;
wire[3:0] Tile_X4Y21_to_EC;
wire[3:0] Tile_X4Y21_to_ED;
wire[3:0] Tile_X4Y21_to_EF;
wire[7:0] Tile_X4Y21_to_EG;
wire[7:0] Tile_X4Y21_to_EH;
wire[11:0] Tile_X4Y21_to_EI;
wire[3:0] Tile_X4Y21_to_WA;
wire[3:0] Tile_X4Y21_to_WB;
wire[3:0] Tile_X4Y21_to_WC;
wire[3:0] Tile_X4Y21_to_WD;
wire[3:0] Tile_X4Y21_to_WF;
wire[7:0] Tile_X4Y21_to_WG;
wire[7:0] Tile_X4Y21_to_WH;
wire[11:0] Tile_X4Y21_to_WI;
wire[3:0] Tile_X4Y21_to_NA;
wire[3:0] Tile_X4Y21_to_NB;
wire[3:0] Tile_X4Y21_to_NC;
wire[3:0] Tile_X4Y21_to_ND;
wire[3:0] Tile_X4Y21_to_NF;
wire[7:0] Tile_X4Y21_to_NG;
wire[7:0] Tile_X4Y21_to_NH;
wire[11:0] Tile_X4Y21_to_NI;
wire[3:0] Tile_X4Y21_to_SA;
wire[3:0] Tile_X4Y21_to_SB;
wire[3:0] Tile_X4Y21_to_SC;
wire[3:0] Tile_X4Y21_to_SD;
wire[3:0] Tile_X4Y21_to_SF;
wire[7:0] Tile_X4Y21_to_SG;
wire[7:0] Tile_X4Y21_to_SH;
wire[11:0] Tile_X4Y21_to_SI;
wire[3:0] Tile_X5Y21_to_EA;
wire[3:0] Tile_X5Y21_to_EB;
wire[3:0] Tile_X5Y21_to_EC;
wire[3:0] Tile_X5Y21_to_ED;
wire[3:0] Tile_X5Y21_to_EF;
wire[7:0] Tile_X5Y21_to_EG;
wire[7:0] Tile_X5Y21_to_EH;
wire[11:0] Tile_X5Y21_to_EI;
wire[3:0] Tile_X5Y21_to_WA;
wire[3:0] Tile_X5Y21_to_WB;
wire[3:0] Tile_X5Y21_to_WC;
wire[3:0] Tile_X5Y21_to_WD;
wire[3:0] Tile_X5Y21_to_WF;
wire[7:0] Tile_X5Y21_to_WG;
wire[7:0] Tile_X5Y21_to_WH;
wire[11:0] Tile_X5Y21_to_WI;
wire[3:0] Tile_X5Y21_to_NA;
wire[3:0] Tile_X5Y21_to_NB;
wire[3:0] Tile_X5Y21_to_NC;
wire[3:0] Tile_X5Y21_to_ND;
wire[3:0] Tile_X5Y21_to_NF;
wire[7:0] Tile_X5Y21_to_NG;
wire[7:0] Tile_X5Y21_to_NH;
wire[11:0] Tile_X5Y21_to_NI;
wire[3:0] Tile_X5Y21_to_SA;
wire[3:0] Tile_X5Y21_to_SB;
wire[3:0] Tile_X5Y21_to_SC;
wire[3:0] Tile_X5Y21_to_SD;
wire[3:0] Tile_X5Y21_to_SF;
wire[7:0] Tile_X5Y21_to_SG;
wire[7:0] Tile_X5Y21_to_SH;
wire[11:0] Tile_X5Y21_to_SI;
wire[3:0] Tile_X6Y21_to_EA;
wire[3:0] Tile_X6Y21_to_EB;
wire[3:0] Tile_X6Y21_to_EC;
wire[3:0] Tile_X6Y21_to_ED;
wire[3:0] Tile_X6Y21_to_EF;
wire[7:0] Tile_X6Y21_to_EG;
wire[7:0] Tile_X6Y21_to_EH;
wire[11:0] Tile_X6Y21_to_EI;
wire[3:0] Tile_X6Y21_to_WA;
wire[3:0] Tile_X6Y21_to_WB;
wire[3:0] Tile_X6Y21_to_WC;
wire[3:0] Tile_X6Y21_to_WD;
wire[3:0] Tile_X6Y21_to_WF;
wire[7:0] Tile_X6Y21_to_WG;
wire[7:0] Tile_X6Y21_to_WH;
wire[11:0] Tile_X6Y21_to_WI;
wire[3:0] Tile_X6Y21_to_NA;
wire[3:0] Tile_X6Y21_to_NB;
wire[3:0] Tile_X6Y21_to_NC;
wire[3:0] Tile_X6Y21_to_ND;
wire[3:0] Tile_X6Y21_to_NF;
wire[7:0] Tile_X6Y21_to_NG;
wire[7:0] Tile_X6Y21_to_NH;
wire[11:0] Tile_X6Y21_to_NI;
wire[3:0] Tile_X6Y21_to_SA;
wire[3:0] Tile_X6Y21_to_SB;
wire[3:0] Tile_X6Y21_to_SC;
wire[3:0] Tile_X6Y21_to_SD;
wire[3:0] Tile_X6Y21_to_SF;
wire[7:0] Tile_X6Y21_to_SG;
wire[7:0] Tile_X6Y21_to_SH;
wire[11:0] Tile_X6Y21_to_SI;
wire[3:0] Tile_X7Y21_to_EA;
wire[3:0] Tile_X7Y21_to_EB;
wire[3:0] Tile_X7Y21_to_EC;
wire[3:0] Tile_X7Y21_to_ED;
wire[3:0] Tile_X7Y21_to_EF;
wire[7:0] Tile_X7Y21_to_EG;
wire[7:0] Tile_X7Y21_to_EH;
wire[11:0] Tile_X7Y21_to_EI;
wire[3:0] Tile_X7Y21_to_WA;
wire[3:0] Tile_X7Y21_to_WB;
wire[3:0] Tile_X7Y21_to_WC;
wire[3:0] Tile_X7Y21_to_WD;
wire[3:0] Tile_X7Y21_to_WF;
wire[7:0] Tile_X7Y21_to_WG;
wire[7:0] Tile_X7Y21_to_WH;
wire[11:0] Tile_X7Y21_to_WI;
wire[3:0] Tile_X7Y21_to_NA;
wire[3:0] Tile_X7Y21_to_NB;
wire[3:0] Tile_X7Y21_to_NC;
wire[3:0] Tile_X7Y21_to_ND;
wire[3:0] Tile_X7Y21_to_NF;
wire[7:0] Tile_X7Y21_to_NG;
wire[7:0] Tile_X7Y21_to_NH;
wire[11:0] Tile_X7Y21_to_NI;
wire[3:0] Tile_X7Y21_to_SA;
wire[3:0] Tile_X7Y21_to_SB;
wire[3:0] Tile_X7Y21_to_SC;
wire[3:0] Tile_X7Y21_to_SD;
wire[3:0] Tile_X7Y21_to_SF;
wire[7:0] Tile_X7Y21_to_SG;
wire[7:0] Tile_X7Y21_to_SH;
wire[11:0] Tile_X7Y21_to_SI;
wire[3:0] Tile_X8Y21_to_WA;
wire[3:0] Tile_X8Y21_to_WB;
wire[3:0] Tile_X8Y21_to_WC;
wire[3:0] Tile_X8Y21_to_WD;
wire[3:0] Tile_X8Y21_to_WF;
wire[7:0] Tile_X8Y21_to_WG;
wire[7:0] Tile_X8Y21_to_WH;
wire[11:0] Tile_X8Y21_to_WI;
wire[3:0] Tile_X8Y21_to_NA;
wire[3:0] Tile_X8Y21_to_NB;
wire[3:0] Tile_X8Y21_to_NC;
wire[3:0] Tile_X8Y21_to_ND;
wire[3:0] Tile_X8Y21_to_NF;
wire[7:0] Tile_X8Y21_to_NG;
wire[7:0] Tile_X8Y21_to_NH;
wire[11:0] Tile_X8Y21_to_NI;
wire[3:0] Tile_X8Y21_to_SA;
wire[3:0] Tile_X8Y21_to_SB;
wire[3:0] Tile_X8Y21_to_SC;
wire[3:0] Tile_X8Y21_to_SD;
wire[3:0] Tile_X8Y21_to_SF;
wire[7:0] Tile_X8Y21_to_SG;
wire[7:0] Tile_X8Y21_to_SH;
wire[11:0] Tile_X8Y21_to_SI;
wire[1:0] Tile_X9Y21_to_EA_1s;
wire[1:0] Tile_X9Y21_to_EB_1s;
wire[1:0] Tile_X9Y21_to_EC_1s;
wire[1:0] Tile_X9Y21_to_ED_1s;
wire[1:0] Tile_X9Y21_to_EF_1s;
wire[1:0] Tile_X9Y21_to_EG_1s;
wire[1:0] Tile_X9Y21_to_EH_1s;
wire[1:0] Tile_X9Y21_to_EI_1s;
wire[1:0] Tile_X9Y21_to_WA_1s;
wire[1:0] Tile_X9Y21_to_WB_1s;
wire[1:0] Tile_X9Y21_to_WC_1s;
wire[1:0] Tile_X9Y21_to_WD_1s;
wire[1:0] Tile_X9Y21_to_WF_1s;
wire[1:0] Tile_X9Y21_to_WG_1s;
wire[1:0] Tile_X9Y21_to_WH_1s;
wire[1:0] Tile_X9Y21_to_WI_1s;
wire[1:0] Tile_X9Y21_to_NA_1s;
wire[1:0] Tile_X9Y21_to_NB_1s;
wire[1:0] Tile_X9Y21_to_NC_1s;
wire[1:0] Tile_X9Y21_to_ND_1s;
wire[1:0] Tile_X9Y21_to_NF_1s;
wire[1:0] Tile_X9Y21_to_NG_1s;
wire[1:0] Tile_X9Y21_to_NH_1s;
wire[1:0] Tile_X9Y21_to_NI_1s;
wire[1:0] Tile_X9Y21_to_SA_1s;
wire[1:0] Tile_X9Y21_to_SB_1s;
wire[1:0] Tile_X9Y21_to_SC_1s;
wire[1:0] Tile_X9Y21_to_SD_1s;
wire[1:0] Tile_X9Y21_to_SF_1s;
wire[1:0] Tile_X9Y21_to_SG_1s;
wire[1:0] Tile_X9Y21_to_SH_1s;
wire[1:0] Tile_X9Y21_to_SI_1s;
wire[1:0] Tile_X10Y21_to_WA_1s;
wire[1:0] Tile_X10Y21_to_WB_1s;
wire[1:0] Tile_X10Y21_to_WC_1s;
wire[1:0] Tile_X10Y21_to_WD_1s;
wire[1:0] Tile_X10Y21_to_WF_1s;
wire[1:0] Tile_X10Y21_to_WG_1s;
wire[1:0] Tile_X10Y21_to_WH_1s;
wire[1:0] Tile_X10Y21_to_WI_1s;
wire[3:0] Tile_X0Y22_to_EA;
wire[3:0] Tile_X0Y22_to_EB;
wire[3:0] Tile_X0Y22_to_EC;
wire[3:0] Tile_X0Y22_to_ED;
wire[3:0] Tile_X0Y22_to_EF;
wire[7:0] Tile_X0Y22_to_EG;
wire[7:0] Tile_X0Y22_to_EH;
wire[11:0] Tile_X0Y22_to_EI;
wire[3:0] Tile_X0Y22_to_NA;
wire[3:0] Tile_X0Y22_to_NB;
wire[3:0] Tile_X0Y22_to_NC;
wire[3:0] Tile_X0Y22_to_ND;
wire[3:0] Tile_X0Y22_to_NF;
wire[7:0] Tile_X0Y22_to_NG;
wire[7:0] Tile_X0Y22_to_NH;
wire[11:0] Tile_X0Y22_to_NI;
wire[3:0] Tile_X0Y22_to_SA;
wire[3:0] Tile_X0Y22_to_SB;
wire[3:0] Tile_X0Y22_to_SC;
wire[3:0] Tile_X0Y22_to_SD;
wire[3:0] Tile_X0Y22_to_SF;
wire[7:0] Tile_X0Y22_to_SG;
wire[7:0] Tile_X0Y22_to_SH;
wire[11:0] Tile_X0Y22_to_SI;
wire[3:0] Tile_X1Y22_to_EA;
wire[3:0] Tile_X1Y22_to_EB;
wire[3:0] Tile_X1Y22_to_EC;
wire[3:0] Tile_X1Y22_to_ED;
wire[3:0] Tile_X1Y22_to_EF;
wire[7:0] Tile_X1Y22_to_EG;
wire[7:0] Tile_X1Y22_to_EH;
wire[11:0] Tile_X1Y22_to_EI;
wire[3:0] Tile_X1Y22_to_WA;
wire[3:0] Tile_X1Y22_to_WB;
wire[3:0] Tile_X1Y22_to_WC;
wire[3:0] Tile_X1Y22_to_WD;
wire[3:0] Tile_X1Y22_to_WF;
wire[7:0] Tile_X1Y22_to_WG;
wire[7:0] Tile_X1Y22_to_WH;
wire[11:0] Tile_X1Y22_to_WI;
wire[3:0] Tile_X1Y22_to_NA;
wire[3:0] Tile_X1Y22_to_NB;
wire[3:0] Tile_X1Y22_to_NC;
wire[3:0] Tile_X1Y22_to_ND;
wire[3:0] Tile_X1Y22_to_NF;
wire[7:0] Tile_X1Y22_to_NG;
wire[7:0] Tile_X1Y22_to_NH;
wire[11:0] Tile_X1Y22_to_NI;
wire[3:0] Tile_X1Y22_to_SA;
wire[3:0] Tile_X1Y22_to_SB;
wire[3:0] Tile_X1Y22_to_SC;
wire[3:0] Tile_X1Y22_to_SD;
wire[3:0] Tile_X1Y22_to_SF;
wire[7:0] Tile_X1Y22_to_SG;
wire[7:0] Tile_X1Y22_to_SH;
wire[11:0] Tile_X1Y22_to_SI;
wire[3:0] Tile_X2Y22_to_EA;
wire[3:0] Tile_X2Y22_to_EB;
wire[3:0] Tile_X2Y22_to_EC;
wire[3:0] Tile_X2Y22_to_ED;
wire[3:0] Tile_X2Y22_to_EF;
wire[7:0] Tile_X2Y22_to_EG;
wire[7:0] Tile_X2Y22_to_EH;
wire[11:0] Tile_X2Y22_to_EI;
wire[3:0] Tile_X2Y22_to_WA;
wire[3:0] Tile_X2Y22_to_WB;
wire[3:0] Tile_X2Y22_to_WC;
wire[3:0] Tile_X2Y22_to_WD;
wire[3:0] Tile_X2Y22_to_WF;
wire[7:0] Tile_X2Y22_to_WG;
wire[7:0] Tile_X2Y22_to_WH;
wire[11:0] Tile_X2Y22_to_WI;
wire[3:0] Tile_X2Y22_to_NA;
wire[3:0] Tile_X2Y22_to_NB;
wire[3:0] Tile_X2Y22_to_NC;
wire[3:0] Tile_X2Y22_to_ND;
wire[3:0] Tile_X2Y22_to_NF;
wire[7:0] Tile_X2Y22_to_NG;
wire[7:0] Tile_X2Y22_to_NH;
wire[11:0] Tile_X2Y22_to_NI;
wire[3:0] Tile_X2Y22_to_SA;
wire[3:0] Tile_X2Y22_to_SB;
wire[3:0] Tile_X2Y22_to_SC;
wire[3:0] Tile_X2Y22_to_SD;
wire[3:0] Tile_X2Y22_to_SF;
wire[7:0] Tile_X2Y22_to_SG;
wire[7:0] Tile_X2Y22_to_SH;
wire[11:0] Tile_X2Y22_to_SI;
wire[3:0] Tile_X3Y22_to_EA;
wire[3:0] Tile_X3Y22_to_EB;
wire[3:0] Tile_X3Y22_to_EC;
wire[3:0] Tile_X3Y22_to_ED;
wire[3:0] Tile_X3Y22_to_EF;
wire[7:0] Tile_X3Y22_to_EG;
wire[7:0] Tile_X3Y22_to_EH;
wire[11:0] Tile_X3Y22_to_EI;
wire[3:0] Tile_X3Y22_to_WA;
wire[3:0] Tile_X3Y22_to_WB;
wire[3:0] Tile_X3Y22_to_WC;
wire[3:0] Tile_X3Y22_to_WD;
wire[3:0] Tile_X3Y22_to_WF;
wire[7:0] Tile_X3Y22_to_WG;
wire[7:0] Tile_X3Y22_to_WH;
wire[11:0] Tile_X3Y22_to_WI;
wire[3:0] Tile_X3Y22_to_NA;
wire[3:0] Tile_X3Y22_to_NB;
wire[3:0] Tile_X3Y22_to_NC;
wire[3:0] Tile_X3Y22_to_ND;
wire[3:0] Tile_X3Y22_to_NF;
wire[7:0] Tile_X3Y22_to_NG;
wire[7:0] Tile_X3Y22_to_NH;
wire[11:0] Tile_X3Y22_to_NI;
wire[3:0] Tile_X3Y22_to_SA;
wire[3:0] Tile_X3Y22_to_SB;
wire[3:0] Tile_X3Y22_to_SC;
wire[3:0] Tile_X3Y22_to_SD;
wire[3:0] Tile_X3Y22_to_SF;
wire[7:0] Tile_X3Y22_to_SG;
wire[7:0] Tile_X3Y22_to_SH;
wire[11:0] Tile_X3Y22_to_SI;
wire[3:0] Tile_X4Y22_to_EA;
wire[3:0] Tile_X4Y22_to_EB;
wire[3:0] Tile_X4Y22_to_EC;
wire[3:0] Tile_X4Y22_to_ED;
wire[3:0] Tile_X4Y22_to_EF;
wire[7:0] Tile_X4Y22_to_EG;
wire[7:0] Tile_X4Y22_to_EH;
wire[11:0] Tile_X4Y22_to_EI;
wire[3:0] Tile_X4Y22_to_WA;
wire[3:0] Tile_X4Y22_to_WB;
wire[3:0] Tile_X4Y22_to_WC;
wire[3:0] Tile_X4Y22_to_WD;
wire[3:0] Tile_X4Y22_to_WF;
wire[7:0] Tile_X4Y22_to_WG;
wire[7:0] Tile_X4Y22_to_WH;
wire[11:0] Tile_X4Y22_to_WI;
wire[3:0] Tile_X4Y22_to_NA;
wire[3:0] Tile_X4Y22_to_NB;
wire[3:0] Tile_X4Y22_to_NC;
wire[3:0] Tile_X4Y22_to_ND;
wire[3:0] Tile_X4Y22_to_NF;
wire[7:0] Tile_X4Y22_to_NG;
wire[7:0] Tile_X4Y22_to_NH;
wire[11:0] Tile_X4Y22_to_NI;
wire[3:0] Tile_X4Y22_to_SA;
wire[3:0] Tile_X4Y22_to_SB;
wire[3:0] Tile_X4Y22_to_SC;
wire[3:0] Tile_X4Y22_to_SD;
wire[3:0] Tile_X4Y22_to_SF;
wire[7:0] Tile_X4Y22_to_SG;
wire[7:0] Tile_X4Y22_to_SH;
wire[11:0] Tile_X4Y22_to_SI;
wire[3:0] Tile_X5Y22_to_EA;
wire[3:0] Tile_X5Y22_to_EB;
wire[3:0] Tile_X5Y22_to_EC;
wire[3:0] Tile_X5Y22_to_ED;
wire[3:0] Tile_X5Y22_to_EF;
wire[7:0] Tile_X5Y22_to_EG;
wire[7:0] Tile_X5Y22_to_EH;
wire[11:0] Tile_X5Y22_to_EI;
wire[3:0] Tile_X5Y22_to_WA;
wire[3:0] Tile_X5Y22_to_WB;
wire[3:0] Tile_X5Y22_to_WC;
wire[3:0] Tile_X5Y22_to_WD;
wire[3:0] Tile_X5Y22_to_WF;
wire[7:0] Tile_X5Y22_to_WG;
wire[7:0] Tile_X5Y22_to_WH;
wire[11:0] Tile_X5Y22_to_WI;
wire[3:0] Tile_X5Y22_to_NA;
wire[3:0] Tile_X5Y22_to_NB;
wire[3:0] Tile_X5Y22_to_NC;
wire[3:0] Tile_X5Y22_to_ND;
wire[3:0] Tile_X5Y22_to_NF;
wire[7:0] Tile_X5Y22_to_NG;
wire[7:0] Tile_X5Y22_to_NH;
wire[11:0] Tile_X5Y22_to_NI;
wire[3:0] Tile_X5Y22_to_SA;
wire[3:0] Tile_X5Y22_to_SB;
wire[3:0] Tile_X5Y22_to_SC;
wire[3:0] Tile_X5Y22_to_SD;
wire[3:0] Tile_X5Y22_to_SF;
wire[7:0] Tile_X5Y22_to_SG;
wire[7:0] Tile_X5Y22_to_SH;
wire[11:0] Tile_X5Y22_to_SI;
wire[3:0] Tile_X6Y22_to_EA;
wire[3:0] Tile_X6Y22_to_EB;
wire[3:0] Tile_X6Y22_to_EC;
wire[3:0] Tile_X6Y22_to_ED;
wire[3:0] Tile_X6Y22_to_EF;
wire[7:0] Tile_X6Y22_to_EG;
wire[7:0] Tile_X6Y22_to_EH;
wire[11:0] Tile_X6Y22_to_EI;
wire[3:0] Tile_X6Y22_to_WA;
wire[3:0] Tile_X6Y22_to_WB;
wire[3:0] Tile_X6Y22_to_WC;
wire[3:0] Tile_X6Y22_to_WD;
wire[3:0] Tile_X6Y22_to_WF;
wire[7:0] Tile_X6Y22_to_WG;
wire[7:0] Tile_X6Y22_to_WH;
wire[11:0] Tile_X6Y22_to_WI;
wire[3:0] Tile_X6Y22_to_NA;
wire[3:0] Tile_X6Y22_to_NB;
wire[3:0] Tile_X6Y22_to_NC;
wire[3:0] Tile_X6Y22_to_ND;
wire[3:0] Tile_X6Y22_to_NF;
wire[7:0] Tile_X6Y22_to_NG;
wire[7:0] Tile_X6Y22_to_NH;
wire[11:0] Tile_X6Y22_to_NI;
wire[3:0] Tile_X6Y22_to_SA;
wire[3:0] Tile_X6Y22_to_SB;
wire[3:0] Tile_X6Y22_to_SC;
wire[3:0] Tile_X6Y22_to_SD;
wire[3:0] Tile_X6Y22_to_SF;
wire[7:0] Tile_X6Y22_to_SG;
wire[7:0] Tile_X6Y22_to_SH;
wire[11:0] Tile_X6Y22_to_SI;
wire[3:0] Tile_X7Y22_to_EA;
wire[3:0] Tile_X7Y22_to_EB;
wire[3:0] Tile_X7Y22_to_EC;
wire[3:0] Tile_X7Y22_to_ED;
wire[3:0] Tile_X7Y22_to_EF;
wire[7:0] Tile_X7Y22_to_EG;
wire[7:0] Tile_X7Y22_to_EH;
wire[11:0] Tile_X7Y22_to_EI;
wire[3:0] Tile_X7Y22_to_WA;
wire[3:0] Tile_X7Y22_to_WB;
wire[3:0] Tile_X7Y22_to_WC;
wire[3:0] Tile_X7Y22_to_WD;
wire[3:0] Tile_X7Y22_to_WF;
wire[7:0] Tile_X7Y22_to_WG;
wire[7:0] Tile_X7Y22_to_WH;
wire[11:0] Tile_X7Y22_to_WI;
wire[3:0] Tile_X7Y22_to_NA;
wire[3:0] Tile_X7Y22_to_NB;
wire[3:0] Tile_X7Y22_to_NC;
wire[3:0] Tile_X7Y22_to_ND;
wire[3:0] Tile_X7Y22_to_NF;
wire[7:0] Tile_X7Y22_to_NG;
wire[7:0] Tile_X7Y22_to_NH;
wire[11:0] Tile_X7Y22_to_NI;
wire[3:0] Tile_X7Y22_to_SA;
wire[3:0] Tile_X7Y22_to_SB;
wire[3:0] Tile_X7Y22_to_SC;
wire[3:0] Tile_X7Y22_to_SD;
wire[3:0] Tile_X7Y22_to_SF;
wire[7:0] Tile_X7Y22_to_SG;
wire[7:0] Tile_X7Y22_to_SH;
wire[11:0] Tile_X7Y22_to_SI;
wire[3:0] Tile_X8Y22_to_WA;
wire[3:0] Tile_X8Y22_to_WB;
wire[3:0] Tile_X8Y22_to_WC;
wire[3:0] Tile_X8Y22_to_WD;
wire[3:0] Tile_X8Y22_to_WF;
wire[7:0] Tile_X8Y22_to_WG;
wire[7:0] Tile_X8Y22_to_WH;
wire[11:0] Tile_X8Y22_to_WI;
wire[3:0] Tile_X8Y22_to_NA;
wire[3:0] Tile_X8Y22_to_NB;
wire[3:0] Tile_X8Y22_to_NC;
wire[3:0] Tile_X8Y22_to_ND;
wire[3:0] Tile_X8Y22_to_NF;
wire[7:0] Tile_X8Y22_to_NG;
wire[7:0] Tile_X8Y22_to_NH;
wire[11:0] Tile_X8Y22_to_NI;
wire[3:0] Tile_X8Y22_to_SA;
wire[3:0] Tile_X8Y22_to_SB;
wire[3:0] Tile_X8Y22_to_SC;
wire[3:0] Tile_X8Y22_to_SD;
wire[3:0] Tile_X8Y22_to_SF;
wire[7:0] Tile_X8Y22_to_SG;
wire[7:0] Tile_X8Y22_to_SH;
wire[11:0] Tile_X8Y22_to_SI;
wire[1:0] Tile_X9Y22_to_EA_1s;
wire[1:0] Tile_X9Y22_to_EB_1s;
wire[1:0] Tile_X9Y22_to_EC_1s;
wire[1:0] Tile_X9Y22_to_ED_1s;
wire[1:0] Tile_X9Y22_to_EF_1s;
wire[1:0] Tile_X9Y22_to_EG_1s;
wire[1:0] Tile_X9Y22_to_EH_1s;
wire[1:0] Tile_X9Y22_to_EI_1s;
wire[1:0] Tile_X9Y22_to_WA_1s;
wire[1:0] Tile_X9Y22_to_WB_1s;
wire[1:0] Tile_X9Y22_to_WC_1s;
wire[1:0] Tile_X9Y22_to_WD_1s;
wire[1:0] Tile_X9Y22_to_WF_1s;
wire[1:0] Tile_X9Y22_to_WG_1s;
wire[1:0] Tile_X9Y22_to_WH_1s;
wire[1:0] Tile_X9Y22_to_WI_1s;
wire[1:0] Tile_X9Y22_to_NA_1s;
wire[1:0] Tile_X9Y22_to_NB_1s;
wire[1:0] Tile_X9Y22_to_NC_1s;
wire[1:0] Tile_X9Y22_to_ND_1s;
wire[1:0] Tile_X9Y22_to_NF_1s;
wire[1:0] Tile_X9Y22_to_NG_1s;
wire[1:0] Tile_X9Y22_to_NH_1s;
wire[1:0] Tile_X9Y22_to_NI_1s;
wire[1:0] Tile_X9Y22_to_SA_1s;
wire[1:0] Tile_X9Y22_to_SB_1s;
wire[1:0] Tile_X9Y22_to_SC_1s;
wire[1:0] Tile_X9Y22_to_SD_1s;
wire[1:0] Tile_X9Y22_to_SF_1s;
wire[1:0] Tile_X9Y22_to_SG_1s;
wire[1:0] Tile_X9Y22_to_SH_1s;
wire[1:0] Tile_X9Y22_to_SI_1s;
wire[1:0] Tile_X10Y22_to_WA_1s;
wire[1:0] Tile_X10Y22_to_WB_1s;
wire[1:0] Tile_X10Y22_to_WC_1s;
wire[1:0] Tile_X10Y22_to_WD_1s;
wire[1:0] Tile_X10Y22_to_WF_1s;
wire[1:0] Tile_X10Y22_to_WG_1s;
wire[1:0] Tile_X10Y22_to_WH_1s;
wire[1:0] Tile_X10Y22_to_WI_1s;
wire[3:0] Tile_X0Y23_to_EA;
wire[3:0] Tile_X0Y23_to_EB;
wire[3:0] Tile_X0Y23_to_EC;
wire[3:0] Tile_X0Y23_to_ED;
wire[3:0] Tile_X0Y23_to_EF;
wire[7:0] Tile_X0Y23_to_EG;
wire[7:0] Tile_X0Y23_to_EH;
wire[11:0] Tile_X0Y23_to_EI;
wire[3:0] Tile_X0Y23_to_NA;
wire[3:0] Tile_X0Y23_to_NB;
wire[3:0] Tile_X0Y23_to_NC;
wire[3:0] Tile_X0Y23_to_ND;
wire[3:0] Tile_X0Y23_to_NF;
wire[7:0] Tile_X0Y23_to_NG;
wire[7:0] Tile_X0Y23_to_NH;
wire[11:0] Tile_X0Y23_to_NI;
wire[3:0] Tile_X0Y23_to_SA;
wire[3:0] Tile_X0Y23_to_SB;
wire[3:0] Tile_X0Y23_to_SC;
wire[3:0] Tile_X0Y23_to_SD;
wire[3:0] Tile_X0Y23_to_SF;
wire[7:0] Tile_X0Y23_to_SG;
wire[7:0] Tile_X0Y23_to_SH;
wire[11:0] Tile_X0Y23_to_SI;
wire[3:0] Tile_X1Y23_to_EA;
wire[3:0] Tile_X1Y23_to_EB;
wire[3:0] Tile_X1Y23_to_EC;
wire[3:0] Tile_X1Y23_to_ED;
wire[3:0] Tile_X1Y23_to_EF;
wire[7:0] Tile_X1Y23_to_EG;
wire[7:0] Tile_X1Y23_to_EH;
wire[11:0] Tile_X1Y23_to_EI;
wire[3:0] Tile_X1Y23_to_WA;
wire[3:0] Tile_X1Y23_to_WB;
wire[3:0] Tile_X1Y23_to_WC;
wire[3:0] Tile_X1Y23_to_WD;
wire[3:0] Tile_X1Y23_to_WF;
wire[7:0] Tile_X1Y23_to_WG;
wire[7:0] Tile_X1Y23_to_WH;
wire[11:0] Tile_X1Y23_to_WI;
wire[3:0] Tile_X1Y23_to_NA;
wire[3:0] Tile_X1Y23_to_NB;
wire[3:0] Tile_X1Y23_to_NC;
wire[3:0] Tile_X1Y23_to_ND;
wire[3:0] Tile_X1Y23_to_NF;
wire[7:0] Tile_X1Y23_to_NG;
wire[7:0] Tile_X1Y23_to_NH;
wire[11:0] Tile_X1Y23_to_NI;
wire[3:0] Tile_X1Y23_to_SA;
wire[3:0] Tile_X1Y23_to_SB;
wire[3:0] Tile_X1Y23_to_SC;
wire[3:0] Tile_X1Y23_to_SD;
wire[3:0] Tile_X1Y23_to_SF;
wire[7:0] Tile_X1Y23_to_SG;
wire[7:0] Tile_X1Y23_to_SH;
wire[11:0] Tile_X1Y23_to_SI;
wire[3:0] Tile_X2Y23_to_EA;
wire[3:0] Tile_X2Y23_to_EB;
wire[3:0] Tile_X2Y23_to_EC;
wire[3:0] Tile_X2Y23_to_ED;
wire[3:0] Tile_X2Y23_to_EF;
wire[7:0] Tile_X2Y23_to_EG;
wire[7:0] Tile_X2Y23_to_EH;
wire[11:0] Tile_X2Y23_to_EI;
wire[3:0] Tile_X2Y23_to_WA;
wire[3:0] Tile_X2Y23_to_WB;
wire[3:0] Tile_X2Y23_to_WC;
wire[3:0] Tile_X2Y23_to_WD;
wire[3:0] Tile_X2Y23_to_WF;
wire[7:0] Tile_X2Y23_to_WG;
wire[7:0] Tile_X2Y23_to_WH;
wire[11:0] Tile_X2Y23_to_WI;
wire[3:0] Tile_X2Y23_to_NA;
wire[3:0] Tile_X2Y23_to_NB;
wire[3:0] Tile_X2Y23_to_NC;
wire[3:0] Tile_X2Y23_to_ND;
wire[3:0] Tile_X2Y23_to_NF;
wire[7:0] Tile_X2Y23_to_NG;
wire[7:0] Tile_X2Y23_to_NH;
wire[11:0] Tile_X2Y23_to_NI;
wire[3:0] Tile_X2Y23_to_SA;
wire[3:0] Tile_X2Y23_to_SB;
wire[3:0] Tile_X2Y23_to_SC;
wire[3:0] Tile_X2Y23_to_SD;
wire[3:0] Tile_X2Y23_to_SF;
wire[7:0] Tile_X2Y23_to_SG;
wire[7:0] Tile_X2Y23_to_SH;
wire[11:0] Tile_X2Y23_to_SI;
wire[3:0] Tile_X3Y23_to_EA;
wire[3:0] Tile_X3Y23_to_EB;
wire[3:0] Tile_X3Y23_to_EC;
wire[3:0] Tile_X3Y23_to_ED;
wire[3:0] Tile_X3Y23_to_EF;
wire[7:0] Tile_X3Y23_to_EG;
wire[7:0] Tile_X3Y23_to_EH;
wire[11:0] Tile_X3Y23_to_EI;
wire[3:0] Tile_X3Y23_to_WA;
wire[3:0] Tile_X3Y23_to_WB;
wire[3:0] Tile_X3Y23_to_WC;
wire[3:0] Tile_X3Y23_to_WD;
wire[3:0] Tile_X3Y23_to_WF;
wire[7:0] Tile_X3Y23_to_WG;
wire[7:0] Tile_X3Y23_to_WH;
wire[11:0] Tile_X3Y23_to_WI;
wire[3:0] Tile_X3Y23_to_NA;
wire[3:0] Tile_X3Y23_to_NB;
wire[3:0] Tile_X3Y23_to_NC;
wire[3:0] Tile_X3Y23_to_ND;
wire[3:0] Tile_X3Y23_to_NF;
wire[7:0] Tile_X3Y23_to_NG;
wire[7:0] Tile_X3Y23_to_NH;
wire[11:0] Tile_X3Y23_to_NI;
wire[3:0] Tile_X3Y23_to_SA;
wire[3:0] Tile_X3Y23_to_SB;
wire[3:0] Tile_X3Y23_to_SC;
wire[3:0] Tile_X3Y23_to_SD;
wire[3:0] Tile_X3Y23_to_SF;
wire[7:0] Tile_X3Y23_to_SG;
wire[7:0] Tile_X3Y23_to_SH;
wire[11:0] Tile_X3Y23_to_SI;
wire[3:0] Tile_X4Y23_to_EA;
wire[3:0] Tile_X4Y23_to_EB;
wire[3:0] Tile_X4Y23_to_EC;
wire[3:0] Tile_X4Y23_to_ED;
wire[3:0] Tile_X4Y23_to_EF;
wire[7:0] Tile_X4Y23_to_EG;
wire[7:0] Tile_X4Y23_to_EH;
wire[11:0] Tile_X4Y23_to_EI;
wire[3:0] Tile_X4Y23_to_WA;
wire[3:0] Tile_X4Y23_to_WB;
wire[3:0] Tile_X4Y23_to_WC;
wire[3:0] Tile_X4Y23_to_WD;
wire[3:0] Tile_X4Y23_to_WF;
wire[7:0] Tile_X4Y23_to_WG;
wire[7:0] Tile_X4Y23_to_WH;
wire[11:0] Tile_X4Y23_to_WI;
wire[3:0] Tile_X4Y23_to_NA;
wire[3:0] Tile_X4Y23_to_NB;
wire[3:0] Tile_X4Y23_to_NC;
wire[3:0] Tile_X4Y23_to_ND;
wire[3:0] Tile_X4Y23_to_NF;
wire[7:0] Tile_X4Y23_to_NG;
wire[7:0] Tile_X4Y23_to_NH;
wire[11:0] Tile_X4Y23_to_NI;
wire[3:0] Tile_X4Y23_to_SA;
wire[3:0] Tile_X4Y23_to_SB;
wire[3:0] Tile_X4Y23_to_SC;
wire[3:0] Tile_X4Y23_to_SD;
wire[3:0] Tile_X4Y23_to_SF;
wire[7:0] Tile_X4Y23_to_SG;
wire[7:0] Tile_X4Y23_to_SH;
wire[11:0] Tile_X4Y23_to_SI;
wire[3:0] Tile_X5Y23_to_EA;
wire[3:0] Tile_X5Y23_to_EB;
wire[3:0] Tile_X5Y23_to_EC;
wire[3:0] Tile_X5Y23_to_ED;
wire[3:0] Tile_X5Y23_to_EF;
wire[7:0] Tile_X5Y23_to_EG;
wire[7:0] Tile_X5Y23_to_EH;
wire[11:0] Tile_X5Y23_to_EI;
wire[3:0] Tile_X5Y23_to_WA;
wire[3:0] Tile_X5Y23_to_WB;
wire[3:0] Tile_X5Y23_to_WC;
wire[3:0] Tile_X5Y23_to_WD;
wire[3:0] Tile_X5Y23_to_WF;
wire[7:0] Tile_X5Y23_to_WG;
wire[7:0] Tile_X5Y23_to_WH;
wire[11:0] Tile_X5Y23_to_WI;
wire[3:0] Tile_X5Y23_to_NA;
wire[3:0] Tile_X5Y23_to_NB;
wire[3:0] Tile_X5Y23_to_NC;
wire[3:0] Tile_X5Y23_to_ND;
wire[3:0] Tile_X5Y23_to_NF;
wire[7:0] Tile_X5Y23_to_NG;
wire[7:0] Tile_X5Y23_to_NH;
wire[11:0] Tile_X5Y23_to_NI;
wire[3:0] Tile_X5Y23_to_SA;
wire[3:0] Tile_X5Y23_to_SB;
wire[3:0] Tile_X5Y23_to_SC;
wire[3:0] Tile_X5Y23_to_SD;
wire[3:0] Tile_X5Y23_to_SF;
wire[7:0] Tile_X5Y23_to_SG;
wire[7:0] Tile_X5Y23_to_SH;
wire[11:0] Tile_X5Y23_to_SI;
wire[3:0] Tile_X6Y23_to_EA;
wire[3:0] Tile_X6Y23_to_EB;
wire[3:0] Tile_X6Y23_to_EC;
wire[3:0] Tile_X6Y23_to_ED;
wire[3:0] Tile_X6Y23_to_EF;
wire[7:0] Tile_X6Y23_to_EG;
wire[7:0] Tile_X6Y23_to_EH;
wire[11:0] Tile_X6Y23_to_EI;
wire[3:0] Tile_X6Y23_to_WA;
wire[3:0] Tile_X6Y23_to_WB;
wire[3:0] Tile_X6Y23_to_WC;
wire[3:0] Tile_X6Y23_to_WD;
wire[3:0] Tile_X6Y23_to_WF;
wire[7:0] Tile_X6Y23_to_WG;
wire[7:0] Tile_X6Y23_to_WH;
wire[11:0] Tile_X6Y23_to_WI;
wire[3:0] Tile_X6Y23_to_NA;
wire[3:0] Tile_X6Y23_to_NB;
wire[3:0] Tile_X6Y23_to_NC;
wire[3:0] Tile_X6Y23_to_ND;
wire[3:0] Tile_X6Y23_to_NF;
wire[7:0] Tile_X6Y23_to_NG;
wire[7:0] Tile_X6Y23_to_NH;
wire[11:0] Tile_X6Y23_to_NI;
wire[3:0] Tile_X6Y23_to_SA;
wire[3:0] Tile_X6Y23_to_SB;
wire[3:0] Tile_X6Y23_to_SC;
wire[3:0] Tile_X6Y23_to_SD;
wire[3:0] Tile_X6Y23_to_SF;
wire[7:0] Tile_X6Y23_to_SG;
wire[7:0] Tile_X6Y23_to_SH;
wire[11:0] Tile_X6Y23_to_SI;
wire[3:0] Tile_X7Y23_to_EA;
wire[3:0] Tile_X7Y23_to_EB;
wire[3:0] Tile_X7Y23_to_EC;
wire[3:0] Tile_X7Y23_to_ED;
wire[3:0] Tile_X7Y23_to_EF;
wire[7:0] Tile_X7Y23_to_EG;
wire[7:0] Tile_X7Y23_to_EH;
wire[11:0] Tile_X7Y23_to_EI;
wire[3:0] Tile_X7Y23_to_WA;
wire[3:0] Tile_X7Y23_to_WB;
wire[3:0] Tile_X7Y23_to_WC;
wire[3:0] Tile_X7Y23_to_WD;
wire[3:0] Tile_X7Y23_to_WF;
wire[7:0] Tile_X7Y23_to_WG;
wire[7:0] Tile_X7Y23_to_WH;
wire[11:0] Tile_X7Y23_to_WI;
wire[3:0] Tile_X7Y23_to_NA;
wire[3:0] Tile_X7Y23_to_NB;
wire[3:0] Tile_X7Y23_to_NC;
wire[3:0] Tile_X7Y23_to_ND;
wire[3:0] Tile_X7Y23_to_NF;
wire[7:0] Tile_X7Y23_to_NG;
wire[7:0] Tile_X7Y23_to_NH;
wire[11:0] Tile_X7Y23_to_NI;
wire[3:0] Tile_X7Y23_to_SA;
wire[3:0] Tile_X7Y23_to_SB;
wire[3:0] Tile_X7Y23_to_SC;
wire[3:0] Tile_X7Y23_to_SD;
wire[3:0] Tile_X7Y23_to_SF;
wire[7:0] Tile_X7Y23_to_SG;
wire[7:0] Tile_X7Y23_to_SH;
wire[11:0] Tile_X7Y23_to_SI;
wire[3:0] Tile_X8Y23_to_WA;
wire[3:0] Tile_X8Y23_to_WB;
wire[3:0] Tile_X8Y23_to_WC;
wire[3:0] Tile_X8Y23_to_WD;
wire[3:0] Tile_X8Y23_to_WF;
wire[7:0] Tile_X8Y23_to_WG;
wire[7:0] Tile_X8Y23_to_WH;
wire[11:0] Tile_X8Y23_to_WI;
wire[3:0] Tile_X8Y23_to_NA;
wire[3:0] Tile_X8Y23_to_NB;
wire[3:0] Tile_X8Y23_to_NC;
wire[3:0] Tile_X8Y23_to_ND;
wire[3:0] Tile_X8Y23_to_NF;
wire[7:0] Tile_X8Y23_to_NG;
wire[7:0] Tile_X8Y23_to_NH;
wire[11:0] Tile_X8Y23_to_NI;
wire[3:0] Tile_X8Y23_to_SA;
wire[3:0] Tile_X8Y23_to_SB;
wire[3:0] Tile_X8Y23_to_SC;
wire[3:0] Tile_X8Y23_to_SD;
wire[3:0] Tile_X8Y23_to_SF;
wire[7:0] Tile_X8Y23_to_SG;
wire[7:0] Tile_X8Y23_to_SH;
wire[11:0] Tile_X8Y23_to_SI;
wire[1:0] Tile_X9Y23_to_EA_1s;
wire[1:0] Tile_X9Y23_to_EB_1s;
wire[1:0] Tile_X9Y23_to_EC_1s;
wire[1:0] Tile_X9Y23_to_ED_1s;
wire[1:0] Tile_X9Y23_to_EF_1s;
wire[1:0] Tile_X9Y23_to_EG_1s;
wire[1:0] Tile_X9Y23_to_EH_1s;
wire[1:0] Tile_X9Y23_to_EI_1s;
wire[1:0] Tile_X9Y23_to_WA_1s;
wire[1:0] Tile_X9Y23_to_WB_1s;
wire[1:0] Tile_X9Y23_to_WC_1s;
wire[1:0] Tile_X9Y23_to_WD_1s;
wire[1:0] Tile_X9Y23_to_WF_1s;
wire[1:0] Tile_X9Y23_to_WG_1s;
wire[1:0] Tile_X9Y23_to_WH_1s;
wire[1:0] Tile_X9Y23_to_WI_1s;
wire[1:0] Tile_X9Y23_to_NA_1s;
wire[1:0] Tile_X9Y23_to_NB_1s;
wire[1:0] Tile_X9Y23_to_NC_1s;
wire[1:0] Tile_X9Y23_to_ND_1s;
wire[1:0] Tile_X9Y23_to_NF_1s;
wire[1:0] Tile_X9Y23_to_NG_1s;
wire[1:0] Tile_X9Y23_to_NH_1s;
wire[1:0] Tile_X9Y23_to_NI_1s;
wire[1:0] Tile_X9Y23_to_SA_1s;
wire[1:0] Tile_X9Y23_to_SB_1s;
wire[1:0] Tile_X9Y23_to_SC_1s;
wire[1:0] Tile_X9Y23_to_SD_1s;
wire[1:0] Tile_X9Y23_to_SF_1s;
wire[1:0] Tile_X9Y23_to_SG_1s;
wire[1:0] Tile_X9Y23_to_SH_1s;
wire[1:0] Tile_X9Y23_to_SI_1s;
wire[1:0] Tile_X10Y23_to_WA_1s;
wire[1:0] Tile_X10Y23_to_WB_1s;
wire[1:0] Tile_X10Y23_to_WC_1s;
wire[1:0] Tile_X10Y23_to_WD_1s;
wire[1:0] Tile_X10Y23_to_WF_1s;
wire[1:0] Tile_X10Y23_to_WG_1s;
wire[1:0] Tile_X10Y23_to_WH_1s;
wire[1:0] Tile_X10Y23_to_WI_1s;
wire[3:0] Tile_X0Y24_to_NA;
wire[3:0] Tile_X0Y24_to_NB;
wire[3:0] Tile_X0Y24_to_NC;
wire[3:0] Tile_X0Y24_to_ND;
wire[3:0] Tile_X0Y24_to_NF;
wire[7:0] Tile_X0Y24_to_NG;
wire[7:0] Tile_X0Y24_to_NH;
wire[11:0] Tile_X0Y24_to_NI;
wire[3:0] Tile_X1Y24_to_NA;
wire[3:0] Tile_X1Y24_to_NB;
wire[3:0] Tile_X1Y24_to_NC;
wire[3:0] Tile_X1Y24_to_ND;
wire[3:0] Tile_X1Y24_to_NF;
wire[7:0] Tile_X1Y24_to_NG;
wire[7:0] Tile_X1Y24_to_NH;
wire[11:0] Tile_X1Y24_to_NI;
wire[3:0] Tile_X2Y24_to_NA;
wire[3:0] Tile_X2Y24_to_NB;
wire[3:0] Tile_X2Y24_to_NC;
wire[3:0] Tile_X2Y24_to_ND;
wire[3:0] Tile_X2Y24_to_NF;
wire[7:0] Tile_X2Y24_to_NG;
wire[7:0] Tile_X2Y24_to_NH;
wire[11:0] Tile_X2Y24_to_NI;
wire[3:0] Tile_X3Y24_to_NA;
wire[3:0] Tile_X3Y24_to_NB;
wire[3:0] Tile_X3Y24_to_NC;
wire[3:0] Tile_X3Y24_to_ND;
wire[3:0] Tile_X3Y24_to_NF;
wire[7:0] Tile_X3Y24_to_NG;
wire[7:0] Tile_X3Y24_to_NH;
wire[11:0] Tile_X3Y24_to_NI;
wire[3:0] Tile_X4Y24_to_NA;
wire[3:0] Tile_X4Y24_to_NB;
wire[3:0] Tile_X4Y24_to_NC;
wire[3:0] Tile_X4Y24_to_ND;
wire[3:0] Tile_X4Y24_to_NF;
wire[7:0] Tile_X4Y24_to_NG;
wire[7:0] Tile_X4Y24_to_NH;
wire[11:0] Tile_X4Y24_to_NI;
wire[3:0] Tile_X5Y24_to_NA;
wire[3:0] Tile_X5Y24_to_NB;
wire[3:0] Tile_X5Y24_to_NC;
wire[3:0] Tile_X5Y24_to_ND;
wire[3:0] Tile_X5Y24_to_NF;
wire[7:0] Tile_X5Y24_to_NG;
wire[7:0] Tile_X5Y24_to_NH;
wire[11:0] Tile_X5Y24_to_NI;
wire[3:0] Tile_X6Y24_to_NA;
wire[3:0] Tile_X6Y24_to_NB;
wire[3:0] Tile_X6Y24_to_NC;
wire[3:0] Tile_X6Y24_to_ND;
wire[3:0] Tile_X6Y24_to_NF;
wire[7:0] Tile_X6Y24_to_NG;
wire[7:0] Tile_X6Y24_to_NH;
wire[11:0] Tile_X6Y24_to_NI;
wire[3:0] Tile_X7Y24_to_NA;
wire[3:0] Tile_X7Y24_to_NB;
wire[3:0] Tile_X7Y24_to_NC;
wire[3:0] Tile_X7Y24_to_ND;
wire[3:0] Tile_X7Y24_to_NF;
wire[7:0] Tile_X7Y24_to_NG;
wire[7:0] Tile_X7Y24_to_NH;
wire[11:0] Tile_X7Y24_to_NI;
wire[3:0] Tile_X8Y24_to_NA;
wire[3:0] Tile_X8Y24_to_NB;
wire[3:0] Tile_X8Y24_to_NC;
wire[3:0] Tile_X8Y24_to_ND;
wire[3:0] Tile_X8Y24_to_NF;
wire[7:0] Tile_X8Y24_to_NG;
wire[7:0] Tile_X8Y24_to_NH;
wire[11:0] Tile_X8Y24_to_NI;
wire[1:0] Tile_X9Y24_to_NA_1s;
wire[1:0] Tile_X9Y24_to_NB_1s;
wire[1:0] Tile_X9Y24_to_NC_1s;
wire[1:0] Tile_X9Y24_to_ND_1s;
wire[1:0] Tile_X9Y24_to_NF_1s;
wire[1:0] Tile_X9Y24_to_NG_1s;
wire[1:0] Tile_X9Y24_to_NH_1s;
wire[1:0] Tile_X9Y24_to_NI_1s;
wire[1:0] Tile_X10Y24_to_NA_1s;
wire[1:0] Tile_X10Y24_to_NB_1s;
wire[1:0] Tile_X10Y24_to_NC_1s;
wire[1:0] Tile_X10Y24_to_ND_1s;
wire[1:0] Tile_X10Y24_to_NF_1s;
wire[1:0] Tile_X10Y24_to_NG_1s;
wire[1:0] Tile_X10Y24_to_NH_1s;
wire[1:0] Tile_X10Y24_to_NI_1s;

assign Tile_Y1_FrameData = FrameData[FrameBitsPerRow*(1+1)-1:FrameBitsPerRow*1];
assign Tile_Y2_FrameData = FrameData[FrameBitsPerRow*(2+1)-1:FrameBitsPerRow*2];
assign Tile_Y3_FrameData = FrameData[FrameBitsPerRow*(3+1)-1:FrameBitsPerRow*3];
assign Tile_Y4_FrameData = FrameData[FrameBitsPerRow*(4+1)-1:FrameBitsPerRow*4];
assign Tile_Y5_FrameData = FrameData[FrameBitsPerRow*(5+1)-1:FrameBitsPerRow*5];
assign Tile_Y6_FrameData = FrameData[FrameBitsPerRow*(6+1)-1:FrameBitsPerRow*6];
assign Tile_Y7_FrameData = FrameData[FrameBitsPerRow*(7+1)-1:FrameBitsPerRow*7];
assign Tile_Y8_FrameData = FrameData[FrameBitsPerRow*(8+1)-1:FrameBitsPerRow*8];
assign Tile_Y9_FrameData = FrameData[FrameBitsPerRow*(9+1)-1:FrameBitsPerRow*9];
assign Tile_Y10_FrameData = FrameData[FrameBitsPerRow*(10+1)-1:FrameBitsPerRow*10];
assign Tile_Y11_FrameData = FrameData[FrameBitsPerRow*(11+1)-1:FrameBitsPerRow*11];
assign Tile_Y12_FrameData = FrameData[FrameBitsPerRow*(12+1)-1:FrameBitsPerRow*12];
assign Tile_Y13_FrameData = FrameData[FrameBitsPerRow*(13+1)-1:FrameBitsPerRow*13];
assign Tile_Y14_FrameData = FrameData[FrameBitsPerRow*(14+1)-1:FrameBitsPerRow*14];
assign Tile_Y15_FrameData = FrameData[FrameBitsPerRow*(15+1)-1:FrameBitsPerRow*15];
assign Tile_Y16_FrameData = FrameData[FrameBitsPerRow*(16+1)-1:FrameBitsPerRow*16];
assign Tile_Y17_FrameData = FrameData[FrameBitsPerRow*(17+1)-1:FrameBitsPerRow*17];
assign Tile_Y18_FrameData = FrameData[FrameBitsPerRow*(18+1)-1:FrameBitsPerRow*18];
assign Tile_Y19_FrameData = FrameData[FrameBitsPerRow*(19+1)-1:FrameBitsPerRow*19];
assign Tile_Y20_FrameData = FrameData[FrameBitsPerRow*(20+1)-1:FrameBitsPerRow*20];
assign Tile_Y21_FrameData = FrameData[FrameBitsPerRow*(21+1)-1:FrameBitsPerRow*21];
assign Tile_Y22_FrameData = FrameData[FrameBitsPerRow*(22+1)-1:FrameBitsPerRow*22];
assign Tile_Y23_FrameData = FrameData[FrameBitsPerRow*(23+1)-1:FrameBitsPerRow*23];
assign Tile_X0_FrameStrobe = FrameStrobe[MaxFramesPerCol*(0+1)-1:MaxFramesPerCol*0];
assign Tile_X1_FrameStrobe = FrameStrobe[MaxFramesPerCol*(1+1)-1:MaxFramesPerCol*1];
assign Tile_X2_FrameStrobe = FrameStrobe[MaxFramesPerCol*(2+1)-1:MaxFramesPerCol*2];
assign Tile_X3_FrameStrobe = FrameStrobe[MaxFramesPerCol*(3+1)-1:MaxFramesPerCol*3];
assign Tile_X4_FrameStrobe = FrameStrobe[MaxFramesPerCol*(4+1)-1:MaxFramesPerCol*4];
assign Tile_X5_FrameStrobe = FrameStrobe[MaxFramesPerCol*(5+1)-1:MaxFramesPerCol*5];
assign Tile_X6_FrameStrobe = FrameStrobe[MaxFramesPerCol*(6+1)-1:MaxFramesPerCol*6];
assign Tile_X7_FrameStrobe = FrameStrobe[MaxFramesPerCol*(7+1)-1:MaxFramesPerCol*7];
assign Tile_X8_FrameStrobe = FrameStrobe[MaxFramesPerCol*(8+1)-1:MaxFramesPerCol*8];
assign Tile_X9_FrameStrobe = FrameStrobe[MaxFramesPerCol*(9+1)-1:MaxFramesPerCol*9];
assign Tile_X10_FrameStrobe = FrameStrobe[MaxFramesPerCol*(10+1)-1:MaxFramesPerCol*10];

 //tile IO port will get directly connected to top-level tile module
N_term_custom Tile_X0Y0_N_term_custom (
    .from_NA(Tile_X0Y1_to_NA),
    .from_NB(Tile_X0Y1_to_NB),
    .from_NC(Tile_X0Y1_to_NC),
    .from_ND(Tile_X0Y1_to_ND),
    .from_NF(Tile_X0Y1_to_NF),
    .from_NG(Tile_X0Y1_to_NG),
    .from_NH(Tile_X0Y1_to_NH),
    .from_NI(Tile_X0Y1_to_NI),
    .to_SA(Tile_X0Y0_to_SA),
    .to_SB(Tile_X0Y0_to_SB),
    .to_SC(Tile_X0Y0_to_SC),
    .to_SD(Tile_X0Y0_to_SD),
    .to_SF(Tile_X0Y0_to_SF),
    .to_SG(Tile_X0Y0_to_SG),
    .to_SH(Tile_X0Y0_to_SH),
    .to_SI(Tile_X0Y0_to_SI),
    .UserCLK(Tile_X0Y1_UserCLKo),
    .UserCLKo(Tile_X0Y0_UserCLKo),
    .rst(Tile_X0Y1_rsto),
    .rsto(Tile_X0Y0_rsto),
    .FrameStrobe(Tile_X0Y1_FrameStrobe_O),
    .FrameStrobe_O(Tile_X0Y0_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
N_term_custom Tile_X1Y0_N_term_custom (
    .from_NA(Tile_X1Y1_to_NA),
    .from_NB(Tile_X1Y1_to_NB),
    .from_NC(Tile_X1Y1_to_NC),
    .from_ND(Tile_X1Y1_to_ND),
    .from_NF(Tile_X1Y1_to_NF),
    .from_NG(Tile_X1Y1_to_NG),
    .from_NH(Tile_X1Y1_to_NH),
    .from_NI(Tile_X1Y1_to_NI),
    .to_SA(Tile_X1Y0_to_SA),
    .to_SB(Tile_X1Y0_to_SB),
    .to_SC(Tile_X1Y0_to_SC),
    .to_SD(Tile_X1Y0_to_SD),
    .to_SF(Tile_X1Y0_to_SF),
    .to_SG(Tile_X1Y0_to_SG),
    .to_SH(Tile_X1Y0_to_SH),
    .to_SI(Tile_X1Y0_to_SI),
    .UserCLK(Tile_X1Y1_UserCLKo),
    .UserCLKo(Tile_X1Y0_UserCLKo),
    .rst(Tile_X1Y1_rsto),
    .rsto(Tile_X1Y0_rsto),
    .FrameStrobe(Tile_X1Y1_FrameStrobe_O),
    .FrameStrobe_O(Tile_X1Y0_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
N_term_custom Tile_X2Y0_N_term_custom (
    .from_NA(Tile_X2Y1_to_NA),
    .from_NB(Tile_X2Y1_to_NB),
    .from_NC(Tile_X2Y1_to_NC),
    .from_ND(Tile_X2Y1_to_ND),
    .from_NF(Tile_X2Y1_to_NF),
    .from_NG(Tile_X2Y1_to_NG),
    .from_NH(Tile_X2Y1_to_NH),
    .from_NI(Tile_X2Y1_to_NI),
    .to_SA(Tile_X2Y0_to_SA),
    .to_SB(Tile_X2Y0_to_SB),
    .to_SC(Tile_X2Y0_to_SC),
    .to_SD(Tile_X2Y0_to_SD),
    .to_SF(Tile_X2Y0_to_SF),
    .to_SG(Tile_X2Y0_to_SG),
    .to_SH(Tile_X2Y0_to_SH),
    .to_SI(Tile_X2Y0_to_SI),
    .UserCLK(Tile_X2Y1_UserCLKo),
    .UserCLKo(Tile_X2Y0_UserCLKo),
    .rst(Tile_X2Y1_rsto),
    .rsto(Tile_X2Y0_rsto),
    .FrameStrobe(Tile_X2Y1_FrameStrobe_O),
    .FrameStrobe_O(Tile_X2Y0_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
N_term_custom Tile_X3Y0_N_term_custom (
    .from_NA(Tile_X3Y1_to_NA),
    .from_NB(Tile_X3Y1_to_NB),
    .from_NC(Tile_X3Y1_to_NC),
    .from_ND(Tile_X3Y1_to_ND),
    .from_NF(Tile_X3Y1_to_NF),
    .from_NG(Tile_X3Y1_to_NG),
    .from_NH(Tile_X3Y1_to_NH),
    .from_NI(Tile_X3Y1_to_NI),
    .to_SA(Tile_X3Y0_to_SA),
    .to_SB(Tile_X3Y0_to_SB),
    .to_SC(Tile_X3Y0_to_SC),
    .to_SD(Tile_X3Y0_to_SD),
    .to_SF(Tile_X3Y0_to_SF),
    .to_SG(Tile_X3Y0_to_SG),
    .to_SH(Tile_X3Y0_to_SH),
    .to_SI(Tile_X3Y0_to_SI),
    .UserCLK(Tile_X3Y1_UserCLKo),
    .UserCLKo(Tile_X3Y0_UserCLKo),
    .rst(Tile_X3Y1_rsto),
    .rsto(Tile_X3Y0_rsto),
    .FrameStrobe(Tile_X3Y1_FrameStrobe_O),
    .FrameStrobe_O(Tile_X3Y0_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
N_term_custom Tile_X4Y0_N_term_custom (
    .from_NA(Tile_X4Y1_to_NA),
    .from_NB(Tile_X4Y1_to_NB),
    .from_NC(Tile_X4Y1_to_NC),
    .from_ND(Tile_X4Y1_to_ND),
    .from_NF(Tile_X4Y1_to_NF),
    .from_NG(Tile_X4Y1_to_NG),
    .from_NH(Tile_X4Y1_to_NH),
    .from_NI(Tile_X4Y1_to_NI),
    .to_SA(Tile_X4Y0_to_SA),
    .to_SB(Tile_X4Y0_to_SB),
    .to_SC(Tile_X4Y0_to_SC),
    .to_SD(Tile_X4Y0_to_SD),
    .to_SF(Tile_X4Y0_to_SF),
    .to_SG(Tile_X4Y0_to_SG),
    .to_SH(Tile_X4Y0_to_SH),
    .to_SI(Tile_X4Y0_to_SI),
    .UserCLK(Tile_X4Y1_UserCLKo),
    .UserCLKo(Tile_X4Y0_UserCLKo),
    .rst(Tile_X4Y1_rsto),
    .rsto(Tile_X4Y0_rsto),
    .FrameStrobe(Tile_X4Y1_FrameStrobe_O),
    .FrameStrobe_O(Tile_X4Y0_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
N_term_custom Tile_X5Y0_N_term_custom (
    .from_NA(Tile_X5Y1_to_NA),
    .from_NB(Tile_X5Y1_to_NB),
    .from_NC(Tile_X5Y1_to_NC),
    .from_ND(Tile_X5Y1_to_ND),
    .from_NF(Tile_X5Y1_to_NF),
    .from_NG(Tile_X5Y1_to_NG),
    .from_NH(Tile_X5Y1_to_NH),
    .from_NI(Tile_X5Y1_to_NI),
    .to_SA(Tile_X5Y0_to_SA),
    .to_SB(Tile_X5Y0_to_SB),
    .to_SC(Tile_X5Y0_to_SC),
    .to_SD(Tile_X5Y0_to_SD),
    .to_SF(Tile_X5Y0_to_SF),
    .to_SG(Tile_X5Y0_to_SG),
    .to_SH(Tile_X5Y0_to_SH),
    .to_SI(Tile_X5Y0_to_SI),
    .UserCLK(Tile_X5Y1_UserCLKo),
    .UserCLKo(Tile_X5Y0_UserCLKo),
    .rst(Tile_X5Y1_rsto),
    .rsto(Tile_X5Y0_rsto),
    .FrameStrobe(Tile_X5Y1_FrameStrobe_O),
    .FrameStrobe_O(Tile_X5Y0_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
N_term_custom Tile_X6Y0_N_term_custom (
    .from_NA(Tile_X6Y1_to_NA),
    .from_NB(Tile_X6Y1_to_NB),
    .from_NC(Tile_X6Y1_to_NC),
    .from_ND(Tile_X6Y1_to_ND),
    .from_NF(Tile_X6Y1_to_NF),
    .from_NG(Tile_X6Y1_to_NG),
    .from_NH(Tile_X6Y1_to_NH),
    .from_NI(Tile_X6Y1_to_NI),
    .to_SA(Tile_X6Y0_to_SA),
    .to_SB(Tile_X6Y0_to_SB),
    .to_SC(Tile_X6Y0_to_SC),
    .to_SD(Tile_X6Y0_to_SD),
    .to_SF(Tile_X6Y0_to_SF),
    .to_SG(Tile_X6Y0_to_SG),
    .to_SH(Tile_X6Y0_to_SH),
    .to_SI(Tile_X6Y0_to_SI),
    .UserCLK(Tile_X6Y1_UserCLKo),
    .UserCLKo(Tile_X6Y0_UserCLKo),
    .rst(Tile_X6Y1_rsto),
    .rsto(Tile_X6Y0_rsto),
    .FrameStrobe(Tile_X6Y1_FrameStrobe_O),
    .FrameStrobe_O(Tile_X6Y0_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
N_term_custom Tile_X7Y0_N_term_custom (
    .from_NA(Tile_X7Y1_to_NA),
    .from_NB(Tile_X7Y1_to_NB),
    .from_NC(Tile_X7Y1_to_NC),
    .from_ND(Tile_X7Y1_to_ND),
    .from_NF(Tile_X7Y1_to_NF),
    .from_NG(Tile_X7Y1_to_NG),
    .from_NH(Tile_X7Y1_to_NH),
    .from_NI(Tile_X7Y1_to_NI),
    .to_SA(Tile_X7Y0_to_SA),
    .to_SB(Tile_X7Y0_to_SB),
    .to_SC(Tile_X7Y0_to_SC),
    .to_SD(Tile_X7Y0_to_SD),
    .to_SF(Tile_X7Y0_to_SF),
    .to_SG(Tile_X7Y0_to_SG),
    .to_SH(Tile_X7Y0_to_SH),
    .to_SI(Tile_X7Y0_to_SI),
    .UserCLK(Tile_X7Y1_UserCLKo),
    .UserCLKo(Tile_X7Y0_UserCLKo),
    .rst(Tile_X7Y1_rsto),
    .rsto(Tile_X7Y0_rsto),
    .FrameStrobe(Tile_X7Y1_FrameStrobe_O),
    .FrameStrobe_O(Tile_X7Y0_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
N_term_custom Tile_X8Y0_N_term_custom (
    .from_NA(Tile_X8Y1_to_NA),
    .from_NB(Tile_X8Y1_to_NB),
    .from_NC(Tile_X8Y1_to_NC),
    .from_ND(Tile_X8Y1_to_ND),
    .from_NF(Tile_X8Y1_to_NF),
    .from_NG(Tile_X8Y1_to_NG),
    .from_NH(Tile_X8Y1_to_NH),
    .from_NI(Tile_X8Y1_to_NI),
    .to_SA(Tile_X8Y0_to_SA),
    .to_SB(Tile_X8Y0_to_SB),
    .to_SC(Tile_X8Y0_to_SC),
    .to_SD(Tile_X8Y0_to_SD),
    .to_SF(Tile_X8Y0_to_SF),
    .to_SG(Tile_X8Y0_to_SG),
    .to_SH(Tile_X8Y0_to_SH),
    .to_SI(Tile_X8Y0_to_SI),
    .UserCLK(Tile_X8Y1_UserCLKo),
    .UserCLKo(Tile_X8Y0_UserCLKo),
    .rst(Tile_X8Y1_rsto),
    .rsto(Tile_X8Y0_rsto),
    .FrameStrobe(Tile_X8Y1_FrameStrobe_O),
    .FrameStrobe_O(Tile_X8Y0_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
N_term_s1 Tile_X9Y0_N_term_s1 (
    .from_NA_1s(Tile_X9Y1_to_NA_1s),
    .from_NB_1s(Tile_X9Y1_to_NB_1s),
    .from_NC_1s(Tile_X9Y1_to_NC_1s),
    .from_ND_1s(Tile_X9Y1_to_ND_1s),
    .from_NF_1s(Tile_X9Y1_to_NF_1s),
    .from_NG_1s(Tile_X9Y1_to_NG_1s),
    .from_NH_1s(Tile_X9Y1_to_NH_1s),
    .from_NI_1s(Tile_X9Y1_to_NI_1s),
    .to_SA_1s(Tile_X9Y0_to_SA_1s),
    .to_SB_1s(Tile_X9Y0_to_SB_1s),
    .to_SC_1s(Tile_X9Y0_to_SC_1s),
    .to_SD_1s(Tile_X9Y0_to_SD_1s),
    .to_SF_1s(Tile_X9Y0_to_SF_1s),
    .to_SG_1s(Tile_X9Y0_to_SG_1s),
    .to_SH_1s(Tile_X9Y0_to_SH_1s),
    .to_SI_1s(Tile_X9Y0_to_SI_1s),
    .UserCLK(Tile_X9Y1_UserCLKo),
    .UserCLKo(Tile_X9Y0_UserCLKo),
    .rst(Tile_X9Y1_rsto),
    .rsto(Tile_X9Y0_rsto),
    .FrameStrobe(Tile_X9Y1_FrameStrobe_O),
    .FrameStrobe_O(Tile_X9Y0_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
N_term_s1 Tile_X10Y0_N_term_s1 (
    .to_SA_1s(Tile_X10Y0_to_SA_1s),
    .to_SB_1s(Tile_X10Y0_to_SB_1s),
    .to_SC_1s(Tile_X10Y0_to_SC_1s),
    .to_SD_1s(Tile_X10Y0_to_SD_1s),
    .to_SF_1s(Tile_X10Y0_to_SF_1s),
    .to_SG_1s(Tile_X10Y0_to_SG_1s),
    .to_SH_1s(Tile_X10Y0_to_SH_1s),
    .to_SI_1s(Tile_X10Y0_to_SI_1s),
    .UserCLK(Tile_X10Y1_UserCLKo),
    .UserCLKo(Tile_X10Y0_UserCLKo),
    .rst(Tile_X10Y1_rsto),
    .rsto(Tile_X10Y0_rsto),
    .FrameStrobe(Tile_X10Y1_FrameStrobe_O),
    .FrameStrobe_O(Tile_X10Y0_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
W_IO_custom
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X0Y1_Emulate_Bitstream)
    )
`endif
    Tile_X0Y1_W_IO_custom
    (
    .from_NA(Tile_X0Y2_to_NA),
    .from_NB(Tile_X0Y2_to_NB),
    .from_NC(Tile_X0Y2_to_NC),
    .from_ND(Tile_X0Y2_to_ND),
    .from_NF(Tile_X0Y2_to_NF),
    .from_NG(Tile_X0Y2_to_NG),
    .from_NH(Tile_X0Y2_to_NH),
    .from_NI(Tile_X0Y2_to_NI),
    .from_SA(Tile_X0Y0_to_SA),
    .from_SB(Tile_X0Y0_to_SB),
    .from_SC(Tile_X0Y0_to_SC),
    .from_SD(Tile_X0Y0_to_SD),
    .from_SF(Tile_X0Y0_to_SF),
    .from_SG(Tile_X0Y0_to_SG),
    .from_SH(Tile_X0Y0_to_SH),
    .from_SI(Tile_X0Y0_to_SI),
    .from_WA(Tile_X1Y1_to_WA),
    .from_WB(Tile_X1Y1_to_WB),
    .from_WC(Tile_X1Y1_to_WC),
    .from_WD(Tile_X1Y1_to_WD),
    .from_WF(Tile_X1Y1_to_WF),
    .from_WG(Tile_X1Y1_to_WG),
    .from_WH(Tile_X1Y1_to_WH),
    .from_WI(Tile_X1Y1_to_WI),
    .to_EA(Tile_X0Y1_to_EA),
    .to_EB(Tile_X0Y1_to_EB),
    .to_EC(Tile_X0Y1_to_EC),
    .to_ED(Tile_X0Y1_to_ED),
    .to_EF(Tile_X0Y1_to_EF),
    .to_EG(Tile_X0Y1_to_EG),
    .to_EH(Tile_X0Y1_to_EH),
    .to_EI(Tile_X0Y1_to_EI),
    .to_NA(Tile_X0Y1_to_NA),
    .to_NB(Tile_X0Y1_to_NB),
    .to_NC(Tile_X0Y1_to_NC),
    .to_ND(Tile_X0Y1_to_ND),
    .to_NF(Tile_X0Y1_to_NF),
    .to_NG(Tile_X0Y1_to_NG),
    .to_NH(Tile_X0Y1_to_NH),
    .to_NI(Tile_X0Y1_to_NI),
    .to_SA(Tile_X0Y1_to_SA),
    .to_SB(Tile_X0Y1_to_SB),
    .to_SC(Tile_X0Y1_to_SC),
    .to_SD(Tile_X0Y1_to_SD),
    .to_SF(Tile_X0Y1_to_SF),
    .to_SG(Tile_X0Y1_to_SG),
    .to_SH(Tile_X0Y1_to_SH),
    .to_SI(Tile_X0Y1_to_SI),
    .A_O_top_0_t(Tile_X0Y1_A_O_top_0_t),
    .A_O_top_0_f(Tile_X0Y1_A_O_top_0_f),
    .A_O_top_1_t(Tile_X0Y1_A_O_top_1_t),
    .A_O_top_1_f(Tile_X0Y1_A_O_top_1_f),
    .A_prech1(Tile_X0Y1_A_prech1),
    .A_prech2(Tile_X0Y1_A_prech2),
    .A_DR_fault(Tile_X0Y1_A_DR_fault),
    .A_I_top_0_t(Tile_X0Y1_A_I_top_0_t),
    .A_I_top_0_f(Tile_X0Y1_A_I_top_0_f),
    .A_I_top_1_t(Tile_X0Y1_A_I_top_1_t),
    .A_I_top_1_f(Tile_X0Y1_A_I_top_1_f),
    .A_T_top(Tile_X0Y1_A_T_top),
    .A_F_masked1(Tile_X0Y1_A_F_masked1),
    .A_F_masked2(Tile_X0Y1_A_F_masked2),
    .A_config_C_bit0(Tile_X0Y1_A_config_C_bit0),
    .A_config_C_bit1(Tile_X0Y1_A_config_C_bit1),
    .A_config_C_bit2(Tile_X0Y1_A_config_C_bit2),
    .A_config_C_bit3(Tile_X0Y1_A_config_C_bit3),
    .B_config_C_bit0(Tile_X0Y1_B_config_C_bit0),
    .B_config_C_bit1(Tile_X0Y1_B_config_C_bit1),
    .B_config_C_bit2(Tile_X0Y1_B_config_C_bit2),
    .B_config_C_bit3(Tile_X0Y1_B_config_C_bit3),
    .UserCLK(Tile_X0Y2_UserCLKo),
    .UserCLKo(Tile_X0Y1_UserCLKo),
    .rst(Tile_X0Y2_rsto),
    .rsto(Tile_X0Y1_rsto),
    .FrameData(Tile_Y1_FrameData),
    .FrameData_O(Tile_X0Y1_FrameData_O),
    .FrameStrobe(Tile_X0Y2_FrameStrobe_O),
    .FrameStrobe_O(Tile_X0Y1_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X1Y1_Emulate_Bitstream)
    )
`endif
    Tile_X1Y1_linear_LMDPL
    (
    .from_NA(Tile_X1Y2_to_NA),
    .from_NB(Tile_X1Y2_to_NB),
    .from_NC(Tile_X1Y2_to_NC),
    .from_ND(Tile_X1Y2_to_ND),
    .from_NF(Tile_X1Y2_to_NF),
    .from_NG(Tile_X1Y2_to_NG),
    .from_NH(Tile_X1Y2_to_NH),
    .from_NI(Tile_X1Y2_to_NI),
    .from_EA(Tile_X0Y1_to_EA),
    .from_EB(Tile_X0Y1_to_EB),
    .from_EC(Tile_X0Y1_to_EC),
    .from_ED(Tile_X0Y1_to_ED),
    .from_EF(Tile_X0Y1_to_EF),
    .from_EG(Tile_X0Y1_to_EG),
    .from_EH(Tile_X0Y1_to_EH),
    .from_EI(Tile_X0Y1_to_EI),
    .from_SA(Tile_X1Y0_to_SA),
    .from_SB(Tile_X1Y0_to_SB),
    .from_SC(Tile_X1Y0_to_SC),
    .from_SD(Tile_X1Y0_to_SD),
    .from_SF(Tile_X1Y0_to_SF),
    .from_SG(Tile_X1Y0_to_SG),
    .from_SH(Tile_X1Y0_to_SH),
    .from_SI(Tile_X1Y0_to_SI),
    .from_WA(Tile_X2Y1_to_WA),
    .from_WB(Tile_X2Y1_to_WB),
    .from_WC(Tile_X2Y1_to_WC),
    .from_WD(Tile_X2Y1_to_WD),
    .from_WF(Tile_X2Y1_to_WF),
    .from_WG(Tile_X2Y1_to_WG),
    .from_WH(Tile_X2Y1_to_WH),
    .from_WI(Tile_X2Y1_to_WI),
    .to_EA(Tile_X1Y1_to_EA),
    .to_EB(Tile_X1Y1_to_EB),
    .to_EC(Tile_X1Y1_to_EC),
    .to_ED(Tile_X1Y1_to_ED),
    .to_EF(Tile_X1Y1_to_EF),
    .to_EG(Tile_X1Y1_to_EG),
    .to_EH(Tile_X1Y1_to_EH),
    .to_EI(Tile_X1Y1_to_EI),
    .to_WA(Tile_X1Y1_to_WA),
    .to_WB(Tile_X1Y1_to_WB),
    .to_WC(Tile_X1Y1_to_WC),
    .to_WD(Tile_X1Y1_to_WD),
    .to_WF(Tile_X1Y1_to_WF),
    .to_WG(Tile_X1Y1_to_WG),
    .to_WH(Tile_X1Y1_to_WH),
    .to_WI(Tile_X1Y1_to_WI),
    .to_NA(Tile_X1Y1_to_NA),
    .to_NB(Tile_X1Y1_to_NB),
    .to_NC(Tile_X1Y1_to_NC),
    .to_ND(Tile_X1Y1_to_ND),
    .to_NF(Tile_X1Y1_to_NF),
    .to_NG(Tile_X1Y1_to_NG),
    .to_NH(Tile_X1Y1_to_NH),
    .to_NI(Tile_X1Y1_to_NI),
    .to_SA(Tile_X1Y1_to_SA),
    .to_SB(Tile_X1Y1_to_SB),
    .to_SC(Tile_X1Y1_to_SC),
    .to_SD(Tile_X1Y1_to_SD),
    .to_SF(Tile_X1Y1_to_SF),
    .to_SG(Tile_X1Y1_to_SG),
    .to_SH(Tile_X1Y1_to_SH),
    .to_SI(Tile_X1Y1_to_SI),
    .F_masked1(Tile_X1Y1_F_masked1),
    .F_masked2(Tile_X1Y1_F_masked2),
    .UserCLK(Tile_X1Y2_UserCLKo),
    .UserCLKo(Tile_X1Y1_UserCLKo),
    .rst(Tile_X1Y2_rsto),
    .rsto(Tile_X1Y1_rsto),
    .FrameData(Tile_X0Y1_FrameData_O),
    .FrameData_O(Tile_X1Y1_FrameData_O),
    .FrameStrobe(Tile_X1Y2_FrameStrobe_O),
    .FrameStrobe_O(Tile_X1Y1_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X2Y1_Emulate_Bitstream)
    )
`endif
    Tile_X2Y1_linear_LMDPL
    (
    .from_NA(Tile_X2Y2_to_NA),
    .from_NB(Tile_X2Y2_to_NB),
    .from_NC(Tile_X2Y2_to_NC),
    .from_ND(Tile_X2Y2_to_ND),
    .from_NF(Tile_X2Y2_to_NF),
    .from_NG(Tile_X2Y2_to_NG),
    .from_NH(Tile_X2Y2_to_NH),
    .from_NI(Tile_X2Y2_to_NI),
    .from_EA(Tile_X1Y1_to_EA),
    .from_EB(Tile_X1Y1_to_EB),
    .from_EC(Tile_X1Y1_to_EC),
    .from_ED(Tile_X1Y1_to_ED),
    .from_EF(Tile_X1Y1_to_EF),
    .from_EG(Tile_X1Y1_to_EG),
    .from_EH(Tile_X1Y1_to_EH),
    .from_EI(Tile_X1Y1_to_EI),
    .from_SA(Tile_X2Y0_to_SA),
    .from_SB(Tile_X2Y0_to_SB),
    .from_SC(Tile_X2Y0_to_SC),
    .from_SD(Tile_X2Y0_to_SD),
    .from_SF(Tile_X2Y0_to_SF),
    .from_SG(Tile_X2Y0_to_SG),
    .from_SH(Tile_X2Y0_to_SH),
    .from_SI(Tile_X2Y0_to_SI),
    .from_WA(Tile_X3Y1_to_WA),
    .from_WB(Tile_X3Y1_to_WB),
    .from_WC(Tile_X3Y1_to_WC),
    .from_WD(Tile_X3Y1_to_WD),
    .from_WF(Tile_X3Y1_to_WF),
    .from_WG(Tile_X3Y1_to_WG),
    .from_WH(Tile_X3Y1_to_WH),
    .from_WI(Tile_X3Y1_to_WI),
    .to_EA(Tile_X2Y1_to_EA),
    .to_EB(Tile_X2Y1_to_EB),
    .to_EC(Tile_X2Y1_to_EC),
    .to_ED(Tile_X2Y1_to_ED),
    .to_EF(Tile_X2Y1_to_EF),
    .to_EG(Tile_X2Y1_to_EG),
    .to_EH(Tile_X2Y1_to_EH),
    .to_EI(Tile_X2Y1_to_EI),
    .to_WA(Tile_X2Y1_to_WA),
    .to_WB(Tile_X2Y1_to_WB),
    .to_WC(Tile_X2Y1_to_WC),
    .to_WD(Tile_X2Y1_to_WD),
    .to_WF(Tile_X2Y1_to_WF),
    .to_WG(Tile_X2Y1_to_WG),
    .to_WH(Tile_X2Y1_to_WH),
    .to_WI(Tile_X2Y1_to_WI),
    .to_NA(Tile_X2Y1_to_NA),
    .to_NB(Tile_X2Y1_to_NB),
    .to_NC(Tile_X2Y1_to_NC),
    .to_ND(Tile_X2Y1_to_ND),
    .to_NF(Tile_X2Y1_to_NF),
    .to_NG(Tile_X2Y1_to_NG),
    .to_NH(Tile_X2Y1_to_NH),
    .to_NI(Tile_X2Y1_to_NI),
    .to_SA(Tile_X2Y1_to_SA),
    .to_SB(Tile_X2Y1_to_SB),
    .to_SC(Tile_X2Y1_to_SC),
    .to_SD(Tile_X2Y1_to_SD),
    .to_SF(Tile_X2Y1_to_SF),
    .to_SG(Tile_X2Y1_to_SG),
    .to_SH(Tile_X2Y1_to_SH),
    .to_SI(Tile_X2Y1_to_SI),
    .F_masked1(Tile_X2Y1_F_masked1),
    .F_masked2(Tile_X2Y1_F_masked2),
    .UserCLK(Tile_X2Y2_UserCLKo),
    .UserCLKo(Tile_X2Y1_UserCLKo),
    .rst(Tile_X2Y2_rsto),
    .rsto(Tile_X2Y1_rsto),
    .FrameData(Tile_X1Y1_FrameData_O),
    .FrameData_O(Tile_X2Y1_FrameData_O),
    .FrameStrobe(Tile_X2Y2_FrameStrobe_O),
    .FrameStrobe_O(Tile_X2Y1_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
nonlinear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X3Y1_Emulate_Bitstream)
    )
`endif
    Tile_X3Y1_nonlinear_LMDPL
    (
    .from_NA(Tile_X3Y2_to_NA),
    .from_NB(Tile_X3Y2_to_NB),
    .from_NC(Tile_X3Y2_to_NC),
    .from_ND(Tile_X3Y2_to_ND),
    .from_NF(Tile_X3Y2_to_NF),
    .from_NG(Tile_X3Y2_to_NG),
    .from_NH(Tile_X3Y2_to_NH),
    .from_NI(Tile_X3Y2_to_NI),
    .from_EA(Tile_X2Y1_to_EA),
    .from_EB(Tile_X2Y1_to_EB),
    .from_EC(Tile_X2Y1_to_EC),
    .from_ED(Tile_X2Y1_to_ED),
    .from_EF(Tile_X2Y1_to_EF),
    .from_EG(Tile_X2Y1_to_EG),
    .from_EH(Tile_X2Y1_to_EH),
    .from_EI(Tile_X2Y1_to_EI),
    .from_SA(Tile_X3Y0_to_SA),
    .from_SB(Tile_X3Y0_to_SB),
    .from_SC(Tile_X3Y0_to_SC),
    .from_SD(Tile_X3Y0_to_SD),
    .from_SF(Tile_X3Y0_to_SF),
    .from_SG(Tile_X3Y0_to_SG),
    .from_SH(Tile_X3Y0_to_SH),
    .from_SI(Tile_X3Y0_to_SI),
    .from_WA(Tile_X4Y1_to_WA),
    .from_WB(Tile_X4Y1_to_WB),
    .from_WC(Tile_X4Y1_to_WC),
    .from_WD(Tile_X4Y1_to_WD),
    .from_WF(Tile_X4Y1_to_WF),
    .from_WG(Tile_X4Y1_to_WG),
    .from_WH(Tile_X4Y1_to_WH),
    .from_WI(Tile_X4Y1_to_WI),
    .to_EA(Tile_X3Y1_to_EA),
    .to_EB(Tile_X3Y1_to_EB),
    .to_EC(Tile_X3Y1_to_EC),
    .to_ED(Tile_X3Y1_to_ED),
    .to_EF(Tile_X3Y1_to_EF),
    .to_EG(Tile_X3Y1_to_EG),
    .to_EH(Tile_X3Y1_to_EH),
    .to_EI(Tile_X3Y1_to_EI),
    .to_WA(Tile_X3Y1_to_WA),
    .to_WB(Tile_X3Y1_to_WB),
    .to_WC(Tile_X3Y1_to_WC),
    .to_WD(Tile_X3Y1_to_WD),
    .to_WF(Tile_X3Y1_to_WF),
    .to_WG(Tile_X3Y1_to_WG),
    .to_WH(Tile_X3Y1_to_WH),
    .to_WI(Tile_X3Y1_to_WI),
    .to_NA(Tile_X3Y1_to_NA),
    .to_NB(Tile_X3Y1_to_NB),
    .to_NC(Tile_X3Y1_to_NC),
    .to_ND(Tile_X3Y1_to_ND),
    .to_NF(Tile_X3Y1_to_NF),
    .to_NG(Tile_X3Y1_to_NG),
    .to_NH(Tile_X3Y1_to_NH),
    .to_NI(Tile_X3Y1_to_NI),
    .to_SA(Tile_X3Y1_to_SA),
    .to_SB(Tile_X3Y1_to_SB),
    .to_SC(Tile_X3Y1_to_SC),
    .to_SD(Tile_X3Y1_to_SD),
    .to_SF(Tile_X3Y1_to_SF),
    .to_SG(Tile_X3Y1_to_SG),
    .to_SH(Tile_X3Y1_to_SH),
    .to_SI(Tile_X3Y1_to_SI),
    .R_t(Tile_X3Y1_R_t),
    .R_f(Tile_X3Y1_R_f),
    .F_masked1(Tile_X3Y1_F_masked1),
    .F_masked2(Tile_X3Y1_F_masked2),
    .UserCLK(Tile_X3Y2_UserCLKo),
    .UserCLKo(Tile_X3Y1_UserCLKo),
    .rst(Tile_X3Y2_rsto),
    .rsto(Tile_X3Y1_rsto),
    .FrameData(Tile_X2Y1_FrameData_O),
    .FrameData_O(Tile_X3Y1_FrameData_O),
    .FrameStrobe(Tile_X3Y2_FrameStrobe_O),
    .FrameStrobe_O(Tile_X3Y1_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X4Y1_Emulate_Bitstream)
    )
`endif
    Tile_X4Y1_linear_LMDPL
    (
    .from_NA(Tile_X4Y2_to_NA),
    .from_NB(Tile_X4Y2_to_NB),
    .from_NC(Tile_X4Y2_to_NC),
    .from_ND(Tile_X4Y2_to_ND),
    .from_NF(Tile_X4Y2_to_NF),
    .from_NG(Tile_X4Y2_to_NG),
    .from_NH(Tile_X4Y2_to_NH),
    .from_NI(Tile_X4Y2_to_NI),
    .from_EA(Tile_X3Y1_to_EA),
    .from_EB(Tile_X3Y1_to_EB),
    .from_EC(Tile_X3Y1_to_EC),
    .from_ED(Tile_X3Y1_to_ED),
    .from_EF(Tile_X3Y1_to_EF),
    .from_EG(Tile_X3Y1_to_EG),
    .from_EH(Tile_X3Y1_to_EH),
    .from_EI(Tile_X3Y1_to_EI),
    .from_SA(Tile_X4Y0_to_SA),
    .from_SB(Tile_X4Y0_to_SB),
    .from_SC(Tile_X4Y0_to_SC),
    .from_SD(Tile_X4Y0_to_SD),
    .from_SF(Tile_X4Y0_to_SF),
    .from_SG(Tile_X4Y0_to_SG),
    .from_SH(Tile_X4Y0_to_SH),
    .from_SI(Tile_X4Y0_to_SI),
    .from_WA(Tile_X5Y1_to_WA),
    .from_WB(Tile_X5Y1_to_WB),
    .from_WC(Tile_X5Y1_to_WC),
    .from_WD(Tile_X5Y1_to_WD),
    .from_WF(Tile_X5Y1_to_WF),
    .from_WG(Tile_X5Y1_to_WG),
    .from_WH(Tile_X5Y1_to_WH),
    .from_WI(Tile_X5Y1_to_WI),
    .to_EA(Tile_X4Y1_to_EA),
    .to_EB(Tile_X4Y1_to_EB),
    .to_EC(Tile_X4Y1_to_EC),
    .to_ED(Tile_X4Y1_to_ED),
    .to_EF(Tile_X4Y1_to_EF),
    .to_EG(Tile_X4Y1_to_EG),
    .to_EH(Tile_X4Y1_to_EH),
    .to_EI(Tile_X4Y1_to_EI),
    .to_WA(Tile_X4Y1_to_WA),
    .to_WB(Tile_X4Y1_to_WB),
    .to_WC(Tile_X4Y1_to_WC),
    .to_WD(Tile_X4Y1_to_WD),
    .to_WF(Tile_X4Y1_to_WF),
    .to_WG(Tile_X4Y1_to_WG),
    .to_WH(Tile_X4Y1_to_WH),
    .to_WI(Tile_X4Y1_to_WI),
    .to_NA(Tile_X4Y1_to_NA),
    .to_NB(Tile_X4Y1_to_NB),
    .to_NC(Tile_X4Y1_to_NC),
    .to_ND(Tile_X4Y1_to_ND),
    .to_NF(Tile_X4Y1_to_NF),
    .to_NG(Tile_X4Y1_to_NG),
    .to_NH(Tile_X4Y1_to_NH),
    .to_NI(Tile_X4Y1_to_NI),
    .to_SA(Tile_X4Y1_to_SA),
    .to_SB(Tile_X4Y1_to_SB),
    .to_SC(Tile_X4Y1_to_SC),
    .to_SD(Tile_X4Y1_to_SD),
    .to_SF(Tile_X4Y1_to_SF),
    .to_SG(Tile_X4Y1_to_SG),
    .to_SH(Tile_X4Y1_to_SH),
    .to_SI(Tile_X4Y1_to_SI),
    .F_masked1(Tile_X4Y1_F_masked1),
    .F_masked2(Tile_X4Y1_F_masked2),
    .UserCLK(Tile_X4Y2_UserCLKo),
    .UserCLKo(Tile_X4Y1_UserCLKo),
    .rst(Tile_X4Y2_rsto),
    .rsto(Tile_X4Y1_rsto),
    .FrameData(Tile_X3Y1_FrameData_O),
    .FrameData_O(Tile_X4Y1_FrameData_O),
    .FrameStrobe(Tile_X4Y2_FrameStrobe_O),
    .FrameStrobe_O(Tile_X4Y1_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X5Y1_Emulate_Bitstream)
    )
`endif
    Tile_X5Y1_linear_LMDPL
    (
    .from_NA(Tile_X5Y2_to_NA),
    .from_NB(Tile_X5Y2_to_NB),
    .from_NC(Tile_X5Y2_to_NC),
    .from_ND(Tile_X5Y2_to_ND),
    .from_NF(Tile_X5Y2_to_NF),
    .from_NG(Tile_X5Y2_to_NG),
    .from_NH(Tile_X5Y2_to_NH),
    .from_NI(Tile_X5Y2_to_NI),
    .from_EA(Tile_X4Y1_to_EA),
    .from_EB(Tile_X4Y1_to_EB),
    .from_EC(Tile_X4Y1_to_EC),
    .from_ED(Tile_X4Y1_to_ED),
    .from_EF(Tile_X4Y1_to_EF),
    .from_EG(Tile_X4Y1_to_EG),
    .from_EH(Tile_X4Y1_to_EH),
    .from_EI(Tile_X4Y1_to_EI),
    .from_SA(Tile_X5Y0_to_SA),
    .from_SB(Tile_X5Y0_to_SB),
    .from_SC(Tile_X5Y0_to_SC),
    .from_SD(Tile_X5Y0_to_SD),
    .from_SF(Tile_X5Y0_to_SF),
    .from_SG(Tile_X5Y0_to_SG),
    .from_SH(Tile_X5Y0_to_SH),
    .from_SI(Tile_X5Y0_to_SI),
    .from_WA(Tile_X6Y1_to_WA),
    .from_WB(Tile_X6Y1_to_WB),
    .from_WC(Tile_X6Y1_to_WC),
    .from_WD(Tile_X6Y1_to_WD),
    .from_WF(Tile_X6Y1_to_WF),
    .from_WG(Tile_X6Y1_to_WG),
    .from_WH(Tile_X6Y1_to_WH),
    .from_WI(Tile_X6Y1_to_WI),
    .to_EA(Tile_X5Y1_to_EA),
    .to_EB(Tile_X5Y1_to_EB),
    .to_EC(Tile_X5Y1_to_EC),
    .to_ED(Tile_X5Y1_to_ED),
    .to_EF(Tile_X5Y1_to_EF),
    .to_EG(Tile_X5Y1_to_EG),
    .to_EH(Tile_X5Y1_to_EH),
    .to_EI(Tile_X5Y1_to_EI),
    .to_WA(Tile_X5Y1_to_WA),
    .to_WB(Tile_X5Y1_to_WB),
    .to_WC(Tile_X5Y1_to_WC),
    .to_WD(Tile_X5Y1_to_WD),
    .to_WF(Tile_X5Y1_to_WF),
    .to_WG(Tile_X5Y1_to_WG),
    .to_WH(Tile_X5Y1_to_WH),
    .to_WI(Tile_X5Y1_to_WI),
    .to_NA(Tile_X5Y1_to_NA),
    .to_NB(Tile_X5Y1_to_NB),
    .to_NC(Tile_X5Y1_to_NC),
    .to_ND(Tile_X5Y1_to_ND),
    .to_NF(Tile_X5Y1_to_NF),
    .to_NG(Tile_X5Y1_to_NG),
    .to_NH(Tile_X5Y1_to_NH),
    .to_NI(Tile_X5Y1_to_NI),
    .to_SA(Tile_X5Y1_to_SA),
    .to_SB(Tile_X5Y1_to_SB),
    .to_SC(Tile_X5Y1_to_SC),
    .to_SD(Tile_X5Y1_to_SD),
    .to_SF(Tile_X5Y1_to_SF),
    .to_SG(Tile_X5Y1_to_SG),
    .to_SH(Tile_X5Y1_to_SH),
    .to_SI(Tile_X5Y1_to_SI),
    .F_masked1(Tile_X5Y1_F_masked1),
    .F_masked2(Tile_X5Y1_F_masked2),
    .UserCLK(Tile_X5Y2_UserCLKo),
    .UserCLKo(Tile_X5Y1_UserCLKo),
    .rst(Tile_X5Y2_rsto),
    .rsto(Tile_X5Y1_rsto),
    .FrameData(Tile_X4Y1_FrameData_O),
    .FrameData_O(Tile_X5Y1_FrameData_O),
    .FrameStrobe(Tile_X5Y2_FrameStrobe_O),
    .FrameStrobe_O(Tile_X5Y1_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
nonlinear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X6Y1_Emulate_Bitstream)
    )
`endif
    Tile_X6Y1_nonlinear_LMDPL
    (
    .from_NA(Tile_X6Y2_to_NA),
    .from_NB(Tile_X6Y2_to_NB),
    .from_NC(Tile_X6Y2_to_NC),
    .from_ND(Tile_X6Y2_to_ND),
    .from_NF(Tile_X6Y2_to_NF),
    .from_NG(Tile_X6Y2_to_NG),
    .from_NH(Tile_X6Y2_to_NH),
    .from_NI(Tile_X6Y2_to_NI),
    .from_EA(Tile_X5Y1_to_EA),
    .from_EB(Tile_X5Y1_to_EB),
    .from_EC(Tile_X5Y1_to_EC),
    .from_ED(Tile_X5Y1_to_ED),
    .from_EF(Tile_X5Y1_to_EF),
    .from_EG(Tile_X5Y1_to_EG),
    .from_EH(Tile_X5Y1_to_EH),
    .from_EI(Tile_X5Y1_to_EI),
    .from_SA(Tile_X6Y0_to_SA),
    .from_SB(Tile_X6Y0_to_SB),
    .from_SC(Tile_X6Y0_to_SC),
    .from_SD(Tile_X6Y0_to_SD),
    .from_SF(Tile_X6Y0_to_SF),
    .from_SG(Tile_X6Y0_to_SG),
    .from_SH(Tile_X6Y0_to_SH),
    .from_SI(Tile_X6Y0_to_SI),
    .from_WA(Tile_X7Y1_to_WA),
    .from_WB(Tile_X7Y1_to_WB),
    .from_WC(Tile_X7Y1_to_WC),
    .from_WD(Tile_X7Y1_to_WD),
    .from_WF(Tile_X7Y1_to_WF),
    .from_WG(Tile_X7Y1_to_WG),
    .from_WH(Tile_X7Y1_to_WH),
    .from_WI(Tile_X7Y1_to_WI),
    .to_EA(Tile_X6Y1_to_EA),
    .to_EB(Tile_X6Y1_to_EB),
    .to_EC(Tile_X6Y1_to_EC),
    .to_ED(Tile_X6Y1_to_ED),
    .to_EF(Tile_X6Y1_to_EF),
    .to_EG(Tile_X6Y1_to_EG),
    .to_EH(Tile_X6Y1_to_EH),
    .to_EI(Tile_X6Y1_to_EI),
    .to_WA(Tile_X6Y1_to_WA),
    .to_WB(Tile_X6Y1_to_WB),
    .to_WC(Tile_X6Y1_to_WC),
    .to_WD(Tile_X6Y1_to_WD),
    .to_WF(Tile_X6Y1_to_WF),
    .to_WG(Tile_X6Y1_to_WG),
    .to_WH(Tile_X6Y1_to_WH),
    .to_WI(Tile_X6Y1_to_WI),
    .to_NA(Tile_X6Y1_to_NA),
    .to_NB(Tile_X6Y1_to_NB),
    .to_NC(Tile_X6Y1_to_NC),
    .to_ND(Tile_X6Y1_to_ND),
    .to_NF(Tile_X6Y1_to_NF),
    .to_NG(Tile_X6Y1_to_NG),
    .to_NH(Tile_X6Y1_to_NH),
    .to_NI(Tile_X6Y1_to_NI),
    .to_SA(Tile_X6Y1_to_SA),
    .to_SB(Tile_X6Y1_to_SB),
    .to_SC(Tile_X6Y1_to_SC),
    .to_SD(Tile_X6Y1_to_SD),
    .to_SF(Tile_X6Y1_to_SF),
    .to_SG(Tile_X6Y1_to_SG),
    .to_SH(Tile_X6Y1_to_SH),
    .to_SI(Tile_X6Y1_to_SI),
    .R_t(Tile_X6Y1_R_t),
    .R_f(Tile_X6Y1_R_f),
    .F_masked1(Tile_X6Y1_F_masked1),
    .F_masked2(Tile_X6Y1_F_masked2),
    .UserCLK(Tile_X6Y2_UserCLKo),
    .UserCLKo(Tile_X6Y1_UserCLKo),
    .rst(Tile_X6Y2_rsto),
    .rsto(Tile_X6Y1_rsto),
    .FrameData(Tile_X5Y1_FrameData_O),
    .FrameData_O(Tile_X6Y1_FrameData_O),
    .FrameStrobe(Tile_X6Y2_FrameStrobe_O),
    .FrameStrobe_O(Tile_X6Y1_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X7Y1_Emulate_Bitstream)
    )
`endif
    Tile_X7Y1_linear_LMDPL
    (
    .from_NA(Tile_X7Y2_to_NA),
    .from_NB(Tile_X7Y2_to_NB),
    .from_NC(Tile_X7Y2_to_NC),
    .from_ND(Tile_X7Y2_to_ND),
    .from_NF(Tile_X7Y2_to_NF),
    .from_NG(Tile_X7Y2_to_NG),
    .from_NH(Tile_X7Y2_to_NH),
    .from_NI(Tile_X7Y2_to_NI),
    .from_EA(Tile_X6Y1_to_EA),
    .from_EB(Tile_X6Y1_to_EB),
    .from_EC(Tile_X6Y1_to_EC),
    .from_ED(Tile_X6Y1_to_ED),
    .from_EF(Tile_X6Y1_to_EF),
    .from_EG(Tile_X6Y1_to_EG),
    .from_EH(Tile_X6Y1_to_EH),
    .from_EI(Tile_X6Y1_to_EI),
    .from_SA(Tile_X7Y0_to_SA),
    .from_SB(Tile_X7Y0_to_SB),
    .from_SC(Tile_X7Y0_to_SC),
    .from_SD(Tile_X7Y0_to_SD),
    .from_SF(Tile_X7Y0_to_SF),
    .from_SG(Tile_X7Y0_to_SG),
    .from_SH(Tile_X7Y0_to_SH),
    .from_SI(Tile_X7Y0_to_SI),
    .from_WA(Tile_X8Y1_to_WA),
    .from_WB(Tile_X8Y1_to_WB),
    .from_WC(Tile_X8Y1_to_WC),
    .from_WD(Tile_X8Y1_to_WD),
    .from_WF(Tile_X8Y1_to_WF),
    .from_WG(Tile_X8Y1_to_WG),
    .from_WH(Tile_X8Y1_to_WH),
    .from_WI(Tile_X8Y1_to_WI),
    .to_EA(Tile_X7Y1_to_EA),
    .to_EB(Tile_X7Y1_to_EB),
    .to_EC(Tile_X7Y1_to_EC),
    .to_ED(Tile_X7Y1_to_ED),
    .to_EF(Tile_X7Y1_to_EF),
    .to_EG(Tile_X7Y1_to_EG),
    .to_EH(Tile_X7Y1_to_EH),
    .to_EI(Tile_X7Y1_to_EI),
    .to_WA(Tile_X7Y1_to_WA),
    .to_WB(Tile_X7Y1_to_WB),
    .to_WC(Tile_X7Y1_to_WC),
    .to_WD(Tile_X7Y1_to_WD),
    .to_WF(Tile_X7Y1_to_WF),
    .to_WG(Tile_X7Y1_to_WG),
    .to_WH(Tile_X7Y1_to_WH),
    .to_WI(Tile_X7Y1_to_WI),
    .to_NA(Tile_X7Y1_to_NA),
    .to_NB(Tile_X7Y1_to_NB),
    .to_NC(Tile_X7Y1_to_NC),
    .to_ND(Tile_X7Y1_to_ND),
    .to_NF(Tile_X7Y1_to_NF),
    .to_NG(Tile_X7Y1_to_NG),
    .to_NH(Tile_X7Y1_to_NH),
    .to_NI(Tile_X7Y1_to_NI),
    .to_SA(Tile_X7Y1_to_SA),
    .to_SB(Tile_X7Y1_to_SB),
    .to_SC(Tile_X7Y1_to_SC),
    .to_SD(Tile_X7Y1_to_SD),
    .to_SF(Tile_X7Y1_to_SF),
    .to_SG(Tile_X7Y1_to_SG),
    .to_SH(Tile_X7Y1_to_SH),
    .to_SI(Tile_X7Y1_to_SI),
    .F_masked1(Tile_X7Y1_F_masked1),
    .F_masked2(Tile_X7Y1_F_masked2),
    .UserCLK(Tile_X7Y2_UserCLKo),
    .UserCLKo(Tile_X7Y1_UserCLKo),
    .rst(Tile_X7Y2_rsto),
    .rsto(Tile_X7Y1_rsto),
    .FrameData(Tile_X6Y1_FrameData_O),
    .FrameData_O(Tile_X7Y1_FrameData_O),
    .FrameStrobe(Tile_X7Y2_FrameStrobe_O),
    .FrameStrobe_O(Tile_X7Y1_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
ctrl_to_sec
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X8Y1_Emulate_Bitstream)
    )
`endif
    Tile_X8Y1_ctrl_to_sec
    (
    .from_NA(Tile_X8Y2_to_NA),
    .from_NB(Tile_X8Y2_to_NB),
    .from_NC(Tile_X8Y2_to_NC),
    .from_ND(Tile_X8Y2_to_ND),
    .from_NF(Tile_X8Y2_to_NF),
    .from_NG(Tile_X8Y2_to_NG),
    .from_NH(Tile_X8Y2_to_NH),
    .from_NI(Tile_X8Y2_to_NI),
    .from_EA(Tile_X7Y1_to_EA),
    .from_EB(Tile_X7Y1_to_EB),
    .from_EC(Tile_X7Y1_to_EC),
    .from_ED(Tile_X7Y1_to_ED),
    .from_EF(Tile_X7Y1_to_EF),
    .from_EG(Tile_X7Y1_to_EG),
    .from_EH(Tile_X7Y1_to_EH),
    .from_EI(Tile_X7Y1_to_EI),
    .from_SA(Tile_X8Y0_to_SA),
    .from_SB(Tile_X8Y0_to_SB),
    .from_SC(Tile_X8Y0_to_SC),
    .from_SD(Tile_X8Y0_to_SD),
    .from_SF(Tile_X8Y0_to_SF),
    .from_SG(Tile_X8Y0_to_SG),
    .from_SH(Tile_X8Y0_to_SH),
    .from_SI(Tile_X8Y0_to_SI),
    .from_WA_1s(Tile_X9Y1_to_WA_1s),
    .from_WB_1s(Tile_X9Y1_to_WB_1s),
    .from_WC_1s(Tile_X9Y1_to_WC_1s),
    .from_WD_1s(Tile_X9Y1_to_WD_1s),
    .from_WF_1s(Tile_X9Y1_to_WF_1s),
    .from_WG_1s(Tile_X9Y1_to_WG_1s),
    .from_WH_1s(Tile_X9Y1_to_WH_1s),
    .from_WI_1s(Tile_X9Y1_to_WI_1s),
    .to_WA(Tile_X8Y1_to_WA),
    .to_WB(Tile_X8Y1_to_WB),
    .to_WC(Tile_X8Y1_to_WC),
    .to_WD(Tile_X8Y1_to_WD),
    .to_WF(Tile_X8Y1_to_WF),
    .to_WG(Tile_X8Y1_to_WG),
    .to_WH(Tile_X8Y1_to_WH),
    .to_WI(Tile_X8Y1_to_WI),
    .to_NA(Tile_X8Y1_to_NA),
    .to_NB(Tile_X8Y1_to_NB),
    .to_NC(Tile_X8Y1_to_NC),
    .to_ND(Tile_X8Y1_to_ND),
    .to_NF(Tile_X8Y1_to_NF),
    .to_NG(Tile_X8Y1_to_NG),
    .to_NH(Tile_X8Y1_to_NH),
    .to_NI(Tile_X8Y1_to_NI),
    .to_SA(Tile_X8Y1_to_SA),
    .to_SB(Tile_X8Y1_to_SB),
    .to_SC(Tile_X8Y1_to_SC),
    .to_SD(Tile_X8Y1_to_SD),
    .to_SF(Tile_X8Y1_to_SF),
    .to_SG(Tile_X8Y1_to_SG),
    .to_SH(Tile_X8Y1_to_SH),
    .to_SI(Tile_X8Y1_to_SI),
    .UserCLK(Tile_X8Y2_UserCLKo),
    .UserCLKo(Tile_X8Y1_UserCLKo),
    .rst(Tile_X8Y2_rsto),
    .rsto(Tile_X8Y1_rsto),
    .FrameData(Tile_X7Y1_FrameData_O),
    .FrameData_O(Tile_X8Y1_FrameData_O),
    .FrameStrobe(Tile_X8Y2_FrameStrobe_O),
    .FrameStrobe_O(Tile_X8Y1_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
combined_WDDL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X9Y1_Emulate_Bitstream)
    )
`endif
    Tile_X9Y1_combined_WDDL
    (
    .from_NA_1s(Tile_X9Y2_to_NA_1s),
    .from_NB_1s(Tile_X9Y2_to_NB_1s),
    .from_NC_1s(Tile_X9Y2_to_NC_1s),
    .from_ND_1s(Tile_X9Y2_to_ND_1s),
    .from_NF_1s(Tile_X9Y2_to_NF_1s),
    .from_NG_1s(Tile_X9Y2_to_NG_1s),
    .from_NH_1s(Tile_X9Y2_to_NH_1s),
    .from_NI_1s(Tile_X9Y2_to_NI_1s),
    .from_SA_1s(Tile_X9Y0_to_SA_1s),
    .from_SB_1s(Tile_X9Y0_to_SB_1s),
    .from_SC_1s(Tile_X9Y0_to_SC_1s),
    .from_SD_1s(Tile_X9Y0_to_SD_1s),
    .from_SF_1s(Tile_X9Y0_to_SF_1s),
    .from_SG_1s(Tile_X9Y0_to_SG_1s),
    .from_SH_1s(Tile_X9Y0_to_SH_1s),
    .from_SI_1s(Tile_X9Y0_to_SI_1s),
    .from_WA_1s(Tile_X10Y1_to_WA_1s),
    .from_WB_1s(Tile_X10Y1_to_WB_1s),
    .from_WC_1s(Tile_X10Y1_to_WC_1s),
    .from_WD_1s(Tile_X10Y1_to_WD_1s),
    .from_WF_1s(Tile_X10Y1_to_WF_1s),
    .from_WG_1s(Tile_X10Y1_to_WG_1s),
    .from_WH_1s(Tile_X10Y1_to_WH_1s),
    .from_WI_1s(Tile_X10Y1_to_WI_1s),
    .to_EA_1s(Tile_X9Y1_to_EA_1s),
    .to_EB_1s(Tile_X9Y1_to_EB_1s),
    .to_EC_1s(Tile_X9Y1_to_EC_1s),
    .to_ED_1s(Tile_X9Y1_to_ED_1s),
    .to_EF_1s(Tile_X9Y1_to_EF_1s),
    .to_EG_1s(Tile_X9Y1_to_EG_1s),
    .to_EH_1s(Tile_X9Y1_to_EH_1s),
    .to_EI_1s(Tile_X9Y1_to_EI_1s),
    .to_WA_1s(Tile_X9Y1_to_WA_1s),
    .to_WB_1s(Tile_X9Y1_to_WB_1s),
    .to_WC_1s(Tile_X9Y1_to_WC_1s),
    .to_WD_1s(Tile_X9Y1_to_WD_1s),
    .to_WF_1s(Tile_X9Y1_to_WF_1s),
    .to_WG_1s(Tile_X9Y1_to_WG_1s),
    .to_WH_1s(Tile_X9Y1_to_WH_1s),
    .to_WI_1s(Tile_X9Y1_to_WI_1s),
    .to_NA_1s(Tile_X9Y1_to_NA_1s),
    .to_NB_1s(Tile_X9Y1_to_NB_1s),
    .to_NC_1s(Tile_X9Y1_to_NC_1s),
    .to_ND_1s(Tile_X9Y1_to_ND_1s),
    .to_NF_1s(Tile_X9Y1_to_NF_1s),
    .to_NG_1s(Tile_X9Y1_to_NG_1s),
    .to_NH_1s(Tile_X9Y1_to_NH_1s),
    .to_NI_1s(Tile_X9Y1_to_NI_1s),
    .to_SA_1s(Tile_X9Y1_to_SA_1s),
    .to_SB_1s(Tile_X9Y1_to_SB_1s),
    .to_SC_1s(Tile_X9Y1_to_SC_1s),
    .to_SD_1s(Tile_X9Y1_to_SD_1s),
    .to_SF_1s(Tile_X9Y1_to_SF_1s),
    .to_SG_1s(Tile_X9Y1_to_SG_1s),
    .to_SH_1s(Tile_X9Y1_to_SH_1s),
    .to_SI_1s(Tile_X9Y1_to_SI_1s),
    .F_ctrl(Tile_X9Y1_F_ctrl),
    .UserCLK(Tile_X9Y2_UserCLKo),
    .UserCLKo(Tile_X9Y1_UserCLKo),
    .rst(Tile_X9Y2_rsto),
    .rsto(Tile_X9Y1_rsto),
    .FrameData(Tile_X8Y1_FrameData_O),
    .FrameData_O(Tile_X9Y1_FrameData_O),
    .FrameStrobe(Tile_X9Y2_FrameStrobe_O),
    .FrameStrobe_O(Tile_X9Y1_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
ctrl_IO
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X10Y1_Emulate_Bitstream)
    )
`endif
    Tile_X10Y1_ctrl_IO
    (
    .from_EA_1s(Tile_X9Y1_to_EA_1s),
    .from_EB_1s(Tile_X9Y1_to_EB_1s),
    .from_EC_1s(Tile_X9Y1_to_EC_1s),
    .from_ED_1s(Tile_X9Y1_to_ED_1s),
    .from_EF_1s(Tile_X9Y1_to_EF_1s),
    .from_EG_1s(Tile_X9Y1_to_EG_1s),
    .from_EH_1s(Tile_X9Y1_to_EH_1s),
    .from_EI_1s(Tile_X9Y1_to_EI_1s),
    .to_WA_1s(Tile_X10Y1_to_WA_1s),
    .to_WB_1s(Tile_X10Y1_to_WB_1s),
    .to_WC_1s(Tile_X10Y1_to_WC_1s),
    .to_WD_1s(Tile_X10Y1_to_WD_1s),
    .to_WF_1s(Tile_X10Y1_to_WF_1s),
    .to_WG_1s(Tile_X10Y1_to_WG_1s),
    .to_WH_1s(Tile_X10Y1_to_WH_1s),
    .to_WI_1s(Tile_X10Y1_to_WI_1s),
    .A_O_top_0_t(Tile_X10Y1_A_O_top_0_t),
    .A_O_top_0_f(Tile_X10Y1_A_O_top_0_f),
    .A_prech2(Tile_X10Y1_A_prech2),
    .A_DR_fault(Tile_X10Y1_A_DR_fault),
    .A_I_top_0_t(Tile_X10Y1_A_I_top_0_t),
    .A_I_top_0_f(Tile_X10Y1_A_I_top_0_f),
    .A_T_top(Tile_X10Y1_A_T_top),
    .A_F_ctrl(Tile_X10Y1_A_F_ctrl),
    .UserCLK(Tile_X10Y2_UserCLKo),
    .UserCLKo(Tile_X10Y1_UserCLKo),
    .rst(Tile_X10Y2_rsto),
    .rsto(Tile_X10Y1_rsto),
    .FrameData(Tile_X9Y1_FrameData_O),
    .FrameData_O(Tile_X10Y1_FrameData_O),
    .FrameStrobe(Tile_X10Y2_FrameStrobe_O),
    .FrameStrobe_O(Tile_X10Y1_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
W_IO_custom
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X0Y2_Emulate_Bitstream)
    )
`endif
    Tile_X0Y2_W_IO_custom
    (
    .from_NA(Tile_X0Y3_to_NA),
    .from_NB(Tile_X0Y3_to_NB),
    .from_NC(Tile_X0Y3_to_NC),
    .from_ND(Tile_X0Y3_to_ND),
    .from_NF(Tile_X0Y3_to_NF),
    .from_NG(Tile_X0Y3_to_NG),
    .from_NH(Tile_X0Y3_to_NH),
    .from_NI(Tile_X0Y3_to_NI),
    .from_SA(Tile_X0Y1_to_SA),
    .from_SB(Tile_X0Y1_to_SB),
    .from_SC(Tile_X0Y1_to_SC),
    .from_SD(Tile_X0Y1_to_SD),
    .from_SF(Tile_X0Y1_to_SF),
    .from_SG(Tile_X0Y1_to_SG),
    .from_SH(Tile_X0Y1_to_SH),
    .from_SI(Tile_X0Y1_to_SI),
    .from_WA(Tile_X1Y2_to_WA),
    .from_WB(Tile_X1Y2_to_WB),
    .from_WC(Tile_X1Y2_to_WC),
    .from_WD(Tile_X1Y2_to_WD),
    .from_WF(Tile_X1Y2_to_WF),
    .from_WG(Tile_X1Y2_to_WG),
    .from_WH(Tile_X1Y2_to_WH),
    .from_WI(Tile_X1Y2_to_WI),
    .to_EA(Tile_X0Y2_to_EA),
    .to_EB(Tile_X0Y2_to_EB),
    .to_EC(Tile_X0Y2_to_EC),
    .to_ED(Tile_X0Y2_to_ED),
    .to_EF(Tile_X0Y2_to_EF),
    .to_EG(Tile_X0Y2_to_EG),
    .to_EH(Tile_X0Y2_to_EH),
    .to_EI(Tile_X0Y2_to_EI),
    .to_NA(Tile_X0Y2_to_NA),
    .to_NB(Tile_X0Y2_to_NB),
    .to_NC(Tile_X0Y2_to_NC),
    .to_ND(Tile_X0Y2_to_ND),
    .to_NF(Tile_X0Y2_to_NF),
    .to_NG(Tile_X0Y2_to_NG),
    .to_NH(Tile_X0Y2_to_NH),
    .to_NI(Tile_X0Y2_to_NI),
    .to_SA(Tile_X0Y2_to_SA),
    .to_SB(Tile_X0Y2_to_SB),
    .to_SC(Tile_X0Y2_to_SC),
    .to_SD(Tile_X0Y2_to_SD),
    .to_SF(Tile_X0Y2_to_SF),
    .to_SG(Tile_X0Y2_to_SG),
    .to_SH(Tile_X0Y2_to_SH),
    .to_SI(Tile_X0Y2_to_SI),
    .A_O_top_0_t(Tile_X0Y2_A_O_top_0_t),
    .A_O_top_0_f(Tile_X0Y2_A_O_top_0_f),
    .A_O_top_1_t(Tile_X0Y2_A_O_top_1_t),
    .A_O_top_1_f(Tile_X0Y2_A_O_top_1_f),
    .A_prech1(Tile_X0Y2_A_prech1),
    .A_prech2(Tile_X0Y2_A_prech2),
    .A_DR_fault(Tile_X0Y2_A_DR_fault),
    .A_I_top_0_t(Tile_X0Y2_A_I_top_0_t),
    .A_I_top_0_f(Tile_X0Y2_A_I_top_0_f),
    .A_I_top_1_t(Tile_X0Y2_A_I_top_1_t),
    .A_I_top_1_f(Tile_X0Y2_A_I_top_1_f),
    .A_T_top(Tile_X0Y2_A_T_top),
    .A_F_masked1(Tile_X0Y2_A_F_masked1),
    .A_F_masked2(Tile_X0Y2_A_F_masked2),
    .A_config_C_bit0(Tile_X0Y2_A_config_C_bit0),
    .A_config_C_bit1(Tile_X0Y2_A_config_C_bit1),
    .A_config_C_bit2(Tile_X0Y2_A_config_C_bit2),
    .A_config_C_bit3(Tile_X0Y2_A_config_C_bit3),
    .B_config_C_bit0(Tile_X0Y2_B_config_C_bit0),
    .B_config_C_bit1(Tile_X0Y2_B_config_C_bit1),
    .B_config_C_bit2(Tile_X0Y2_B_config_C_bit2),
    .B_config_C_bit3(Tile_X0Y2_B_config_C_bit3),
    .UserCLK(Tile_X0Y3_UserCLKo),
    .UserCLKo(Tile_X0Y2_UserCLKo),
    .rst(Tile_X0Y3_rsto),
    .rsto(Tile_X0Y2_rsto),
    .FrameData(Tile_Y2_FrameData),
    .FrameData_O(Tile_X0Y2_FrameData_O),
    .FrameStrobe(Tile_X0Y3_FrameStrobe_O),
    .FrameStrobe_O(Tile_X0Y2_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X1Y2_Emulate_Bitstream)
    )
`endif
    Tile_X1Y2_linear_LMDPL
    (
    .from_NA(Tile_X1Y3_to_NA),
    .from_NB(Tile_X1Y3_to_NB),
    .from_NC(Tile_X1Y3_to_NC),
    .from_ND(Tile_X1Y3_to_ND),
    .from_NF(Tile_X1Y3_to_NF),
    .from_NG(Tile_X1Y3_to_NG),
    .from_NH(Tile_X1Y3_to_NH),
    .from_NI(Tile_X1Y3_to_NI),
    .from_EA(Tile_X0Y2_to_EA),
    .from_EB(Tile_X0Y2_to_EB),
    .from_EC(Tile_X0Y2_to_EC),
    .from_ED(Tile_X0Y2_to_ED),
    .from_EF(Tile_X0Y2_to_EF),
    .from_EG(Tile_X0Y2_to_EG),
    .from_EH(Tile_X0Y2_to_EH),
    .from_EI(Tile_X0Y2_to_EI),
    .from_SA(Tile_X1Y1_to_SA),
    .from_SB(Tile_X1Y1_to_SB),
    .from_SC(Tile_X1Y1_to_SC),
    .from_SD(Tile_X1Y1_to_SD),
    .from_SF(Tile_X1Y1_to_SF),
    .from_SG(Tile_X1Y1_to_SG),
    .from_SH(Tile_X1Y1_to_SH),
    .from_SI(Tile_X1Y1_to_SI),
    .from_WA(Tile_X2Y2_to_WA),
    .from_WB(Tile_X2Y2_to_WB),
    .from_WC(Tile_X2Y2_to_WC),
    .from_WD(Tile_X2Y2_to_WD),
    .from_WF(Tile_X2Y2_to_WF),
    .from_WG(Tile_X2Y2_to_WG),
    .from_WH(Tile_X2Y2_to_WH),
    .from_WI(Tile_X2Y2_to_WI),
    .to_EA(Tile_X1Y2_to_EA),
    .to_EB(Tile_X1Y2_to_EB),
    .to_EC(Tile_X1Y2_to_EC),
    .to_ED(Tile_X1Y2_to_ED),
    .to_EF(Tile_X1Y2_to_EF),
    .to_EG(Tile_X1Y2_to_EG),
    .to_EH(Tile_X1Y2_to_EH),
    .to_EI(Tile_X1Y2_to_EI),
    .to_WA(Tile_X1Y2_to_WA),
    .to_WB(Tile_X1Y2_to_WB),
    .to_WC(Tile_X1Y2_to_WC),
    .to_WD(Tile_X1Y2_to_WD),
    .to_WF(Tile_X1Y2_to_WF),
    .to_WG(Tile_X1Y2_to_WG),
    .to_WH(Tile_X1Y2_to_WH),
    .to_WI(Tile_X1Y2_to_WI),
    .to_NA(Tile_X1Y2_to_NA),
    .to_NB(Tile_X1Y2_to_NB),
    .to_NC(Tile_X1Y2_to_NC),
    .to_ND(Tile_X1Y2_to_ND),
    .to_NF(Tile_X1Y2_to_NF),
    .to_NG(Tile_X1Y2_to_NG),
    .to_NH(Tile_X1Y2_to_NH),
    .to_NI(Tile_X1Y2_to_NI),
    .to_SA(Tile_X1Y2_to_SA),
    .to_SB(Tile_X1Y2_to_SB),
    .to_SC(Tile_X1Y2_to_SC),
    .to_SD(Tile_X1Y2_to_SD),
    .to_SF(Tile_X1Y2_to_SF),
    .to_SG(Tile_X1Y2_to_SG),
    .to_SH(Tile_X1Y2_to_SH),
    .to_SI(Tile_X1Y2_to_SI),
    .F_masked1(Tile_X1Y2_F_masked1),
    .F_masked2(Tile_X1Y2_F_masked2),
    .UserCLK(Tile_X1Y3_UserCLKo),
    .UserCLKo(Tile_X1Y2_UserCLKo),
    .rst(Tile_X1Y3_rsto),
    .rsto(Tile_X1Y2_rsto),
    .FrameData(Tile_X0Y2_FrameData_O),
    .FrameData_O(Tile_X1Y2_FrameData_O),
    .FrameStrobe(Tile_X1Y3_FrameStrobe_O),
    .FrameStrobe_O(Tile_X1Y2_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X2Y2_Emulate_Bitstream)
    )
`endif
    Tile_X2Y2_linear_LMDPL
    (
    .from_NA(Tile_X2Y3_to_NA),
    .from_NB(Tile_X2Y3_to_NB),
    .from_NC(Tile_X2Y3_to_NC),
    .from_ND(Tile_X2Y3_to_ND),
    .from_NF(Tile_X2Y3_to_NF),
    .from_NG(Tile_X2Y3_to_NG),
    .from_NH(Tile_X2Y3_to_NH),
    .from_NI(Tile_X2Y3_to_NI),
    .from_EA(Tile_X1Y2_to_EA),
    .from_EB(Tile_X1Y2_to_EB),
    .from_EC(Tile_X1Y2_to_EC),
    .from_ED(Tile_X1Y2_to_ED),
    .from_EF(Tile_X1Y2_to_EF),
    .from_EG(Tile_X1Y2_to_EG),
    .from_EH(Tile_X1Y2_to_EH),
    .from_EI(Tile_X1Y2_to_EI),
    .from_SA(Tile_X2Y1_to_SA),
    .from_SB(Tile_X2Y1_to_SB),
    .from_SC(Tile_X2Y1_to_SC),
    .from_SD(Tile_X2Y1_to_SD),
    .from_SF(Tile_X2Y1_to_SF),
    .from_SG(Tile_X2Y1_to_SG),
    .from_SH(Tile_X2Y1_to_SH),
    .from_SI(Tile_X2Y1_to_SI),
    .from_WA(Tile_X3Y2_to_WA),
    .from_WB(Tile_X3Y2_to_WB),
    .from_WC(Tile_X3Y2_to_WC),
    .from_WD(Tile_X3Y2_to_WD),
    .from_WF(Tile_X3Y2_to_WF),
    .from_WG(Tile_X3Y2_to_WG),
    .from_WH(Tile_X3Y2_to_WH),
    .from_WI(Tile_X3Y2_to_WI),
    .to_EA(Tile_X2Y2_to_EA),
    .to_EB(Tile_X2Y2_to_EB),
    .to_EC(Tile_X2Y2_to_EC),
    .to_ED(Tile_X2Y2_to_ED),
    .to_EF(Tile_X2Y2_to_EF),
    .to_EG(Tile_X2Y2_to_EG),
    .to_EH(Tile_X2Y2_to_EH),
    .to_EI(Tile_X2Y2_to_EI),
    .to_WA(Tile_X2Y2_to_WA),
    .to_WB(Tile_X2Y2_to_WB),
    .to_WC(Tile_X2Y2_to_WC),
    .to_WD(Tile_X2Y2_to_WD),
    .to_WF(Tile_X2Y2_to_WF),
    .to_WG(Tile_X2Y2_to_WG),
    .to_WH(Tile_X2Y2_to_WH),
    .to_WI(Tile_X2Y2_to_WI),
    .to_NA(Tile_X2Y2_to_NA),
    .to_NB(Tile_X2Y2_to_NB),
    .to_NC(Tile_X2Y2_to_NC),
    .to_ND(Tile_X2Y2_to_ND),
    .to_NF(Tile_X2Y2_to_NF),
    .to_NG(Tile_X2Y2_to_NG),
    .to_NH(Tile_X2Y2_to_NH),
    .to_NI(Tile_X2Y2_to_NI),
    .to_SA(Tile_X2Y2_to_SA),
    .to_SB(Tile_X2Y2_to_SB),
    .to_SC(Tile_X2Y2_to_SC),
    .to_SD(Tile_X2Y2_to_SD),
    .to_SF(Tile_X2Y2_to_SF),
    .to_SG(Tile_X2Y2_to_SG),
    .to_SH(Tile_X2Y2_to_SH),
    .to_SI(Tile_X2Y2_to_SI),
    .F_masked1(Tile_X2Y2_F_masked1),
    .F_masked2(Tile_X2Y2_F_masked2),
    .UserCLK(Tile_X2Y3_UserCLKo),
    .UserCLKo(Tile_X2Y2_UserCLKo),
    .rst(Tile_X2Y3_rsto),
    .rsto(Tile_X2Y2_rsto),
    .FrameData(Tile_X1Y2_FrameData_O),
    .FrameData_O(Tile_X2Y2_FrameData_O),
    .FrameStrobe(Tile_X2Y3_FrameStrobe_O),
    .FrameStrobe_O(Tile_X2Y2_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
nonlinear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X3Y2_Emulate_Bitstream)
    )
`endif
    Tile_X3Y2_nonlinear_LMDPL
    (
    .from_NA(Tile_X3Y3_to_NA),
    .from_NB(Tile_X3Y3_to_NB),
    .from_NC(Tile_X3Y3_to_NC),
    .from_ND(Tile_X3Y3_to_ND),
    .from_NF(Tile_X3Y3_to_NF),
    .from_NG(Tile_X3Y3_to_NG),
    .from_NH(Tile_X3Y3_to_NH),
    .from_NI(Tile_X3Y3_to_NI),
    .from_EA(Tile_X2Y2_to_EA),
    .from_EB(Tile_X2Y2_to_EB),
    .from_EC(Tile_X2Y2_to_EC),
    .from_ED(Tile_X2Y2_to_ED),
    .from_EF(Tile_X2Y2_to_EF),
    .from_EG(Tile_X2Y2_to_EG),
    .from_EH(Tile_X2Y2_to_EH),
    .from_EI(Tile_X2Y2_to_EI),
    .from_SA(Tile_X3Y1_to_SA),
    .from_SB(Tile_X3Y1_to_SB),
    .from_SC(Tile_X3Y1_to_SC),
    .from_SD(Tile_X3Y1_to_SD),
    .from_SF(Tile_X3Y1_to_SF),
    .from_SG(Tile_X3Y1_to_SG),
    .from_SH(Tile_X3Y1_to_SH),
    .from_SI(Tile_X3Y1_to_SI),
    .from_WA(Tile_X4Y2_to_WA),
    .from_WB(Tile_X4Y2_to_WB),
    .from_WC(Tile_X4Y2_to_WC),
    .from_WD(Tile_X4Y2_to_WD),
    .from_WF(Tile_X4Y2_to_WF),
    .from_WG(Tile_X4Y2_to_WG),
    .from_WH(Tile_X4Y2_to_WH),
    .from_WI(Tile_X4Y2_to_WI),
    .to_EA(Tile_X3Y2_to_EA),
    .to_EB(Tile_X3Y2_to_EB),
    .to_EC(Tile_X3Y2_to_EC),
    .to_ED(Tile_X3Y2_to_ED),
    .to_EF(Tile_X3Y2_to_EF),
    .to_EG(Tile_X3Y2_to_EG),
    .to_EH(Tile_X3Y2_to_EH),
    .to_EI(Tile_X3Y2_to_EI),
    .to_WA(Tile_X3Y2_to_WA),
    .to_WB(Tile_X3Y2_to_WB),
    .to_WC(Tile_X3Y2_to_WC),
    .to_WD(Tile_X3Y2_to_WD),
    .to_WF(Tile_X3Y2_to_WF),
    .to_WG(Tile_X3Y2_to_WG),
    .to_WH(Tile_X3Y2_to_WH),
    .to_WI(Tile_X3Y2_to_WI),
    .to_NA(Tile_X3Y2_to_NA),
    .to_NB(Tile_X3Y2_to_NB),
    .to_NC(Tile_X3Y2_to_NC),
    .to_ND(Tile_X3Y2_to_ND),
    .to_NF(Tile_X3Y2_to_NF),
    .to_NG(Tile_X3Y2_to_NG),
    .to_NH(Tile_X3Y2_to_NH),
    .to_NI(Tile_X3Y2_to_NI),
    .to_SA(Tile_X3Y2_to_SA),
    .to_SB(Tile_X3Y2_to_SB),
    .to_SC(Tile_X3Y2_to_SC),
    .to_SD(Tile_X3Y2_to_SD),
    .to_SF(Tile_X3Y2_to_SF),
    .to_SG(Tile_X3Y2_to_SG),
    .to_SH(Tile_X3Y2_to_SH),
    .to_SI(Tile_X3Y2_to_SI),
    .R_t(Tile_X3Y2_R_t),
    .R_f(Tile_X3Y2_R_f),
    .F_masked1(Tile_X3Y2_F_masked1),
    .F_masked2(Tile_X3Y2_F_masked2),
    .UserCLK(Tile_X3Y3_UserCLKo),
    .UserCLKo(Tile_X3Y2_UserCLKo),
    .rst(Tile_X3Y3_rsto),
    .rsto(Tile_X3Y2_rsto),
    .FrameData(Tile_X2Y2_FrameData_O),
    .FrameData_O(Tile_X3Y2_FrameData_O),
    .FrameStrobe(Tile_X3Y3_FrameStrobe_O),
    .FrameStrobe_O(Tile_X3Y2_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X4Y2_Emulate_Bitstream)
    )
`endif
    Tile_X4Y2_linear_LMDPL
    (
    .from_NA(Tile_X4Y3_to_NA),
    .from_NB(Tile_X4Y3_to_NB),
    .from_NC(Tile_X4Y3_to_NC),
    .from_ND(Tile_X4Y3_to_ND),
    .from_NF(Tile_X4Y3_to_NF),
    .from_NG(Tile_X4Y3_to_NG),
    .from_NH(Tile_X4Y3_to_NH),
    .from_NI(Tile_X4Y3_to_NI),
    .from_EA(Tile_X3Y2_to_EA),
    .from_EB(Tile_X3Y2_to_EB),
    .from_EC(Tile_X3Y2_to_EC),
    .from_ED(Tile_X3Y2_to_ED),
    .from_EF(Tile_X3Y2_to_EF),
    .from_EG(Tile_X3Y2_to_EG),
    .from_EH(Tile_X3Y2_to_EH),
    .from_EI(Tile_X3Y2_to_EI),
    .from_SA(Tile_X4Y1_to_SA),
    .from_SB(Tile_X4Y1_to_SB),
    .from_SC(Tile_X4Y1_to_SC),
    .from_SD(Tile_X4Y1_to_SD),
    .from_SF(Tile_X4Y1_to_SF),
    .from_SG(Tile_X4Y1_to_SG),
    .from_SH(Tile_X4Y1_to_SH),
    .from_SI(Tile_X4Y1_to_SI),
    .from_WA(Tile_X5Y2_to_WA),
    .from_WB(Tile_X5Y2_to_WB),
    .from_WC(Tile_X5Y2_to_WC),
    .from_WD(Tile_X5Y2_to_WD),
    .from_WF(Tile_X5Y2_to_WF),
    .from_WG(Tile_X5Y2_to_WG),
    .from_WH(Tile_X5Y2_to_WH),
    .from_WI(Tile_X5Y2_to_WI),
    .to_EA(Tile_X4Y2_to_EA),
    .to_EB(Tile_X4Y2_to_EB),
    .to_EC(Tile_X4Y2_to_EC),
    .to_ED(Tile_X4Y2_to_ED),
    .to_EF(Tile_X4Y2_to_EF),
    .to_EG(Tile_X4Y2_to_EG),
    .to_EH(Tile_X4Y2_to_EH),
    .to_EI(Tile_X4Y2_to_EI),
    .to_WA(Tile_X4Y2_to_WA),
    .to_WB(Tile_X4Y2_to_WB),
    .to_WC(Tile_X4Y2_to_WC),
    .to_WD(Tile_X4Y2_to_WD),
    .to_WF(Tile_X4Y2_to_WF),
    .to_WG(Tile_X4Y2_to_WG),
    .to_WH(Tile_X4Y2_to_WH),
    .to_WI(Tile_X4Y2_to_WI),
    .to_NA(Tile_X4Y2_to_NA),
    .to_NB(Tile_X4Y2_to_NB),
    .to_NC(Tile_X4Y2_to_NC),
    .to_ND(Tile_X4Y2_to_ND),
    .to_NF(Tile_X4Y2_to_NF),
    .to_NG(Tile_X4Y2_to_NG),
    .to_NH(Tile_X4Y2_to_NH),
    .to_NI(Tile_X4Y2_to_NI),
    .to_SA(Tile_X4Y2_to_SA),
    .to_SB(Tile_X4Y2_to_SB),
    .to_SC(Tile_X4Y2_to_SC),
    .to_SD(Tile_X4Y2_to_SD),
    .to_SF(Tile_X4Y2_to_SF),
    .to_SG(Tile_X4Y2_to_SG),
    .to_SH(Tile_X4Y2_to_SH),
    .to_SI(Tile_X4Y2_to_SI),
    .F_masked1(Tile_X4Y2_F_masked1),
    .F_masked2(Tile_X4Y2_F_masked2),
    .UserCLK(Tile_X4Y3_UserCLKo),
    .UserCLKo(Tile_X4Y2_UserCLKo),
    .rst(Tile_X4Y3_rsto),
    .rsto(Tile_X4Y2_rsto),
    .FrameData(Tile_X3Y2_FrameData_O),
    .FrameData_O(Tile_X4Y2_FrameData_O),
    .FrameStrobe(Tile_X4Y3_FrameStrobe_O),
    .FrameStrobe_O(Tile_X4Y2_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X5Y2_Emulate_Bitstream)
    )
`endif
    Tile_X5Y2_linear_LMDPL
    (
    .from_NA(Tile_X5Y3_to_NA),
    .from_NB(Tile_X5Y3_to_NB),
    .from_NC(Tile_X5Y3_to_NC),
    .from_ND(Tile_X5Y3_to_ND),
    .from_NF(Tile_X5Y3_to_NF),
    .from_NG(Tile_X5Y3_to_NG),
    .from_NH(Tile_X5Y3_to_NH),
    .from_NI(Tile_X5Y3_to_NI),
    .from_EA(Tile_X4Y2_to_EA),
    .from_EB(Tile_X4Y2_to_EB),
    .from_EC(Tile_X4Y2_to_EC),
    .from_ED(Tile_X4Y2_to_ED),
    .from_EF(Tile_X4Y2_to_EF),
    .from_EG(Tile_X4Y2_to_EG),
    .from_EH(Tile_X4Y2_to_EH),
    .from_EI(Tile_X4Y2_to_EI),
    .from_SA(Tile_X5Y1_to_SA),
    .from_SB(Tile_X5Y1_to_SB),
    .from_SC(Tile_X5Y1_to_SC),
    .from_SD(Tile_X5Y1_to_SD),
    .from_SF(Tile_X5Y1_to_SF),
    .from_SG(Tile_X5Y1_to_SG),
    .from_SH(Tile_X5Y1_to_SH),
    .from_SI(Tile_X5Y1_to_SI),
    .from_WA(Tile_X6Y2_to_WA),
    .from_WB(Tile_X6Y2_to_WB),
    .from_WC(Tile_X6Y2_to_WC),
    .from_WD(Tile_X6Y2_to_WD),
    .from_WF(Tile_X6Y2_to_WF),
    .from_WG(Tile_X6Y2_to_WG),
    .from_WH(Tile_X6Y2_to_WH),
    .from_WI(Tile_X6Y2_to_WI),
    .to_EA(Tile_X5Y2_to_EA),
    .to_EB(Tile_X5Y2_to_EB),
    .to_EC(Tile_X5Y2_to_EC),
    .to_ED(Tile_X5Y2_to_ED),
    .to_EF(Tile_X5Y2_to_EF),
    .to_EG(Tile_X5Y2_to_EG),
    .to_EH(Tile_X5Y2_to_EH),
    .to_EI(Tile_X5Y2_to_EI),
    .to_WA(Tile_X5Y2_to_WA),
    .to_WB(Tile_X5Y2_to_WB),
    .to_WC(Tile_X5Y2_to_WC),
    .to_WD(Tile_X5Y2_to_WD),
    .to_WF(Tile_X5Y2_to_WF),
    .to_WG(Tile_X5Y2_to_WG),
    .to_WH(Tile_X5Y2_to_WH),
    .to_WI(Tile_X5Y2_to_WI),
    .to_NA(Tile_X5Y2_to_NA),
    .to_NB(Tile_X5Y2_to_NB),
    .to_NC(Tile_X5Y2_to_NC),
    .to_ND(Tile_X5Y2_to_ND),
    .to_NF(Tile_X5Y2_to_NF),
    .to_NG(Tile_X5Y2_to_NG),
    .to_NH(Tile_X5Y2_to_NH),
    .to_NI(Tile_X5Y2_to_NI),
    .to_SA(Tile_X5Y2_to_SA),
    .to_SB(Tile_X5Y2_to_SB),
    .to_SC(Tile_X5Y2_to_SC),
    .to_SD(Tile_X5Y2_to_SD),
    .to_SF(Tile_X5Y2_to_SF),
    .to_SG(Tile_X5Y2_to_SG),
    .to_SH(Tile_X5Y2_to_SH),
    .to_SI(Tile_X5Y2_to_SI),
    .F_masked1(Tile_X5Y2_F_masked1),
    .F_masked2(Tile_X5Y2_F_masked2),
    .UserCLK(Tile_X5Y3_UserCLKo),
    .UserCLKo(Tile_X5Y2_UserCLKo),
    .rst(Tile_X5Y3_rsto),
    .rsto(Tile_X5Y2_rsto),
    .FrameData(Tile_X4Y2_FrameData_O),
    .FrameData_O(Tile_X5Y2_FrameData_O),
    .FrameStrobe(Tile_X5Y3_FrameStrobe_O),
    .FrameStrobe_O(Tile_X5Y2_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
nonlinear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X6Y2_Emulate_Bitstream)
    )
`endif
    Tile_X6Y2_nonlinear_LMDPL
    (
    .from_NA(Tile_X6Y3_to_NA),
    .from_NB(Tile_X6Y3_to_NB),
    .from_NC(Tile_X6Y3_to_NC),
    .from_ND(Tile_X6Y3_to_ND),
    .from_NF(Tile_X6Y3_to_NF),
    .from_NG(Tile_X6Y3_to_NG),
    .from_NH(Tile_X6Y3_to_NH),
    .from_NI(Tile_X6Y3_to_NI),
    .from_EA(Tile_X5Y2_to_EA),
    .from_EB(Tile_X5Y2_to_EB),
    .from_EC(Tile_X5Y2_to_EC),
    .from_ED(Tile_X5Y2_to_ED),
    .from_EF(Tile_X5Y2_to_EF),
    .from_EG(Tile_X5Y2_to_EG),
    .from_EH(Tile_X5Y2_to_EH),
    .from_EI(Tile_X5Y2_to_EI),
    .from_SA(Tile_X6Y1_to_SA),
    .from_SB(Tile_X6Y1_to_SB),
    .from_SC(Tile_X6Y1_to_SC),
    .from_SD(Tile_X6Y1_to_SD),
    .from_SF(Tile_X6Y1_to_SF),
    .from_SG(Tile_X6Y1_to_SG),
    .from_SH(Tile_X6Y1_to_SH),
    .from_SI(Tile_X6Y1_to_SI),
    .from_WA(Tile_X7Y2_to_WA),
    .from_WB(Tile_X7Y2_to_WB),
    .from_WC(Tile_X7Y2_to_WC),
    .from_WD(Tile_X7Y2_to_WD),
    .from_WF(Tile_X7Y2_to_WF),
    .from_WG(Tile_X7Y2_to_WG),
    .from_WH(Tile_X7Y2_to_WH),
    .from_WI(Tile_X7Y2_to_WI),
    .to_EA(Tile_X6Y2_to_EA),
    .to_EB(Tile_X6Y2_to_EB),
    .to_EC(Tile_X6Y2_to_EC),
    .to_ED(Tile_X6Y2_to_ED),
    .to_EF(Tile_X6Y2_to_EF),
    .to_EG(Tile_X6Y2_to_EG),
    .to_EH(Tile_X6Y2_to_EH),
    .to_EI(Tile_X6Y2_to_EI),
    .to_WA(Tile_X6Y2_to_WA),
    .to_WB(Tile_X6Y2_to_WB),
    .to_WC(Tile_X6Y2_to_WC),
    .to_WD(Tile_X6Y2_to_WD),
    .to_WF(Tile_X6Y2_to_WF),
    .to_WG(Tile_X6Y2_to_WG),
    .to_WH(Tile_X6Y2_to_WH),
    .to_WI(Tile_X6Y2_to_WI),
    .to_NA(Tile_X6Y2_to_NA),
    .to_NB(Tile_X6Y2_to_NB),
    .to_NC(Tile_X6Y2_to_NC),
    .to_ND(Tile_X6Y2_to_ND),
    .to_NF(Tile_X6Y2_to_NF),
    .to_NG(Tile_X6Y2_to_NG),
    .to_NH(Tile_X6Y2_to_NH),
    .to_NI(Tile_X6Y2_to_NI),
    .to_SA(Tile_X6Y2_to_SA),
    .to_SB(Tile_X6Y2_to_SB),
    .to_SC(Tile_X6Y2_to_SC),
    .to_SD(Tile_X6Y2_to_SD),
    .to_SF(Tile_X6Y2_to_SF),
    .to_SG(Tile_X6Y2_to_SG),
    .to_SH(Tile_X6Y2_to_SH),
    .to_SI(Tile_X6Y2_to_SI),
    .R_t(Tile_X6Y2_R_t),
    .R_f(Tile_X6Y2_R_f),
    .F_masked1(Tile_X6Y2_F_masked1),
    .F_masked2(Tile_X6Y2_F_masked2),
    .UserCLK(Tile_X6Y3_UserCLKo),
    .UserCLKo(Tile_X6Y2_UserCLKo),
    .rst(Tile_X6Y3_rsto),
    .rsto(Tile_X6Y2_rsto),
    .FrameData(Tile_X5Y2_FrameData_O),
    .FrameData_O(Tile_X6Y2_FrameData_O),
    .FrameStrobe(Tile_X6Y3_FrameStrobe_O),
    .FrameStrobe_O(Tile_X6Y2_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X7Y2_Emulate_Bitstream)
    )
`endif
    Tile_X7Y2_linear_LMDPL
    (
    .from_NA(Tile_X7Y3_to_NA),
    .from_NB(Tile_X7Y3_to_NB),
    .from_NC(Tile_X7Y3_to_NC),
    .from_ND(Tile_X7Y3_to_ND),
    .from_NF(Tile_X7Y3_to_NF),
    .from_NG(Tile_X7Y3_to_NG),
    .from_NH(Tile_X7Y3_to_NH),
    .from_NI(Tile_X7Y3_to_NI),
    .from_EA(Tile_X6Y2_to_EA),
    .from_EB(Tile_X6Y2_to_EB),
    .from_EC(Tile_X6Y2_to_EC),
    .from_ED(Tile_X6Y2_to_ED),
    .from_EF(Tile_X6Y2_to_EF),
    .from_EG(Tile_X6Y2_to_EG),
    .from_EH(Tile_X6Y2_to_EH),
    .from_EI(Tile_X6Y2_to_EI),
    .from_SA(Tile_X7Y1_to_SA),
    .from_SB(Tile_X7Y1_to_SB),
    .from_SC(Tile_X7Y1_to_SC),
    .from_SD(Tile_X7Y1_to_SD),
    .from_SF(Tile_X7Y1_to_SF),
    .from_SG(Tile_X7Y1_to_SG),
    .from_SH(Tile_X7Y1_to_SH),
    .from_SI(Tile_X7Y1_to_SI),
    .from_WA(Tile_X8Y2_to_WA),
    .from_WB(Tile_X8Y2_to_WB),
    .from_WC(Tile_X8Y2_to_WC),
    .from_WD(Tile_X8Y2_to_WD),
    .from_WF(Tile_X8Y2_to_WF),
    .from_WG(Tile_X8Y2_to_WG),
    .from_WH(Tile_X8Y2_to_WH),
    .from_WI(Tile_X8Y2_to_WI),
    .to_EA(Tile_X7Y2_to_EA),
    .to_EB(Tile_X7Y2_to_EB),
    .to_EC(Tile_X7Y2_to_EC),
    .to_ED(Tile_X7Y2_to_ED),
    .to_EF(Tile_X7Y2_to_EF),
    .to_EG(Tile_X7Y2_to_EG),
    .to_EH(Tile_X7Y2_to_EH),
    .to_EI(Tile_X7Y2_to_EI),
    .to_WA(Tile_X7Y2_to_WA),
    .to_WB(Tile_X7Y2_to_WB),
    .to_WC(Tile_X7Y2_to_WC),
    .to_WD(Tile_X7Y2_to_WD),
    .to_WF(Tile_X7Y2_to_WF),
    .to_WG(Tile_X7Y2_to_WG),
    .to_WH(Tile_X7Y2_to_WH),
    .to_WI(Tile_X7Y2_to_WI),
    .to_NA(Tile_X7Y2_to_NA),
    .to_NB(Tile_X7Y2_to_NB),
    .to_NC(Tile_X7Y2_to_NC),
    .to_ND(Tile_X7Y2_to_ND),
    .to_NF(Tile_X7Y2_to_NF),
    .to_NG(Tile_X7Y2_to_NG),
    .to_NH(Tile_X7Y2_to_NH),
    .to_NI(Tile_X7Y2_to_NI),
    .to_SA(Tile_X7Y2_to_SA),
    .to_SB(Tile_X7Y2_to_SB),
    .to_SC(Tile_X7Y2_to_SC),
    .to_SD(Tile_X7Y2_to_SD),
    .to_SF(Tile_X7Y2_to_SF),
    .to_SG(Tile_X7Y2_to_SG),
    .to_SH(Tile_X7Y2_to_SH),
    .to_SI(Tile_X7Y2_to_SI),
    .F_masked1(Tile_X7Y2_F_masked1),
    .F_masked2(Tile_X7Y2_F_masked2),
    .UserCLK(Tile_X7Y3_UserCLKo),
    .UserCLKo(Tile_X7Y2_UserCLKo),
    .rst(Tile_X7Y3_rsto),
    .rsto(Tile_X7Y2_rsto),
    .FrameData(Tile_X6Y2_FrameData_O),
    .FrameData_O(Tile_X7Y2_FrameData_O),
    .FrameStrobe(Tile_X7Y3_FrameStrobe_O),
    .FrameStrobe_O(Tile_X7Y2_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
ctrl_to_sec
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X8Y2_Emulate_Bitstream)
    )
`endif
    Tile_X8Y2_ctrl_to_sec
    (
    .from_NA(Tile_X8Y3_to_NA),
    .from_NB(Tile_X8Y3_to_NB),
    .from_NC(Tile_X8Y3_to_NC),
    .from_ND(Tile_X8Y3_to_ND),
    .from_NF(Tile_X8Y3_to_NF),
    .from_NG(Tile_X8Y3_to_NG),
    .from_NH(Tile_X8Y3_to_NH),
    .from_NI(Tile_X8Y3_to_NI),
    .from_EA(Tile_X7Y2_to_EA),
    .from_EB(Tile_X7Y2_to_EB),
    .from_EC(Tile_X7Y2_to_EC),
    .from_ED(Tile_X7Y2_to_ED),
    .from_EF(Tile_X7Y2_to_EF),
    .from_EG(Tile_X7Y2_to_EG),
    .from_EH(Tile_X7Y2_to_EH),
    .from_EI(Tile_X7Y2_to_EI),
    .from_SA(Tile_X8Y1_to_SA),
    .from_SB(Tile_X8Y1_to_SB),
    .from_SC(Tile_X8Y1_to_SC),
    .from_SD(Tile_X8Y1_to_SD),
    .from_SF(Tile_X8Y1_to_SF),
    .from_SG(Tile_X8Y1_to_SG),
    .from_SH(Tile_X8Y1_to_SH),
    .from_SI(Tile_X8Y1_to_SI),
    .from_WA_1s(Tile_X9Y2_to_WA_1s),
    .from_WB_1s(Tile_X9Y2_to_WB_1s),
    .from_WC_1s(Tile_X9Y2_to_WC_1s),
    .from_WD_1s(Tile_X9Y2_to_WD_1s),
    .from_WF_1s(Tile_X9Y2_to_WF_1s),
    .from_WG_1s(Tile_X9Y2_to_WG_1s),
    .from_WH_1s(Tile_X9Y2_to_WH_1s),
    .from_WI_1s(Tile_X9Y2_to_WI_1s),
    .to_WA(Tile_X8Y2_to_WA),
    .to_WB(Tile_X8Y2_to_WB),
    .to_WC(Tile_X8Y2_to_WC),
    .to_WD(Tile_X8Y2_to_WD),
    .to_WF(Tile_X8Y2_to_WF),
    .to_WG(Tile_X8Y2_to_WG),
    .to_WH(Tile_X8Y2_to_WH),
    .to_WI(Tile_X8Y2_to_WI),
    .to_NA(Tile_X8Y2_to_NA),
    .to_NB(Tile_X8Y2_to_NB),
    .to_NC(Tile_X8Y2_to_NC),
    .to_ND(Tile_X8Y2_to_ND),
    .to_NF(Tile_X8Y2_to_NF),
    .to_NG(Tile_X8Y2_to_NG),
    .to_NH(Tile_X8Y2_to_NH),
    .to_NI(Tile_X8Y2_to_NI),
    .to_SA(Tile_X8Y2_to_SA),
    .to_SB(Tile_X8Y2_to_SB),
    .to_SC(Tile_X8Y2_to_SC),
    .to_SD(Tile_X8Y2_to_SD),
    .to_SF(Tile_X8Y2_to_SF),
    .to_SG(Tile_X8Y2_to_SG),
    .to_SH(Tile_X8Y2_to_SH),
    .to_SI(Tile_X8Y2_to_SI),
    .UserCLK(Tile_X8Y3_UserCLKo),
    .UserCLKo(Tile_X8Y2_UserCLKo),
    .rst(Tile_X8Y3_rsto),
    .rsto(Tile_X8Y2_rsto),
    .FrameData(Tile_X7Y2_FrameData_O),
    .FrameData_O(Tile_X8Y2_FrameData_O),
    .FrameStrobe(Tile_X8Y3_FrameStrobe_O),
    .FrameStrobe_O(Tile_X8Y2_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
combined_WDDL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X9Y2_Emulate_Bitstream)
    )
`endif
    Tile_X9Y2_combined_WDDL
    (
    .from_NA_1s(Tile_X9Y3_to_NA_1s),
    .from_NB_1s(Tile_X9Y3_to_NB_1s),
    .from_NC_1s(Tile_X9Y3_to_NC_1s),
    .from_ND_1s(Tile_X9Y3_to_ND_1s),
    .from_NF_1s(Tile_X9Y3_to_NF_1s),
    .from_NG_1s(Tile_X9Y3_to_NG_1s),
    .from_NH_1s(Tile_X9Y3_to_NH_1s),
    .from_NI_1s(Tile_X9Y3_to_NI_1s),
    .from_SA_1s(Tile_X9Y1_to_SA_1s),
    .from_SB_1s(Tile_X9Y1_to_SB_1s),
    .from_SC_1s(Tile_X9Y1_to_SC_1s),
    .from_SD_1s(Tile_X9Y1_to_SD_1s),
    .from_SF_1s(Tile_X9Y1_to_SF_1s),
    .from_SG_1s(Tile_X9Y1_to_SG_1s),
    .from_SH_1s(Tile_X9Y1_to_SH_1s),
    .from_SI_1s(Tile_X9Y1_to_SI_1s),
    .from_WA_1s(Tile_X10Y2_to_WA_1s),
    .from_WB_1s(Tile_X10Y2_to_WB_1s),
    .from_WC_1s(Tile_X10Y2_to_WC_1s),
    .from_WD_1s(Tile_X10Y2_to_WD_1s),
    .from_WF_1s(Tile_X10Y2_to_WF_1s),
    .from_WG_1s(Tile_X10Y2_to_WG_1s),
    .from_WH_1s(Tile_X10Y2_to_WH_1s),
    .from_WI_1s(Tile_X10Y2_to_WI_1s),
    .to_EA_1s(Tile_X9Y2_to_EA_1s),
    .to_EB_1s(Tile_X9Y2_to_EB_1s),
    .to_EC_1s(Tile_X9Y2_to_EC_1s),
    .to_ED_1s(Tile_X9Y2_to_ED_1s),
    .to_EF_1s(Tile_X9Y2_to_EF_1s),
    .to_EG_1s(Tile_X9Y2_to_EG_1s),
    .to_EH_1s(Tile_X9Y2_to_EH_1s),
    .to_EI_1s(Tile_X9Y2_to_EI_1s),
    .to_WA_1s(Tile_X9Y2_to_WA_1s),
    .to_WB_1s(Tile_X9Y2_to_WB_1s),
    .to_WC_1s(Tile_X9Y2_to_WC_1s),
    .to_WD_1s(Tile_X9Y2_to_WD_1s),
    .to_WF_1s(Tile_X9Y2_to_WF_1s),
    .to_WG_1s(Tile_X9Y2_to_WG_1s),
    .to_WH_1s(Tile_X9Y2_to_WH_1s),
    .to_WI_1s(Tile_X9Y2_to_WI_1s),
    .to_NA_1s(Tile_X9Y2_to_NA_1s),
    .to_NB_1s(Tile_X9Y2_to_NB_1s),
    .to_NC_1s(Tile_X9Y2_to_NC_1s),
    .to_ND_1s(Tile_X9Y2_to_ND_1s),
    .to_NF_1s(Tile_X9Y2_to_NF_1s),
    .to_NG_1s(Tile_X9Y2_to_NG_1s),
    .to_NH_1s(Tile_X9Y2_to_NH_1s),
    .to_NI_1s(Tile_X9Y2_to_NI_1s),
    .to_SA_1s(Tile_X9Y2_to_SA_1s),
    .to_SB_1s(Tile_X9Y2_to_SB_1s),
    .to_SC_1s(Tile_X9Y2_to_SC_1s),
    .to_SD_1s(Tile_X9Y2_to_SD_1s),
    .to_SF_1s(Tile_X9Y2_to_SF_1s),
    .to_SG_1s(Tile_X9Y2_to_SG_1s),
    .to_SH_1s(Tile_X9Y2_to_SH_1s),
    .to_SI_1s(Tile_X9Y2_to_SI_1s),
    .F_ctrl(Tile_X9Y2_F_ctrl),
    .UserCLK(Tile_X9Y3_UserCLKo),
    .UserCLKo(Tile_X9Y2_UserCLKo),
    .rst(Tile_X9Y3_rsto),
    .rsto(Tile_X9Y2_rsto),
    .FrameData(Tile_X8Y2_FrameData_O),
    .FrameData_O(Tile_X9Y2_FrameData_O),
    .FrameStrobe(Tile_X9Y3_FrameStrobe_O),
    .FrameStrobe_O(Tile_X9Y2_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
ctrl_IO
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X10Y2_Emulate_Bitstream)
    )
`endif
    Tile_X10Y2_ctrl_IO
    (
    .from_EA_1s(Tile_X9Y2_to_EA_1s),
    .from_EB_1s(Tile_X9Y2_to_EB_1s),
    .from_EC_1s(Tile_X9Y2_to_EC_1s),
    .from_ED_1s(Tile_X9Y2_to_ED_1s),
    .from_EF_1s(Tile_X9Y2_to_EF_1s),
    .from_EG_1s(Tile_X9Y2_to_EG_1s),
    .from_EH_1s(Tile_X9Y2_to_EH_1s),
    .from_EI_1s(Tile_X9Y2_to_EI_1s),
    .to_WA_1s(Tile_X10Y2_to_WA_1s),
    .to_WB_1s(Tile_X10Y2_to_WB_1s),
    .to_WC_1s(Tile_X10Y2_to_WC_1s),
    .to_WD_1s(Tile_X10Y2_to_WD_1s),
    .to_WF_1s(Tile_X10Y2_to_WF_1s),
    .to_WG_1s(Tile_X10Y2_to_WG_1s),
    .to_WH_1s(Tile_X10Y2_to_WH_1s),
    .to_WI_1s(Tile_X10Y2_to_WI_1s),
    .A_O_top_0_t(Tile_X10Y2_A_O_top_0_t),
    .A_O_top_0_f(Tile_X10Y2_A_O_top_0_f),
    .A_prech2(Tile_X10Y2_A_prech2),
    .A_DR_fault(Tile_X10Y2_A_DR_fault),
    .A_I_top_0_t(Tile_X10Y2_A_I_top_0_t),
    .A_I_top_0_f(Tile_X10Y2_A_I_top_0_f),
    .A_T_top(Tile_X10Y2_A_T_top),
    .A_F_ctrl(Tile_X10Y2_A_F_ctrl),
    .UserCLK(Tile_X10Y3_UserCLKo),
    .UserCLKo(Tile_X10Y2_UserCLKo),
    .rst(Tile_X10Y3_rsto),
    .rsto(Tile_X10Y2_rsto),
    .FrameData(Tile_X9Y2_FrameData_O),
    .FrameData_O(Tile_X10Y2_FrameData_O),
    .FrameStrobe(Tile_X10Y3_FrameStrobe_O),
    .FrameStrobe_O(Tile_X10Y2_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
W_IO_custom
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X0Y3_Emulate_Bitstream)
    )
`endif
    Tile_X0Y3_W_IO_custom
    (
    .from_NA(Tile_X0Y4_to_NA),
    .from_NB(Tile_X0Y4_to_NB),
    .from_NC(Tile_X0Y4_to_NC),
    .from_ND(Tile_X0Y4_to_ND),
    .from_NF(Tile_X0Y4_to_NF),
    .from_NG(Tile_X0Y4_to_NG),
    .from_NH(Tile_X0Y4_to_NH),
    .from_NI(Tile_X0Y4_to_NI),
    .from_SA(Tile_X0Y2_to_SA),
    .from_SB(Tile_X0Y2_to_SB),
    .from_SC(Tile_X0Y2_to_SC),
    .from_SD(Tile_X0Y2_to_SD),
    .from_SF(Tile_X0Y2_to_SF),
    .from_SG(Tile_X0Y2_to_SG),
    .from_SH(Tile_X0Y2_to_SH),
    .from_SI(Tile_X0Y2_to_SI),
    .from_WA(Tile_X1Y3_to_WA),
    .from_WB(Tile_X1Y3_to_WB),
    .from_WC(Tile_X1Y3_to_WC),
    .from_WD(Tile_X1Y3_to_WD),
    .from_WF(Tile_X1Y3_to_WF),
    .from_WG(Tile_X1Y3_to_WG),
    .from_WH(Tile_X1Y3_to_WH),
    .from_WI(Tile_X1Y3_to_WI),
    .to_EA(Tile_X0Y3_to_EA),
    .to_EB(Tile_X0Y3_to_EB),
    .to_EC(Tile_X0Y3_to_EC),
    .to_ED(Tile_X0Y3_to_ED),
    .to_EF(Tile_X0Y3_to_EF),
    .to_EG(Tile_X0Y3_to_EG),
    .to_EH(Tile_X0Y3_to_EH),
    .to_EI(Tile_X0Y3_to_EI),
    .to_NA(Tile_X0Y3_to_NA),
    .to_NB(Tile_X0Y3_to_NB),
    .to_NC(Tile_X0Y3_to_NC),
    .to_ND(Tile_X0Y3_to_ND),
    .to_NF(Tile_X0Y3_to_NF),
    .to_NG(Tile_X0Y3_to_NG),
    .to_NH(Tile_X0Y3_to_NH),
    .to_NI(Tile_X0Y3_to_NI),
    .to_SA(Tile_X0Y3_to_SA),
    .to_SB(Tile_X0Y3_to_SB),
    .to_SC(Tile_X0Y3_to_SC),
    .to_SD(Tile_X0Y3_to_SD),
    .to_SF(Tile_X0Y3_to_SF),
    .to_SG(Tile_X0Y3_to_SG),
    .to_SH(Tile_X0Y3_to_SH),
    .to_SI(Tile_X0Y3_to_SI),
    .A_O_top_0_t(Tile_X0Y3_A_O_top_0_t),
    .A_O_top_0_f(Tile_X0Y3_A_O_top_0_f),
    .A_O_top_1_t(Tile_X0Y3_A_O_top_1_t),
    .A_O_top_1_f(Tile_X0Y3_A_O_top_1_f),
    .A_prech1(Tile_X0Y3_A_prech1),
    .A_prech2(Tile_X0Y3_A_prech2),
    .A_DR_fault(Tile_X0Y3_A_DR_fault),
    .A_I_top_0_t(Tile_X0Y3_A_I_top_0_t),
    .A_I_top_0_f(Tile_X0Y3_A_I_top_0_f),
    .A_I_top_1_t(Tile_X0Y3_A_I_top_1_t),
    .A_I_top_1_f(Tile_X0Y3_A_I_top_1_f),
    .A_T_top(Tile_X0Y3_A_T_top),
    .A_F_masked1(Tile_X0Y3_A_F_masked1),
    .A_F_masked2(Tile_X0Y3_A_F_masked2),
    .A_config_C_bit0(Tile_X0Y3_A_config_C_bit0),
    .A_config_C_bit1(Tile_X0Y3_A_config_C_bit1),
    .A_config_C_bit2(Tile_X0Y3_A_config_C_bit2),
    .A_config_C_bit3(Tile_X0Y3_A_config_C_bit3),
    .B_config_C_bit0(Tile_X0Y3_B_config_C_bit0),
    .B_config_C_bit1(Tile_X0Y3_B_config_C_bit1),
    .B_config_C_bit2(Tile_X0Y3_B_config_C_bit2),
    .B_config_C_bit3(Tile_X0Y3_B_config_C_bit3),
    .UserCLK(Tile_X0Y4_UserCLKo),
    .UserCLKo(Tile_X0Y3_UserCLKo),
    .rst(Tile_X0Y4_rsto),
    .rsto(Tile_X0Y3_rsto),
    .FrameData(Tile_Y3_FrameData),
    .FrameData_O(Tile_X0Y3_FrameData_O),
    .FrameStrobe(Tile_X0Y4_FrameStrobe_O),
    .FrameStrobe_O(Tile_X0Y3_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X1Y3_Emulate_Bitstream)
    )
`endif
    Tile_X1Y3_linear_LMDPL
    (
    .from_NA(Tile_X1Y4_to_NA),
    .from_NB(Tile_X1Y4_to_NB),
    .from_NC(Tile_X1Y4_to_NC),
    .from_ND(Tile_X1Y4_to_ND),
    .from_NF(Tile_X1Y4_to_NF),
    .from_NG(Tile_X1Y4_to_NG),
    .from_NH(Tile_X1Y4_to_NH),
    .from_NI(Tile_X1Y4_to_NI),
    .from_EA(Tile_X0Y3_to_EA),
    .from_EB(Tile_X0Y3_to_EB),
    .from_EC(Tile_X0Y3_to_EC),
    .from_ED(Tile_X0Y3_to_ED),
    .from_EF(Tile_X0Y3_to_EF),
    .from_EG(Tile_X0Y3_to_EG),
    .from_EH(Tile_X0Y3_to_EH),
    .from_EI(Tile_X0Y3_to_EI),
    .from_SA(Tile_X1Y2_to_SA),
    .from_SB(Tile_X1Y2_to_SB),
    .from_SC(Tile_X1Y2_to_SC),
    .from_SD(Tile_X1Y2_to_SD),
    .from_SF(Tile_X1Y2_to_SF),
    .from_SG(Tile_X1Y2_to_SG),
    .from_SH(Tile_X1Y2_to_SH),
    .from_SI(Tile_X1Y2_to_SI),
    .from_WA(Tile_X2Y3_to_WA),
    .from_WB(Tile_X2Y3_to_WB),
    .from_WC(Tile_X2Y3_to_WC),
    .from_WD(Tile_X2Y3_to_WD),
    .from_WF(Tile_X2Y3_to_WF),
    .from_WG(Tile_X2Y3_to_WG),
    .from_WH(Tile_X2Y3_to_WH),
    .from_WI(Tile_X2Y3_to_WI),
    .to_EA(Tile_X1Y3_to_EA),
    .to_EB(Tile_X1Y3_to_EB),
    .to_EC(Tile_X1Y3_to_EC),
    .to_ED(Tile_X1Y3_to_ED),
    .to_EF(Tile_X1Y3_to_EF),
    .to_EG(Tile_X1Y3_to_EG),
    .to_EH(Tile_X1Y3_to_EH),
    .to_EI(Tile_X1Y3_to_EI),
    .to_WA(Tile_X1Y3_to_WA),
    .to_WB(Tile_X1Y3_to_WB),
    .to_WC(Tile_X1Y3_to_WC),
    .to_WD(Tile_X1Y3_to_WD),
    .to_WF(Tile_X1Y3_to_WF),
    .to_WG(Tile_X1Y3_to_WG),
    .to_WH(Tile_X1Y3_to_WH),
    .to_WI(Tile_X1Y3_to_WI),
    .to_NA(Tile_X1Y3_to_NA),
    .to_NB(Tile_X1Y3_to_NB),
    .to_NC(Tile_X1Y3_to_NC),
    .to_ND(Tile_X1Y3_to_ND),
    .to_NF(Tile_X1Y3_to_NF),
    .to_NG(Tile_X1Y3_to_NG),
    .to_NH(Tile_X1Y3_to_NH),
    .to_NI(Tile_X1Y3_to_NI),
    .to_SA(Tile_X1Y3_to_SA),
    .to_SB(Tile_X1Y3_to_SB),
    .to_SC(Tile_X1Y3_to_SC),
    .to_SD(Tile_X1Y3_to_SD),
    .to_SF(Tile_X1Y3_to_SF),
    .to_SG(Tile_X1Y3_to_SG),
    .to_SH(Tile_X1Y3_to_SH),
    .to_SI(Tile_X1Y3_to_SI),
    .F_masked1(Tile_X1Y3_F_masked1),
    .F_masked2(Tile_X1Y3_F_masked2),
    .UserCLK(Tile_X1Y4_UserCLKo),
    .UserCLKo(Tile_X1Y3_UserCLKo),
    .rst(Tile_X1Y4_rsto),
    .rsto(Tile_X1Y3_rsto),
    .FrameData(Tile_X0Y3_FrameData_O),
    .FrameData_O(Tile_X1Y3_FrameData_O),
    .FrameStrobe(Tile_X1Y4_FrameStrobe_O),
    .FrameStrobe_O(Tile_X1Y3_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X2Y3_Emulate_Bitstream)
    )
`endif
    Tile_X2Y3_linear_LMDPL
    (
    .from_NA(Tile_X2Y4_to_NA),
    .from_NB(Tile_X2Y4_to_NB),
    .from_NC(Tile_X2Y4_to_NC),
    .from_ND(Tile_X2Y4_to_ND),
    .from_NF(Tile_X2Y4_to_NF),
    .from_NG(Tile_X2Y4_to_NG),
    .from_NH(Tile_X2Y4_to_NH),
    .from_NI(Tile_X2Y4_to_NI),
    .from_EA(Tile_X1Y3_to_EA),
    .from_EB(Tile_X1Y3_to_EB),
    .from_EC(Tile_X1Y3_to_EC),
    .from_ED(Tile_X1Y3_to_ED),
    .from_EF(Tile_X1Y3_to_EF),
    .from_EG(Tile_X1Y3_to_EG),
    .from_EH(Tile_X1Y3_to_EH),
    .from_EI(Tile_X1Y3_to_EI),
    .from_SA(Tile_X2Y2_to_SA),
    .from_SB(Tile_X2Y2_to_SB),
    .from_SC(Tile_X2Y2_to_SC),
    .from_SD(Tile_X2Y2_to_SD),
    .from_SF(Tile_X2Y2_to_SF),
    .from_SG(Tile_X2Y2_to_SG),
    .from_SH(Tile_X2Y2_to_SH),
    .from_SI(Tile_X2Y2_to_SI),
    .from_WA(Tile_X3Y3_to_WA),
    .from_WB(Tile_X3Y3_to_WB),
    .from_WC(Tile_X3Y3_to_WC),
    .from_WD(Tile_X3Y3_to_WD),
    .from_WF(Tile_X3Y3_to_WF),
    .from_WG(Tile_X3Y3_to_WG),
    .from_WH(Tile_X3Y3_to_WH),
    .from_WI(Tile_X3Y3_to_WI),
    .to_EA(Tile_X2Y3_to_EA),
    .to_EB(Tile_X2Y3_to_EB),
    .to_EC(Tile_X2Y3_to_EC),
    .to_ED(Tile_X2Y3_to_ED),
    .to_EF(Tile_X2Y3_to_EF),
    .to_EG(Tile_X2Y3_to_EG),
    .to_EH(Tile_X2Y3_to_EH),
    .to_EI(Tile_X2Y3_to_EI),
    .to_WA(Tile_X2Y3_to_WA),
    .to_WB(Tile_X2Y3_to_WB),
    .to_WC(Tile_X2Y3_to_WC),
    .to_WD(Tile_X2Y3_to_WD),
    .to_WF(Tile_X2Y3_to_WF),
    .to_WG(Tile_X2Y3_to_WG),
    .to_WH(Tile_X2Y3_to_WH),
    .to_WI(Tile_X2Y3_to_WI),
    .to_NA(Tile_X2Y3_to_NA),
    .to_NB(Tile_X2Y3_to_NB),
    .to_NC(Tile_X2Y3_to_NC),
    .to_ND(Tile_X2Y3_to_ND),
    .to_NF(Tile_X2Y3_to_NF),
    .to_NG(Tile_X2Y3_to_NG),
    .to_NH(Tile_X2Y3_to_NH),
    .to_NI(Tile_X2Y3_to_NI),
    .to_SA(Tile_X2Y3_to_SA),
    .to_SB(Tile_X2Y3_to_SB),
    .to_SC(Tile_X2Y3_to_SC),
    .to_SD(Tile_X2Y3_to_SD),
    .to_SF(Tile_X2Y3_to_SF),
    .to_SG(Tile_X2Y3_to_SG),
    .to_SH(Tile_X2Y3_to_SH),
    .to_SI(Tile_X2Y3_to_SI),
    .F_masked1(Tile_X2Y3_F_masked1),
    .F_masked2(Tile_X2Y3_F_masked2),
    .UserCLK(Tile_X2Y4_UserCLKo),
    .UserCLKo(Tile_X2Y3_UserCLKo),
    .rst(Tile_X2Y4_rsto),
    .rsto(Tile_X2Y3_rsto),
    .FrameData(Tile_X1Y3_FrameData_O),
    .FrameData_O(Tile_X2Y3_FrameData_O),
    .FrameStrobe(Tile_X2Y4_FrameStrobe_O),
    .FrameStrobe_O(Tile_X2Y3_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
nonlinear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X3Y3_Emulate_Bitstream)
    )
`endif
    Tile_X3Y3_nonlinear_LMDPL
    (
    .from_NA(Tile_X3Y4_to_NA),
    .from_NB(Tile_X3Y4_to_NB),
    .from_NC(Tile_X3Y4_to_NC),
    .from_ND(Tile_X3Y4_to_ND),
    .from_NF(Tile_X3Y4_to_NF),
    .from_NG(Tile_X3Y4_to_NG),
    .from_NH(Tile_X3Y4_to_NH),
    .from_NI(Tile_X3Y4_to_NI),
    .from_EA(Tile_X2Y3_to_EA),
    .from_EB(Tile_X2Y3_to_EB),
    .from_EC(Tile_X2Y3_to_EC),
    .from_ED(Tile_X2Y3_to_ED),
    .from_EF(Tile_X2Y3_to_EF),
    .from_EG(Tile_X2Y3_to_EG),
    .from_EH(Tile_X2Y3_to_EH),
    .from_EI(Tile_X2Y3_to_EI),
    .from_SA(Tile_X3Y2_to_SA),
    .from_SB(Tile_X3Y2_to_SB),
    .from_SC(Tile_X3Y2_to_SC),
    .from_SD(Tile_X3Y2_to_SD),
    .from_SF(Tile_X3Y2_to_SF),
    .from_SG(Tile_X3Y2_to_SG),
    .from_SH(Tile_X3Y2_to_SH),
    .from_SI(Tile_X3Y2_to_SI),
    .from_WA(Tile_X4Y3_to_WA),
    .from_WB(Tile_X4Y3_to_WB),
    .from_WC(Tile_X4Y3_to_WC),
    .from_WD(Tile_X4Y3_to_WD),
    .from_WF(Tile_X4Y3_to_WF),
    .from_WG(Tile_X4Y3_to_WG),
    .from_WH(Tile_X4Y3_to_WH),
    .from_WI(Tile_X4Y3_to_WI),
    .to_EA(Tile_X3Y3_to_EA),
    .to_EB(Tile_X3Y3_to_EB),
    .to_EC(Tile_X3Y3_to_EC),
    .to_ED(Tile_X3Y3_to_ED),
    .to_EF(Tile_X3Y3_to_EF),
    .to_EG(Tile_X3Y3_to_EG),
    .to_EH(Tile_X3Y3_to_EH),
    .to_EI(Tile_X3Y3_to_EI),
    .to_WA(Tile_X3Y3_to_WA),
    .to_WB(Tile_X3Y3_to_WB),
    .to_WC(Tile_X3Y3_to_WC),
    .to_WD(Tile_X3Y3_to_WD),
    .to_WF(Tile_X3Y3_to_WF),
    .to_WG(Tile_X3Y3_to_WG),
    .to_WH(Tile_X3Y3_to_WH),
    .to_WI(Tile_X3Y3_to_WI),
    .to_NA(Tile_X3Y3_to_NA),
    .to_NB(Tile_X3Y3_to_NB),
    .to_NC(Tile_X3Y3_to_NC),
    .to_ND(Tile_X3Y3_to_ND),
    .to_NF(Tile_X3Y3_to_NF),
    .to_NG(Tile_X3Y3_to_NG),
    .to_NH(Tile_X3Y3_to_NH),
    .to_NI(Tile_X3Y3_to_NI),
    .to_SA(Tile_X3Y3_to_SA),
    .to_SB(Tile_X3Y3_to_SB),
    .to_SC(Tile_X3Y3_to_SC),
    .to_SD(Tile_X3Y3_to_SD),
    .to_SF(Tile_X3Y3_to_SF),
    .to_SG(Tile_X3Y3_to_SG),
    .to_SH(Tile_X3Y3_to_SH),
    .to_SI(Tile_X3Y3_to_SI),
    .R_t(Tile_X3Y3_R_t),
    .R_f(Tile_X3Y3_R_f),
    .F_masked1(Tile_X3Y3_F_masked1),
    .F_masked2(Tile_X3Y3_F_masked2),
    .UserCLK(Tile_X3Y4_UserCLKo),
    .UserCLKo(Tile_X3Y3_UserCLKo),
    .rst(Tile_X3Y4_rsto),
    .rsto(Tile_X3Y3_rsto),
    .FrameData(Tile_X2Y3_FrameData_O),
    .FrameData_O(Tile_X3Y3_FrameData_O),
    .FrameStrobe(Tile_X3Y4_FrameStrobe_O),
    .FrameStrobe_O(Tile_X3Y3_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X4Y3_Emulate_Bitstream)
    )
`endif
    Tile_X4Y3_linear_LMDPL
    (
    .from_NA(Tile_X4Y4_to_NA),
    .from_NB(Tile_X4Y4_to_NB),
    .from_NC(Tile_X4Y4_to_NC),
    .from_ND(Tile_X4Y4_to_ND),
    .from_NF(Tile_X4Y4_to_NF),
    .from_NG(Tile_X4Y4_to_NG),
    .from_NH(Tile_X4Y4_to_NH),
    .from_NI(Tile_X4Y4_to_NI),
    .from_EA(Tile_X3Y3_to_EA),
    .from_EB(Tile_X3Y3_to_EB),
    .from_EC(Tile_X3Y3_to_EC),
    .from_ED(Tile_X3Y3_to_ED),
    .from_EF(Tile_X3Y3_to_EF),
    .from_EG(Tile_X3Y3_to_EG),
    .from_EH(Tile_X3Y3_to_EH),
    .from_EI(Tile_X3Y3_to_EI),
    .from_SA(Tile_X4Y2_to_SA),
    .from_SB(Tile_X4Y2_to_SB),
    .from_SC(Tile_X4Y2_to_SC),
    .from_SD(Tile_X4Y2_to_SD),
    .from_SF(Tile_X4Y2_to_SF),
    .from_SG(Tile_X4Y2_to_SG),
    .from_SH(Tile_X4Y2_to_SH),
    .from_SI(Tile_X4Y2_to_SI),
    .from_WA(Tile_X5Y3_to_WA),
    .from_WB(Tile_X5Y3_to_WB),
    .from_WC(Tile_X5Y3_to_WC),
    .from_WD(Tile_X5Y3_to_WD),
    .from_WF(Tile_X5Y3_to_WF),
    .from_WG(Tile_X5Y3_to_WG),
    .from_WH(Tile_X5Y3_to_WH),
    .from_WI(Tile_X5Y3_to_WI),
    .to_EA(Tile_X4Y3_to_EA),
    .to_EB(Tile_X4Y3_to_EB),
    .to_EC(Tile_X4Y3_to_EC),
    .to_ED(Tile_X4Y3_to_ED),
    .to_EF(Tile_X4Y3_to_EF),
    .to_EG(Tile_X4Y3_to_EG),
    .to_EH(Tile_X4Y3_to_EH),
    .to_EI(Tile_X4Y3_to_EI),
    .to_WA(Tile_X4Y3_to_WA),
    .to_WB(Tile_X4Y3_to_WB),
    .to_WC(Tile_X4Y3_to_WC),
    .to_WD(Tile_X4Y3_to_WD),
    .to_WF(Tile_X4Y3_to_WF),
    .to_WG(Tile_X4Y3_to_WG),
    .to_WH(Tile_X4Y3_to_WH),
    .to_WI(Tile_X4Y3_to_WI),
    .to_NA(Tile_X4Y3_to_NA),
    .to_NB(Tile_X4Y3_to_NB),
    .to_NC(Tile_X4Y3_to_NC),
    .to_ND(Tile_X4Y3_to_ND),
    .to_NF(Tile_X4Y3_to_NF),
    .to_NG(Tile_X4Y3_to_NG),
    .to_NH(Tile_X4Y3_to_NH),
    .to_NI(Tile_X4Y3_to_NI),
    .to_SA(Tile_X4Y3_to_SA),
    .to_SB(Tile_X4Y3_to_SB),
    .to_SC(Tile_X4Y3_to_SC),
    .to_SD(Tile_X4Y3_to_SD),
    .to_SF(Tile_X4Y3_to_SF),
    .to_SG(Tile_X4Y3_to_SG),
    .to_SH(Tile_X4Y3_to_SH),
    .to_SI(Tile_X4Y3_to_SI),
    .F_masked1(Tile_X4Y3_F_masked1),
    .F_masked2(Tile_X4Y3_F_masked2),
    .UserCLK(Tile_X4Y4_UserCLKo),
    .UserCLKo(Tile_X4Y3_UserCLKo),
    .rst(Tile_X4Y4_rsto),
    .rsto(Tile_X4Y3_rsto),
    .FrameData(Tile_X3Y3_FrameData_O),
    .FrameData_O(Tile_X4Y3_FrameData_O),
    .FrameStrobe(Tile_X4Y4_FrameStrobe_O),
    .FrameStrobe_O(Tile_X4Y3_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X5Y3_Emulate_Bitstream)
    )
`endif
    Tile_X5Y3_linear_LMDPL
    (
    .from_NA(Tile_X5Y4_to_NA),
    .from_NB(Tile_X5Y4_to_NB),
    .from_NC(Tile_X5Y4_to_NC),
    .from_ND(Tile_X5Y4_to_ND),
    .from_NF(Tile_X5Y4_to_NF),
    .from_NG(Tile_X5Y4_to_NG),
    .from_NH(Tile_X5Y4_to_NH),
    .from_NI(Tile_X5Y4_to_NI),
    .from_EA(Tile_X4Y3_to_EA),
    .from_EB(Tile_X4Y3_to_EB),
    .from_EC(Tile_X4Y3_to_EC),
    .from_ED(Tile_X4Y3_to_ED),
    .from_EF(Tile_X4Y3_to_EF),
    .from_EG(Tile_X4Y3_to_EG),
    .from_EH(Tile_X4Y3_to_EH),
    .from_EI(Tile_X4Y3_to_EI),
    .from_SA(Tile_X5Y2_to_SA),
    .from_SB(Tile_X5Y2_to_SB),
    .from_SC(Tile_X5Y2_to_SC),
    .from_SD(Tile_X5Y2_to_SD),
    .from_SF(Tile_X5Y2_to_SF),
    .from_SG(Tile_X5Y2_to_SG),
    .from_SH(Tile_X5Y2_to_SH),
    .from_SI(Tile_X5Y2_to_SI),
    .from_WA(Tile_X6Y3_to_WA),
    .from_WB(Tile_X6Y3_to_WB),
    .from_WC(Tile_X6Y3_to_WC),
    .from_WD(Tile_X6Y3_to_WD),
    .from_WF(Tile_X6Y3_to_WF),
    .from_WG(Tile_X6Y3_to_WG),
    .from_WH(Tile_X6Y3_to_WH),
    .from_WI(Tile_X6Y3_to_WI),
    .to_EA(Tile_X5Y3_to_EA),
    .to_EB(Tile_X5Y3_to_EB),
    .to_EC(Tile_X5Y3_to_EC),
    .to_ED(Tile_X5Y3_to_ED),
    .to_EF(Tile_X5Y3_to_EF),
    .to_EG(Tile_X5Y3_to_EG),
    .to_EH(Tile_X5Y3_to_EH),
    .to_EI(Tile_X5Y3_to_EI),
    .to_WA(Tile_X5Y3_to_WA),
    .to_WB(Tile_X5Y3_to_WB),
    .to_WC(Tile_X5Y3_to_WC),
    .to_WD(Tile_X5Y3_to_WD),
    .to_WF(Tile_X5Y3_to_WF),
    .to_WG(Tile_X5Y3_to_WG),
    .to_WH(Tile_X5Y3_to_WH),
    .to_WI(Tile_X5Y3_to_WI),
    .to_NA(Tile_X5Y3_to_NA),
    .to_NB(Tile_X5Y3_to_NB),
    .to_NC(Tile_X5Y3_to_NC),
    .to_ND(Tile_X5Y3_to_ND),
    .to_NF(Tile_X5Y3_to_NF),
    .to_NG(Tile_X5Y3_to_NG),
    .to_NH(Tile_X5Y3_to_NH),
    .to_NI(Tile_X5Y3_to_NI),
    .to_SA(Tile_X5Y3_to_SA),
    .to_SB(Tile_X5Y3_to_SB),
    .to_SC(Tile_X5Y3_to_SC),
    .to_SD(Tile_X5Y3_to_SD),
    .to_SF(Tile_X5Y3_to_SF),
    .to_SG(Tile_X5Y3_to_SG),
    .to_SH(Tile_X5Y3_to_SH),
    .to_SI(Tile_X5Y3_to_SI),
    .F_masked1(Tile_X5Y3_F_masked1),
    .F_masked2(Tile_X5Y3_F_masked2),
    .UserCLK(Tile_X5Y4_UserCLKo),
    .UserCLKo(Tile_X5Y3_UserCLKo),
    .rst(Tile_X5Y4_rsto),
    .rsto(Tile_X5Y3_rsto),
    .FrameData(Tile_X4Y3_FrameData_O),
    .FrameData_O(Tile_X5Y3_FrameData_O),
    .FrameStrobe(Tile_X5Y4_FrameStrobe_O),
    .FrameStrobe_O(Tile_X5Y3_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
nonlinear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X6Y3_Emulate_Bitstream)
    )
`endif
    Tile_X6Y3_nonlinear_LMDPL
    (
    .from_NA(Tile_X6Y4_to_NA),
    .from_NB(Tile_X6Y4_to_NB),
    .from_NC(Tile_X6Y4_to_NC),
    .from_ND(Tile_X6Y4_to_ND),
    .from_NF(Tile_X6Y4_to_NF),
    .from_NG(Tile_X6Y4_to_NG),
    .from_NH(Tile_X6Y4_to_NH),
    .from_NI(Tile_X6Y4_to_NI),
    .from_EA(Tile_X5Y3_to_EA),
    .from_EB(Tile_X5Y3_to_EB),
    .from_EC(Tile_X5Y3_to_EC),
    .from_ED(Tile_X5Y3_to_ED),
    .from_EF(Tile_X5Y3_to_EF),
    .from_EG(Tile_X5Y3_to_EG),
    .from_EH(Tile_X5Y3_to_EH),
    .from_EI(Tile_X5Y3_to_EI),
    .from_SA(Tile_X6Y2_to_SA),
    .from_SB(Tile_X6Y2_to_SB),
    .from_SC(Tile_X6Y2_to_SC),
    .from_SD(Tile_X6Y2_to_SD),
    .from_SF(Tile_X6Y2_to_SF),
    .from_SG(Tile_X6Y2_to_SG),
    .from_SH(Tile_X6Y2_to_SH),
    .from_SI(Tile_X6Y2_to_SI),
    .from_WA(Tile_X7Y3_to_WA),
    .from_WB(Tile_X7Y3_to_WB),
    .from_WC(Tile_X7Y3_to_WC),
    .from_WD(Tile_X7Y3_to_WD),
    .from_WF(Tile_X7Y3_to_WF),
    .from_WG(Tile_X7Y3_to_WG),
    .from_WH(Tile_X7Y3_to_WH),
    .from_WI(Tile_X7Y3_to_WI),
    .to_EA(Tile_X6Y3_to_EA),
    .to_EB(Tile_X6Y3_to_EB),
    .to_EC(Tile_X6Y3_to_EC),
    .to_ED(Tile_X6Y3_to_ED),
    .to_EF(Tile_X6Y3_to_EF),
    .to_EG(Tile_X6Y3_to_EG),
    .to_EH(Tile_X6Y3_to_EH),
    .to_EI(Tile_X6Y3_to_EI),
    .to_WA(Tile_X6Y3_to_WA),
    .to_WB(Tile_X6Y3_to_WB),
    .to_WC(Tile_X6Y3_to_WC),
    .to_WD(Tile_X6Y3_to_WD),
    .to_WF(Tile_X6Y3_to_WF),
    .to_WG(Tile_X6Y3_to_WG),
    .to_WH(Tile_X6Y3_to_WH),
    .to_WI(Tile_X6Y3_to_WI),
    .to_NA(Tile_X6Y3_to_NA),
    .to_NB(Tile_X6Y3_to_NB),
    .to_NC(Tile_X6Y3_to_NC),
    .to_ND(Tile_X6Y3_to_ND),
    .to_NF(Tile_X6Y3_to_NF),
    .to_NG(Tile_X6Y3_to_NG),
    .to_NH(Tile_X6Y3_to_NH),
    .to_NI(Tile_X6Y3_to_NI),
    .to_SA(Tile_X6Y3_to_SA),
    .to_SB(Tile_X6Y3_to_SB),
    .to_SC(Tile_X6Y3_to_SC),
    .to_SD(Tile_X6Y3_to_SD),
    .to_SF(Tile_X6Y3_to_SF),
    .to_SG(Tile_X6Y3_to_SG),
    .to_SH(Tile_X6Y3_to_SH),
    .to_SI(Tile_X6Y3_to_SI),
    .R_t(Tile_X6Y3_R_t),
    .R_f(Tile_X6Y3_R_f),
    .F_masked1(Tile_X6Y3_F_masked1),
    .F_masked2(Tile_X6Y3_F_masked2),
    .UserCLK(Tile_X6Y4_UserCLKo),
    .UserCLKo(Tile_X6Y3_UserCLKo),
    .rst(Tile_X6Y4_rsto),
    .rsto(Tile_X6Y3_rsto),
    .FrameData(Tile_X5Y3_FrameData_O),
    .FrameData_O(Tile_X6Y3_FrameData_O),
    .FrameStrobe(Tile_X6Y4_FrameStrobe_O),
    .FrameStrobe_O(Tile_X6Y3_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X7Y3_Emulate_Bitstream)
    )
`endif
    Tile_X7Y3_linear_LMDPL
    (
    .from_NA(Tile_X7Y4_to_NA),
    .from_NB(Tile_X7Y4_to_NB),
    .from_NC(Tile_X7Y4_to_NC),
    .from_ND(Tile_X7Y4_to_ND),
    .from_NF(Tile_X7Y4_to_NF),
    .from_NG(Tile_X7Y4_to_NG),
    .from_NH(Tile_X7Y4_to_NH),
    .from_NI(Tile_X7Y4_to_NI),
    .from_EA(Tile_X6Y3_to_EA),
    .from_EB(Tile_X6Y3_to_EB),
    .from_EC(Tile_X6Y3_to_EC),
    .from_ED(Tile_X6Y3_to_ED),
    .from_EF(Tile_X6Y3_to_EF),
    .from_EG(Tile_X6Y3_to_EG),
    .from_EH(Tile_X6Y3_to_EH),
    .from_EI(Tile_X6Y3_to_EI),
    .from_SA(Tile_X7Y2_to_SA),
    .from_SB(Tile_X7Y2_to_SB),
    .from_SC(Tile_X7Y2_to_SC),
    .from_SD(Tile_X7Y2_to_SD),
    .from_SF(Tile_X7Y2_to_SF),
    .from_SG(Tile_X7Y2_to_SG),
    .from_SH(Tile_X7Y2_to_SH),
    .from_SI(Tile_X7Y2_to_SI),
    .from_WA(Tile_X8Y3_to_WA),
    .from_WB(Tile_X8Y3_to_WB),
    .from_WC(Tile_X8Y3_to_WC),
    .from_WD(Tile_X8Y3_to_WD),
    .from_WF(Tile_X8Y3_to_WF),
    .from_WG(Tile_X8Y3_to_WG),
    .from_WH(Tile_X8Y3_to_WH),
    .from_WI(Tile_X8Y3_to_WI),
    .to_EA(Tile_X7Y3_to_EA),
    .to_EB(Tile_X7Y3_to_EB),
    .to_EC(Tile_X7Y3_to_EC),
    .to_ED(Tile_X7Y3_to_ED),
    .to_EF(Tile_X7Y3_to_EF),
    .to_EG(Tile_X7Y3_to_EG),
    .to_EH(Tile_X7Y3_to_EH),
    .to_EI(Tile_X7Y3_to_EI),
    .to_WA(Tile_X7Y3_to_WA),
    .to_WB(Tile_X7Y3_to_WB),
    .to_WC(Tile_X7Y3_to_WC),
    .to_WD(Tile_X7Y3_to_WD),
    .to_WF(Tile_X7Y3_to_WF),
    .to_WG(Tile_X7Y3_to_WG),
    .to_WH(Tile_X7Y3_to_WH),
    .to_WI(Tile_X7Y3_to_WI),
    .to_NA(Tile_X7Y3_to_NA),
    .to_NB(Tile_X7Y3_to_NB),
    .to_NC(Tile_X7Y3_to_NC),
    .to_ND(Tile_X7Y3_to_ND),
    .to_NF(Tile_X7Y3_to_NF),
    .to_NG(Tile_X7Y3_to_NG),
    .to_NH(Tile_X7Y3_to_NH),
    .to_NI(Tile_X7Y3_to_NI),
    .to_SA(Tile_X7Y3_to_SA),
    .to_SB(Tile_X7Y3_to_SB),
    .to_SC(Tile_X7Y3_to_SC),
    .to_SD(Tile_X7Y3_to_SD),
    .to_SF(Tile_X7Y3_to_SF),
    .to_SG(Tile_X7Y3_to_SG),
    .to_SH(Tile_X7Y3_to_SH),
    .to_SI(Tile_X7Y3_to_SI),
    .F_masked1(Tile_X7Y3_F_masked1),
    .F_masked2(Tile_X7Y3_F_masked2),
    .UserCLK(Tile_X7Y4_UserCLKo),
    .UserCLKo(Tile_X7Y3_UserCLKo),
    .rst(Tile_X7Y4_rsto),
    .rsto(Tile_X7Y3_rsto),
    .FrameData(Tile_X6Y3_FrameData_O),
    .FrameData_O(Tile_X7Y3_FrameData_O),
    .FrameStrobe(Tile_X7Y4_FrameStrobe_O),
    .FrameStrobe_O(Tile_X7Y3_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
ctrl_to_sec
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X8Y3_Emulate_Bitstream)
    )
`endif
    Tile_X8Y3_ctrl_to_sec
    (
    .from_NA(Tile_X8Y4_to_NA),
    .from_NB(Tile_X8Y4_to_NB),
    .from_NC(Tile_X8Y4_to_NC),
    .from_ND(Tile_X8Y4_to_ND),
    .from_NF(Tile_X8Y4_to_NF),
    .from_NG(Tile_X8Y4_to_NG),
    .from_NH(Tile_X8Y4_to_NH),
    .from_NI(Tile_X8Y4_to_NI),
    .from_EA(Tile_X7Y3_to_EA),
    .from_EB(Tile_X7Y3_to_EB),
    .from_EC(Tile_X7Y3_to_EC),
    .from_ED(Tile_X7Y3_to_ED),
    .from_EF(Tile_X7Y3_to_EF),
    .from_EG(Tile_X7Y3_to_EG),
    .from_EH(Tile_X7Y3_to_EH),
    .from_EI(Tile_X7Y3_to_EI),
    .from_SA(Tile_X8Y2_to_SA),
    .from_SB(Tile_X8Y2_to_SB),
    .from_SC(Tile_X8Y2_to_SC),
    .from_SD(Tile_X8Y2_to_SD),
    .from_SF(Tile_X8Y2_to_SF),
    .from_SG(Tile_X8Y2_to_SG),
    .from_SH(Tile_X8Y2_to_SH),
    .from_SI(Tile_X8Y2_to_SI),
    .from_WA_1s(Tile_X9Y3_to_WA_1s),
    .from_WB_1s(Tile_X9Y3_to_WB_1s),
    .from_WC_1s(Tile_X9Y3_to_WC_1s),
    .from_WD_1s(Tile_X9Y3_to_WD_1s),
    .from_WF_1s(Tile_X9Y3_to_WF_1s),
    .from_WG_1s(Tile_X9Y3_to_WG_1s),
    .from_WH_1s(Tile_X9Y3_to_WH_1s),
    .from_WI_1s(Tile_X9Y3_to_WI_1s),
    .to_WA(Tile_X8Y3_to_WA),
    .to_WB(Tile_X8Y3_to_WB),
    .to_WC(Tile_X8Y3_to_WC),
    .to_WD(Tile_X8Y3_to_WD),
    .to_WF(Tile_X8Y3_to_WF),
    .to_WG(Tile_X8Y3_to_WG),
    .to_WH(Tile_X8Y3_to_WH),
    .to_WI(Tile_X8Y3_to_WI),
    .to_NA(Tile_X8Y3_to_NA),
    .to_NB(Tile_X8Y3_to_NB),
    .to_NC(Tile_X8Y3_to_NC),
    .to_ND(Tile_X8Y3_to_ND),
    .to_NF(Tile_X8Y3_to_NF),
    .to_NG(Tile_X8Y3_to_NG),
    .to_NH(Tile_X8Y3_to_NH),
    .to_NI(Tile_X8Y3_to_NI),
    .to_SA(Tile_X8Y3_to_SA),
    .to_SB(Tile_X8Y3_to_SB),
    .to_SC(Tile_X8Y3_to_SC),
    .to_SD(Tile_X8Y3_to_SD),
    .to_SF(Tile_X8Y3_to_SF),
    .to_SG(Tile_X8Y3_to_SG),
    .to_SH(Tile_X8Y3_to_SH),
    .to_SI(Tile_X8Y3_to_SI),
    .UserCLK(Tile_X8Y4_UserCLKo),
    .UserCLKo(Tile_X8Y3_UserCLKo),
    .rst(Tile_X8Y4_rsto),
    .rsto(Tile_X8Y3_rsto),
    .FrameData(Tile_X7Y3_FrameData_O),
    .FrameData_O(Tile_X8Y3_FrameData_O),
    .FrameStrobe(Tile_X8Y4_FrameStrobe_O),
    .FrameStrobe_O(Tile_X8Y3_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
combined_WDDL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X9Y3_Emulate_Bitstream)
    )
`endif
    Tile_X9Y3_combined_WDDL
    (
    .from_NA_1s(Tile_X9Y4_to_NA_1s),
    .from_NB_1s(Tile_X9Y4_to_NB_1s),
    .from_NC_1s(Tile_X9Y4_to_NC_1s),
    .from_ND_1s(Tile_X9Y4_to_ND_1s),
    .from_NF_1s(Tile_X9Y4_to_NF_1s),
    .from_NG_1s(Tile_X9Y4_to_NG_1s),
    .from_NH_1s(Tile_X9Y4_to_NH_1s),
    .from_NI_1s(Tile_X9Y4_to_NI_1s),
    .from_SA_1s(Tile_X9Y2_to_SA_1s),
    .from_SB_1s(Tile_X9Y2_to_SB_1s),
    .from_SC_1s(Tile_X9Y2_to_SC_1s),
    .from_SD_1s(Tile_X9Y2_to_SD_1s),
    .from_SF_1s(Tile_X9Y2_to_SF_1s),
    .from_SG_1s(Tile_X9Y2_to_SG_1s),
    .from_SH_1s(Tile_X9Y2_to_SH_1s),
    .from_SI_1s(Tile_X9Y2_to_SI_1s),
    .from_WA_1s(Tile_X10Y3_to_WA_1s),
    .from_WB_1s(Tile_X10Y3_to_WB_1s),
    .from_WC_1s(Tile_X10Y3_to_WC_1s),
    .from_WD_1s(Tile_X10Y3_to_WD_1s),
    .from_WF_1s(Tile_X10Y3_to_WF_1s),
    .from_WG_1s(Tile_X10Y3_to_WG_1s),
    .from_WH_1s(Tile_X10Y3_to_WH_1s),
    .from_WI_1s(Tile_X10Y3_to_WI_1s),
    .to_EA_1s(Tile_X9Y3_to_EA_1s),
    .to_EB_1s(Tile_X9Y3_to_EB_1s),
    .to_EC_1s(Tile_X9Y3_to_EC_1s),
    .to_ED_1s(Tile_X9Y3_to_ED_1s),
    .to_EF_1s(Tile_X9Y3_to_EF_1s),
    .to_EG_1s(Tile_X9Y3_to_EG_1s),
    .to_EH_1s(Tile_X9Y3_to_EH_1s),
    .to_EI_1s(Tile_X9Y3_to_EI_1s),
    .to_WA_1s(Tile_X9Y3_to_WA_1s),
    .to_WB_1s(Tile_X9Y3_to_WB_1s),
    .to_WC_1s(Tile_X9Y3_to_WC_1s),
    .to_WD_1s(Tile_X9Y3_to_WD_1s),
    .to_WF_1s(Tile_X9Y3_to_WF_1s),
    .to_WG_1s(Tile_X9Y3_to_WG_1s),
    .to_WH_1s(Tile_X9Y3_to_WH_1s),
    .to_WI_1s(Tile_X9Y3_to_WI_1s),
    .to_NA_1s(Tile_X9Y3_to_NA_1s),
    .to_NB_1s(Tile_X9Y3_to_NB_1s),
    .to_NC_1s(Tile_X9Y3_to_NC_1s),
    .to_ND_1s(Tile_X9Y3_to_ND_1s),
    .to_NF_1s(Tile_X9Y3_to_NF_1s),
    .to_NG_1s(Tile_X9Y3_to_NG_1s),
    .to_NH_1s(Tile_X9Y3_to_NH_1s),
    .to_NI_1s(Tile_X9Y3_to_NI_1s),
    .to_SA_1s(Tile_X9Y3_to_SA_1s),
    .to_SB_1s(Tile_X9Y3_to_SB_1s),
    .to_SC_1s(Tile_X9Y3_to_SC_1s),
    .to_SD_1s(Tile_X9Y3_to_SD_1s),
    .to_SF_1s(Tile_X9Y3_to_SF_1s),
    .to_SG_1s(Tile_X9Y3_to_SG_1s),
    .to_SH_1s(Tile_X9Y3_to_SH_1s),
    .to_SI_1s(Tile_X9Y3_to_SI_1s),
    .F_ctrl(Tile_X9Y3_F_ctrl),
    .UserCLK(Tile_X9Y4_UserCLKo),
    .UserCLKo(Tile_X9Y3_UserCLKo),
    .rst(Tile_X9Y4_rsto),
    .rsto(Tile_X9Y3_rsto),
    .FrameData(Tile_X8Y3_FrameData_O),
    .FrameData_O(Tile_X9Y3_FrameData_O),
    .FrameStrobe(Tile_X9Y4_FrameStrobe_O),
    .FrameStrobe_O(Tile_X9Y3_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
ctrl_IO
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X10Y3_Emulate_Bitstream)
    )
`endif
    Tile_X10Y3_ctrl_IO
    (
    .from_EA_1s(Tile_X9Y3_to_EA_1s),
    .from_EB_1s(Tile_X9Y3_to_EB_1s),
    .from_EC_1s(Tile_X9Y3_to_EC_1s),
    .from_ED_1s(Tile_X9Y3_to_ED_1s),
    .from_EF_1s(Tile_X9Y3_to_EF_1s),
    .from_EG_1s(Tile_X9Y3_to_EG_1s),
    .from_EH_1s(Tile_X9Y3_to_EH_1s),
    .from_EI_1s(Tile_X9Y3_to_EI_1s),
    .to_WA_1s(Tile_X10Y3_to_WA_1s),
    .to_WB_1s(Tile_X10Y3_to_WB_1s),
    .to_WC_1s(Tile_X10Y3_to_WC_1s),
    .to_WD_1s(Tile_X10Y3_to_WD_1s),
    .to_WF_1s(Tile_X10Y3_to_WF_1s),
    .to_WG_1s(Tile_X10Y3_to_WG_1s),
    .to_WH_1s(Tile_X10Y3_to_WH_1s),
    .to_WI_1s(Tile_X10Y3_to_WI_1s),
    .A_O_top_0_t(Tile_X10Y3_A_O_top_0_t),
    .A_O_top_0_f(Tile_X10Y3_A_O_top_0_f),
    .A_prech2(Tile_X10Y3_A_prech2),
    .A_DR_fault(Tile_X10Y3_A_DR_fault),
    .A_I_top_0_t(Tile_X10Y3_A_I_top_0_t),
    .A_I_top_0_f(Tile_X10Y3_A_I_top_0_f),
    .A_T_top(Tile_X10Y3_A_T_top),
    .A_F_ctrl(Tile_X10Y3_A_F_ctrl),
    .UserCLK(Tile_X10Y4_UserCLKo),
    .UserCLKo(Tile_X10Y3_UserCLKo),
    .rst(Tile_X10Y4_rsto),
    .rsto(Tile_X10Y3_rsto),
    .FrameData(Tile_X9Y3_FrameData_O),
    .FrameData_O(Tile_X10Y3_FrameData_O),
    .FrameStrobe(Tile_X10Y4_FrameStrobe_O),
    .FrameStrobe_O(Tile_X10Y3_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
W_IO_custom
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X0Y4_Emulate_Bitstream)
    )
`endif
    Tile_X0Y4_W_IO_custom
    (
    .from_NA(Tile_X0Y5_to_NA),
    .from_NB(Tile_X0Y5_to_NB),
    .from_NC(Tile_X0Y5_to_NC),
    .from_ND(Tile_X0Y5_to_ND),
    .from_NF(Tile_X0Y5_to_NF),
    .from_NG(Tile_X0Y5_to_NG),
    .from_NH(Tile_X0Y5_to_NH),
    .from_NI(Tile_X0Y5_to_NI),
    .from_SA(Tile_X0Y3_to_SA),
    .from_SB(Tile_X0Y3_to_SB),
    .from_SC(Tile_X0Y3_to_SC),
    .from_SD(Tile_X0Y3_to_SD),
    .from_SF(Tile_X0Y3_to_SF),
    .from_SG(Tile_X0Y3_to_SG),
    .from_SH(Tile_X0Y3_to_SH),
    .from_SI(Tile_X0Y3_to_SI),
    .from_WA(Tile_X1Y4_to_WA),
    .from_WB(Tile_X1Y4_to_WB),
    .from_WC(Tile_X1Y4_to_WC),
    .from_WD(Tile_X1Y4_to_WD),
    .from_WF(Tile_X1Y4_to_WF),
    .from_WG(Tile_X1Y4_to_WG),
    .from_WH(Tile_X1Y4_to_WH),
    .from_WI(Tile_X1Y4_to_WI),
    .to_EA(Tile_X0Y4_to_EA),
    .to_EB(Tile_X0Y4_to_EB),
    .to_EC(Tile_X0Y4_to_EC),
    .to_ED(Tile_X0Y4_to_ED),
    .to_EF(Tile_X0Y4_to_EF),
    .to_EG(Tile_X0Y4_to_EG),
    .to_EH(Tile_X0Y4_to_EH),
    .to_EI(Tile_X0Y4_to_EI),
    .to_NA(Tile_X0Y4_to_NA),
    .to_NB(Tile_X0Y4_to_NB),
    .to_NC(Tile_X0Y4_to_NC),
    .to_ND(Tile_X0Y4_to_ND),
    .to_NF(Tile_X0Y4_to_NF),
    .to_NG(Tile_X0Y4_to_NG),
    .to_NH(Tile_X0Y4_to_NH),
    .to_NI(Tile_X0Y4_to_NI),
    .to_SA(Tile_X0Y4_to_SA),
    .to_SB(Tile_X0Y4_to_SB),
    .to_SC(Tile_X0Y4_to_SC),
    .to_SD(Tile_X0Y4_to_SD),
    .to_SF(Tile_X0Y4_to_SF),
    .to_SG(Tile_X0Y4_to_SG),
    .to_SH(Tile_X0Y4_to_SH),
    .to_SI(Tile_X0Y4_to_SI),
    .A_O_top_0_t(Tile_X0Y4_A_O_top_0_t),
    .A_O_top_0_f(Tile_X0Y4_A_O_top_0_f),
    .A_O_top_1_t(Tile_X0Y4_A_O_top_1_t),
    .A_O_top_1_f(Tile_X0Y4_A_O_top_1_f),
    .A_prech1(Tile_X0Y4_A_prech1),
    .A_prech2(Tile_X0Y4_A_prech2),
    .A_DR_fault(Tile_X0Y4_A_DR_fault),
    .A_I_top_0_t(Tile_X0Y4_A_I_top_0_t),
    .A_I_top_0_f(Tile_X0Y4_A_I_top_0_f),
    .A_I_top_1_t(Tile_X0Y4_A_I_top_1_t),
    .A_I_top_1_f(Tile_X0Y4_A_I_top_1_f),
    .A_T_top(Tile_X0Y4_A_T_top),
    .A_F_masked1(Tile_X0Y4_A_F_masked1),
    .A_F_masked2(Tile_X0Y4_A_F_masked2),
    .A_config_C_bit0(Tile_X0Y4_A_config_C_bit0),
    .A_config_C_bit1(Tile_X0Y4_A_config_C_bit1),
    .A_config_C_bit2(Tile_X0Y4_A_config_C_bit2),
    .A_config_C_bit3(Tile_X0Y4_A_config_C_bit3),
    .B_config_C_bit0(Tile_X0Y4_B_config_C_bit0),
    .B_config_C_bit1(Tile_X0Y4_B_config_C_bit1),
    .B_config_C_bit2(Tile_X0Y4_B_config_C_bit2),
    .B_config_C_bit3(Tile_X0Y4_B_config_C_bit3),
    .UserCLK(Tile_X0Y5_UserCLKo),
    .UserCLKo(Tile_X0Y4_UserCLKo),
    .rst(Tile_X0Y5_rsto),
    .rsto(Tile_X0Y4_rsto),
    .FrameData(Tile_Y4_FrameData),
    .FrameData_O(Tile_X0Y4_FrameData_O),
    .FrameStrobe(Tile_X0Y5_FrameStrobe_O),
    .FrameStrobe_O(Tile_X0Y4_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X1Y4_Emulate_Bitstream)
    )
`endif
    Tile_X1Y4_linear_LMDPL
    (
    .from_NA(Tile_X1Y5_to_NA),
    .from_NB(Tile_X1Y5_to_NB),
    .from_NC(Tile_X1Y5_to_NC),
    .from_ND(Tile_X1Y5_to_ND),
    .from_NF(Tile_X1Y5_to_NF),
    .from_NG(Tile_X1Y5_to_NG),
    .from_NH(Tile_X1Y5_to_NH),
    .from_NI(Tile_X1Y5_to_NI),
    .from_EA(Tile_X0Y4_to_EA),
    .from_EB(Tile_X0Y4_to_EB),
    .from_EC(Tile_X0Y4_to_EC),
    .from_ED(Tile_X0Y4_to_ED),
    .from_EF(Tile_X0Y4_to_EF),
    .from_EG(Tile_X0Y4_to_EG),
    .from_EH(Tile_X0Y4_to_EH),
    .from_EI(Tile_X0Y4_to_EI),
    .from_SA(Tile_X1Y3_to_SA),
    .from_SB(Tile_X1Y3_to_SB),
    .from_SC(Tile_X1Y3_to_SC),
    .from_SD(Tile_X1Y3_to_SD),
    .from_SF(Tile_X1Y3_to_SF),
    .from_SG(Tile_X1Y3_to_SG),
    .from_SH(Tile_X1Y3_to_SH),
    .from_SI(Tile_X1Y3_to_SI),
    .from_WA(Tile_X2Y4_to_WA),
    .from_WB(Tile_X2Y4_to_WB),
    .from_WC(Tile_X2Y4_to_WC),
    .from_WD(Tile_X2Y4_to_WD),
    .from_WF(Tile_X2Y4_to_WF),
    .from_WG(Tile_X2Y4_to_WG),
    .from_WH(Tile_X2Y4_to_WH),
    .from_WI(Tile_X2Y4_to_WI),
    .to_EA(Tile_X1Y4_to_EA),
    .to_EB(Tile_X1Y4_to_EB),
    .to_EC(Tile_X1Y4_to_EC),
    .to_ED(Tile_X1Y4_to_ED),
    .to_EF(Tile_X1Y4_to_EF),
    .to_EG(Tile_X1Y4_to_EG),
    .to_EH(Tile_X1Y4_to_EH),
    .to_EI(Tile_X1Y4_to_EI),
    .to_WA(Tile_X1Y4_to_WA),
    .to_WB(Tile_X1Y4_to_WB),
    .to_WC(Tile_X1Y4_to_WC),
    .to_WD(Tile_X1Y4_to_WD),
    .to_WF(Tile_X1Y4_to_WF),
    .to_WG(Tile_X1Y4_to_WG),
    .to_WH(Tile_X1Y4_to_WH),
    .to_WI(Tile_X1Y4_to_WI),
    .to_NA(Tile_X1Y4_to_NA),
    .to_NB(Tile_X1Y4_to_NB),
    .to_NC(Tile_X1Y4_to_NC),
    .to_ND(Tile_X1Y4_to_ND),
    .to_NF(Tile_X1Y4_to_NF),
    .to_NG(Tile_X1Y4_to_NG),
    .to_NH(Tile_X1Y4_to_NH),
    .to_NI(Tile_X1Y4_to_NI),
    .to_SA(Tile_X1Y4_to_SA),
    .to_SB(Tile_X1Y4_to_SB),
    .to_SC(Tile_X1Y4_to_SC),
    .to_SD(Tile_X1Y4_to_SD),
    .to_SF(Tile_X1Y4_to_SF),
    .to_SG(Tile_X1Y4_to_SG),
    .to_SH(Tile_X1Y4_to_SH),
    .to_SI(Tile_X1Y4_to_SI),
    .F_masked1(Tile_X1Y4_F_masked1),
    .F_masked2(Tile_X1Y4_F_masked2),
    .UserCLK(Tile_X1Y5_UserCLKo),
    .UserCLKo(Tile_X1Y4_UserCLKo),
    .rst(Tile_X1Y5_rsto),
    .rsto(Tile_X1Y4_rsto),
    .FrameData(Tile_X0Y4_FrameData_O),
    .FrameData_O(Tile_X1Y4_FrameData_O),
    .FrameStrobe(Tile_X1Y5_FrameStrobe_O),
    .FrameStrobe_O(Tile_X1Y4_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X2Y4_Emulate_Bitstream)
    )
`endif
    Tile_X2Y4_linear_LMDPL
    (
    .from_NA(Tile_X2Y5_to_NA),
    .from_NB(Tile_X2Y5_to_NB),
    .from_NC(Tile_X2Y5_to_NC),
    .from_ND(Tile_X2Y5_to_ND),
    .from_NF(Tile_X2Y5_to_NF),
    .from_NG(Tile_X2Y5_to_NG),
    .from_NH(Tile_X2Y5_to_NH),
    .from_NI(Tile_X2Y5_to_NI),
    .from_EA(Tile_X1Y4_to_EA),
    .from_EB(Tile_X1Y4_to_EB),
    .from_EC(Tile_X1Y4_to_EC),
    .from_ED(Tile_X1Y4_to_ED),
    .from_EF(Tile_X1Y4_to_EF),
    .from_EG(Tile_X1Y4_to_EG),
    .from_EH(Tile_X1Y4_to_EH),
    .from_EI(Tile_X1Y4_to_EI),
    .from_SA(Tile_X2Y3_to_SA),
    .from_SB(Tile_X2Y3_to_SB),
    .from_SC(Tile_X2Y3_to_SC),
    .from_SD(Tile_X2Y3_to_SD),
    .from_SF(Tile_X2Y3_to_SF),
    .from_SG(Tile_X2Y3_to_SG),
    .from_SH(Tile_X2Y3_to_SH),
    .from_SI(Tile_X2Y3_to_SI),
    .from_WA(Tile_X3Y4_to_WA),
    .from_WB(Tile_X3Y4_to_WB),
    .from_WC(Tile_X3Y4_to_WC),
    .from_WD(Tile_X3Y4_to_WD),
    .from_WF(Tile_X3Y4_to_WF),
    .from_WG(Tile_X3Y4_to_WG),
    .from_WH(Tile_X3Y4_to_WH),
    .from_WI(Tile_X3Y4_to_WI),
    .to_EA(Tile_X2Y4_to_EA),
    .to_EB(Tile_X2Y4_to_EB),
    .to_EC(Tile_X2Y4_to_EC),
    .to_ED(Tile_X2Y4_to_ED),
    .to_EF(Tile_X2Y4_to_EF),
    .to_EG(Tile_X2Y4_to_EG),
    .to_EH(Tile_X2Y4_to_EH),
    .to_EI(Tile_X2Y4_to_EI),
    .to_WA(Tile_X2Y4_to_WA),
    .to_WB(Tile_X2Y4_to_WB),
    .to_WC(Tile_X2Y4_to_WC),
    .to_WD(Tile_X2Y4_to_WD),
    .to_WF(Tile_X2Y4_to_WF),
    .to_WG(Tile_X2Y4_to_WG),
    .to_WH(Tile_X2Y4_to_WH),
    .to_WI(Tile_X2Y4_to_WI),
    .to_NA(Tile_X2Y4_to_NA),
    .to_NB(Tile_X2Y4_to_NB),
    .to_NC(Tile_X2Y4_to_NC),
    .to_ND(Tile_X2Y4_to_ND),
    .to_NF(Tile_X2Y4_to_NF),
    .to_NG(Tile_X2Y4_to_NG),
    .to_NH(Tile_X2Y4_to_NH),
    .to_NI(Tile_X2Y4_to_NI),
    .to_SA(Tile_X2Y4_to_SA),
    .to_SB(Tile_X2Y4_to_SB),
    .to_SC(Tile_X2Y4_to_SC),
    .to_SD(Tile_X2Y4_to_SD),
    .to_SF(Tile_X2Y4_to_SF),
    .to_SG(Tile_X2Y4_to_SG),
    .to_SH(Tile_X2Y4_to_SH),
    .to_SI(Tile_X2Y4_to_SI),
    .F_masked1(Tile_X2Y4_F_masked1),
    .F_masked2(Tile_X2Y4_F_masked2),
    .UserCLK(Tile_X2Y5_UserCLKo),
    .UserCLKo(Tile_X2Y4_UserCLKo),
    .rst(Tile_X2Y5_rsto),
    .rsto(Tile_X2Y4_rsto),
    .FrameData(Tile_X1Y4_FrameData_O),
    .FrameData_O(Tile_X2Y4_FrameData_O),
    .FrameStrobe(Tile_X2Y5_FrameStrobe_O),
    .FrameStrobe_O(Tile_X2Y4_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
nonlinear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X3Y4_Emulate_Bitstream)
    )
`endif
    Tile_X3Y4_nonlinear_LMDPL
    (
    .from_NA(Tile_X3Y5_to_NA),
    .from_NB(Tile_X3Y5_to_NB),
    .from_NC(Tile_X3Y5_to_NC),
    .from_ND(Tile_X3Y5_to_ND),
    .from_NF(Tile_X3Y5_to_NF),
    .from_NG(Tile_X3Y5_to_NG),
    .from_NH(Tile_X3Y5_to_NH),
    .from_NI(Tile_X3Y5_to_NI),
    .from_EA(Tile_X2Y4_to_EA),
    .from_EB(Tile_X2Y4_to_EB),
    .from_EC(Tile_X2Y4_to_EC),
    .from_ED(Tile_X2Y4_to_ED),
    .from_EF(Tile_X2Y4_to_EF),
    .from_EG(Tile_X2Y4_to_EG),
    .from_EH(Tile_X2Y4_to_EH),
    .from_EI(Tile_X2Y4_to_EI),
    .from_SA(Tile_X3Y3_to_SA),
    .from_SB(Tile_X3Y3_to_SB),
    .from_SC(Tile_X3Y3_to_SC),
    .from_SD(Tile_X3Y3_to_SD),
    .from_SF(Tile_X3Y3_to_SF),
    .from_SG(Tile_X3Y3_to_SG),
    .from_SH(Tile_X3Y3_to_SH),
    .from_SI(Tile_X3Y3_to_SI),
    .from_WA(Tile_X4Y4_to_WA),
    .from_WB(Tile_X4Y4_to_WB),
    .from_WC(Tile_X4Y4_to_WC),
    .from_WD(Tile_X4Y4_to_WD),
    .from_WF(Tile_X4Y4_to_WF),
    .from_WG(Tile_X4Y4_to_WG),
    .from_WH(Tile_X4Y4_to_WH),
    .from_WI(Tile_X4Y4_to_WI),
    .to_EA(Tile_X3Y4_to_EA),
    .to_EB(Tile_X3Y4_to_EB),
    .to_EC(Tile_X3Y4_to_EC),
    .to_ED(Tile_X3Y4_to_ED),
    .to_EF(Tile_X3Y4_to_EF),
    .to_EG(Tile_X3Y4_to_EG),
    .to_EH(Tile_X3Y4_to_EH),
    .to_EI(Tile_X3Y4_to_EI),
    .to_WA(Tile_X3Y4_to_WA),
    .to_WB(Tile_X3Y4_to_WB),
    .to_WC(Tile_X3Y4_to_WC),
    .to_WD(Tile_X3Y4_to_WD),
    .to_WF(Tile_X3Y4_to_WF),
    .to_WG(Tile_X3Y4_to_WG),
    .to_WH(Tile_X3Y4_to_WH),
    .to_WI(Tile_X3Y4_to_WI),
    .to_NA(Tile_X3Y4_to_NA),
    .to_NB(Tile_X3Y4_to_NB),
    .to_NC(Tile_X3Y4_to_NC),
    .to_ND(Tile_X3Y4_to_ND),
    .to_NF(Tile_X3Y4_to_NF),
    .to_NG(Tile_X3Y4_to_NG),
    .to_NH(Tile_X3Y4_to_NH),
    .to_NI(Tile_X3Y4_to_NI),
    .to_SA(Tile_X3Y4_to_SA),
    .to_SB(Tile_X3Y4_to_SB),
    .to_SC(Tile_X3Y4_to_SC),
    .to_SD(Tile_X3Y4_to_SD),
    .to_SF(Tile_X3Y4_to_SF),
    .to_SG(Tile_X3Y4_to_SG),
    .to_SH(Tile_X3Y4_to_SH),
    .to_SI(Tile_X3Y4_to_SI),
    .R_t(Tile_X3Y4_R_t),
    .R_f(Tile_X3Y4_R_f),
    .F_masked1(Tile_X3Y4_F_masked1),
    .F_masked2(Tile_X3Y4_F_masked2),
    .UserCLK(Tile_X3Y5_UserCLKo),
    .UserCLKo(Tile_X3Y4_UserCLKo),
    .rst(Tile_X3Y5_rsto),
    .rsto(Tile_X3Y4_rsto),
    .FrameData(Tile_X2Y4_FrameData_O),
    .FrameData_O(Tile_X3Y4_FrameData_O),
    .FrameStrobe(Tile_X3Y5_FrameStrobe_O),
    .FrameStrobe_O(Tile_X3Y4_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X4Y4_Emulate_Bitstream)
    )
`endif
    Tile_X4Y4_linear_LMDPL
    (
    .from_NA(Tile_X4Y5_to_NA),
    .from_NB(Tile_X4Y5_to_NB),
    .from_NC(Tile_X4Y5_to_NC),
    .from_ND(Tile_X4Y5_to_ND),
    .from_NF(Tile_X4Y5_to_NF),
    .from_NG(Tile_X4Y5_to_NG),
    .from_NH(Tile_X4Y5_to_NH),
    .from_NI(Tile_X4Y5_to_NI),
    .from_EA(Tile_X3Y4_to_EA),
    .from_EB(Tile_X3Y4_to_EB),
    .from_EC(Tile_X3Y4_to_EC),
    .from_ED(Tile_X3Y4_to_ED),
    .from_EF(Tile_X3Y4_to_EF),
    .from_EG(Tile_X3Y4_to_EG),
    .from_EH(Tile_X3Y4_to_EH),
    .from_EI(Tile_X3Y4_to_EI),
    .from_SA(Tile_X4Y3_to_SA),
    .from_SB(Tile_X4Y3_to_SB),
    .from_SC(Tile_X4Y3_to_SC),
    .from_SD(Tile_X4Y3_to_SD),
    .from_SF(Tile_X4Y3_to_SF),
    .from_SG(Tile_X4Y3_to_SG),
    .from_SH(Tile_X4Y3_to_SH),
    .from_SI(Tile_X4Y3_to_SI),
    .from_WA(Tile_X5Y4_to_WA),
    .from_WB(Tile_X5Y4_to_WB),
    .from_WC(Tile_X5Y4_to_WC),
    .from_WD(Tile_X5Y4_to_WD),
    .from_WF(Tile_X5Y4_to_WF),
    .from_WG(Tile_X5Y4_to_WG),
    .from_WH(Tile_X5Y4_to_WH),
    .from_WI(Tile_X5Y4_to_WI),
    .to_EA(Tile_X4Y4_to_EA),
    .to_EB(Tile_X4Y4_to_EB),
    .to_EC(Tile_X4Y4_to_EC),
    .to_ED(Tile_X4Y4_to_ED),
    .to_EF(Tile_X4Y4_to_EF),
    .to_EG(Tile_X4Y4_to_EG),
    .to_EH(Tile_X4Y4_to_EH),
    .to_EI(Tile_X4Y4_to_EI),
    .to_WA(Tile_X4Y4_to_WA),
    .to_WB(Tile_X4Y4_to_WB),
    .to_WC(Tile_X4Y4_to_WC),
    .to_WD(Tile_X4Y4_to_WD),
    .to_WF(Tile_X4Y4_to_WF),
    .to_WG(Tile_X4Y4_to_WG),
    .to_WH(Tile_X4Y4_to_WH),
    .to_WI(Tile_X4Y4_to_WI),
    .to_NA(Tile_X4Y4_to_NA),
    .to_NB(Tile_X4Y4_to_NB),
    .to_NC(Tile_X4Y4_to_NC),
    .to_ND(Tile_X4Y4_to_ND),
    .to_NF(Tile_X4Y4_to_NF),
    .to_NG(Tile_X4Y4_to_NG),
    .to_NH(Tile_X4Y4_to_NH),
    .to_NI(Tile_X4Y4_to_NI),
    .to_SA(Tile_X4Y4_to_SA),
    .to_SB(Tile_X4Y4_to_SB),
    .to_SC(Tile_X4Y4_to_SC),
    .to_SD(Tile_X4Y4_to_SD),
    .to_SF(Tile_X4Y4_to_SF),
    .to_SG(Tile_X4Y4_to_SG),
    .to_SH(Tile_X4Y4_to_SH),
    .to_SI(Tile_X4Y4_to_SI),
    .F_masked1(Tile_X4Y4_F_masked1),
    .F_masked2(Tile_X4Y4_F_masked2),
    .UserCLK(Tile_X4Y5_UserCLKo),
    .UserCLKo(Tile_X4Y4_UserCLKo),
    .rst(Tile_X4Y5_rsto),
    .rsto(Tile_X4Y4_rsto),
    .FrameData(Tile_X3Y4_FrameData_O),
    .FrameData_O(Tile_X4Y4_FrameData_O),
    .FrameStrobe(Tile_X4Y5_FrameStrobe_O),
    .FrameStrobe_O(Tile_X4Y4_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X5Y4_Emulate_Bitstream)
    )
`endif
    Tile_X5Y4_linear_LMDPL
    (
    .from_NA(Tile_X5Y5_to_NA),
    .from_NB(Tile_X5Y5_to_NB),
    .from_NC(Tile_X5Y5_to_NC),
    .from_ND(Tile_X5Y5_to_ND),
    .from_NF(Tile_X5Y5_to_NF),
    .from_NG(Tile_X5Y5_to_NG),
    .from_NH(Tile_X5Y5_to_NH),
    .from_NI(Tile_X5Y5_to_NI),
    .from_EA(Tile_X4Y4_to_EA),
    .from_EB(Tile_X4Y4_to_EB),
    .from_EC(Tile_X4Y4_to_EC),
    .from_ED(Tile_X4Y4_to_ED),
    .from_EF(Tile_X4Y4_to_EF),
    .from_EG(Tile_X4Y4_to_EG),
    .from_EH(Tile_X4Y4_to_EH),
    .from_EI(Tile_X4Y4_to_EI),
    .from_SA(Tile_X5Y3_to_SA),
    .from_SB(Tile_X5Y3_to_SB),
    .from_SC(Tile_X5Y3_to_SC),
    .from_SD(Tile_X5Y3_to_SD),
    .from_SF(Tile_X5Y3_to_SF),
    .from_SG(Tile_X5Y3_to_SG),
    .from_SH(Tile_X5Y3_to_SH),
    .from_SI(Tile_X5Y3_to_SI),
    .from_WA(Tile_X6Y4_to_WA),
    .from_WB(Tile_X6Y4_to_WB),
    .from_WC(Tile_X6Y4_to_WC),
    .from_WD(Tile_X6Y4_to_WD),
    .from_WF(Tile_X6Y4_to_WF),
    .from_WG(Tile_X6Y4_to_WG),
    .from_WH(Tile_X6Y4_to_WH),
    .from_WI(Tile_X6Y4_to_WI),
    .to_EA(Tile_X5Y4_to_EA),
    .to_EB(Tile_X5Y4_to_EB),
    .to_EC(Tile_X5Y4_to_EC),
    .to_ED(Tile_X5Y4_to_ED),
    .to_EF(Tile_X5Y4_to_EF),
    .to_EG(Tile_X5Y4_to_EG),
    .to_EH(Tile_X5Y4_to_EH),
    .to_EI(Tile_X5Y4_to_EI),
    .to_WA(Tile_X5Y4_to_WA),
    .to_WB(Tile_X5Y4_to_WB),
    .to_WC(Tile_X5Y4_to_WC),
    .to_WD(Tile_X5Y4_to_WD),
    .to_WF(Tile_X5Y4_to_WF),
    .to_WG(Tile_X5Y4_to_WG),
    .to_WH(Tile_X5Y4_to_WH),
    .to_WI(Tile_X5Y4_to_WI),
    .to_NA(Tile_X5Y4_to_NA),
    .to_NB(Tile_X5Y4_to_NB),
    .to_NC(Tile_X5Y4_to_NC),
    .to_ND(Tile_X5Y4_to_ND),
    .to_NF(Tile_X5Y4_to_NF),
    .to_NG(Tile_X5Y4_to_NG),
    .to_NH(Tile_X5Y4_to_NH),
    .to_NI(Tile_X5Y4_to_NI),
    .to_SA(Tile_X5Y4_to_SA),
    .to_SB(Tile_X5Y4_to_SB),
    .to_SC(Tile_X5Y4_to_SC),
    .to_SD(Tile_X5Y4_to_SD),
    .to_SF(Tile_X5Y4_to_SF),
    .to_SG(Tile_X5Y4_to_SG),
    .to_SH(Tile_X5Y4_to_SH),
    .to_SI(Tile_X5Y4_to_SI),
    .F_masked1(Tile_X5Y4_F_masked1),
    .F_masked2(Tile_X5Y4_F_masked2),
    .UserCLK(Tile_X5Y5_UserCLKo),
    .UserCLKo(Tile_X5Y4_UserCLKo),
    .rst(Tile_X5Y5_rsto),
    .rsto(Tile_X5Y4_rsto),
    .FrameData(Tile_X4Y4_FrameData_O),
    .FrameData_O(Tile_X5Y4_FrameData_O),
    .FrameStrobe(Tile_X5Y5_FrameStrobe_O),
    .FrameStrobe_O(Tile_X5Y4_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
nonlinear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X6Y4_Emulate_Bitstream)
    )
`endif
    Tile_X6Y4_nonlinear_LMDPL
    (
    .from_NA(Tile_X6Y5_to_NA),
    .from_NB(Tile_X6Y5_to_NB),
    .from_NC(Tile_X6Y5_to_NC),
    .from_ND(Tile_X6Y5_to_ND),
    .from_NF(Tile_X6Y5_to_NF),
    .from_NG(Tile_X6Y5_to_NG),
    .from_NH(Tile_X6Y5_to_NH),
    .from_NI(Tile_X6Y5_to_NI),
    .from_EA(Tile_X5Y4_to_EA),
    .from_EB(Tile_X5Y4_to_EB),
    .from_EC(Tile_X5Y4_to_EC),
    .from_ED(Tile_X5Y4_to_ED),
    .from_EF(Tile_X5Y4_to_EF),
    .from_EG(Tile_X5Y4_to_EG),
    .from_EH(Tile_X5Y4_to_EH),
    .from_EI(Tile_X5Y4_to_EI),
    .from_SA(Tile_X6Y3_to_SA),
    .from_SB(Tile_X6Y3_to_SB),
    .from_SC(Tile_X6Y3_to_SC),
    .from_SD(Tile_X6Y3_to_SD),
    .from_SF(Tile_X6Y3_to_SF),
    .from_SG(Tile_X6Y3_to_SG),
    .from_SH(Tile_X6Y3_to_SH),
    .from_SI(Tile_X6Y3_to_SI),
    .from_WA(Tile_X7Y4_to_WA),
    .from_WB(Tile_X7Y4_to_WB),
    .from_WC(Tile_X7Y4_to_WC),
    .from_WD(Tile_X7Y4_to_WD),
    .from_WF(Tile_X7Y4_to_WF),
    .from_WG(Tile_X7Y4_to_WG),
    .from_WH(Tile_X7Y4_to_WH),
    .from_WI(Tile_X7Y4_to_WI),
    .to_EA(Tile_X6Y4_to_EA),
    .to_EB(Tile_X6Y4_to_EB),
    .to_EC(Tile_X6Y4_to_EC),
    .to_ED(Tile_X6Y4_to_ED),
    .to_EF(Tile_X6Y4_to_EF),
    .to_EG(Tile_X6Y4_to_EG),
    .to_EH(Tile_X6Y4_to_EH),
    .to_EI(Tile_X6Y4_to_EI),
    .to_WA(Tile_X6Y4_to_WA),
    .to_WB(Tile_X6Y4_to_WB),
    .to_WC(Tile_X6Y4_to_WC),
    .to_WD(Tile_X6Y4_to_WD),
    .to_WF(Tile_X6Y4_to_WF),
    .to_WG(Tile_X6Y4_to_WG),
    .to_WH(Tile_X6Y4_to_WH),
    .to_WI(Tile_X6Y4_to_WI),
    .to_NA(Tile_X6Y4_to_NA),
    .to_NB(Tile_X6Y4_to_NB),
    .to_NC(Tile_X6Y4_to_NC),
    .to_ND(Tile_X6Y4_to_ND),
    .to_NF(Tile_X6Y4_to_NF),
    .to_NG(Tile_X6Y4_to_NG),
    .to_NH(Tile_X6Y4_to_NH),
    .to_NI(Tile_X6Y4_to_NI),
    .to_SA(Tile_X6Y4_to_SA),
    .to_SB(Tile_X6Y4_to_SB),
    .to_SC(Tile_X6Y4_to_SC),
    .to_SD(Tile_X6Y4_to_SD),
    .to_SF(Tile_X6Y4_to_SF),
    .to_SG(Tile_X6Y4_to_SG),
    .to_SH(Tile_X6Y4_to_SH),
    .to_SI(Tile_X6Y4_to_SI),
    .R_t(Tile_X6Y4_R_t),
    .R_f(Tile_X6Y4_R_f),
    .F_masked1(Tile_X6Y4_F_masked1),
    .F_masked2(Tile_X6Y4_F_masked2),
    .UserCLK(Tile_X6Y5_UserCLKo),
    .UserCLKo(Tile_X6Y4_UserCLKo),
    .rst(Tile_X6Y5_rsto),
    .rsto(Tile_X6Y4_rsto),
    .FrameData(Tile_X5Y4_FrameData_O),
    .FrameData_O(Tile_X6Y4_FrameData_O),
    .FrameStrobe(Tile_X6Y5_FrameStrobe_O),
    .FrameStrobe_O(Tile_X6Y4_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X7Y4_Emulate_Bitstream)
    )
`endif
    Tile_X7Y4_linear_LMDPL
    (
    .from_NA(Tile_X7Y5_to_NA),
    .from_NB(Tile_X7Y5_to_NB),
    .from_NC(Tile_X7Y5_to_NC),
    .from_ND(Tile_X7Y5_to_ND),
    .from_NF(Tile_X7Y5_to_NF),
    .from_NG(Tile_X7Y5_to_NG),
    .from_NH(Tile_X7Y5_to_NH),
    .from_NI(Tile_X7Y5_to_NI),
    .from_EA(Tile_X6Y4_to_EA),
    .from_EB(Tile_X6Y4_to_EB),
    .from_EC(Tile_X6Y4_to_EC),
    .from_ED(Tile_X6Y4_to_ED),
    .from_EF(Tile_X6Y4_to_EF),
    .from_EG(Tile_X6Y4_to_EG),
    .from_EH(Tile_X6Y4_to_EH),
    .from_EI(Tile_X6Y4_to_EI),
    .from_SA(Tile_X7Y3_to_SA),
    .from_SB(Tile_X7Y3_to_SB),
    .from_SC(Tile_X7Y3_to_SC),
    .from_SD(Tile_X7Y3_to_SD),
    .from_SF(Tile_X7Y3_to_SF),
    .from_SG(Tile_X7Y3_to_SG),
    .from_SH(Tile_X7Y3_to_SH),
    .from_SI(Tile_X7Y3_to_SI),
    .from_WA(Tile_X8Y4_to_WA),
    .from_WB(Tile_X8Y4_to_WB),
    .from_WC(Tile_X8Y4_to_WC),
    .from_WD(Tile_X8Y4_to_WD),
    .from_WF(Tile_X8Y4_to_WF),
    .from_WG(Tile_X8Y4_to_WG),
    .from_WH(Tile_X8Y4_to_WH),
    .from_WI(Tile_X8Y4_to_WI),
    .to_EA(Tile_X7Y4_to_EA),
    .to_EB(Tile_X7Y4_to_EB),
    .to_EC(Tile_X7Y4_to_EC),
    .to_ED(Tile_X7Y4_to_ED),
    .to_EF(Tile_X7Y4_to_EF),
    .to_EG(Tile_X7Y4_to_EG),
    .to_EH(Tile_X7Y4_to_EH),
    .to_EI(Tile_X7Y4_to_EI),
    .to_WA(Tile_X7Y4_to_WA),
    .to_WB(Tile_X7Y4_to_WB),
    .to_WC(Tile_X7Y4_to_WC),
    .to_WD(Tile_X7Y4_to_WD),
    .to_WF(Tile_X7Y4_to_WF),
    .to_WG(Tile_X7Y4_to_WG),
    .to_WH(Tile_X7Y4_to_WH),
    .to_WI(Tile_X7Y4_to_WI),
    .to_NA(Tile_X7Y4_to_NA),
    .to_NB(Tile_X7Y4_to_NB),
    .to_NC(Tile_X7Y4_to_NC),
    .to_ND(Tile_X7Y4_to_ND),
    .to_NF(Tile_X7Y4_to_NF),
    .to_NG(Tile_X7Y4_to_NG),
    .to_NH(Tile_X7Y4_to_NH),
    .to_NI(Tile_X7Y4_to_NI),
    .to_SA(Tile_X7Y4_to_SA),
    .to_SB(Tile_X7Y4_to_SB),
    .to_SC(Tile_X7Y4_to_SC),
    .to_SD(Tile_X7Y4_to_SD),
    .to_SF(Tile_X7Y4_to_SF),
    .to_SG(Tile_X7Y4_to_SG),
    .to_SH(Tile_X7Y4_to_SH),
    .to_SI(Tile_X7Y4_to_SI),
    .F_masked1(Tile_X7Y4_F_masked1),
    .F_masked2(Tile_X7Y4_F_masked2),
    .UserCLK(Tile_X7Y5_UserCLKo),
    .UserCLKo(Tile_X7Y4_UserCLKo),
    .rst(Tile_X7Y5_rsto),
    .rsto(Tile_X7Y4_rsto),
    .FrameData(Tile_X6Y4_FrameData_O),
    .FrameData_O(Tile_X7Y4_FrameData_O),
    .FrameStrobe(Tile_X7Y5_FrameStrobe_O),
    .FrameStrobe_O(Tile_X7Y4_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
ctrl_to_sec
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X8Y4_Emulate_Bitstream)
    )
`endif
    Tile_X8Y4_ctrl_to_sec
    (
    .from_NA(Tile_X8Y5_to_NA),
    .from_NB(Tile_X8Y5_to_NB),
    .from_NC(Tile_X8Y5_to_NC),
    .from_ND(Tile_X8Y5_to_ND),
    .from_NF(Tile_X8Y5_to_NF),
    .from_NG(Tile_X8Y5_to_NG),
    .from_NH(Tile_X8Y5_to_NH),
    .from_NI(Tile_X8Y5_to_NI),
    .from_EA(Tile_X7Y4_to_EA),
    .from_EB(Tile_X7Y4_to_EB),
    .from_EC(Tile_X7Y4_to_EC),
    .from_ED(Tile_X7Y4_to_ED),
    .from_EF(Tile_X7Y4_to_EF),
    .from_EG(Tile_X7Y4_to_EG),
    .from_EH(Tile_X7Y4_to_EH),
    .from_EI(Tile_X7Y4_to_EI),
    .from_SA(Tile_X8Y3_to_SA),
    .from_SB(Tile_X8Y3_to_SB),
    .from_SC(Tile_X8Y3_to_SC),
    .from_SD(Tile_X8Y3_to_SD),
    .from_SF(Tile_X8Y3_to_SF),
    .from_SG(Tile_X8Y3_to_SG),
    .from_SH(Tile_X8Y3_to_SH),
    .from_SI(Tile_X8Y3_to_SI),
    .from_WA_1s(Tile_X9Y4_to_WA_1s),
    .from_WB_1s(Tile_X9Y4_to_WB_1s),
    .from_WC_1s(Tile_X9Y4_to_WC_1s),
    .from_WD_1s(Tile_X9Y4_to_WD_1s),
    .from_WF_1s(Tile_X9Y4_to_WF_1s),
    .from_WG_1s(Tile_X9Y4_to_WG_1s),
    .from_WH_1s(Tile_X9Y4_to_WH_1s),
    .from_WI_1s(Tile_X9Y4_to_WI_1s),
    .to_WA(Tile_X8Y4_to_WA),
    .to_WB(Tile_X8Y4_to_WB),
    .to_WC(Tile_X8Y4_to_WC),
    .to_WD(Tile_X8Y4_to_WD),
    .to_WF(Tile_X8Y4_to_WF),
    .to_WG(Tile_X8Y4_to_WG),
    .to_WH(Tile_X8Y4_to_WH),
    .to_WI(Tile_X8Y4_to_WI),
    .to_NA(Tile_X8Y4_to_NA),
    .to_NB(Tile_X8Y4_to_NB),
    .to_NC(Tile_X8Y4_to_NC),
    .to_ND(Tile_X8Y4_to_ND),
    .to_NF(Tile_X8Y4_to_NF),
    .to_NG(Tile_X8Y4_to_NG),
    .to_NH(Tile_X8Y4_to_NH),
    .to_NI(Tile_X8Y4_to_NI),
    .to_SA(Tile_X8Y4_to_SA),
    .to_SB(Tile_X8Y4_to_SB),
    .to_SC(Tile_X8Y4_to_SC),
    .to_SD(Tile_X8Y4_to_SD),
    .to_SF(Tile_X8Y4_to_SF),
    .to_SG(Tile_X8Y4_to_SG),
    .to_SH(Tile_X8Y4_to_SH),
    .to_SI(Tile_X8Y4_to_SI),
    .UserCLK(Tile_X8Y5_UserCLKo),
    .UserCLKo(Tile_X8Y4_UserCLKo),
    .rst(Tile_X8Y5_rsto),
    .rsto(Tile_X8Y4_rsto),
    .FrameData(Tile_X7Y4_FrameData_O),
    .FrameData_O(Tile_X8Y4_FrameData_O),
    .FrameStrobe(Tile_X8Y5_FrameStrobe_O),
    .FrameStrobe_O(Tile_X8Y4_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
combined_WDDL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X9Y4_Emulate_Bitstream)
    )
`endif
    Tile_X9Y4_combined_WDDL
    (
    .from_NA_1s(Tile_X9Y5_to_NA_1s),
    .from_NB_1s(Tile_X9Y5_to_NB_1s),
    .from_NC_1s(Tile_X9Y5_to_NC_1s),
    .from_ND_1s(Tile_X9Y5_to_ND_1s),
    .from_NF_1s(Tile_X9Y5_to_NF_1s),
    .from_NG_1s(Tile_X9Y5_to_NG_1s),
    .from_NH_1s(Tile_X9Y5_to_NH_1s),
    .from_NI_1s(Tile_X9Y5_to_NI_1s),
    .from_SA_1s(Tile_X9Y3_to_SA_1s),
    .from_SB_1s(Tile_X9Y3_to_SB_1s),
    .from_SC_1s(Tile_X9Y3_to_SC_1s),
    .from_SD_1s(Tile_X9Y3_to_SD_1s),
    .from_SF_1s(Tile_X9Y3_to_SF_1s),
    .from_SG_1s(Tile_X9Y3_to_SG_1s),
    .from_SH_1s(Tile_X9Y3_to_SH_1s),
    .from_SI_1s(Tile_X9Y3_to_SI_1s),
    .from_WA_1s(Tile_X10Y4_to_WA_1s),
    .from_WB_1s(Tile_X10Y4_to_WB_1s),
    .from_WC_1s(Tile_X10Y4_to_WC_1s),
    .from_WD_1s(Tile_X10Y4_to_WD_1s),
    .from_WF_1s(Tile_X10Y4_to_WF_1s),
    .from_WG_1s(Tile_X10Y4_to_WG_1s),
    .from_WH_1s(Tile_X10Y4_to_WH_1s),
    .from_WI_1s(Tile_X10Y4_to_WI_1s),
    .to_EA_1s(Tile_X9Y4_to_EA_1s),
    .to_EB_1s(Tile_X9Y4_to_EB_1s),
    .to_EC_1s(Tile_X9Y4_to_EC_1s),
    .to_ED_1s(Tile_X9Y4_to_ED_1s),
    .to_EF_1s(Tile_X9Y4_to_EF_1s),
    .to_EG_1s(Tile_X9Y4_to_EG_1s),
    .to_EH_1s(Tile_X9Y4_to_EH_1s),
    .to_EI_1s(Tile_X9Y4_to_EI_1s),
    .to_WA_1s(Tile_X9Y4_to_WA_1s),
    .to_WB_1s(Tile_X9Y4_to_WB_1s),
    .to_WC_1s(Tile_X9Y4_to_WC_1s),
    .to_WD_1s(Tile_X9Y4_to_WD_1s),
    .to_WF_1s(Tile_X9Y4_to_WF_1s),
    .to_WG_1s(Tile_X9Y4_to_WG_1s),
    .to_WH_1s(Tile_X9Y4_to_WH_1s),
    .to_WI_1s(Tile_X9Y4_to_WI_1s),
    .to_NA_1s(Tile_X9Y4_to_NA_1s),
    .to_NB_1s(Tile_X9Y4_to_NB_1s),
    .to_NC_1s(Tile_X9Y4_to_NC_1s),
    .to_ND_1s(Tile_X9Y4_to_ND_1s),
    .to_NF_1s(Tile_X9Y4_to_NF_1s),
    .to_NG_1s(Tile_X9Y4_to_NG_1s),
    .to_NH_1s(Tile_X9Y4_to_NH_1s),
    .to_NI_1s(Tile_X9Y4_to_NI_1s),
    .to_SA_1s(Tile_X9Y4_to_SA_1s),
    .to_SB_1s(Tile_X9Y4_to_SB_1s),
    .to_SC_1s(Tile_X9Y4_to_SC_1s),
    .to_SD_1s(Tile_X9Y4_to_SD_1s),
    .to_SF_1s(Tile_X9Y4_to_SF_1s),
    .to_SG_1s(Tile_X9Y4_to_SG_1s),
    .to_SH_1s(Tile_X9Y4_to_SH_1s),
    .to_SI_1s(Tile_X9Y4_to_SI_1s),
    .F_ctrl(Tile_X9Y4_F_ctrl),
    .UserCLK(Tile_X9Y5_UserCLKo),
    .UserCLKo(Tile_X9Y4_UserCLKo),
    .rst(Tile_X9Y5_rsto),
    .rsto(Tile_X9Y4_rsto),
    .FrameData(Tile_X8Y4_FrameData_O),
    .FrameData_O(Tile_X9Y4_FrameData_O),
    .FrameStrobe(Tile_X9Y5_FrameStrobe_O),
    .FrameStrobe_O(Tile_X9Y4_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
ctrl_IO
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X10Y4_Emulate_Bitstream)
    )
`endif
    Tile_X10Y4_ctrl_IO
    (
    .from_EA_1s(Tile_X9Y4_to_EA_1s),
    .from_EB_1s(Tile_X9Y4_to_EB_1s),
    .from_EC_1s(Tile_X9Y4_to_EC_1s),
    .from_ED_1s(Tile_X9Y4_to_ED_1s),
    .from_EF_1s(Tile_X9Y4_to_EF_1s),
    .from_EG_1s(Tile_X9Y4_to_EG_1s),
    .from_EH_1s(Tile_X9Y4_to_EH_1s),
    .from_EI_1s(Tile_X9Y4_to_EI_1s),
    .to_WA_1s(Tile_X10Y4_to_WA_1s),
    .to_WB_1s(Tile_X10Y4_to_WB_1s),
    .to_WC_1s(Tile_X10Y4_to_WC_1s),
    .to_WD_1s(Tile_X10Y4_to_WD_1s),
    .to_WF_1s(Tile_X10Y4_to_WF_1s),
    .to_WG_1s(Tile_X10Y4_to_WG_1s),
    .to_WH_1s(Tile_X10Y4_to_WH_1s),
    .to_WI_1s(Tile_X10Y4_to_WI_1s),
    .A_O_top_0_t(Tile_X10Y4_A_O_top_0_t),
    .A_O_top_0_f(Tile_X10Y4_A_O_top_0_f),
    .A_prech2(Tile_X10Y4_A_prech2),
    .A_DR_fault(Tile_X10Y4_A_DR_fault),
    .A_I_top_0_t(Tile_X10Y4_A_I_top_0_t),
    .A_I_top_0_f(Tile_X10Y4_A_I_top_0_f),
    .A_T_top(Tile_X10Y4_A_T_top),
    .A_F_ctrl(Tile_X10Y4_A_F_ctrl),
    .UserCLK(Tile_X10Y5_UserCLKo),
    .UserCLKo(Tile_X10Y4_UserCLKo),
    .rst(Tile_X10Y5_rsto),
    .rsto(Tile_X10Y4_rsto),
    .FrameData(Tile_X9Y4_FrameData_O),
    .FrameData_O(Tile_X10Y4_FrameData_O),
    .FrameStrobe(Tile_X10Y5_FrameStrobe_O),
    .FrameStrobe_O(Tile_X10Y4_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
W_IO_custom
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X0Y5_Emulate_Bitstream)
    )
`endif
    Tile_X0Y5_W_IO_custom
    (
    .from_NA(Tile_X0Y6_to_NA),
    .from_NB(Tile_X0Y6_to_NB),
    .from_NC(Tile_X0Y6_to_NC),
    .from_ND(Tile_X0Y6_to_ND),
    .from_NF(Tile_X0Y6_to_NF),
    .from_NG(Tile_X0Y6_to_NG),
    .from_NH(Tile_X0Y6_to_NH),
    .from_NI(Tile_X0Y6_to_NI),
    .from_SA(Tile_X0Y4_to_SA),
    .from_SB(Tile_X0Y4_to_SB),
    .from_SC(Tile_X0Y4_to_SC),
    .from_SD(Tile_X0Y4_to_SD),
    .from_SF(Tile_X0Y4_to_SF),
    .from_SG(Tile_X0Y4_to_SG),
    .from_SH(Tile_X0Y4_to_SH),
    .from_SI(Tile_X0Y4_to_SI),
    .from_WA(Tile_X1Y5_to_WA),
    .from_WB(Tile_X1Y5_to_WB),
    .from_WC(Tile_X1Y5_to_WC),
    .from_WD(Tile_X1Y5_to_WD),
    .from_WF(Tile_X1Y5_to_WF),
    .from_WG(Tile_X1Y5_to_WG),
    .from_WH(Tile_X1Y5_to_WH),
    .from_WI(Tile_X1Y5_to_WI),
    .to_EA(Tile_X0Y5_to_EA),
    .to_EB(Tile_X0Y5_to_EB),
    .to_EC(Tile_X0Y5_to_EC),
    .to_ED(Tile_X0Y5_to_ED),
    .to_EF(Tile_X0Y5_to_EF),
    .to_EG(Tile_X0Y5_to_EG),
    .to_EH(Tile_X0Y5_to_EH),
    .to_EI(Tile_X0Y5_to_EI),
    .to_NA(Tile_X0Y5_to_NA),
    .to_NB(Tile_X0Y5_to_NB),
    .to_NC(Tile_X0Y5_to_NC),
    .to_ND(Tile_X0Y5_to_ND),
    .to_NF(Tile_X0Y5_to_NF),
    .to_NG(Tile_X0Y5_to_NG),
    .to_NH(Tile_X0Y5_to_NH),
    .to_NI(Tile_X0Y5_to_NI),
    .to_SA(Tile_X0Y5_to_SA),
    .to_SB(Tile_X0Y5_to_SB),
    .to_SC(Tile_X0Y5_to_SC),
    .to_SD(Tile_X0Y5_to_SD),
    .to_SF(Tile_X0Y5_to_SF),
    .to_SG(Tile_X0Y5_to_SG),
    .to_SH(Tile_X0Y5_to_SH),
    .to_SI(Tile_X0Y5_to_SI),
    .A_O_top_0_t(Tile_X0Y5_A_O_top_0_t),
    .A_O_top_0_f(Tile_X0Y5_A_O_top_0_f),
    .A_O_top_1_t(Tile_X0Y5_A_O_top_1_t),
    .A_O_top_1_f(Tile_X0Y5_A_O_top_1_f),
    .A_prech1(Tile_X0Y5_A_prech1),
    .A_prech2(Tile_X0Y5_A_prech2),
    .A_DR_fault(Tile_X0Y5_A_DR_fault),
    .A_I_top_0_t(Tile_X0Y5_A_I_top_0_t),
    .A_I_top_0_f(Tile_X0Y5_A_I_top_0_f),
    .A_I_top_1_t(Tile_X0Y5_A_I_top_1_t),
    .A_I_top_1_f(Tile_X0Y5_A_I_top_1_f),
    .A_T_top(Tile_X0Y5_A_T_top),
    .A_F_masked1(Tile_X0Y5_A_F_masked1),
    .A_F_masked2(Tile_X0Y5_A_F_masked2),
    .A_config_C_bit0(Tile_X0Y5_A_config_C_bit0),
    .A_config_C_bit1(Tile_X0Y5_A_config_C_bit1),
    .A_config_C_bit2(Tile_X0Y5_A_config_C_bit2),
    .A_config_C_bit3(Tile_X0Y5_A_config_C_bit3),
    .B_config_C_bit0(Tile_X0Y5_B_config_C_bit0),
    .B_config_C_bit1(Tile_X0Y5_B_config_C_bit1),
    .B_config_C_bit2(Tile_X0Y5_B_config_C_bit2),
    .B_config_C_bit3(Tile_X0Y5_B_config_C_bit3),
    .UserCLK(Tile_X0Y6_UserCLKo),
    .UserCLKo(Tile_X0Y5_UserCLKo),
    .rst(Tile_X0Y6_rsto),
    .rsto(Tile_X0Y5_rsto),
    .FrameData(Tile_Y5_FrameData),
    .FrameData_O(Tile_X0Y5_FrameData_O),
    .FrameStrobe(Tile_X0Y6_FrameStrobe_O),
    .FrameStrobe_O(Tile_X0Y5_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X1Y5_Emulate_Bitstream)
    )
`endif
    Tile_X1Y5_linear_LMDPL
    (
    .from_NA(Tile_X1Y6_to_NA),
    .from_NB(Tile_X1Y6_to_NB),
    .from_NC(Tile_X1Y6_to_NC),
    .from_ND(Tile_X1Y6_to_ND),
    .from_NF(Tile_X1Y6_to_NF),
    .from_NG(Tile_X1Y6_to_NG),
    .from_NH(Tile_X1Y6_to_NH),
    .from_NI(Tile_X1Y6_to_NI),
    .from_EA(Tile_X0Y5_to_EA),
    .from_EB(Tile_X0Y5_to_EB),
    .from_EC(Tile_X0Y5_to_EC),
    .from_ED(Tile_X0Y5_to_ED),
    .from_EF(Tile_X0Y5_to_EF),
    .from_EG(Tile_X0Y5_to_EG),
    .from_EH(Tile_X0Y5_to_EH),
    .from_EI(Tile_X0Y5_to_EI),
    .from_SA(Tile_X1Y4_to_SA),
    .from_SB(Tile_X1Y4_to_SB),
    .from_SC(Tile_X1Y4_to_SC),
    .from_SD(Tile_X1Y4_to_SD),
    .from_SF(Tile_X1Y4_to_SF),
    .from_SG(Tile_X1Y4_to_SG),
    .from_SH(Tile_X1Y4_to_SH),
    .from_SI(Tile_X1Y4_to_SI),
    .from_WA(Tile_X2Y5_to_WA),
    .from_WB(Tile_X2Y5_to_WB),
    .from_WC(Tile_X2Y5_to_WC),
    .from_WD(Tile_X2Y5_to_WD),
    .from_WF(Tile_X2Y5_to_WF),
    .from_WG(Tile_X2Y5_to_WG),
    .from_WH(Tile_X2Y5_to_WH),
    .from_WI(Tile_X2Y5_to_WI),
    .to_EA(Tile_X1Y5_to_EA),
    .to_EB(Tile_X1Y5_to_EB),
    .to_EC(Tile_X1Y5_to_EC),
    .to_ED(Tile_X1Y5_to_ED),
    .to_EF(Tile_X1Y5_to_EF),
    .to_EG(Tile_X1Y5_to_EG),
    .to_EH(Tile_X1Y5_to_EH),
    .to_EI(Tile_X1Y5_to_EI),
    .to_WA(Tile_X1Y5_to_WA),
    .to_WB(Tile_X1Y5_to_WB),
    .to_WC(Tile_X1Y5_to_WC),
    .to_WD(Tile_X1Y5_to_WD),
    .to_WF(Tile_X1Y5_to_WF),
    .to_WG(Tile_X1Y5_to_WG),
    .to_WH(Tile_X1Y5_to_WH),
    .to_WI(Tile_X1Y5_to_WI),
    .to_NA(Tile_X1Y5_to_NA),
    .to_NB(Tile_X1Y5_to_NB),
    .to_NC(Tile_X1Y5_to_NC),
    .to_ND(Tile_X1Y5_to_ND),
    .to_NF(Tile_X1Y5_to_NF),
    .to_NG(Tile_X1Y5_to_NG),
    .to_NH(Tile_X1Y5_to_NH),
    .to_NI(Tile_X1Y5_to_NI),
    .to_SA(Tile_X1Y5_to_SA),
    .to_SB(Tile_X1Y5_to_SB),
    .to_SC(Tile_X1Y5_to_SC),
    .to_SD(Tile_X1Y5_to_SD),
    .to_SF(Tile_X1Y5_to_SF),
    .to_SG(Tile_X1Y5_to_SG),
    .to_SH(Tile_X1Y5_to_SH),
    .to_SI(Tile_X1Y5_to_SI),
    .F_masked1(Tile_X1Y5_F_masked1),
    .F_masked2(Tile_X1Y5_F_masked2),
    .UserCLK(Tile_X1Y6_UserCLKo),
    .UserCLKo(Tile_X1Y5_UserCLKo),
    .rst(Tile_X1Y6_rsto),
    .rsto(Tile_X1Y5_rsto),
    .FrameData(Tile_X0Y5_FrameData_O),
    .FrameData_O(Tile_X1Y5_FrameData_O),
    .FrameStrobe(Tile_X1Y6_FrameStrobe_O),
    .FrameStrobe_O(Tile_X1Y5_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X2Y5_Emulate_Bitstream)
    )
`endif
    Tile_X2Y5_linear_LMDPL
    (
    .from_NA(Tile_X2Y6_to_NA),
    .from_NB(Tile_X2Y6_to_NB),
    .from_NC(Tile_X2Y6_to_NC),
    .from_ND(Tile_X2Y6_to_ND),
    .from_NF(Tile_X2Y6_to_NF),
    .from_NG(Tile_X2Y6_to_NG),
    .from_NH(Tile_X2Y6_to_NH),
    .from_NI(Tile_X2Y6_to_NI),
    .from_EA(Tile_X1Y5_to_EA),
    .from_EB(Tile_X1Y5_to_EB),
    .from_EC(Tile_X1Y5_to_EC),
    .from_ED(Tile_X1Y5_to_ED),
    .from_EF(Tile_X1Y5_to_EF),
    .from_EG(Tile_X1Y5_to_EG),
    .from_EH(Tile_X1Y5_to_EH),
    .from_EI(Tile_X1Y5_to_EI),
    .from_SA(Tile_X2Y4_to_SA),
    .from_SB(Tile_X2Y4_to_SB),
    .from_SC(Tile_X2Y4_to_SC),
    .from_SD(Tile_X2Y4_to_SD),
    .from_SF(Tile_X2Y4_to_SF),
    .from_SG(Tile_X2Y4_to_SG),
    .from_SH(Tile_X2Y4_to_SH),
    .from_SI(Tile_X2Y4_to_SI),
    .from_WA(Tile_X3Y5_to_WA),
    .from_WB(Tile_X3Y5_to_WB),
    .from_WC(Tile_X3Y5_to_WC),
    .from_WD(Tile_X3Y5_to_WD),
    .from_WF(Tile_X3Y5_to_WF),
    .from_WG(Tile_X3Y5_to_WG),
    .from_WH(Tile_X3Y5_to_WH),
    .from_WI(Tile_X3Y5_to_WI),
    .to_EA(Tile_X2Y5_to_EA),
    .to_EB(Tile_X2Y5_to_EB),
    .to_EC(Tile_X2Y5_to_EC),
    .to_ED(Tile_X2Y5_to_ED),
    .to_EF(Tile_X2Y5_to_EF),
    .to_EG(Tile_X2Y5_to_EG),
    .to_EH(Tile_X2Y5_to_EH),
    .to_EI(Tile_X2Y5_to_EI),
    .to_WA(Tile_X2Y5_to_WA),
    .to_WB(Tile_X2Y5_to_WB),
    .to_WC(Tile_X2Y5_to_WC),
    .to_WD(Tile_X2Y5_to_WD),
    .to_WF(Tile_X2Y5_to_WF),
    .to_WG(Tile_X2Y5_to_WG),
    .to_WH(Tile_X2Y5_to_WH),
    .to_WI(Tile_X2Y5_to_WI),
    .to_NA(Tile_X2Y5_to_NA),
    .to_NB(Tile_X2Y5_to_NB),
    .to_NC(Tile_X2Y5_to_NC),
    .to_ND(Tile_X2Y5_to_ND),
    .to_NF(Tile_X2Y5_to_NF),
    .to_NG(Tile_X2Y5_to_NG),
    .to_NH(Tile_X2Y5_to_NH),
    .to_NI(Tile_X2Y5_to_NI),
    .to_SA(Tile_X2Y5_to_SA),
    .to_SB(Tile_X2Y5_to_SB),
    .to_SC(Tile_X2Y5_to_SC),
    .to_SD(Tile_X2Y5_to_SD),
    .to_SF(Tile_X2Y5_to_SF),
    .to_SG(Tile_X2Y5_to_SG),
    .to_SH(Tile_X2Y5_to_SH),
    .to_SI(Tile_X2Y5_to_SI),
    .F_masked1(Tile_X2Y5_F_masked1),
    .F_masked2(Tile_X2Y5_F_masked2),
    .UserCLK(Tile_X2Y6_UserCLKo),
    .UserCLKo(Tile_X2Y5_UserCLKo),
    .rst(Tile_X2Y6_rsto),
    .rsto(Tile_X2Y5_rsto),
    .FrameData(Tile_X1Y5_FrameData_O),
    .FrameData_O(Tile_X2Y5_FrameData_O),
    .FrameStrobe(Tile_X2Y6_FrameStrobe_O),
    .FrameStrobe_O(Tile_X2Y5_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
nonlinear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X3Y5_Emulate_Bitstream)
    )
`endif
    Tile_X3Y5_nonlinear_LMDPL
    (
    .from_NA(Tile_X3Y6_to_NA),
    .from_NB(Tile_X3Y6_to_NB),
    .from_NC(Tile_X3Y6_to_NC),
    .from_ND(Tile_X3Y6_to_ND),
    .from_NF(Tile_X3Y6_to_NF),
    .from_NG(Tile_X3Y6_to_NG),
    .from_NH(Tile_X3Y6_to_NH),
    .from_NI(Tile_X3Y6_to_NI),
    .from_EA(Tile_X2Y5_to_EA),
    .from_EB(Tile_X2Y5_to_EB),
    .from_EC(Tile_X2Y5_to_EC),
    .from_ED(Tile_X2Y5_to_ED),
    .from_EF(Tile_X2Y5_to_EF),
    .from_EG(Tile_X2Y5_to_EG),
    .from_EH(Tile_X2Y5_to_EH),
    .from_EI(Tile_X2Y5_to_EI),
    .from_SA(Tile_X3Y4_to_SA),
    .from_SB(Tile_X3Y4_to_SB),
    .from_SC(Tile_X3Y4_to_SC),
    .from_SD(Tile_X3Y4_to_SD),
    .from_SF(Tile_X3Y4_to_SF),
    .from_SG(Tile_X3Y4_to_SG),
    .from_SH(Tile_X3Y4_to_SH),
    .from_SI(Tile_X3Y4_to_SI),
    .from_WA(Tile_X4Y5_to_WA),
    .from_WB(Tile_X4Y5_to_WB),
    .from_WC(Tile_X4Y5_to_WC),
    .from_WD(Tile_X4Y5_to_WD),
    .from_WF(Tile_X4Y5_to_WF),
    .from_WG(Tile_X4Y5_to_WG),
    .from_WH(Tile_X4Y5_to_WH),
    .from_WI(Tile_X4Y5_to_WI),
    .to_EA(Tile_X3Y5_to_EA),
    .to_EB(Tile_X3Y5_to_EB),
    .to_EC(Tile_X3Y5_to_EC),
    .to_ED(Tile_X3Y5_to_ED),
    .to_EF(Tile_X3Y5_to_EF),
    .to_EG(Tile_X3Y5_to_EG),
    .to_EH(Tile_X3Y5_to_EH),
    .to_EI(Tile_X3Y5_to_EI),
    .to_WA(Tile_X3Y5_to_WA),
    .to_WB(Tile_X3Y5_to_WB),
    .to_WC(Tile_X3Y5_to_WC),
    .to_WD(Tile_X3Y5_to_WD),
    .to_WF(Tile_X3Y5_to_WF),
    .to_WG(Tile_X3Y5_to_WG),
    .to_WH(Tile_X3Y5_to_WH),
    .to_WI(Tile_X3Y5_to_WI),
    .to_NA(Tile_X3Y5_to_NA),
    .to_NB(Tile_X3Y5_to_NB),
    .to_NC(Tile_X3Y5_to_NC),
    .to_ND(Tile_X3Y5_to_ND),
    .to_NF(Tile_X3Y5_to_NF),
    .to_NG(Tile_X3Y5_to_NG),
    .to_NH(Tile_X3Y5_to_NH),
    .to_NI(Tile_X3Y5_to_NI),
    .to_SA(Tile_X3Y5_to_SA),
    .to_SB(Tile_X3Y5_to_SB),
    .to_SC(Tile_X3Y5_to_SC),
    .to_SD(Tile_X3Y5_to_SD),
    .to_SF(Tile_X3Y5_to_SF),
    .to_SG(Tile_X3Y5_to_SG),
    .to_SH(Tile_X3Y5_to_SH),
    .to_SI(Tile_X3Y5_to_SI),
    .R_t(Tile_X3Y5_R_t),
    .R_f(Tile_X3Y5_R_f),
    .F_masked1(Tile_X3Y5_F_masked1),
    .F_masked2(Tile_X3Y5_F_masked2),
    .UserCLK(Tile_X3Y6_UserCLKo),
    .UserCLKo(Tile_X3Y5_UserCLKo),
    .rst(Tile_X3Y6_rsto),
    .rsto(Tile_X3Y5_rsto),
    .FrameData(Tile_X2Y5_FrameData_O),
    .FrameData_O(Tile_X3Y5_FrameData_O),
    .FrameStrobe(Tile_X3Y6_FrameStrobe_O),
    .FrameStrobe_O(Tile_X3Y5_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X4Y5_Emulate_Bitstream)
    )
`endif
    Tile_X4Y5_linear_LMDPL
    (
    .from_NA(Tile_X4Y6_to_NA),
    .from_NB(Tile_X4Y6_to_NB),
    .from_NC(Tile_X4Y6_to_NC),
    .from_ND(Tile_X4Y6_to_ND),
    .from_NF(Tile_X4Y6_to_NF),
    .from_NG(Tile_X4Y6_to_NG),
    .from_NH(Tile_X4Y6_to_NH),
    .from_NI(Tile_X4Y6_to_NI),
    .from_EA(Tile_X3Y5_to_EA),
    .from_EB(Tile_X3Y5_to_EB),
    .from_EC(Tile_X3Y5_to_EC),
    .from_ED(Tile_X3Y5_to_ED),
    .from_EF(Tile_X3Y5_to_EF),
    .from_EG(Tile_X3Y5_to_EG),
    .from_EH(Tile_X3Y5_to_EH),
    .from_EI(Tile_X3Y5_to_EI),
    .from_SA(Tile_X4Y4_to_SA),
    .from_SB(Tile_X4Y4_to_SB),
    .from_SC(Tile_X4Y4_to_SC),
    .from_SD(Tile_X4Y4_to_SD),
    .from_SF(Tile_X4Y4_to_SF),
    .from_SG(Tile_X4Y4_to_SG),
    .from_SH(Tile_X4Y4_to_SH),
    .from_SI(Tile_X4Y4_to_SI),
    .from_WA(Tile_X5Y5_to_WA),
    .from_WB(Tile_X5Y5_to_WB),
    .from_WC(Tile_X5Y5_to_WC),
    .from_WD(Tile_X5Y5_to_WD),
    .from_WF(Tile_X5Y5_to_WF),
    .from_WG(Tile_X5Y5_to_WG),
    .from_WH(Tile_X5Y5_to_WH),
    .from_WI(Tile_X5Y5_to_WI),
    .to_EA(Tile_X4Y5_to_EA),
    .to_EB(Tile_X4Y5_to_EB),
    .to_EC(Tile_X4Y5_to_EC),
    .to_ED(Tile_X4Y5_to_ED),
    .to_EF(Tile_X4Y5_to_EF),
    .to_EG(Tile_X4Y5_to_EG),
    .to_EH(Tile_X4Y5_to_EH),
    .to_EI(Tile_X4Y5_to_EI),
    .to_WA(Tile_X4Y5_to_WA),
    .to_WB(Tile_X4Y5_to_WB),
    .to_WC(Tile_X4Y5_to_WC),
    .to_WD(Tile_X4Y5_to_WD),
    .to_WF(Tile_X4Y5_to_WF),
    .to_WG(Tile_X4Y5_to_WG),
    .to_WH(Tile_X4Y5_to_WH),
    .to_WI(Tile_X4Y5_to_WI),
    .to_NA(Tile_X4Y5_to_NA),
    .to_NB(Tile_X4Y5_to_NB),
    .to_NC(Tile_X4Y5_to_NC),
    .to_ND(Tile_X4Y5_to_ND),
    .to_NF(Tile_X4Y5_to_NF),
    .to_NG(Tile_X4Y5_to_NG),
    .to_NH(Tile_X4Y5_to_NH),
    .to_NI(Tile_X4Y5_to_NI),
    .to_SA(Tile_X4Y5_to_SA),
    .to_SB(Tile_X4Y5_to_SB),
    .to_SC(Tile_X4Y5_to_SC),
    .to_SD(Tile_X4Y5_to_SD),
    .to_SF(Tile_X4Y5_to_SF),
    .to_SG(Tile_X4Y5_to_SG),
    .to_SH(Tile_X4Y5_to_SH),
    .to_SI(Tile_X4Y5_to_SI),
    .F_masked1(Tile_X4Y5_F_masked1),
    .F_masked2(Tile_X4Y5_F_masked2),
    .UserCLK(Tile_X4Y6_UserCLKo),
    .UserCLKo(Tile_X4Y5_UserCLKo),
    .rst(Tile_X4Y6_rsto),
    .rsto(Tile_X4Y5_rsto),
    .FrameData(Tile_X3Y5_FrameData_O),
    .FrameData_O(Tile_X4Y5_FrameData_O),
    .FrameStrobe(Tile_X4Y6_FrameStrobe_O),
    .FrameStrobe_O(Tile_X4Y5_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X5Y5_Emulate_Bitstream)
    )
`endif
    Tile_X5Y5_linear_LMDPL
    (
    .from_NA(Tile_X5Y6_to_NA),
    .from_NB(Tile_X5Y6_to_NB),
    .from_NC(Tile_X5Y6_to_NC),
    .from_ND(Tile_X5Y6_to_ND),
    .from_NF(Tile_X5Y6_to_NF),
    .from_NG(Tile_X5Y6_to_NG),
    .from_NH(Tile_X5Y6_to_NH),
    .from_NI(Tile_X5Y6_to_NI),
    .from_EA(Tile_X4Y5_to_EA),
    .from_EB(Tile_X4Y5_to_EB),
    .from_EC(Tile_X4Y5_to_EC),
    .from_ED(Tile_X4Y5_to_ED),
    .from_EF(Tile_X4Y5_to_EF),
    .from_EG(Tile_X4Y5_to_EG),
    .from_EH(Tile_X4Y5_to_EH),
    .from_EI(Tile_X4Y5_to_EI),
    .from_SA(Tile_X5Y4_to_SA),
    .from_SB(Tile_X5Y4_to_SB),
    .from_SC(Tile_X5Y4_to_SC),
    .from_SD(Tile_X5Y4_to_SD),
    .from_SF(Tile_X5Y4_to_SF),
    .from_SG(Tile_X5Y4_to_SG),
    .from_SH(Tile_X5Y4_to_SH),
    .from_SI(Tile_X5Y4_to_SI),
    .from_WA(Tile_X6Y5_to_WA),
    .from_WB(Tile_X6Y5_to_WB),
    .from_WC(Tile_X6Y5_to_WC),
    .from_WD(Tile_X6Y5_to_WD),
    .from_WF(Tile_X6Y5_to_WF),
    .from_WG(Tile_X6Y5_to_WG),
    .from_WH(Tile_X6Y5_to_WH),
    .from_WI(Tile_X6Y5_to_WI),
    .to_EA(Tile_X5Y5_to_EA),
    .to_EB(Tile_X5Y5_to_EB),
    .to_EC(Tile_X5Y5_to_EC),
    .to_ED(Tile_X5Y5_to_ED),
    .to_EF(Tile_X5Y5_to_EF),
    .to_EG(Tile_X5Y5_to_EG),
    .to_EH(Tile_X5Y5_to_EH),
    .to_EI(Tile_X5Y5_to_EI),
    .to_WA(Tile_X5Y5_to_WA),
    .to_WB(Tile_X5Y5_to_WB),
    .to_WC(Tile_X5Y5_to_WC),
    .to_WD(Tile_X5Y5_to_WD),
    .to_WF(Tile_X5Y5_to_WF),
    .to_WG(Tile_X5Y5_to_WG),
    .to_WH(Tile_X5Y5_to_WH),
    .to_WI(Tile_X5Y5_to_WI),
    .to_NA(Tile_X5Y5_to_NA),
    .to_NB(Tile_X5Y5_to_NB),
    .to_NC(Tile_X5Y5_to_NC),
    .to_ND(Tile_X5Y5_to_ND),
    .to_NF(Tile_X5Y5_to_NF),
    .to_NG(Tile_X5Y5_to_NG),
    .to_NH(Tile_X5Y5_to_NH),
    .to_NI(Tile_X5Y5_to_NI),
    .to_SA(Tile_X5Y5_to_SA),
    .to_SB(Tile_X5Y5_to_SB),
    .to_SC(Tile_X5Y5_to_SC),
    .to_SD(Tile_X5Y5_to_SD),
    .to_SF(Tile_X5Y5_to_SF),
    .to_SG(Tile_X5Y5_to_SG),
    .to_SH(Tile_X5Y5_to_SH),
    .to_SI(Tile_X5Y5_to_SI),
    .F_masked1(Tile_X5Y5_F_masked1),
    .F_masked2(Tile_X5Y5_F_masked2),
    .UserCLK(Tile_X5Y6_UserCLKo),
    .UserCLKo(Tile_X5Y5_UserCLKo),
    .rst(Tile_X5Y6_rsto),
    .rsto(Tile_X5Y5_rsto),
    .FrameData(Tile_X4Y5_FrameData_O),
    .FrameData_O(Tile_X5Y5_FrameData_O),
    .FrameStrobe(Tile_X5Y6_FrameStrobe_O),
    .FrameStrobe_O(Tile_X5Y5_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
nonlinear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X6Y5_Emulate_Bitstream)
    )
`endif
    Tile_X6Y5_nonlinear_LMDPL
    (
    .from_NA(Tile_X6Y6_to_NA),
    .from_NB(Tile_X6Y6_to_NB),
    .from_NC(Tile_X6Y6_to_NC),
    .from_ND(Tile_X6Y6_to_ND),
    .from_NF(Tile_X6Y6_to_NF),
    .from_NG(Tile_X6Y6_to_NG),
    .from_NH(Tile_X6Y6_to_NH),
    .from_NI(Tile_X6Y6_to_NI),
    .from_EA(Tile_X5Y5_to_EA),
    .from_EB(Tile_X5Y5_to_EB),
    .from_EC(Tile_X5Y5_to_EC),
    .from_ED(Tile_X5Y5_to_ED),
    .from_EF(Tile_X5Y5_to_EF),
    .from_EG(Tile_X5Y5_to_EG),
    .from_EH(Tile_X5Y5_to_EH),
    .from_EI(Tile_X5Y5_to_EI),
    .from_SA(Tile_X6Y4_to_SA),
    .from_SB(Tile_X6Y4_to_SB),
    .from_SC(Tile_X6Y4_to_SC),
    .from_SD(Tile_X6Y4_to_SD),
    .from_SF(Tile_X6Y4_to_SF),
    .from_SG(Tile_X6Y4_to_SG),
    .from_SH(Tile_X6Y4_to_SH),
    .from_SI(Tile_X6Y4_to_SI),
    .from_WA(Tile_X7Y5_to_WA),
    .from_WB(Tile_X7Y5_to_WB),
    .from_WC(Tile_X7Y5_to_WC),
    .from_WD(Tile_X7Y5_to_WD),
    .from_WF(Tile_X7Y5_to_WF),
    .from_WG(Tile_X7Y5_to_WG),
    .from_WH(Tile_X7Y5_to_WH),
    .from_WI(Tile_X7Y5_to_WI),
    .to_EA(Tile_X6Y5_to_EA),
    .to_EB(Tile_X6Y5_to_EB),
    .to_EC(Tile_X6Y5_to_EC),
    .to_ED(Tile_X6Y5_to_ED),
    .to_EF(Tile_X6Y5_to_EF),
    .to_EG(Tile_X6Y5_to_EG),
    .to_EH(Tile_X6Y5_to_EH),
    .to_EI(Tile_X6Y5_to_EI),
    .to_WA(Tile_X6Y5_to_WA),
    .to_WB(Tile_X6Y5_to_WB),
    .to_WC(Tile_X6Y5_to_WC),
    .to_WD(Tile_X6Y5_to_WD),
    .to_WF(Tile_X6Y5_to_WF),
    .to_WG(Tile_X6Y5_to_WG),
    .to_WH(Tile_X6Y5_to_WH),
    .to_WI(Tile_X6Y5_to_WI),
    .to_NA(Tile_X6Y5_to_NA),
    .to_NB(Tile_X6Y5_to_NB),
    .to_NC(Tile_X6Y5_to_NC),
    .to_ND(Tile_X6Y5_to_ND),
    .to_NF(Tile_X6Y5_to_NF),
    .to_NG(Tile_X6Y5_to_NG),
    .to_NH(Tile_X6Y5_to_NH),
    .to_NI(Tile_X6Y5_to_NI),
    .to_SA(Tile_X6Y5_to_SA),
    .to_SB(Tile_X6Y5_to_SB),
    .to_SC(Tile_X6Y5_to_SC),
    .to_SD(Tile_X6Y5_to_SD),
    .to_SF(Tile_X6Y5_to_SF),
    .to_SG(Tile_X6Y5_to_SG),
    .to_SH(Tile_X6Y5_to_SH),
    .to_SI(Tile_X6Y5_to_SI),
    .R_t(Tile_X6Y5_R_t),
    .R_f(Tile_X6Y5_R_f),
    .F_masked1(Tile_X6Y5_F_masked1),
    .F_masked2(Tile_X6Y5_F_masked2),
    .UserCLK(Tile_X6Y6_UserCLKo),
    .UserCLKo(Tile_X6Y5_UserCLKo),
    .rst(Tile_X6Y6_rsto),
    .rsto(Tile_X6Y5_rsto),
    .FrameData(Tile_X5Y5_FrameData_O),
    .FrameData_O(Tile_X6Y5_FrameData_O),
    .FrameStrobe(Tile_X6Y6_FrameStrobe_O),
    .FrameStrobe_O(Tile_X6Y5_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X7Y5_Emulate_Bitstream)
    )
`endif
    Tile_X7Y5_linear_LMDPL
    (
    .from_NA(Tile_X7Y6_to_NA),
    .from_NB(Tile_X7Y6_to_NB),
    .from_NC(Tile_X7Y6_to_NC),
    .from_ND(Tile_X7Y6_to_ND),
    .from_NF(Tile_X7Y6_to_NF),
    .from_NG(Tile_X7Y6_to_NG),
    .from_NH(Tile_X7Y6_to_NH),
    .from_NI(Tile_X7Y6_to_NI),
    .from_EA(Tile_X6Y5_to_EA),
    .from_EB(Tile_X6Y5_to_EB),
    .from_EC(Tile_X6Y5_to_EC),
    .from_ED(Tile_X6Y5_to_ED),
    .from_EF(Tile_X6Y5_to_EF),
    .from_EG(Tile_X6Y5_to_EG),
    .from_EH(Tile_X6Y5_to_EH),
    .from_EI(Tile_X6Y5_to_EI),
    .from_SA(Tile_X7Y4_to_SA),
    .from_SB(Tile_X7Y4_to_SB),
    .from_SC(Tile_X7Y4_to_SC),
    .from_SD(Tile_X7Y4_to_SD),
    .from_SF(Tile_X7Y4_to_SF),
    .from_SG(Tile_X7Y4_to_SG),
    .from_SH(Tile_X7Y4_to_SH),
    .from_SI(Tile_X7Y4_to_SI),
    .from_WA(Tile_X8Y5_to_WA),
    .from_WB(Tile_X8Y5_to_WB),
    .from_WC(Tile_X8Y5_to_WC),
    .from_WD(Tile_X8Y5_to_WD),
    .from_WF(Tile_X8Y5_to_WF),
    .from_WG(Tile_X8Y5_to_WG),
    .from_WH(Tile_X8Y5_to_WH),
    .from_WI(Tile_X8Y5_to_WI),
    .to_EA(Tile_X7Y5_to_EA),
    .to_EB(Tile_X7Y5_to_EB),
    .to_EC(Tile_X7Y5_to_EC),
    .to_ED(Tile_X7Y5_to_ED),
    .to_EF(Tile_X7Y5_to_EF),
    .to_EG(Tile_X7Y5_to_EG),
    .to_EH(Tile_X7Y5_to_EH),
    .to_EI(Tile_X7Y5_to_EI),
    .to_WA(Tile_X7Y5_to_WA),
    .to_WB(Tile_X7Y5_to_WB),
    .to_WC(Tile_X7Y5_to_WC),
    .to_WD(Tile_X7Y5_to_WD),
    .to_WF(Tile_X7Y5_to_WF),
    .to_WG(Tile_X7Y5_to_WG),
    .to_WH(Tile_X7Y5_to_WH),
    .to_WI(Tile_X7Y5_to_WI),
    .to_NA(Tile_X7Y5_to_NA),
    .to_NB(Tile_X7Y5_to_NB),
    .to_NC(Tile_X7Y5_to_NC),
    .to_ND(Tile_X7Y5_to_ND),
    .to_NF(Tile_X7Y5_to_NF),
    .to_NG(Tile_X7Y5_to_NG),
    .to_NH(Tile_X7Y5_to_NH),
    .to_NI(Tile_X7Y5_to_NI),
    .to_SA(Tile_X7Y5_to_SA),
    .to_SB(Tile_X7Y5_to_SB),
    .to_SC(Tile_X7Y5_to_SC),
    .to_SD(Tile_X7Y5_to_SD),
    .to_SF(Tile_X7Y5_to_SF),
    .to_SG(Tile_X7Y5_to_SG),
    .to_SH(Tile_X7Y5_to_SH),
    .to_SI(Tile_X7Y5_to_SI),
    .F_masked1(Tile_X7Y5_F_masked1),
    .F_masked2(Tile_X7Y5_F_masked2),
    .UserCLK(Tile_X7Y6_UserCLKo),
    .UserCLKo(Tile_X7Y5_UserCLKo),
    .rst(Tile_X7Y6_rsto),
    .rsto(Tile_X7Y5_rsto),
    .FrameData(Tile_X6Y5_FrameData_O),
    .FrameData_O(Tile_X7Y5_FrameData_O),
    .FrameStrobe(Tile_X7Y6_FrameStrobe_O),
    .FrameStrobe_O(Tile_X7Y5_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
ctrl_to_sec
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X8Y5_Emulate_Bitstream)
    )
`endif
    Tile_X8Y5_ctrl_to_sec
    (
    .from_NA(Tile_X8Y6_to_NA),
    .from_NB(Tile_X8Y6_to_NB),
    .from_NC(Tile_X8Y6_to_NC),
    .from_ND(Tile_X8Y6_to_ND),
    .from_NF(Tile_X8Y6_to_NF),
    .from_NG(Tile_X8Y6_to_NG),
    .from_NH(Tile_X8Y6_to_NH),
    .from_NI(Tile_X8Y6_to_NI),
    .from_EA(Tile_X7Y5_to_EA),
    .from_EB(Tile_X7Y5_to_EB),
    .from_EC(Tile_X7Y5_to_EC),
    .from_ED(Tile_X7Y5_to_ED),
    .from_EF(Tile_X7Y5_to_EF),
    .from_EG(Tile_X7Y5_to_EG),
    .from_EH(Tile_X7Y5_to_EH),
    .from_EI(Tile_X7Y5_to_EI),
    .from_SA(Tile_X8Y4_to_SA),
    .from_SB(Tile_X8Y4_to_SB),
    .from_SC(Tile_X8Y4_to_SC),
    .from_SD(Tile_X8Y4_to_SD),
    .from_SF(Tile_X8Y4_to_SF),
    .from_SG(Tile_X8Y4_to_SG),
    .from_SH(Tile_X8Y4_to_SH),
    .from_SI(Tile_X8Y4_to_SI),
    .from_WA_1s(Tile_X9Y5_to_WA_1s),
    .from_WB_1s(Tile_X9Y5_to_WB_1s),
    .from_WC_1s(Tile_X9Y5_to_WC_1s),
    .from_WD_1s(Tile_X9Y5_to_WD_1s),
    .from_WF_1s(Tile_X9Y5_to_WF_1s),
    .from_WG_1s(Tile_X9Y5_to_WG_1s),
    .from_WH_1s(Tile_X9Y5_to_WH_1s),
    .from_WI_1s(Tile_X9Y5_to_WI_1s),
    .to_WA(Tile_X8Y5_to_WA),
    .to_WB(Tile_X8Y5_to_WB),
    .to_WC(Tile_X8Y5_to_WC),
    .to_WD(Tile_X8Y5_to_WD),
    .to_WF(Tile_X8Y5_to_WF),
    .to_WG(Tile_X8Y5_to_WG),
    .to_WH(Tile_X8Y5_to_WH),
    .to_WI(Tile_X8Y5_to_WI),
    .to_NA(Tile_X8Y5_to_NA),
    .to_NB(Tile_X8Y5_to_NB),
    .to_NC(Tile_X8Y5_to_NC),
    .to_ND(Tile_X8Y5_to_ND),
    .to_NF(Tile_X8Y5_to_NF),
    .to_NG(Tile_X8Y5_to_NG),
    .to_NH(Tile_X8Y5_to_NH),
    .to_NI(Tile_X8Y5_to_NI),
    .to_SA(Tile_X8Y5_to_SA),
    .to_SB(Tile_X8Y5_to_SB),
    .to_SC(Tile_X8Y5_to_SC),
    .to_SD(Tile_X8Y5_to_SD),
    .to_SF(Tile_X8Y5_to_SF),
    .to_SG(Tile_X8Y5_to_SG),
    .to_SH(Tile_X8Y5_to_SH),
    .to_SI(Tile_X8Y5_to_SI),
    .UserCLK(Tile_X8Y6_UserCLKo),
    .UserCLKo(Tile_X8Y5_UserCLKo),
    .rst(Tile_X8Y6_rsto),
    .rsto(Tile_X8Y5_rsto),
    .FrameData(Tile_X7Y5_FrameData_O),
    .FrameData_O(Tile_X8Y5_FrameData_O),
    .FrameStrobe(Tile_X8Y6_FrameStrobe_O),
    .FrameStrobe_O(Tile_X8Y5_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
combined_WDDL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X9Y5_Emulate_Bitstream)
    )
`endif
    Tile_X9Y5_combined_WDDL
    (
    .from_NA_1s(Tile_X9Y6_to_NA_1s),
    .from_NB_1s(Tile_X9Y6_to_NB_1s),
    .from_NC_1s(Tile_X9Y6_to_NC_1s),
    .from_ND_1s(Tile_X9Y6_to_ND_1s),
    .from_NF_1s(Tile_X9Y6_to_NF_1s),
    .from_NG_1s(Tile_X9Y6_to_NG_1s),
    .from_NH_1s(Tile_X9Y6_to_NH_1s),
    .from_NI_1s(Tile_X9Y6_to_NI_1s),
    .from_SA_1s(Tile_X9Y4_to_SA_1s),
    .from_SB_1s(Tile_X9Y4_to_SB_1s),
    .from_SC_1s(Tile_X9Y4_to_SC_1s),
    .from_SD_1s(Tile_X9Y4_to_SD_1s),
    .from_SF_1s(Tile_X9Y4_to_SF_1s),
    .from_SG_1s(Tile_X9Y4_to_SG_1s),
    .from_SH_1s(Tile_X9Y4_to_SH_1s),
    .from_SI_1s(Tile_X9Y4_to_SI_1s),
    .from_WA_1s(Tile_X10Y5_to_WA_1s),
    .from_WB_1s(Tile_X10Y5_to_WB_1s),
    .from_WC_1s(Tile_X10Y5_to_WC_1s),
    .from_WD_1s(Tile_X10Y5_to_WD_1s),
    .from_WF_1s(Tile_X10Y5_to_WF_1s),
    .from_WG_1s(Tile_X10Y5_to_WG_1s),
    .from_WH_1s(Tile_X10Y5_to_WH_1s),
    .from_WI_1s(Tile_X10Y5_to_WI_1s),
    .to_EA_1s(Tile_X9Y5_to_EA_1s),
    .to_EB_1s(Tile_X9Y5_to_EB_1s),
    .to_EC_1s(Tile_X9Y5_to_EC_1s),
    .to_ED_1s(Tile_X9Y5_to_ED_1s),
    .to_EF_1s(Tile_X9Y5_to_EF_1s),
    .to_EG_1s(Tile_X9Y5_to_EG_1s),
    .to_EH_1s(Tile_X9Y5_to_EH_1s),
    .to_EI_1s(Tile_X9Y5_to_EI_1s),
    .to_WA_1s(Tile_X9Y5_to_WA_1s),
    .to_WB_1s(Tile_X9Y5_to_WB_1s),
    .to_WC_1s(Tile_X9Y5_to_WC_1s),
    .to_WD_1s(Tile_X9Y5_to_WD_1s),
    .to_WF_1s(Tile_X9Y5_to_WF_1s),
    .to_WG_1s(Tile_X9Y5_to_WG_1s),
    .to_WH_1s(Tile_X9Y5_to_WH_1s),
    .to_WI_1s(Tile_X9Y5_to_WI_1s),
    .to_NA_1s(Tile_X9Y5_to_NA_1s),
    .to_NB_1s(Tile_X9Y5_to_NB_1s),
    .to_NC_1s(Tile_X9Y5_to_NC_1s),
    .to_ND_1s(Tile_X9Y5_to_ND_1s),
    .to_NF_1s(Tile_X9Y5_to_NF_1s),
    .to_NG_1s(Tile_X9Y5_to_NG_1s),
    .to_NH_1s(Tile_X9Y5_to_NH_1s),
    .to_NI_1s(Tile_X9Y5_to_NI_1s),
    .to_SA_1s(Tile_X9Y5_to_SA_1s),
    .to_SB_1s(Tile_X9Y5_to_SB_1s),
    .to_SC_1s(Tile_X9Y5_to_SC_1s),
    .to_SD_1s(Tile_X9Y5_to_SD_1s),
    .to_SF_1s(Tile_X9Y5_to_SF_1s),
    .to_SG_1s(Tile_X9Y5_to_SG_1s),
    .to_SH_1s(Tile_X9Y5_to_SH_1s),
    .to_SI_1s(Tile_X9Y5_to_SI_1s),
    .F_ctrl(Tile_X9Y5_F_ctrl),
    .UserCLK(Tile_X9Y6_UserCLKo),
    .UserCLKo(Tile_X9Y5_UserCLKo),
    .rst(Tile_X9Y6_rsto),
    .rsto(Tile_X9Y5_rsto),
    .FrameData(Tile_X8Y5_FrameData_O),
    .FrameData_O(Tile_X9Y5_FrameData_O),
    .FrameStrobe(Tile_X9Y6_FrameStrobe_O),
    .FrameStrobe_O(Tile_X9Y5_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
ctrl_IO
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X10Y5_Emulate_Bitstream)
    )
`endif
    Tile_X10Y5_ctrl_IO
    (
    .from_EA_1s(Tile_X9Y5_to_EA_1s),
    .from_EB_1s(Tile_X9Y5_to_EB_1s),
    .from_EC_1s(Tile_X9Y5_to_EC_1s),
    .from_ED_1s(Tile_X9Y5_to_ED_1s),
    .from_EF_1s(Tile_X9Y5_to_EF_1s),
    .from_EG_1s(Tile_X9Y5_to_EG_1s),
    .from_EH_1s(Tile_X9Y5_to_EH_1s),
    .from_EI_1s(Tile_X9Y5_to_EI_1s),
    .to_WA_1s(Tile_X10Y5_to_WA_1s),
    .to_WB_1s(Tile_X10Y5_to_WB_1s),
    .to_WC_1s(Tile_X10Y5_to_WC_1s),
    .to_WD_1s(Tile_X10Y5_to_WD_1s),
    .to_WF_1s(Tile_X10Y5_to_WF_1s),
    .to_WG_1s(Tile_X10Y5_to_WG_1s),
    .to_WH_1s(Tile_X10Y5_to_WH_1s),
    .to_WI_1s(Tile_X10Y5_to_WI_1s),
    .A_O_top_0_t(Tile_X10Y5_A_O_top_0_t),
    .A_O_top_0_f(Tile_X10Y5_A_O_top_0_f),
    .A_prech2(Tile_X10Y5_A_prech2),
    .A_DR_fault(Tile_X10Y5_A_DR_fault),
    .A_I_top_0_t(Tile_X10Y5_A_I_top_0_t),
    .A_I_top_0_f(Tile_X10Y5_A_I_top_0_f),
    .A_T_top(Tile_X10Y5_A_T_top),
    .A_F_ctrl(Tile_X10Y5_A_F_ctrl),
    .UserCLK(Tile_X10Y6_UserCLKo),
    .UserCLKo(Tile_X10Y5_UserCLKo),
    .rst(Tile_X10Y6_rsto),
    .rsto(Tile_X10Y5_rsto),
    .FrameData(Tile_X9Y5_FrameData_O),
    .FrameData_O(Tile_X10Y5_FrameData_O),
    .FrameStrobe(Tile_X10Y6_FrameStrobe_O),
    .FrameStrobe_O(Tile_X10Y5_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
W_IO_custom
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X0Y6_Emulate_Bitstream)
    )
`endif
    Tile_X0Y6_W_IO_custom
    (
    .from_NA(Tile_X0Y7_to_NA),
    .from_NB(Tile_X0Y7_to_NB),
    .from_NC(Tile_X0Y7_to_NC),
    .from_ND(Tile_X0Y7_to_ND),
    .from_NF(Tile_X0Y7_to_NF),
    .from_NG(Tile_X0Y7_to_NG),
    .from_NH(Tile_X0Y7_to_NH),
    .from_NI(Tile_X0Y7_to_NI),
    .from_SA(Tile_X0Y5_to_SA),
    .from_SB(Tile_X0Y5_to_SB),
    .from_SC(Tile_X0Y5_to_SC),
    .from_SD(Tile_X0Y5_to_SD),
    .from_SF(Tile_X0Y5_to_SF),
    .from_SG(Tile_X0Y5_to_SG),
    .from_SH(Tile_X0Y5_to_SH),
    .from_SI(Tile_X0Y5_to_SI),
    .from_WA(Tile_X1Y6_to_WA),
    .from_WB(Tile_X1Y6_to_WB),
    .from_WC(Tile_X1Y6_to_WC),
    .from_WD(Tile_X1Y6_to_WD),
    .from_WF(Tile_X1Y6_to_WF),
    .from_WG(Tile_X1Y6_to_WG),
    .from_WH(Tile_X1Y6_to_WH),
    .from_WI(Tile_X1Y6_to_WI),
    .to_EA(Tile_X0Y6_to_EA),
    .to_EB(Tile_X0Y6_to_EB),
    .to_EC(Tile_X0Y6_to_EC),
    .to_ED(Tile_X0Y6_to_ED),
    .to_EF(Tile_X0Y6_to_EF),
    .to_EG(Tile_X0Y6_to_EG),
    .to_EH(Tile_X0Y6_to_EH),
    .to_EI(Tile_X0Y6_to_EI),
    .to_NA(Tile_X0Y6_to_NA),
    .to_NB(Tile_X0Y6_to_NB),
    .to_NC(Tile_X0Y6_to_NC),
    .to_ND(Tile_X0Y6_to_ND),
    .to_NF(Tile_X0Y6_to_NF),
    .to_NG(Tile_X0Y6_to_NG),
    .to_NH(Tile_X0Y6_to_NH),
    .to_NI(Tile_X0Y6_to_NI),
    .to_SA(Tile_X0Y6_to_SA),
    .to_SB(Tile_X0Y6_to_SB),
    .to_SC(Tile_X0Y6_to_SC),
    .to_SD(Tile_X0Y6_to_SD),
    .to_SF(Tile_X0Y6_to_SF),
    .to_SG(Tile_X0Y6_to_SG),
    .to_SH(Tile_X0Y6_to_SH),
    .to_SI(Tile_X0Y6_to_SI),
    .A_O_top_0_t(Tile_X0Y6_A_O_top_0_t),
    .A_O_top_0_f(Tile_X0Y6_A_O_top_0_f),
    .A_O_top_1_t(Tile_X0Y6_A_O_top_1_t),
    .A_O_top_1_f(Tile_X0Y6_A_O_top_1_f),
    .A_prech1(Tile_X0Y6_A_prech1),
    .A_prech2(Tile_X0Y6_A_prech2),
    .A_DR_fault(Tile_X0Y6_A_DR_fault),
    .A_I_top_0_t(Tile_X0Y6_A_I_top_0_t),
    .A_I_top_0_f(Tile_X0Y6_A_I_top_0_f),
    .A_I_top_1_t(Tile_X0Y6_A_I_top_1_t),
    .A_I_top_1_f(Tile_X0Y6_A_I_top_1_f),
    .A_T_top(Tile_X0Y6_A_T_top),
    .A_F_masked1(Tile_X0Y6_A_F_masked1),
    .A_F_masked2(Tile_X0Y6_A_F_masked2),
    .A_config_C_bit0(Tile_X0Y6_A_config_C_bit0),
    .A_config_C_bit1(Tile_X0Y6_A_config_C_bit1),
    .A_config_C_bit2(Tile_X0Y6_A_config_C_bit2),
    .A_config_C_bit3(Tile_X0Y6_A_config_C_bit3),
    .B_config_C_bit0(Tile_X0Y6_B_config_C_bit0),
    .B_config_C_bit1(Tile_X0Y6_B_config_C_bit1),
    .B_config_C_bit2(Tile_X0Y6_B_config_C_bit2),
    .B_config_C_bit3(Tile_X0Y6_B_config_C_bit3),
    .UserCLK(Tile_X0Y7_UserCLKo),
    .UserCLKo(Tile_X0Y6_UserCLKo),
    .rst(Tile_X0Y7_rsto),
    .rsto(Tile_X0Y6_rsto),
    .FrameData(Tile_Y6_FrameData),
    .FrameData_O(Tile_X0Y6_FrameData_O),
    .FrameStrobe(Tile_X0Y7_FrameStrobe_O),
    .FrameStrobe_O(Tile_X0Y6_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X1Y6_Emulate_Bitstream)
    )
`endif
    Tile_X1Y6_linear_LMDPL
    (
    .from_NA(Tile_X1Y7_to_NA),
    .from_NB(Tile_X1Y7_to_NB),
    .from_NC(Tile_X1Y7_to_NC),
    .from_ND(Tile_X1Y7_to_ND),
    .from_NF(Tile_X1Y7_to_NF),
    .from_NG(Tile_X1Y7_to_NG),
    .from_NH(Tile_X1Y7_to_NH),
    .from_NI(Tile_X1Y7_to_NI),
    .from_EA(Tile_X0Y6_to_EA),
    .from_EB(Tile_X0Y6_to_EB),
    .from_EC(Tile_X0Y6_to_EC),
    .from_ED(Tile_X0Y6_to_ED),
    .from_EF(Tile_X0Y6_to_EF),
    .from_EG(Tile_X0Y6_to_EG),
    .from_EH(Tile_X0Y6_to_EH),
    .from_EI(Tile_X0Y6_to_EI),
    .from_SA(Tile_X1Y5_to_SA),
    .from_SB(Tile_X1Y5_to_SB),
    .from_SC(Tile_X1Y5_to_SC),
    .from_SD(Tile_X1Y5_to_SD),
    .from_SF(Tile_X1Y5_to_SF),
    .from_SG(Tile_X1Y5_to_SG),
    .from_SH(Tile_X1Y5_to_SH),
    .from_SI(Tile_X1Y5_to_SI),
    .from_WA(Tile_X2Y6_to_WA),
    .from_WB(Tile_X2Y6_to_WB),
    .from_WC(Tile_X2Y6_to_WC),
    .from_WD(Tile_X2Y6_to_WD),
    .from_WF(Tile_X2Y6_to_WF),
    .from_WG(Tile_X2Y6_to_WG),
    .from_WH(Tile_X2Y6_to_WH),
    .from_WI(Tile_X2Y6_to_WI),
    .to_EA(Tile_X1Y6_to_EA),
    .to_EB(Tile_X1Y6_to_EB),
    .to_EC(Tile_X1Y6_to_EC),
    .to_ED(Tile_X1Y6_to_ED),
    .to_EF(Tile_X1Y6_to_EF),
    .to_EG(Tile_X1Y6_to_EG),
    .to_EH(Tile_X1Y6_to_EH),
    .to_EI(Tile_X1Y6_to_EI),
    .to_WA(Tile_X1Y6_to_WA),
    .to_WB(Tile_X1Y6_to_WB),
    .to_WC(Tile_X1Y6_to_WC),
    .to_WD(Tile_X1Y6_to_WD),
    .to_WF(Tile_X1Y6_to_WF),
    .to_WG(Tile_X1Y6_to_WG),
    .to_WH(Tile_X1Y6_to_WH),
    .to_WI(Tile_X1Y6_to_WI),
    .to_NA(Tile_X1Y6_to_NA),
    .to_NB(Tile_X1Y6_to_NB),
    .to_NC(Tile_X1Y6_to_NC),
    .to_ND(Tile_X1Y6_to_ND),
    .to_NF(Tile_X1Y6_to_NF),
    .to_NG(Tile_X1Y6_to_NG),
    .to_NH(Tile_X1Y6_to_NH),
    .to_NI(Tile_X1Y6_to_NI),
    .to_SA(Tile_X1Y6_to_SA),
    .to_SB(Tile_X1Y6_to_SB),
    .to_SC(Tile_X1Y6_to_SC),
    .to_SD(Tile_X1Y6_to_SD),
    .to_SF(Tile_X1Y6_to_SF),
    .to_SG(Tile_X1Y6_to_SG),
    .to_SH(Tile_X1Y6_to_SH),
    .to_SI(Tile_X1Y6_to_SI),
    .F_masked1(Tile_X1Y6_F_masked1),
    .F_masked2(Tile_X1Y6_F_masked2),
    .UserCLK(Tile_X1Y7_UserCLKo),
    .UserCLKo(Tile_X1Y6_UserCLKo),
    .rst(Tile_X1Y7_rsto),
    .rsto(Tile_X1Y6_rsto),
    .FrameData(Tile_X0Y6_FrameData_O),
    .FrameData_O(Tile_X1Y6_FrameData_O),
    .FrameStrobe(Tile_X1Y7_FrameStrobe_O),
    .FrameStrobe_O(Tile_X1Y6_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X2Y6_Emulate_Bitstream)
    )
`endif
    Tile_X2Y6_linear_LMDPL
    (
    .from_NA(Tile_X2Y7_to_NA),
    .from_NB(Tile_X2Y7_to_NB),
    .from_NC(Tile_X2Y7_to_NC),
    .from_ND(Tile_X2Y7_to_ND),
    .from_NF(Tile_X2Y7_to_NF),
    .from_NG(Tile_X2Y7_to_NG),
    .from_NH(Tile_X2Y7_to_NH),
    .from_NI(Tile_X2Y7_to_NI),
    .from_EA(Tile_X1Y6_to_EA),
    .from_EB(Tile_X1Y6_to_EB),
    .from_EC(Tile_X1Y6_to_EC),
    .from_ED(Tile_X1Y6_to_ED),
    .from_EF(Tile_X1Y6_to_EF),
    .from_EG(Tile_X1Y6_to_EG),
    .from_EH(Tile_X1Y6_to_EH),
    .from_EI(Tile_X1Y6_to_EI),
    .from_SA(Tile_X2Y5_to_SA),
    .from_SB(Tile_X2Y5_to_SB),
    .from_SC(Tile_X2Y5_to_SC),
    .from_SD(Tile_X2Y5_to_SD),
    .from_SF(Tile_X2Y5_to_SF),
    .from_SG(Tile_X2Y5_to_SG),
    .from_SH(Tile_X2Y5_to_SH),
    .from_SI(Tile_X2Y5_to_SI),
    .from_WA(Tile_X3Y6_to_WA),
    .from_WB(Tile_X3Y6_to_WB),
    .from_WC(Tile_X3Y6_to_WC),
    .from_WD(Tile_X3Y6_to_WD),
    .from_WF(Tile_X3Y6_to_WF),
    .from_WG(Tile_X3Y6_to_WG),
    .from_WH(Tile_X3Y6_to_WH),
    .from_WI(Tile_X3Y6_to_WI),
    .to_EA(Tile_X2Y6_to_EA),
    .to_EB(Tile_X2Y6_to_EB),
    .to_EC(Tile_X2Y6_to_EC),
    .to_ED(Tile_X2Y6_to_ED),
    .to_EF(Tile_X2Y6_to_EF),
    .to_EG(Tile_X2Y6_to_EG),
    .to_EH(Tile_X2Y6_to_EH),
    .to_EI(Tile_X2Y6_to_EI),
    .to_WA(Tile_X2Y6_to_WA),
    .to_WB(Tile_X2Y6_to_WB),
    .to_WC(Tile_X2Y6_to_WC),
    .to_WD(Tile_X2Y6_to_WD),
    .to_WF(Tile_X2Y6_to_WF),
    .to_WG(Tile_X2Y6_to_WG),
    .to_WH(Tile_X2Y6_to_WH),
    .to_WI(Tile_X2Y6_to_WI),
    .to_NA(Tile_X2Y6_to_NA),
    .to_NB(Tile_X2Y6_to_NB),
    .to_NC(Tile_X2Y6_to_NC),
    .to_ND(Tile_X2Y6_to_ND),
    .to_NF(Tile_X2Y6_to_NF),
    .to_NG(Tile_X2Y6_to_NG),
    .to_NH(Tile_X2Y6_to_NH),
    .to_NI(Tile_X2Y6_to_NI),
    .to_SA(Tile_X2Y6_to_SA),
    .to_SB(Tile_X2Y6_to_SB),
    .to_SC(Tile_X2Y6_to_SC),
    .to_SD(Tile_X2Y6_to_SD),
    .to_SF(Tile_X2Y6_to_SF),
    .to_SG(Tile_X2Y6_to_SG),
    .to_SH(Tile_X2Y6_to_SH),
    .to_SI(Tile_X2Y6_to_SI),
    .F_masked1(Tile_X2Y6_F_masked1),
    .F_masked2(Tile_X2Y6_F_masked2),
    .UserCLK(Tile_X2Y7_UserCLKo),
    .UserCLKo(Tile_X2Y6_UserCLKo),
    .rst(Tile_X2Y7_rsto),
    .rsto(Tile_X2Y6_rsto),
    .FrameData(Tile_X1Y6_FrameData_O),
    .FrameData_O(Tile_X2Y6_FrameData_O),
    .FrameStrobe(Tile_X2Y7_FrameStrobe_O),
    .FrameStrobe_O(Tile_X2Y6_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
nonlinear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X3Y6_Emulate_Bitstream)
    )
`endif
    Tile_X3Y6_nonlinear_LMDPL
    (
    .from_NA(Tile_X3Y7_to_NA),
    .from_NB(Tile_X3Y7_to_NB),
    .from_NC(Tile_X3Y7_to_NC),
    .from_ND(Tile_X3Y7_to_ND),
    .from_NF(Tile_X3Y7_to_NF),
    .from_NG(Tile_X3Y7_to_NG),
    .from_NH(Tile_X3Y7_to_NH),
    .from_NI(Tile_X3Y7_to_NI),
    .from_EA(Tile_X2Y6_to_EA),
    .from_EB(Tile_X2Y6_to_EB),
    .from_EC(Tile_X2Y6_to_EC),
    .from_ED(Tile_X2Y6_to_ED),
    .from_EF(Tile_X2Y6_to_EF),
    .from_EG(Tile_X2Y6_to_EG),
    .from_EH(Tile_X2Y6_to_EH),
    .from_EI(Tile_X2Y6_to_EI),
    .from_SA(Tile_X3Y5_to_SA),
    .from_SB(Tile_X3Y5_to_SB),
    .from_SC(Tile_X3Y5_to_SC),
    .from_SD(Tile_X3Y5_to_SD),
    .from_SF(Tile_X3Y5_to_SF),
    .from_SG(Tile_X3Y5_to_SG),
    .from_SH(Tile_X3Y5_to_SH),
    .from_SI(Tile_X3Y5_to_SI),
    .from_WA(Tile_X4Y6_to_WA),
    .from_WB(Tile_X4Y6_to_WB),
    .from_WC(Tile_X4Y6_to_WC),
    .from_WD(Tile_X4Y6_to_WD),
    .from_WF(Tile_X4Y6_to_WF),
    .from_WG(Tile_X4Y6_to_WG),
    .from_WH(Tile_X4Y6_to_WH),
    .from_WI(Tile_X4Y6_to_WI),
    .to_EA(Tile_X3Y6_to_EA),
    .to_EB(Tile_X3Y6_to_EB),
    .to_EC(Tile_X3Y6_to_EC),
    .to_ED(Tile_X3Y6_to_ED),
    .to_EF(Tile_X3Y6_to_EF),
    .to_EG(Tile_X3Y6_to_EG),
    .to_EH(Tile_X3Y6_to_EH),
    .to_EI(Tile_X3Y6_to_EI),
    .to_WA(Tile_X3Y6_to_WA),
    .to_WB(Tile_X3Y6_to_WB),
    .to_WC(Tile_X3Y6_to_WC),
    .to_WD(Tile_X3Y6_to_WD),
    .to_WF(Tile_X3Y6_to_WF),
    .to_WG(Tile_X3Y6_to_WG),
    .to_WH(Tile_X3Y6_to_WH),
    .to_WI(Tile_X3Y6_to_WI),
    .to_NA(Tile_X3Y6_to_NA),
    .to_NB(Tile_X3Y6_to_NB),
    .to_NC(Tile_X3Y6_to_NC),
    .to_ND(Tile_X3Y6_to_ND),
    .to_NF(Tile_X3Y6_to_NF),
    .to_NG(Tile_X3Y6_to_NG),
    .to_NH(Tile_X3Y6_to_NH),
    .to_NI(Tile_X3Y6_to_NI),
    .to_SA(Tile_X3Y6_to_SA),
    .to_SB(Tile_X3Y6_to_SB),
    .to_SC(Tile_X3Y6_to_SC),
    .to_SD(Tile_X3Y6_to_SD),
    .to_SF(Tile_X3Y6_to_SF),
    .to_SG(Tile_X3Y6_to_SG),
    .to_SH(Tile_X3Y6_to_SH),
    .to_SI(Tile_X3Y6_to_SI),
    .R_t(Tile_X3Y6_R_t),
    .R_f(Tile_X3Y6_R_f),
    .F_masked1(Tile_X3Y6_F_masked1),
    .F_masked2(Tile_X3Y6_F_masked2),
    .UserCLK(Tile_X3Y7_UserCLKo),
    .UserCLKo(Tile_X3Y6_UserCLKo),
    .rst(Tile_X3Y7_rsto),
    .rsto(Tile_X3Y6_rsto),
    .FrameData(Tile_X2Y6_FrameData_O),
    .FrameData_O(Tile_X3Y6_FrameData_O),
    .FrameStrobe(Tile_X3Y7_FrameStrobe_O),
    .FrameStrobe_O(Tile_X3Y6_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X4Y6_Emulate_Bitstream)
    )
`endif
    Tile_X4Y6_linear_LMDPL
    (
    .from_NA(Tile_X4Y7_to_NA),
    .from_NB(Tile_X4Y7_to_NB),
    .from_NC(Tile_X4Y7_to_NC),
    .from_ND(Tile_X4Y7_to_ND),
    .from_NF(Tile_X4Y7_to_NF),
    .from_NG(Tile_X4Y7_to_NG),
    .from_NH(Tile_X4Y7_to_NH),
    .from_NI(Tile_X4Y7_to_NI),
    .from_EA(Tile_X3Y6_to_EA),
    .from_EB(Tile_X3Y6_to_EB),
    .from_EC(Tile_X3Y6_to_EC),
    .from_ED(Tile_X3Y6_to_ED),
    .from_EF(Tile_X3Y6_to_EF),
    .from_EG(Tile_X3Y6_to_EG),
    .from_EH(Tile_X3Y6_to_EH),
    .from_EI(Tile_X3Y6_to_EI),
    .from_SA(Tile_X4Y5_to_SA),
    .from_SB(Tile_X4Y5_to_SB),
    .from_SC(Tile_X4Y5_to_SC),
    .from_SD(Tile_X4Y5_to_SD),
    .from_SF(Tile_X4Y5_to_SF),
    .from_SG(Tile_X4Y5_to_SG),
    .from_SH(Tile_X4Y5_to_SH),
    .from_SI(Tile_X4Y5_to_SI),
    .from_WA(Tile_X5Y6_to_WA),
    .from_WB(Tile_X5Y6_to_WB),
    .from_WC(Tile_X5Y6_to_WC),
    .from_WD(Tile_X5Y6_to_WD),
    .from_WF(Tile_X5Y6_to_WF),
    .from_WG(Tile_X5Y6_to_WG),
    .from_WH(Tile_X5Y6_to_WH),
    .from_WI(Tile_X5Y6_to_WI),
    .to_EA(Tile_X4Y6_to_EA),
    .to_EB(Tile_X4Y6_to_EB),
    .to_EC(Tile_X4Y6_to_EC),
    .to_ED(Tile_X4Y6_to_ED),
    .to_EF(Tile_X4Y6_to_EF),
    .to_EG(Tile_X4Y6_to_EG),
    .to_EH(Tile_X4Y6_to_EH),
    .to_EI(Tile_X4Y6_to_EI),
    .to_WA(Tile_X4Y6_to_WA),
    .to_WB(Tile_X4Y6_to_WB),
    .to_WC(Tile_X4Y6_to_WC),
    .to_WD(Tile_X4Y6_to_WD),
    .to_WF(Tile_X4Y6_to_WF),
    .to_WG(Tile_X4Y6_to_WG),
    .to_WH(Tile_X4Y6_to_WH),
    .to_WI(Tile_X4Y6_to_WI),
    .to_NA(Tile_X4Y6_to_NA),
    .to_NB(Tile_X4Y6_to_NB),
    .to_NC(Tile_X4Y6_to_NC),
    .to_ND(Tile_X4Y6_to_ND),
    .to_NF(Tile_X4Y6_to_NF),
    .to_NG(Tile_X4Y6_to_NG),
    .to_NH(Tile_X4Y6_to_NH),
    .to_NI(Tile_X4Y6_to_NI),
    .to_SA(Tile_X4Y6_to_SA),
    .to_SB(Tile_X4Y6_to_SB),
    .to_SC(Tile_X4Y6_to_SC),
    .to_SD(Tile_X4Y6_to_SD),
    .to_SF(Tile_X4Y6_to_SF),
    .to_SG(Tile_X4Y6_to_SG),
    .to_SH(Tile_X4Y6_to_SH),
    .to_SI(Tile_X4Y6_to_SI),
    .F_masked1(Tile_X4Y6_F_masked1),
    .F_masked2(Tile_X4Y6_F_masked2),
    .UserCLK(Tile_X4Y7_UserCLKo),
    .UserCLKo(Tile_X4Y6_UserCLKo),
    .rst(Tile_X4Y7_rsto),
    .rsto(Tile_X4Y6_rsto),
    .FrameData(Tile_X3Y6_FrameData_O),
    .FrameData_O(Tile_X4Y6_FrameData_O),
    .FrameStrobe(Tile_X4Y7_FrameStrobe_O),
    .FrameStrobe_O(Tile_X4Y6_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X5Y6_Emulate_Bitstream)
    )
`endif
    Tile_X5Y6_linear_LMDPL
    (
    .from_NA(Tile_X5Y7_to_NA),
    .from_NB(Tile_X5Y7_to_NB),
    .from_NC(Tile_X5Y7_to_NC),
    .from_ND(Tile_X5Y7_to_ND),
    .from_NF(Tile_X5Y7_to_NF),
    .from_NG(Tile_X5Y7_to_NG),
    .from_NH(Tile_X5Y7_to_NH),
    .from_NI(Tile_X5Y7_to_NI),
    .from_EA(Tile_X4Y6_to_EA),
    .from_EB(Tile_X4Y6_to_EB),
    .from_EC(Tile_X4Y6_to_EC),
    .from_ED(Tile_X4Y6_to_ED),
    .from_EF(Tile_X4Y6_to_EF),
    .from_EG(Tile_X4Y6_to_EG),
    .from_EH(Tile_X4Y6_to_EH),
    .from_EI(Tile_X4Y6_to_EI),
    .from_SA(Tile_X5Y5_to_SA),
    .from_SB(Tile_X5Y5_to_SB),
    .from_SC(Tile_X5Y5_to_SC),
    .from_SD(Tile_X5Y5_to_SD),
    .from_SF(Tile_X5Y5_to_SF),
    .from_SG(Tile_X5Y5_to_SG),
    .from_SH(Tile_X5Y5_to_SH),
    .from_SI(Tile_X5Y5_to_SI),
    .from_WA(Tile_X6Y6_to_WA),
    .from_WB(Tile_X6Y6_to_WB),
    .from_WC(Tile_X6Y6_to_WC),
    .from_WD(Tile_X6Y6_to_WD),
    .from_WF(Tile_X6Y6_to_WF),
    .from_WG(Tile_X6Y6_to_WG),
    .from_WH(Tile_X6Y6_to_WH),
    .from_WI(Tile_X6Y6_to_WI),
    .to_EA(Tile_X5Y6_to_EA),
    .to_EB(Tile_X5Y6_to_EB),
    .to_EC(Tile_X5Y6_to_EC),
    .to_ED(Tile_X5Y6_to_ED),
    .to_EF(Tile_X5Y6_to_EF),
    .to_EG(Tile_X5Y6_to_EG),
    .to_EH(Tile_X5Y6_to_EH),
    .to_EI(Tile_X5Y6_to_EI),
    .to_WA(Tile_X5Y6_to_WA),
    .to_WB(Tile_X5Y6_to_WB),
    .to_WC(Tile_X5Y6_to_WC),
    .to_WD(Tile_X5Y6_to_WD),
    .to_WF(Tile_X5Y6_to_WF),
    .to_WG(Tile_X5Y6_to_WG),
    .to_WH(Tile_X5Y6_to_WH),
    .to_WI(Tile_X5Y6_to_WI),
    .to_NA(Tile_X5Y6_to_NA),
    .to_NB(Tile_X5Y6_to_NB),
    .to_NC(Tile_X5Y6_to_NC),
    .to_ND(Tile_X5Y6_to_ND),
    .to_NF(Tile_X5Y6_to_NF),
    .to_NG(Tile_X5Y6_to_NG),
    .to_NH(Tile_X5Y6_to_NH),
    .to_NI(Tile_X5Y6_to_NI),
    .to_SA(Tile_X5Y6_to_SA),
    .to_SB(Tile_X5Y6_to_SB),
    .to_SC(Tile_X5Y6_to_SC),
    .to_SD(Tile_X5Y6_to_SD),
    .to_SF(Tile_X5Y6_to_SF),
    .to_SG(Tile_X5Y6_to_SG),
    .to_SH(Tile_X5Y6_to_SH),
    .to_SI(Tile_X5Y6_to_SI),
    .F_masked1(Tile_X5Y6_F_masked1),
    .F_masked2(Tile_X5Y6_F_masked2),
    .UserCLK(Tile_X5Y7_UserCLKo),
    .UserCLKo(Tile_X5Y6_UserCLKo),
    .rst(Tile_X5Y7_rsto),
    .rsto(Tile_X5Y6_rsto),
    .FrameData(Tile_X4Y6_FrameData_O),
    .FrameData_O(Tile_X5Y6_FrameData_O),
    .FrameStrobe(Tile_X5Y7_FrameStrobe_O),
    .FrameStrobe_O(Tile_X5Y6_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
nonlinear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X6Y6_Emulate_Bitstream)
    )
`endif
    Tile_X6Y6_nonlinear_LMDPL
    (
    .from_NA(Tile_X6Y7_to_NA),
    .from_NB(Tile_X6Y7_to_NB),
    .from_NC(Tile_X6Y7_to_NC),
    .from_ND(Tile_X6Y7_to_ND),
    .from_NF(Tile_X6Y7_to_NF),
    .from_NG(Tile_X6Y7_to_NG),
    .from_NH(Tile_X6Y7_to_NH),
    .from_NI(Tile_X6Y7_to_NI),
    .from_EA(Tile_X5Y6_to_EA),
    .from_EB(Tile_X5Y6_to_EB),
    .from_EC(Tile_X5Y6_to_EC),
    .from_ED(Tile_X5Y6_to_ED),
    .from_EF(Tile_X5Y6_to_EF),
    .from_EG(Tile_X5Y6_to_EG),
    .from_EH(Tile_X5Y6_to_EH),
    .from_EI(Tile_X5Y6_to_EI),
    .from_SA(Tile_X6Y5_to_SA),
    .from_SB(Tile_X6Y5_to_SB),
    .from_SC(Tile_X6Y5_to_SC),
    .from_SD(Tile_X6Y5_to_SD),
    .from_SF(Tile_X6Y5_to_SF),
    .from_SG(Tile_X6Y5_to_SG),
    .from_SH(Tile_X6Y5_to_SH),
    .from_SI(Tile_X6Y5_to_SI),
    .from_WA(Tile_X7Y6_to_WA),
    .from_WB(Tile_X7Y6_to_WB),
    .from_WC(Tile_X7Y6_to_WC),
    .from_WD(Tile_X7Y6_to_WD),
    .from_WF(Tile_X7Y6_to_WF),
    .from_WG(Tile_X7Y6_to_WG),
    .from_WH(Tile_X7Y6_to_WH),
    .from_WI(Tile_X7Y6_to_WI),
    .to_EA(Tile_X6Y6_to_EA),
    .to_EB(Tile_X6Y6_to_EB),
    .to_EC(Tile_X6Y6_to_EC),
    .to_ED(Tile_X6Y6_to_ED),
    .to_EF(Tile_X6Y6_to_EF),
    .to_EG(Tile_X6Y6_to_EG),
    .to_EH(Tile_X6Y6_to_EH),
    .to_EI(Tile_X6Y6_to_EI),
    .to_WA(Tile_X6Y6_to_WA),
    .to_WB(Tile_X6Y6_to_WB),
    .to_WC(Tile_X6Y6_to_WC),
    .to_WD(Tile_X6Y6_to_WD),
    .to_WF(Tile_X6Y6_to_WF),
    .to_WG(Tile_X6Y6_to_WG),
    .to_WH(Tile_X6Y6_to_WH),
    .to_WI(Tile_X6Y6_to_WI),
    .to_NA(Tile_X6Y6_to_NA),
    .to_NB(Tile_X6Y6_to_NB),
    .to_NC(Tile_X6Y6_to_NC),
    .to_ND(Tile_X6Y6_to_ND),
    .to_NF(Tile_X6Y6_to_NF),
    .to_NG(Tile_X6Y6_to_NG),
    .to_NH(Tile_X6Y6_to_NH),
    .to_NI(Tile_X6Y6_to_NI),
    .to_SA(Tile_X6Y6_to_SA),
    .to_SB(Tile_X6Y6_to_SB),
    .to_SC(Tile_X6Y6_to_SC),
    .to_SD(Tile_X6Y6_to_SD),
    .to_SF(Tile_X6Y6_to_SF),
    .to_SG(Tile_X6Y6_to_SG),
    .to_SH(Tile_X6Y6_to_SH),
    .to_SI(Tile_X6Y6_to_SI),
    .R_t(Tile_X6Y6_R_t),
    .R_f(Tile_X6Y6_R_f),
    .F_masked1(Tile_X6Y6_F_masked1),
    .F_masked2(Tile_X6Y6_F_masked2),
    .UserCLK(Tile_X6Y7_UserCLKo),
    .UserCLKo(Tile_X6Y6_UserCLKo),
    .rst(Tile_X6Y7_rsto),
    .rsto(Tile_X6Y6_rsto),
    .FrameData(Tile_X5Y6_FrameData_O),
    .FrameData_O(Tile_X6Y6_FrameData_O),
    .FrameStrobe(Tile_X6Y7_FrameStrobe_O),
    .FrameStrobe_O(Tile_X6Y6_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X7Y6_Emulate_Bitstream)
    )
`endif
    Tile_X7Y6_linear_LMDPL
    (
    .from_NA(Tile_X7Y7_to_NA),
    .from_NB(Tile_X7Y7_to_NB),
    .from_NC(Tile_X7Y7_to_NC),
    .from_ND(Tile_X7Y7_to_ND),
    .from_NF(Tile_X7Y7_to_NF),
    .from_NG(Tile_X7Y7_to_NG),
    .from_NH(Tile_X7Y7_to_NH),
    .from_NI(Tile_X7Y7_to_NI),
    .from_EA(Tile_X6Y6_to_EA),
    .from_EB(Tile_X6Y6_to_EB),
    .from_EC(Tile_X6Y6_to_EC),
    .from_ED(Tile_X6Y6_to_ED),
    .from_EF(Tile_X6Y6_to_EF),
    .from_EG(Tile_X6Y6_to_EG),
    .from_EH(Tile_X6Y6_to_EH),
    .from_EI(Tile_X6Y6_to_EI),
    .from_SA(Tile_X7Y5_to_SA),
    .from_SB(Tile_X7Y5_to_SB),
    .from_SC(Tile_X7Y5_to_SC),
    .from_SD(Tile_X7Y5_to_SD),
    .from_SF(Tile_X7Y5_to_SF),
    .from_SG(Tile_X7Y5_to_SG),
    .from_SH(Tile_X7Y5_to_SH),
    .from_SI(Tile_X7Y5_to_SI),
    .from_WA(Tile_X8Y6_to_WA),
    .from_WB(Tile_X8Y6_to_WB),
    .from_WC(Tile_X8Y6_to_WC),
    .from_WD(Tile_X8Y6_to_WD),
    .from_WF(Tile_X8Y6_to_WF),
    .from_WG(Tile_X8Y6_to_WG),
    .from_WH(Tile_X8Y6_to_WH),
    .from_WI(Tile_X8Y6_to_WI),
    .to_EA(Tile_X7Y6_to_EA),
    .to_EB(Tile_X7Y6_to_EB),
    .to_EC(Tile_X7Y6_to_EC),
    .to_ED(Tile_X7Y6_to_ED),
    .to_EF(Tile_X7Y6_to_EF),
    .to_EG(Tile_X7Y6_to_EG),
    .to_EH(Tile_X7Y6_to_EH),
    .to_EI(Tile_X7Y6_to_EI),
    .to_WA(Tile_X7Y6_to_WA),
    .to_WB(Tile_X7Y6_to_WB),
    .to_WC(Tile_X7Y6_to_WC),
    .to_WD(Tile_X7Y6_to_WD),
    .to_WF(Tile_X7Y6_to_WF),
    .to_WG(Tile_X7Y6_to_WG),
    .to_WH(Tile_X7Y6_to_WH),
    .to_WI(Tile_X7Y6_to_WI),
    .to_NA(Tile_X7Y6_to_NA),
    .to_NB(Tile_X7Y6_to_NB),
    .to_NC(Tile_X7Y6_to_NC),
    .to_ND(Tile_X7Y6_to_ND),
    .to_NF(Tile_X7Y6_to_NF),
    .to_NG(Tile_X7Y6_to_NG),
    .to_NH(Tile_X7Y6_to_NH),
    .to_NI(Tile_X7Y6_to_NI),
    .to_SA(Tile_X7Y6_to_SA),
    .to_SB(Tile_X7Y6_to_SB),
    .to_SC(Tile_X7Y6_to_SC),
    .to_SD(Tile_X7Y6_to_SD),
    .to_SF(Tile_X7Y6_to_SF),
    .to_SG(Tile_X7Y6_to_SG),
    .to_SH(Tile_X7Y6_to_SH),
    .to_SI(Tile_X7Y6_to_SI),
    .F_masked1(Tile_X7Y6_F_masked1),
    .F_masked2(Tile_X7Y6_F_masked2),
    .UserCLK(Tile_X7Y7_UserCLKo),
    .UserCLKo(Tile_X7Y6_UserCLKo),
    .rst(Tile_X7Y7_rsto),
    .rsto(Tile_X7Y6_rsto),
    .FrameData(Tile_X6Y6_FrameData_O),
    .FrameData_O(Tile_X7Y6_FrameData_O),
    .FrameStrobe(Tile_X7Y7_FrameStrobe_O),
    .FrameStrobe_O(Tile_X7Y6_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
ctrl_to_sec
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X8Y6_Emulate_Bitstream)
    )
`endif
    Tile_X8Y6_ctrl_to_sec
    (
    .from_NA(Tile_X8Y7_to_NA),
    .from_NB(Tile_X8Y7_to_NB),
    .from_NC(Tile_X8Y7_to_NC),
    .from_ND(Tile_X8Y7_to_ND),
    .from_NF(Tile_X8Y7_to_NF),
    .from_NG(Tile_X8Y7_to_NG),
    .from_NH(Tile_X8Y7_to_NH),
    .from_NI(Tile_X8Y7_to_NI),
    .from_EA(Tile_X7Y6_to_EA),
    .from_EB(Tile_X7Y6_to_EB),
    .from_EC(Tile_X7Y6_to_EC),
    .from_ED(Tile_X7Y6_to_ED),
    .from_EF(Tile_X7Y6_to_EF),
    .from_EG(Tile_X7Y6_to_EG),
    .from_EH(Tile_X7Y6_to_EH),
    .from_EI(Tile_X7Y6_to_EI),
    .from_SA(Tile_X8Y5_to_SA),
    .from_SB(Tile_X8Y5_to_SB),
    .from_SC(Tile_X8Y5_to_SC),
    .from_SD(Tile_X8Y5_to_SD),
    .from_SF(Tile_X8Y5_to_SF),
    .from_SG(Tile_X8Y5_to_SG),
    .from_SH(Tile_X8Y5_to_SH),
    .from_SI(Tile_X8Y5_to_SI),
    .from_WA_1s(Tile_X9Y6_to_WA_1s),
    .from_WB_1s(Tile_X9Y6_to_WB_1s),
    .from_WC_1s(Tile_X9Y6_to_WC_1s),
    .from_WD_1s(Tile_X9Y6_to_WD_1s),
    .from_WF_1s(Tile_X9Y6_to_WF_1s),
    .from_WG_1s(Tile_X9Y6_to_WG_1s),
    .from_WH_1s(Tile_X9Y6_to_WH_1s),
    .from_WI_1s(Tile_X9Y6_to_WI_1s),
    .to_WA(Tile_X8Y6_to_WA),
    .to_WB(Tile_X8Y6_to_WB),
    .to_WC(Tile_X8Y6_to_WC),
    .to_WD(Tile_X8Y6_to_WD),
    .to_WF(Tile_X8Y6_to_WF),
    .to_WG(Tile_X8Y6_to_WG),
    .to_WH(Tile_X8Y6_to_WH),
    .to_WI(Tile_X8Y6_to_WI),
    .to_NA(Tile_X8Y6_to_NA),
    .to_NB(Tile_X8Y6_to_NB),
    .to_NC(Tile_X8Y6_to_NC),
    .to_ND(Tile_X8Y6_to_ND),
    .to_NF(Tile_X8Y6_to_NF),
    .to_NG(Tile_X8Y6_to_NG),
    .to_NH(Tile_X8Y6_to_NH),
    .to_NI(Tile_X8Y6_to_NI),
    .to_SA(Tile_X8Y6_to_SA),
    .to_SB(Tile_X8Y6_to_SB),
    .to_SC(Tile_X8Y6_to_SC),
    .to_SD(Tile_X8Y6_to_SD),
    .to_SF(Tile_X8Y6_to_SF),
    .to_SG(Tile_X8Y6_to_SG),
    .to_SH(Tile_X8Y6_to_SH),
    .to_SI(Tile_X8Y6_to_SI),
    .UserCLK(Tile_X8Y7_UserCLKo),
    .UserCLKo(Tile_X8Y6_UserCLKo),
    .rst(Tile_X8Y7_rsto),
    .rsto(Tile_X8Y6_rsto),
    .FrameData(Tile_X7Y6_FrameData_O),
    .FrameData_O(Tile_X8Y6_FrameData_O),
    .FrameStrobe(Tile_X8Y7_FrameStrobe_O),
    .FrameStrobe_O(Tile_X8Y6_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
combined_WDDL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X9Y6_Emulate_Bitstream)
    )
`endif
    Tile_X9Y6_combined_WDDL
    (
    .from_NA_1s(Tile_X9Y7_to_NA_1s),
    .from_NB_1s(Tile_X9Y7_to_NB_1s),
    .from_NC_1s(Tile_X9Y7_to_NC_1s),
    .from_ND_1s(Tile_X9Y7_to_ND_1s),
    .from_NF_1s(Tile_X9Y7_to_NF_1s),
    .from_NG_1s(Tile_X9Y7_to_NG_1s),
    .from_NH_1s(Tile_X9Y7_to_NH_1s),
    .from_NI_1s(Tile_X9Y7_to_NI_1s),
    .from_SA_1s(Tile_X9Y5_to_SA_1s),
    .from_SB_1s(Tile_X9Y5_to_SB_1s),
    .from_SC_1s(Tile_X9Y5_to_SC_1s),
    .from_SD_1s(Tile_X9Y5_to_SD_1s),
    .from_SF_1s(Tile_X9Y5_to_SF_1s),
    .from_SG_1s(Tile_X9Y5_to_SG_1s),
    .from_SH_1s(Tile_X9Y5_to_SH_1s),
    .from_SI_1s(Tile_X9Y5_to_SI_1s),
    .from_WA_1s(Tile_X10Y6_to_WA_1s),
    .from_WB_1s(Tile_X10Y6_to_WB_1s),
    .from_WC_1s(Tile_X10Y6_to_WC_1s),
    .from_WD_1s(Tile_X10Y6_to_WD_1s),
    .from_WF_1s(Tile_X10Y6_to_WF_1s),
    .from_WG_1s(Tile_X10Y6_to_WG_1s),
    .from_WH_1s(Tile_X10Y6_to_WH_1s),
    .from_WI_1s(Tile_X10Y6_to_WI_1s),
    .to_EA_1s(Tile_X9Y6_to_EA_1s),
    .to_EB_1s(Tile_X9Y6_to_EB_1s),
    .to_EC_1s(Tile_X9Y6_to_EC_1s),
    .to_ED_1s(Tile_X9Y6_to_ED_1s),
    .to_EF_1s(Tile_X9Y6_to_EF_1s),
    .to_EG_1s(Tile_X9Y6_to_EG_1s),
    .to_EH_1s(Tile_X9Y6_to_EH_1s),
    .to_EI_1s(Tile_X9Y6_to_EI_1s),
    .to_WA_1s(Tile_X9Y6_to_WA_1s),
    .to_WB_1s(Tile_X9Y6_to_WB_1s),
    .to_WC_1s(Tile_X9Y6_to_WC_1s),
    .to_WD_1s(Tile_X9Y6_to_WD_1s),
    .to_WF_1s(Tile_X9Y6_to_WF_1s),
    .to_WG_1s(Tile_X9Y6_to_WG_1s),
    .to_WH_1s(Tile_X9Y6_to_WH_1s),
    .to_WI_1s(Tile_X9Y6_to_WI_1s),
    .to_NA_1s(Tile_X9Y6_to_NA_1s),
    .to_NB_1s(Tile_X9Y6_to_NB_1s),
    .to_NC_1s(Tile_X9Y6_to_NC_1s),
    .to_ND_1s(Tile_X9Y6_to_ND_1s),
    .to_NF_1s(Tile_X9Y6_to_NF_1s),
    .to_NG_1s(Tile_X9Y6_to_NG_1s),
    .to_NH_1s(Tile_X9Y6_to_NH_1s),
    .to_NI_1s(Tile_X9Y6_to_NI_1s),
    .to_SA_1s(Tile_X9Y6_to_SA_1s),
    .to_SB_1s(Tile_X9Y6_to_SB_1s),
    .to_SC_1s(Tile_X9Y6_to_SC_1s),
    .to_SD_1s(Tile_X9Y6_to_SD_1s),
    .to_SF_1s(Tile_X9Y6_to_SF_1s),
    .to_SG_1s(Tile_X9Y6_to_SG_1s),
    .to_SH_1s(Tile_X9Y6_to_SH_1s),
    .to_SI_1s(Tile_X9Y6_to_SI_1s),
    .F_ctrl(Tile_X9Y6_F_ctrl),
    .UserCLK(Tile_X9Y7_UserCLKo),
    .UserCLKo(Tile_X9Y6_UserCLKo),
    .rst(Tile_X9Y7_rsto),
    .rsto(Tile_X9Y6_rsto),
    .FrameData(Tile_X8Y6_FrameData_O),
    .FrameData_O(Tile_X9Y6_FrameData_O),
    .FrameStrobe(Tile_X9Y7_FrameStrobe_O),
    .FrameStrobe_O(Tile_X9Y6_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
ctrl_IO
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X10Y6_Emulate_Bitstream)
    )
`endif
    Tile_X10Y6_ctrl_IO
    (
    .from_EA_1s(Tile_X9Y6_to_EA_1s),
    .from_EB_1s(Tile_X9Y6_to_EB_1s),
    .from_EC_1s(Tile_X9Y6_to_EC_1s),
    .from_ED_1s(Tile_X9Y6_to_ED_1s),
    .from_EF_1s(Tile_X9Y6_to_EF_1s),
    .from_EG_1s(Tile_X9Y6_to_EG_1s),
    .from_EH_1s(Tile_X9Y6_to_EH_1s),
    .from_EI_1s(Tile_X9Y6_to_EI_1s),
    .to_WA_1s(Tile_X10Y6_to_WA_1s),
    .to_WB_1s(Tile_X10Y6_to_WB_1s),
    .to_WC_1s(Tile_X10Y6_to_WC_1s),
    .to_WD_1s(Tile_X10Y6_to_WD_1s),
    .to_WF_1s(Tile_X10Y6_to_WF_1s),
    .to_WG_1s(Tile_X10Y6_to_WG_1s),
    .to_WH_1s(Tile_X10Y6_to_WH_1s),
    .to_WI_1s(Tile_X10Y6_to_WI_1s),
    .A_O_top_0_t(Tile_X10Y6_A_O_top_0_t),
    .A_O_top_0_f(Tile_X10Y6_A_O_top_0_f),
    .A_prech2(Tile_X10Y6_A_prech2),
    .A_DR_fault(Tile_X10Y6_A_DR_fault),
    .A_I_top_0_t(Tile_X10Y6_A_I_top_0_t),
    .A_I_top_0_f(Tile_X10Y6_A_I_top_0_f),
    .A_T_top(Tile_X10Y6_A_T_top),
    .A_F_ctrl(Tile_X10Y6_A_F_ctrl),
    .UserCLK(Tile_X10Y7_UserCLKo),
    .UserCLKo(Tile_X10Y6_UserCLKo),
    .rst(Tile_X10Y7_rsto),
    .rsto(Tile_X10Y6_rsto),
    .FrameData(Tile_X9Y6_FrameData_O),
    .FrameData_O(Tile_X10Y6_FrameData_O),
    .FrameStrobe(Tile_X10Y7_FrameStrobe_O),
    .FrameStrobe_O(Tile_X10Y6_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
W_IO_custom
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X0Y7_Emulate_Bitstream)
    )
`endif
    Tile_X0Y7_W_IO_custom
    (
    .from_NA(Tile_X0Y8_to_NA),
    .from_NB(Tile_X0Y8_to_NB),
    .from_NC(Tile_X0Y8_to_NC),
    .from_ND(Tile_X0Y8_to_ND),
    .from_NF(Tile_X0Y8_to_NF),
    .from_NG(Tile_X0Y8_to_NG),
    .from_NH(Tile_X0Y8_to_NH),
    .from_NI(Tile_X0Y8_to_NI),
    .from_SA(Tile_X0Y6_to_SA),
    .from_SB(Tile_X0Y6_to_SB),
    .from_SC(Tile_X0Y6_to_SC),
    .from_SD(Tile_X0Y6_to_SD),
    .from_SF(Tile_X0Y6_to_SF),
    .from_SG(Tile_X0Y6_to_SG),
    .from_SH(Tile_X0Y6_to_SH),
    .from_SI(Tile_X0Y6_to_SI),
    .from_WA(Tile_X1Y7_to_WA),
    .from_WB(Tile_X1Y7_to_WB),
    .from_WC(Tile_X1Y7_to_WC),
    .from_WD(Tile_X1Y7_to_WD),
    .from_WF(Tile_X1Y7_to_WF),
    .from_WG(Tile_X1Y7_to_WG),
    .from_WH(Tile_X1Y7_to_WH),
    .from_WI(Tile_X1Y7_to_WI),
    .to_EA(Tile_X0Y7_to_EA),
    .to_EB(Tile_X0Y7_to_EB),
    .to_EC(Tile_X0Y7_to_EC),
    .to_ED(Tile_X0Y7_to_ED),
    .to_EF(Tile_X0Y7_to_EF),
    .to_EG(Tile_X0Y7_to_EG),
    .to_EH(Tile_X0Y7_to_EH),
    .to_EI(Tile_X0Y7_to_EI),
    .to_NA(Tile_X0Y7_to_NA),
    .to_NB(Tile_X0Y7_to_NB),
    .to_NC(Tile_X0Y7_to_NC),
    .to_ND(Tile_X0Y7_to_ND),
    .to_NF(Tile_X0Y7_to_NF),
    .to_NG(Tile_X0Y7_to_NG),
    .to_NH(Tile_X0Y7_to_NH),
    .to_NI(Tile_X0Y7_to_NI),
    .to_SA(Tile_X0Y7_to_SA),
    .to_SB(Tile_X0Y7_to_SB),
    .to_SC(Tile_X0Y7_to_SC),
    .to_SD(Tile_X0Y7_to_SD),
    .to_SF(Tile_X0Y7_to_SF),
    .to_SG(Tile_X0Y7_to_SG),
    .to_SH(Tile_X0Y7_to_SH),
    .to_SI(Tile_X0Y7_to_SI),
    .A_O_top_0_t(Tile_X0Y7_A_O_top_0_t),
    .A_O_top_0_f(Tile_X0Y7_A_O_top_0_f),
    .A_O_top_1_t(Tile_X0Y7_A_O_top_1_t),
    .A_O_top_1_f(Tile_X0Y7_A_O_top_1_f),
    .A_prech1(Tile_X0Y7_A_prech1),
    .A_prech2(Tile_X0Y7_A_prech2),
    .A_DR_fault(Tile_X0Y7_A_DR_fault),
    .A_I_top_0_t(Tile_X0Y7_A_I_top_0_t),
    .A_I_top_0_f(Tile_X0Y7_A_I_top_0_f),
    .A_I_top_1_t(Tile_X0Y7_A_I_top_1_t),
    .A_I_top_1_f(Tile_X0Y7_A_I_top_1_f),
    .A_T_top(Tile_X0Y7_A_T_top),
    .A_F_masked1(Tile_X0Y7_A_F_masked1),
    .A_F_masked2(Tile_X0Y7_A_F_masked2),
    .A_config_C_bit0(Tile_X0Y7_A_config_C_bit0),
    .A_config_C_bit1(Tile_X0Y7_A_config_C_bit1),
    .A_config_C_bit2(Tile_X0Y7_A_config_C_bit2),
    .A_config_C_bit3(Tile_X0Y7_A_config_C_bit3),
    .B_config_C_bit0(Tile_X0Y7_B_config_C_bit0),
    .B_config_C_bit1(Tile_X0Y7_B_config_C_bit1),
    .B_config_C_bit2(Tile_X0Y7_B_config_C_bit2),
    .B_config_C_bit3(Tile_X0Y7_B_config_C_bit3),
    .UserCLK(Tile_X0Y8_UserCLKo),
    .UserCLKo(Tile_X0Y7_UserCLKo),
    .rst(Tile_X0Y8_rsto),
    .rsto(Tile_X0Y7_rsto),
    .FrameData(Tile_Y7_FrameData),
    .FrameData_O(Tile_X0Y7_FrameData_O),
    .FrameStrobe(Tile_X0Y8_FrameStrobe_O),
    .FrameStrobe_O(Tile_X0Y7_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X1Y7_Emulate_Bitstream)
    )
`endif
    Tile_X1Y7_linear_LMDPL
    (
    .from_NA(Tile_X1Y8_to_NA),
    .from_NB(Tile_X1Y8_to_NB),
    .from_NC(Tile_X1Y8_to_NC),
    .from_ND(Tile_X1Y8_to_ND),
    .from_NF(Tile_X1Y8_to_NF),
    .from_NG(Tile_X1Y8_to_NG),
    .from_NH(Tile_X1Y8_to_NH),
    .from_NI(Tile_X1Y8_to_NI),
    .from_EA(Tile_X0Y7_to_EA),
    .from_EB(Tile_X0Y7_to_EB),
    .from_EC(Tile_X0Y7_to_EC),
    .from_ED(Tile_X0Y7_to_ED),
    .from_EF(Tile_X0Y7_to_EF),
    .from_EG(Tile_X0Y7_to_EG),
    .from_EH(Tile_X0Y7_to_EH),
    .from_EI(Tile_X0Y7_to_EI),
    .from_SA(Tile_X1Y6_to_SA),
    .from_SB(Tile_X1Y6_to_SB),
    .from_SC(Tile_X1Y6_to_SC),
    .from_SD(Tile_X1Y6_to_SD),
    .from_SF(Tile_X1Y6_to_SF),
    .from_SG(Tile_X1Y6_to_SG),
    .from_SH(Tile_X1Y6_to_SH),
    .from_SI(Tile_X1Y6_to_SI),
    .from_WA(Tile_X2Y7_to_WA),
    .from_WB(Tile_X2Y7_to_WB),
    .from_WC(Tile_X2Y7_to_WC),
    .from_WD(Tile_X2Y7_to_WD),
    .from_WF(Tile_X2Y7_to_WF),
    .from_WG(Tile_X2Y7_to_WG),
    .from_WH(Tile_X2Y7_to_WH),
    .from_WI(Tile_X2Y7_to_WI),
    .to_EA(Tile_X1Y7_to_EA),
    .to_EB(Tile_X1Y7_to_EB),
    .to_EC(Tile_X1Y7_to_EC),
    .to_ED(Tile_X1Y7_to_ED),
    .to_EF(Tile_X1Y7_to_EF),
    .to_EG(Tile_X1Y7_to_EG),
    .to_EH(Tile_X1Y7_to_EH),
    .to_EI(Tile_X1Y7_to_EI),
    .to_WA(Tile_X1Y7_to_WA),
    .to_WB(Tile_X1Y7_to_WB),
    .to_WC(Tile_X1Y7_to_WC),
    .to_WD(Tile_X1Y7_to_WD),
    .to_WF(Tile_X1Y7_to_WF),
    .to_WG(Tile_X1Y7_to_WG),
    .to_WH(Tile_X1Y7_to_WH),
    .to_WI(Tile_X1Y7_to_WI),
    .to_NA(Tile_X1Y7_to_NA),
    .to_NB(Tile_X1Y7_to_NB),
    .to_NC(Tile_X1Y7_to_NC),
    .to_ND(Tile_X1Y7_to_ND),
    .to_NF(Tile_X1Y7_to_NF),
    .to_NG(Tile_X1Y7_to_NG),
    .to_NH(Tile_X1Y7_to_NH),
    .to_NI(Tile_X1Y7_to_NI),
    .to_SA(Tile_X1Y7_to_SA),
    .to_SB(Tile_X1Y7_to_SB),
    .to_SC(Tile_X1Y7_to_SC),
    .to_SD(Tile_X1Y7_to_SD),
    .to_SF(Tile_X1Y7_to_SF),
    .to_SG(Tile_X1Y7_to_SG),
    .to_SH(Tile_X1Y7_to_SH),
    .to_SI(Tile_X1Y7_to_SI),
    .F_masked1(Tile_X1Y7_F_masked1),
    .F_masked2(Tile_X1Y7_F_masked2),
    .UserCLK(Tile_X1Y8_UserCLKo),
    .UserCLKo(Tile_X1Y7_UserCLKo),
    .rst(Tile_X1Y8_rsto),
    .rsto(Tile_X1Y7_rsto),
    .FrameData(Tile_X0Y7_FrameData_O),
    .FrameData_O(Tile_X1Y7_FrameData_O),
    .FrameStrobe(Tile_X1Y8_FrameStrobe_O),
    .FrameStrobe_O(Tile_X1Y7_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X2Y7_Emulate_Bitstream)
    )
`endif
    Tile_X2Y7_linear_LMDPL
    (
    .from_NA(Tile_X2Y8_to_NA),
    .from_NB(Tile_X2Y8_to_NB),
    .from_NC(Tile_X2Y8_to_NC),
    .from_ND(Tile_X2Y8_to_ND),
    .from_NF(Tile_X2Y8_to_NF),
    .from_NG(Tile_X2Y8_to_NG),
    .from_NH(Tile_X2Y8_to_NH),
    .from_NI(Tile_X2Y8_to_NI),
    .from_EA(Tile_X1Y7_to_EA),
    .from_EB(Tile_X1Y7_to_EB),
    .from_EC(Tile_X1Y7_to_EC),
    .from_ED(Tile_X1Y7_to_ED),
    .from_EF(Tile_X1Y7_to_EF),
    .from_EG(Tile_X1Y7_to_EG),
    .from_EH(Tile_X1Y7_to_EH),
    .from_EI(Tile_X1Y7_to_EI),
    .from_SA(Tile_X2Y6_to_SA),
    .from_SB(Tile_X2Y6_to_SB),
    .from_SC(Tile_X2Y6_to_SC),
    .from_SD(Tile_X2Y6_to_SD),
    .from_SF(Tile_X2Y6_to_SF),
    .from_SG(Tile_X2Y6_to_SG),
    .from_SH(Tile_X2Y6_to_SH),
    .from_SI(Tile_X2Y6_to_SI),
    .from_WA(Tile_X3Y7_to_WA),
    .from_WB(Tile_X3Y7_to_WB),
    .from_WC(Tile_X3Y7_to_WC),
    .from_WD(Tile_X3Y7_to_WD),
    .from_WF(Tile_X3Y7_to_WF),
    .from_WG(Tile_X3Y7_to_WG),
    .from_WH(Tile_X3Y7_to_WH),
    .from_WI(Tile_X3Y7_to_WI),
    .to_EA(Tile_X2Y7_to_EA),
    .to_EB(Tile_X2Y7_to_EB),
    .to_EC(Tile_X2Y7_to_EC),
    .to_ED(Tile_X2Y7_to_ED),
    .to_EF(Tile_X2Y7_to_EF),
    .to_EG(Tile_X2Y7_to_EG),
    .to_EH(Tile_X2Y7_to_EH),
    .to_EI(Tile_X2Y7_to_EI),
    .to_WA(Tile_X2Y7_to_WA),
    .to_WB(Tile_X2Y7_to_WB),
    .to_WC(Tile_X2Y7_to_WC),
    .to_WD(Tile_X2Y7_to_WD),
    .to_WF(Tile_X2Y7_to_WF),
    .to_WG(Tile_X2Y7_to_WG),
    .to_WH(Tile_X2Y7_to_WH),
    .to_WI(Tile_X2Y7_to_WI),
    .to_NA(Tile_X2Y7_to_NA),
    .to_NB(Tile_X2Y7_to_NB),
    .to_NC(Tile_X2Y7_to_NC),
    .to_ND(Tile_X2Y7_to_ND),
    .to_NF(Tile_X2Y7_to_NF),
    .to_NG(Tile_X2Y7_to_NG),
    .to_NH(Tile_X2Y7_to_NH),
    .to_NI(Tile_X2Y7_to_NI),
    .to_SA(Tile_X2Y7_to_SA),
    .to_SB(Tile_X2Y7_to_SB),
    .to_SC(Tile_X2Y7_to_SC),
    .to_SD(Tile_X2Y7_to_SD),
    .to_SF(Tile_X2Y7_to_SF),
    .to_SG(Tile_X2Y7_to_SG),
    .to_SH(Tile_X2Y7_to_SH),
    .to_SI(Tile_X2Y7_to_SI),
    .F_masked1(Tile_X2Y7_F_masked1),
    .F_masked2(Tile_X2Y7_F_masked2),
    .UserCLK(Tile_X2Y8_UserCLKo),
    .UserCLKo(Tile_X2Y7_UserCLKo),
    .rst(Tile_X2Y8_rsto),
    .rsto(Tile_X2Y7_rsto),
    .FrameData(Tile_X1Y7_FrameData_O),
    .FrameData_O(Tile_X2Y7_FrameData_O),
    .FrameStrobe(Tile_X2Y8_FrameStrobe_O),
    .FrameStrobe_O(Tile_X2Y7_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
nonlinear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X3Y7_Emulate_Bitstream)
    )
`endif
    Tile_X3Y7_nonlinear_LMDPL
    (
    .from_NA(Tile_X3Y8_to_NA),
    .from_NB(Tile_X3Y8_to_NB),
    .from_NC(Tile_X3Y8_to_NC),
    .from_ND(Tile_X3Y8_to_ND),
    .from_NF(Tile_X3Y8_to_NF),
    .from_NG(Tile_X3Y8_to_NG),
    .from_NH(Tile_X3Y8_to_NH),
    .from_NI(Tile_X3Y8_to_NI),
    .from_EA(Tile_X2Y7_to_EA),
    .from_EB(Tile_X2Y7_to_EB),
    .from_EC(Tile_X2Y7_to_EC),
    .from_ED(Tile_X2Y7_to_ED),
    .from_EF(Tile_X2Y7_to_EF),
    .from_EG(Tile_X2Y7_to_EG),
    .from_EH(Tile_X2Y7_to_EH),
    .from_EI(Tile_X2Y7_to_EI),
    .from_SA(Tile_X3Y6_to_SA),
    .from_SB(Tile_X3Y6_to_SB),
    .from_SC(Tile_X3Y6_to_SC),
    .from_SD(Tile_X3Y6_to_SD),
    .from_SF(Tile_X3Y6_to_SF),
    .from_SG(Tile_X3Y6_to_SG),
    .from_SH(Tile_X3Y6_to_SH),
    .from_SI(Tile_X3Y6_to_SI),
    .from_WA(Tile_X4Y7_to_WA),
    .from_WB(Tile_X4Y7_to_WB),
    .from_WC(Tile_X4Y7_to_WC),
    .from_WD(Tile_X4Y7_to_WD),
    .from_WF(Tile_X4Y7_to_WF),
    .from_WG(Tile_X4Y7_to_WG),
    .from_WH(Tile_X4Y7_to_WH),
    .from_WI(Tile_X4Y7_to_WI),
    .to_EA(Tile_X3Y7_to_EA),
    .to_EB(Tile_X3Y7_to_EB),
    .to_EC(Tile_X3Y7_to_EC),
    .to_ED(Tile_X3Y7_to_ED),
    .to_EF(Tile_X3Y7_to_EF),
    .to_EG(Tile_X3Y7_to_EG),
    .to_EH(Tile_X3Y7_to_EH),
    .to_EI(Tile_X3Y7_to_EI),
    .to_WA(Tile_X3Y7_to_WA),
    .to_WB(Tile_X3Y7_to_WB),
    .to_WC(Tile_X3Y7_to_WC),
    .to_WD(Tile_X3Y7_to_WD),
    .to_WF(Tile_X3Y7_to_WF),
    .to_WG(Tile_X3Y7_to_WG),
    .to_WH(Tile_X3Y7_to_WH),
    .to_WI(Tile_X3Y7_to_WI),
    .to_NA(Tile_X3Y7_to_NA),
    .to_NB(Tile_X3Y7_to_NB),
    .to_NC(Tile_X3Y7_to_NC),
    .to_ND(Tile_X3Y7_to_ND),
    .to_NF(Tile_X3Y7_to_NF),
    .to_NG(Tile_X3Y7_to_NG),
    .to_NH(Tile_X3Y7_to_NH),
    .to_NI(Tile_X3Y7_to_NI),
    .to_SA(Tile_X3Y7_to_SA),
    .to_SB(Tile_X3Y7_to_SB),
    .to_SC(Tile_X3Y7_to_SC),
    .to_SD(Tile_X3Y7_to_SD),
    .to_SF(Tile_X3Y7_to_SF),
    .to_SG(Tile_X3Y7_to_SG),
    .to_SH(Tile_X3Y7_to_SH),
    .to_SI(Tile_X3Y7_to_SI),
    .R_t(Tile_X3Y7_R_t),
    .R_f(Tile_X3Y7_R_f),
    .F_masked1(Tile_X3Y7_F_masked1),
    .F_masked2(Tile_X3Y7_F_masked2),
    .UserCLK(Tile_X3Y8_UserCLKo),
    .UserCLKo(Tile_X3Y7_UserCLKo),
    .rst(Tile_X3Y8_rsto),
    .rsto(Tile_X3Y7_rsto),
    .FrameData(Tile_X2Y7_FrameData_O),
    .FrameData_O(Tile_X3Y7_FrameData_O),
    .FrameStrobe(Tile_X3Y8_FrameStrobe_O),
    .FrameStrobe_O(Tile_X3Y7_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X4Y7_Emulate_Bitstream)
    )
`endif
    Tile_X4Y7_linear_LMDPL
    (
    .from_NA(Tile_X4Y8_to_NA),
    .from_NB(Tile_X4Y8_to_NB),
    .from_NC(Tile_X4Y8_to_NC),
    .from_ND(Tile_X4Y8_to_ND),
    .from_NF(Tile_X4Y8_to_NF),
    .from_NG(Tile_X4Y8_to_NG),
    .from_NH(Tile_X4Y8_to_NH),
    .from_NI(Tile_X4Y8_to_NI),
    .from_EA(Tile_X3Y7_to_EA),
    .from_EB(Tile_X3Y7_to_EB),
    .from_EC(Tile_X3Y7_to_EC),
    .from_ED(Tile_X3Y7_to_ED),
    .from_EF(Tile_X3Y7_to_EF),
    .from_EG(Tile_X3Y7_to_EG),
    .from_EH(Tile_X3Y7_to_EH),
    .from_EI(Tile_X3Y7_to_EI),
    .from_SA(Tile_X4Y6_to_SA),
    .from_SB(Tile_X4Y6_to_SB),
    .from_SC(Tile_X4Y6_to_SC),
    .from_SD(Tile_X4Y6_to_SD),
    .from_SF(Tile_X4Y6_to_SF),
    .from_SG(Tile_X4Y6_to_SG),
    .from_SH(Tile_X4Y6_to_SH),
    .from_SI(Tile_X4Y6_to_SI),
    .from_WA(Tile_X5Y7_to_WA),
    .from_WB(Tile_X5Y7_to_WB),
    .from_WC(Tile_X5Y7_to_WC),
    .from_WD(Tile_X5Y7_to_WD),
    .from_WF(Tile_X5Y7_to_WF),
    .from_WG(Tile_X5Y7_to_WG),
    .from_WH(Tile_X5Y7_to_WH),
    .from_WI(Tile_X5Y7_to_WI),
    .to_EA(Tile_X4Y7_to_EA),
    .to_EB(Tile_X4Y7_to_EB),
    .to_EC(Tile_X4Y7_to_EC),
    .to_ED(Tile_X4Y7_to_ED),
    .to_EF(Tile_X4Y7_to_EF),
    .to_EG(Tile_X4Y7_to_EG),
    .to_EH(Tile_X4Y7_to_EH),
    .to_EI(Tile_X4Y7_to_EI),
    .to_WA(Tile_X4Y7_to_WA),
    .to_WB(Tile_X4Y7_to_WB),
    .to_WC(Tile_X4Y7_to_WC),
    .to_WD(Tile_X4Y7_to_WD),
    .to_WF(Tile_X4Y7_to_WF),
    .to_WG(Tile_X4Y7_to_WG),
    .to_WH(Tile_X4Y7_to_WH),
    .to_WI(Tile_X4Y7_to_WI),
    .to_NA(Tile_X4Y7_to_NA),
    .to_NB(Tile_X4Y7_to_NB),
    .to_NC(Tile_X4Y7_to_NC),
    .to_ND(Tile_X4Y7_to_ND),
    .to_NF(Tile_X4Y7_to_NF),
    .to_NG(Tile_X4Y7_to_NG),
    .to_NH(Tile_X4Y7_to_NH),
    .to_NI(Tile_X4Y7_to_NI),
    .to_SA(Tile_X4Y7_to_SA),
    .to_SB(Tile_X4Y7_to_SB),
    .to_SC(Tile_X4Y7_to_SC),
    .to_SD(Tile_X4Y7_to_SD),
    .to_SF(Tile_X4Y7_to_SF),
    .to_SG(Tile_X4Y7_to_SG),
    .to_SH(Tile_X4Y7_to_SH),
    .to_SI(Tile_X4Y7_to_SI),
    .F_masked1(Tile_X4Y7_F_masked1),
    .F_masked2(Tile_X4Y7_F_masked2),
    .UserCLK(Tile_X4Y8_UserCLKo),
    .UserCLKo(Tile_X4Y7_UserCLKo),
    .rst(Tile_X4Y8_rsto),
    .rsto(Tile_X4Y7_rsto),
    .FrameData(Tile_X3Y7_FrameData_O),
    .FrameData_O(Tile_X4Y7_FrameData_O),
    .FrameStrobe(Tile_X4Y8_FrameStrobe_O),
    .FrameStrobe_O(Tile_X4Y7_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X5Y7_Emulate_Bitstream)
    )
`endif
    Tile_X5Y7_linear_LMDPL
    (
    .from_NA(Tile_X5Y8_to_NA),
    .from_NB(Tile_X5Y8_to_NB),
    .from_NC(Tile_X5Y8_to_NC),
    .from_ND(Tile_X5Y8_to_ND),
    .from_NF(Tile_X5Y8_to_NF),
    .from_NG(Tile_X5Y8_to_NG),
    .from_NH(Tile_X5Y8_to_NH),
    .from_NI(Tile_X5Y8_to_NI),
    .from_EA(Tile_X4Y7_to_EA),
    .from_EB(Tile_X4Y7_to_EB),
    .from_EC(Tile_X4Y7_to_EC),
    .from_ED(Tile_X4Y7_to_ED),
    .from_EF(Tile_X4Y7_to_EF),
    .from_EG(Tile_X4Y7_to_EG),
    .from_EH(Tile_X4Y7_to_EH),
    .from_EI(Tile_X4Y7_to_EI),
    .from_SA(Tile_X5Y6_to_SA),
    .from_SB(Tile_X5Y6_to_SB),
    .from_SC(Tile_X5Y6_to_SC),
    .from_SD(Tile_X5Y6_to_SD),
    .from_SF(Tile_X5Y6_to_SF),
    .from_SG(Tile_X5Y6_to_SG),
    .from_SH(Tile_X5Y6_to_SH),
    .from_SI(Tile_X5Y6_to_SI),
    .from_WA(Tile_X6Y7_to_WA),
    .from_WB(Tile_X6Y7_to_WB),
    .from_WC(Tile_X6Y7_to_WC),
    .from_WD(Tile_X6Y7_to_WD),
    .from_WF(Tile_X6Y7_to_WF),
    .from_WG(Tile_X6Y7_to_WG),
    .from_WH(Tile_X6Y7_to_WH),
    .from_WI(Tile_X6Y7_to_WI),
    .to_EA(Tile_X5Y7_to_EA),
    .to_EB(Tile_X5Y7_to_EB),
    .to_EC(Tile_X5Y7_to_EC),
    .to_ED(Tile_X5Y7_to_ED),
    .to_EF(Tile_X5Y7_to_EF),
    .to_EG(Tile_X5Y7_to_EG),
    .to_EH(Tile_X5Y7_to_EH),
    .to_EI(Tile_X5Y7_to_EI),
    .to_WA(Tile_X5Y7_to_WA),
    .to_WB(Tile_X5Y7_to_WB),
    .to_WC(Tile_X5Y7_to_WC),
    .to_WD(Tile_X5Y7_to_WD),
    .to_WF(Tile_X5Y7_to_WF),
    .to_WG(Tile_X5Y7_to_WG),
    .to_WH(Tile_X5Y7_to_WH),
    .to_WI(Tile_X5Y7_to_WI),
    .to_NA(Tile_X5Y7_to_NA),
    .to_NB(Tile_X5Y7_to_NB),
    .to_NC(Tile_X5Y7_to_NC),
    .to_ND(Tile_X5Y7_to_ND),
    .to_NF(Tile_X5Y7_to_NF),
    .to_NG(Tile_X5Y7_to_NG),
    .to_NH(Tile_X5Y7_to_NH),
    .to_NI(Tile_X5Y7_to_NI),
    .to_SA(Tile_X5Y7_to_SA),
    .to_SB(Tile_X5Y7_to_SB),
    .to_SC(Tile_X5Y7_to_SC),
    .to_SD(Tile_X5Y7_to_SD),
    .to_SF(Tile_X5Y7_to_SF),
    .to_SG(Tile_X5Y7_to_SG),
    .to_SH(Tile_X5Y7_to_SH),
    .to_SI(Tile_X5Y7_to_SI),
    .F_masked1(Tile_X5Y7_F_masked1),
    .F_masked2(Tile_X5Y7_F_masked2),
    .UserCLK(Tile_X5Y8_UserCLKo),
    .UserCLKo(Tile_X5Y7_UserCLKo),
    .rst(Tile_X5Y8_rsto),
    .rsto(Tile_X5Y7_rsto),
    .FrameData(Tile_X4Y7_FrameData_O),
    .FrameData_O(Tile_X5Y7_FrameData_O),
    .FrameStrobe(Tile_X5Y8_FrameStrobe_O),
    .FrameStrobe_O(Tile_X5Y7_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
nonlinear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X6Y7_Emulate_Bitstream)
    )
`endif
    Tile_X6Y7_nonlinear_LMDPL
    (
    .from_NA(Tile_X6Y8_to_NA),
    .from_NB(Tile_X6Y8_to_NB),
    .from_NC(Tile_X6Y8_to_NC),
    .from_ND(Tile_X6Y8_to_ND),
    .from_NF(Tile_X6Y8_to_NF),
    .from_NG(Tile_X6Y8_to_NG),
    .from_NH(Tile_X6Y8_to_NH),
    .from_NI(Tile_X6Y8_to_NI),
    .from_EA(Tile_X5Y7_to_EA),
    .from_EB(Tile_X5Y7_to_EB),
    .from_EC(Tile_X5Y7_to_EC),
    .from_ED(Tile_X5Y7_to_ED),
    .from_EF(Tile_X5Y7_to_EF),
    .from_EG(Tile_X5Y7_to_EG),
    .from_EH(Tile_X5Y7_to_EH),
    .from_EI(Tile_X5Y7_to_EI),
    .from_SA(Tile_X6Y6_to_SA),
    .from_SB(Tile_X6Y6_to_SB),
    .from_SC(Tile_X6Y6_to_SC),
    .from_SD(Tile_X6Y6_to_SD),
    .from_SF(Tile_X6Y6_to_SF),
    .from_SG(Tile_X6Y6_to_SG),
    .from_SH(Tile_X6Y6_to_SH),
    .from_SI(Tile_X6Y6_to_SI),
    .from_WA(Tile_X7Y7_to_WA),
    .from_WB(Tile_X7Y7_to_WB),
    .from_WC(Tile_X7Y7_to_WC),
    .from_WD(Tile_X7Y7_to_WD),
    .from_WF(Tile_X7Y7_to_WF),
    .from_WG(Tile_X7Y7_to_WG),
    .from_WH(Tile_X7Y7_to_WH),
    .from_WI(Tile_X7Y7_to_WI),
    .to_EA(Tile_X6Y7_to_EA),
    .to_EB(Tile_X6Y7_to_EB),
    .to_EC(Tile_X6Y7_to_EC),
    .to_ED(Tile_X6Y7_to_ED),
    .to_EF(Tile_X6Y7_to_EF),
    .to_EG(Tile_X6Y7_to_EG),
    .to_EH(Tile_X6Y7_to_EH),
    .to_EI(Tile_X6Y7_to_EI),
    .to_WA(Tile_X6Y7_to_WA),
    .to_WB(Tile_X6Y7_to_WB),
    .to_WC(Tile_X6Y7_to_WC),
    .to_WD(Tile_X6Y7_to_WD),
    .to_WF(Tile_X6Y7_to_WF),
    .to_WG(Tile_X6Y7_to_WG),
    .to_WH(Tile_X6Y7_to_WH),
    .to_WI(Tile_X6Y7_to_WI),
    .to_NA(Tile_X6Y7_to_NA),
    .to_NB(Tile_X6Y7_to_NB),
    .to_NC(Tile_X6Y7_to_NC),
    .to_ND(Tile_X6Y7_to_ND),
    .to_NF(Tile_X6Y7_to_NF),
    .to_NG(Tile_X6Y7_to_NG),
    .to_NH(Tile_X6Y7_to_NH),
    .to_NI(Tile_X6Y7_to_NI),
    .to_SA(Tile_X6Y7_to_SA),
    .to_SB(Tile_X6Y7_to_SB),
    .to_SC(Tile_X6Y7_to_SC),
    .to_SD(Tile_X6Y7_to_SD),
    .to_SF(Tile_X6Y7_to_SF),
    .to_SG(Tile_X6Y7_to_SG),
    .to_SH(Tile_X6Y7_to_SH),
    .to_SI(Tile_X6Y7_to_SI),
    .R_t(Tile_X6Y7_R_t),
    .R_f(Tile_X6Y7_R_f),
    .F_masked1(Tile_X6Y7_F_masked1),
    .F_masked2(Tile_X6Y7_F_masked2),
    .UserCLK(Tile_X6Y8_UserCLKo),
    .UserCLKo(Tile_X6Y7_UserCLKo),
    .rst(Tile_X6Y8_rsto),
    .rsto(Tile_X6Y7_rsto),
    .FrameData(Tile_X5Y7_FrameData_O),
    .FrameData_O(Tile_X6Y7_FrameData_O),
    .FrameStrobe(Tile_X6Y8_FrameStrobe_O),
    .FrameStrobe_O(Tile_X6Y7_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X7Y7_Emulate_Bitstream)
    )
`endif
    Tile_X7Y7_linear_LMDPL
    (
    .from_NA(Tile_X7Y8_to_NA),
    .from_NB(Tile_X7Y8_to_NB),
    .from_NC(Tile_X7Y8_to_NC),
    .from_ND(Tile_X7Y8_to_ND),
    .from_NF(Tile_X7Y8_to_NF),
    .from_NG(Tile_X7Y8_to_NG),
    .from_NH(Tile_X7Y8_to_NH),
    .from_NI(Tile_X7Y8_to_NI),
    .from_EA(Tile_X6Y7_to_EA),
    .from_EB(Tile_X6Y7_to_EB),
    .from_EC(Tile_X6Y7_to_EC),
    .from_ED(Tile_X6Y7_to_ED),
    .from_EF(Tile_X6Y7_to_EF),
    .from_EG(Tile_X6Y7_to_EG),
    .from_EH(Tile_X6Y7_to_EH),
    .from_EI(Tile_X6Y7_to_EI),
    .from_SA(Tile_X7Y6_to_SA),
    .from_SB(Tile_X7Y6_to_SB),
    .from_SC(Tile_X7Y6_to_SC),
    .from_SD(Tile_X7Y6_to_SD),
    .from_SF(Tile_X7Y6_to_SF),
    .from_SG(Tile_X7Y6_to_SG),
    .from_SH(Tile_X7Y6_to_SH),
    .from_SI(Tile_X7Y6_to_SI),
    .from_WA(Tile_X8Y7_to_WA),
    .from_WB(Tile_X8Y7_to_WB),
    .from_WC(Tile_X8Y7_to_WC),
    .from_WD(Tile_X8Y7_to_WD),
    .from_WF(Tile_X8Y7_to_WF),
    .from_WG(Tile_X8Y7_to_WG),
    .from_WH(Tile_X8Y7_to_WH),
    .from_WI(Tile_X8Y7_to_WI),
    .to_EA(Tile_X7Y7_to_EA),
    .to_EB(Tile_X7Y7_to_EB),
    .to_EC(Tile_X7Y7_to_EC),
    .to_ED(Tile_X7Y7_to_ED),
    .to_EF(Tile_X7Y7_to_EF),
    .to_EG(Tile_X7Y7_to_EG),
    .to_EH(Tile_X7Y7_to_EH),
    .to_EI(Tile_X7Y7_to_EI),
    .to_WA(Tile_X7Y7_to_WA),
    .to_WB(Tile_X7Y7_to_WB),
    .to_WC(Tile_X7Y7_to_WC),
    .to_WD(Tile_X7Y7_to_WD),
    .to_WF(Tile_X7Y7_to_WF),
    .to_WG(Tile_X7Y7_to_WG),
    .to_WH(Tile_X7Y7_to_WH),
    .to_WI(Tile_X7Y7_to_WI),
    .to_NA(Tile_X7Y7_to_NA),
    .to_NB(Tile_X7Y7_to_NB),
    .to_NC(Tile_X7Y7_to_NC),
    .to_ND(Tile_X7Y7_to_ND),
    .to_NF(Tile_X7Y7_to_NF),
    .to_NG(Tile_X7Y7_to_NG),
    .to_NH(Tile_X7Y7_to_NH),
    .to_NI(Tile_X7Y7_to_NI),
    .to_SA(Tile_X7Y7_to_SA),
    .to_SB(Tile_X7Y7_to_SB),
    .to_SC(Tile_X7Y7_to_SC),
    .to_SD(Tile_X7Y7_to_SD),
    .to_SF(Tile_X7Y7_to_SF),
    .to_SG(Tile_X7Y7_to_SG),
    .to_SH(Tile_X7Y7_to_SH),
    .to_SI(Tile_X7Y7_to_SI),
    .F_masked1(Tile_X7Y7_F_masked1),
    .F_masked2(Tile_X7Y7_F_masked2),
    .UserCLK(Tile_X7Y8_UserCLKo),
    .UserCLKo(Tile_X7Y7_UserCLKo),
    .rst(Tile_X7Y8_rsto),
    .rsto(Tile_X7Y7_rsto),
    .FrameData(Tile_X6Y7_FrameData_O),
    .FrameData_O(Tile_X7Y7_FrameData_O),
    .FrameStrobe(Tile_X7Y8_FrameStrobe_O),
    .FrameStrobe_O(Tile_X7Y7_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
ctrl_to_sec
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X8Y7_Emulate_Bitstream)
    )
`endif
    Tile_X8Y7_ctrl_to_sec
    (
    .from_NA(Tile_X8Y8_to_NA),
    .from_NB(Tile_X8Y8_to_NB),
    .from_NC(Tile_X8Y8_to_NC),
    .from_ND(Tile_X8Y8_to_ND),
    .from_NF(Tile_X8Y8_to_NF),
    .from_NG(Tile_X8Y8_to_NG),
    .from_NH(Tile_X8Y8_to_NH),
    .from_NI(Tile_X8Y8_to_NI),
    .from_EA(Tile_X7Y7_to_EA),
    .from_EB(Tile_X7Y7_to_EB),
    .from_EC(Tile_X7Y7_to_EC),
    .from_ED(Tile_X7Y7_to_ED),
    .from_EF(Tile_X7Y7_to_EF),
    .from_EG(Tile_X7Y7_to_EG),
    .from_EH(Tile_X7Y7_to_EH),
    .from_EI(Tile_X7Y7_to_EI),
    .from_SA(Tile_X8Y6_to_SA),
    .from_SB(Tile_X8Y6_to_SB),
    .from_SC(Tile_X8Y6_to_SC),
    .from_SD(Tile_X8Y6_to_SD),
    .from_SF(Tile_X8Y6_to_SF),
    .from_SG(Tile_X8Y6_to_SG),
    .from_SH(Tile_X8Y6_to_SH),
    .from_SI(Tile_X8Y6_to_SI),
    .from_WA_1s(Tile_X9Y7_to_WA_1s),
    .from_WB_1s(Tile_X9Y7_to_WB_1s),
    .from_WC_1s(Tile_X9Y7_to_WC_1s),
    .from_WD_1s(Tile_X9Y7_to_WD_1s),
    .from_WF_1s(Tile_X9Y7_to_WF_1s),
    .from_WG_1s(Tile_X9Y7_to_WG_1s),
    .from_WH_1s(Tile_X9Y7_to_WH_1s),
    .from_WI_1s(Tile_X9Y7_to_WI_1s),
    .to_WA(Tile_X8Y7_to_WA),
    .to_WB(Tile_X8Y7_to_WB),
    .to_WC(Tile_X8Y7_to_WC),
    .to_WD(Tile_X8Y7_to_WD),
    .to_WF(Tile_X8Y7_to_WF),
    .to_WG(Tile_X8Y7_to_WG),
    .to_WH(Tile_X8Y7_to_WH),
    .to_WI(Tile_X8Y7_to_WI),
    .to_NA(Tile_X8Y7_to_NA),
    .to_NB(Tile_X8Y7_to_NB),
    .to_NC(Tile_X8Y7_to_NC),
    .to_ND(Tile_X8Y7_to_ND),
    .to_NF(Tile_X8Y7_to_NF),
    .to_NG(Tile_X8Y7_to_NG),
    .to_NH(Tile_X8Y7_to_NH),
    .to_NI(Tile_X8Y7_to_NI),
    .to_SA(Tile_X8Y7_to_SA),
    .to_SB(Tile_X8Y7_to_SB),
    .to_SC(Tile_X8Y7_to_SC),
    .to_SD(Tile_X8Y7_to_SD),
    .to_SF(Tile_X8Y7_to_SF),
    .to_SG(Tile_X8Y7_to_SG),
    .to_SH(Tile_X8Y7_to_SH),
    .to_SI(Tile_X8Y7_to_SI),
    .UserCLK(Tile_X8Y8_UserCLKo),
    .UserCLKo(Tile_X8Y7_UserCLKo),
    .rst(Tile_X8Y8_rsto),
    .rsto(Tile_X8Y7_rsto),
    .FrameData(Tile_X7Y7_FrameData_O),
    .FrameData_O(Tile_X8Y7_FrameData_O),
    .FrameStrobe(Tile_X8Y8_FrameStrobe_O),
    .FrameStrobe_O(Tile_X8Y7_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
combined_WDDL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X9Y7_Emulate_Bitstream)
    )
`endif
    Tile_X9Y7_combined_WDDL
    (
    .from_NA_1s(Tile_X9Y8_to_NA_1s),
    .from_NB_1s(Tile_X9Y8_to_NB_1s),
    .from_NC_1s(Tile_X9Y8_to_NC_1s),
    .from_ND_1s(Tile_X9Y8_to_ND_1s),
    .from_NF_1s(Tile_X9Y8_to_NF_1s),
    .from_NG_1s(Tile_X9Y8_to_NG_1s),
    .from_NH_1s(Tile_X9Y8_to_NH_1s),
    .from_NI_1s(Tile_X9Y8_to_NI_1s),
    .from_SA_1s(Tile_X9Y6_to_SA_1s),
    .from_SB_1s(Tile_X9Y6_to_SB_1s),
    .from_SC_1s(Tile_X9Y6_to_SC_1s),
    .from_SD_1s(Tile_X9Y6_to_SD_1s),
    .from_SF_1s(Tile_X9Y6_to_SF_1s),
    .from_SG_1s(Tile_X9Y6_to_SG_1s),
    .from_SH_1s(Tile_X9Y6_to_SH_1s),
    .from_SI_1s(Tile_X9Y6_to_SI_1s),
    .from_WA_1s(Tile_X10Y7_to_WA_1s),
    .from_WB_1s(Tile_X10Y7_to_WB_1s),
    .from_WC_1s(Tile_X10Y7_to_WC_1s),
    .from_WD_1s(Tile_X10Y7_to_WD_1s),
    .from_WF_1s(Tile_X10Y7_to_WF_1s),
    .from_WG_1s(Tile_X10Y7_to_WG_1s),
    .from_WH_1s(Tile_X10Y7_to_WH_1s),
    .from_WI_1s(Tile_X10Y7_to_WI_1s),
    .to_EA_1s(Tile_X9Y7_to_EA_1s),
    .to_EB_1s(Tile_X9Y7_to_EB_1s),
    .to_EC_1s(Tile_X9Y7_to_EC_1s),
    .to_ED_1s(Tile_X9Y7_to_ED_1s),
    .to_EF_1s(Tile_X9Y7_to_EF_1s),
    .to_EG_1s(Tile_X9Y7_to_EG_1s),
    .to_EH_1s(Tile_X9Y7_to_EH_1s),
    .to_EI_1s(Tile_X9Y7_to_EI_1s),
    .to_WA_1s(Tile_X9Y7_to_WA_1s),
    .to_WB_1s(Tile_X9Y7_to_WB_1s),
    .to_WC_1s(Tile_X9Y7_to_WC_1s),
    .to_WD_1s(Tile_X9Y7_to_WD_1s),
    .to_WF_1s(Tile_X9Y7_to_WF_1s),
    .to_WG_1s(Tile_X9Y7_to_WG_1s),
    .to_WH_1s(Tile_X9Y7_to_WH_1s),
    .to_WI_1s(Tile_X9Y7_to_WI_1s),
    .to_NA_1s(Tile_X9Y7_to_NA_1s),
    .to_NB_1s(Tile_X9Y7_to_NB_1s),
    .to_NC_1s(Tile_X9Y7_to_NC_1s),
    .to_ND_1s(Tile_X9Y7_to_ND_1s),
    .to_NF_1s(Tile_X9Y7_to_NF_1s),
    .to_NG_1s(Tile_X9Y7_to_NG_1s),
    .to_NH_1s(Tile_X9Y7_to_NH_1s),
    .to_NI_1s(Tile_X9Y7_to_NI_1s),
    .to_SA_1s(Tile_X9Y7_to_SA_1s),
    .to_SB_1s(Tile_X9Y7_to_SB_1s),
    .to_SC_1s(Tile_X9Y7_to_SC_1s),
    .to_SD_1s(Tile_X9Y7_to_SD_1s),
    .to_SF_1s(Tile_X9Y7_to_SF_1s),
    .to_SG_1s(Tile_X9Y7_to_SG_1s),
    .to_SH_1s(Tile_X9Y7_to_SH_1s),
    .to_SI_1s(Tile_X9Y7_to_SI_1s),
    .F_ctrl(Tile_X9Y7_F_ctrl),
    .UserCLK(Tile_X9Y8_UserCLKo),
    .UserCLKo(Tile_X9Y7_UserCLKo),
    .rst(Tile_X9Y8_rsto),
    .rsto(Tile_X9Y7_rsto),
    .FrameData(Tile_X8Y7_FrameData_O),
    .FrameData_O(Tile_X9Y7_FrameData_O),
    .FrameStrobe(Tile_X9Y8_FrameStrobe_O),
    .FrameStrobe_O(Tile_X9Y7_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
ctrl_IO
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X10Y7_Emulate_Bitstream)
    )
`endif
    Tile_X10Y7_ctrl_IO
    (
    .from_EA_1s(Tile_X9Y7_to_EA_1s),
    .from_EB_1s(Tile_X9Y7_to_EB_1s),
    .from_EC_1s(Tile_X9Y7_to_EC_1s),
    .from_ED_1s(Tile_X9Y7_to_ED_1s),
    .from_EF_1s(Tile_X9Y7_to_EF_1s),
    .from_EG_1s(Tile_X9Y7_to_EG_1s),
    .from_EH_1s(Tile_X9Y7_to_EH_1s),
    .from_EI_1s(Tile_X9Y7_to_EI_1s),
    .to_WA_1s(Tile_X10Y7_to_WA_1s),
    .to_WB_1s(Tile_X10Y7_to_WB_1s),
    .to_WC_1s(Tile_X10Y7_to_WC_1s),
    .to_WD_1s(Tile_X10Y7_to_WD_1s),
    .to_WF_1s(Tile_X10Y7_to_WF_1s),
    .to_WG_1s(Tile_X10Y7_to_WG_1s),
    .to_WH_1s(Tile_X10Y7_to_WH_1s),
    .to_WI_1s(Tile_X10Y7_to_WI_1s),
    .A_O_top_0_t(Tile_X10Y7_A_O_top_0_t),
    .A_O_top_0_f(Tile_X10Y7_A_O_top_0_f),
    .A_prech2(Tile_X10Y7_A_prech2),
    .A_DR_fault(Tile_X10Y7_A_DR_fault),
    .A_I_top_0_t(Tile_X10Y7_A_I_top_0_t),
    .A_I_top_0_f(Tile_X10Y7_A_I_top_0_f),
    .A_T_top(Tile_X10Y7_A_T_top),
    .A_F_ctrl(Tile_X10Y7_A_F_ctrl),
    .UserCLK(Tile_X10Y8_UserCLKo),
    .UserCLKo(Tile_X10Y7_UserCLKo),
    .rst(Tile_X10Y8_rsto),
    .rsto(Tile_X10Y7_rsto),
    .FrameData(Tile_X9Y7_FrameData_O),
    .FrameData_O(Tile_X10Y7_FrameData_O),
    .FrameStrobe(Tile_X10Y8_FrameStrobe_O),
    .FrameStrobe_O(Tile_X10Y7_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
W_IO_custom
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X0Y8_Emulate_Bitstream)
    )
`endif
    Tile_X0Y8_W_IO_custom
    (
    .from_NA(Tile_X0Y9_to_NA),
    .from_NB(Tile_X0Y9_to_NB),
    .from_NC(Tile_X0Y9_to_NC),
    .from_ND(Tile_X0Y9_to_ND),
    .from_NF(Tile_X0Y9_to_NF),
    .from_NG(Tile_X0Y9_to_NG),
    .from_NH(Tile_X0Y9_to_NH),
    .from_NI(Tile_X0Y9_to_NI),
    .from_SA(Tile_X0Y7_to_SA),
    .from_SB(Tile_X0Y7_to_SB),
    .from_SC(Tile_X0Y7_to_SC),
    .from_SD(Tile_X0Y7_to_SD),
    .from_SF(Tile_X0Y7_to_SF),
    .from_SG(Tile_X0Y7_to_SG),
    .from_SH(Tile_X0Y7_to_SH),
    .from_SI(Tile_X0Y7_to_SI),
    .from_WA(Tile_X1Y8_to_WA),
    .from_WB(Tile_X1Y8_to_WB),
    .from_WC(Tile_X1Y8_to_WC),
    .from_WD(Tile_X1Y8_to_WD),
    .from_WF(Tile_X1Y8_to_WF),
    .from_WG(Tile_X1Y8_to_WG),
    .from_WH(Tile_X1Y8_to_WH),
    .from_WI(Tile_X1Y8_to_WI),
    .to_EA(Tile_X0Y8_to_EA),
    .to_EB(Tile_X0Y8_to_EB),
    .to_EC(Tile_X0Y8_to_EC),
    .to_ED(Tile_X0Y8_to_ED),
    .to_EF(Tile_X0Y8_to_EF),
    .to_EG(Tile_X0Y8_to_EG),
    .to_EH(Tile_X0Y8_to_EH),
    .to_EI(Tile_X0Y8_to_EI),
    .to_NA(Tile_X0Y8_to_NA),
    .to_NB(Tile_X0Y8_to_NB),
    .to_NC(Tile_X0Y8_to_NC),
    .to_ND(Tile_X0Y8_to_ND),
    .to_NF(Tile_X0Y8_to_NF),
    .to_NG(Tile_X0Y8_to_NG),
    .to_NH(Tile_X0Y8_to_NH),
    .to_NI(Tile_X0Y8_to_NI),
    .to_SA(Tile_X0Y8_to_SA),
    .to_SB(Tile_X0Y8_to_SB),
    .to_SC(Tile_X0Y8_to_SC),
    .to_SD(Tile_X0Y8_to_SD),
    .to_SF(Tile_X0Y8_to_SF),
    .to_SG(Tile_X0Y8_to_SG),
    .to_SH(Tile_X0Y8_to_SH),
    .to_SI(Tile_X0Y8_to_SI),
    .A_O_top_0_t(Tile_X0Y8_A_O_top_0_t),
    .A_O_top_0_f(Tile_X0Y8_A_O_top_0_f),
    .A_O_top_1_t(Tile_X0Y8_A_O_top_1_t),
    .A_O_top_1_f(Tile_X0Y8_A_O_top_1_f),
    .A_prech1(Tile_X0Y8_A_prech1),
    .A_prech2(Tile_X0Y8_A_prech2),
    .A_DR_fault(Tile_X0Y8_A_DR_fault),
    .A_I_top_0_t(Tile_X0Y8_A_I_top_0_t),
    .A_I_top_0_f(Tile_X0Y8_A_I_top_0_f),
    .A_I_top_1_t(Tile_X0Y8_A_I_top_1_t),
    .A_I_top_1_f(Tile_X0Y8_A_I_top_1_f),
    .A_T_top(Tile_X0Y8_A_T_top),
    .A_F_masked1(Tile_X0Y8_A_F_masked1),
    .A_F_masked2(Tile_X0Y8_A_F_masked2),
    .A_config_C_bit0(Tile_X0Y8_A_config_C_bit0),
    .A_config_C_bit1(Tile_X0Y8_A_config_C_bit1),
    .A_config_C_bit2(Tile_X0Y8_A_config_C_bit2),
    .A_config_C_bit3(Tile_X0Y8_A_config_C_bit3),
    .B_config_C_bit0(Tile_X0Y8_B_config_C_bit0),
    .B_config_C_bit1(Tile_X0Y8_B_config_C_bit1),
    .B_config_C_bit2(Tile_X0Y8_B_config_C_bit2),
    .B_config_C_bit3(Tile_X0Y8_B_config_C_bit3),
    .UserCLK(Tile_X0Y9_UserCLKo),
    .UserCLKo(Tile_X0Y8_UserCLKo),
    .rst(Tile_X0Y9_rsto),
    .rsto(Tile_X0Y8_rsto),
    .FrameData(Tile_Y8_FrameData),
    .FrameData_O(Tile_X0Y8_FrameData_O),
    .FrameStrobe(Tile_X0Y9_FrameStrobe_O),
    .FrameStrobe_O(Tile_X0Y8_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X1Y8_Emulate_Bitstream)
    )
`endif
    Tile_X1Y8_linear_LMDPL
    (
    .from_NA(Tile_X1Y9_to_NA),
    .from_NB(Tile_X1Y9_to_NB),
    .from_NC(Tile_X1Y9_to_NC),
    .from_ND(Tile_X1Y9_to_ND),
    .from_NF(Tile_X1Y9_to_NF),
    .from_NG(Tile_X1Y9_to_NG),
    .from_NH(Tile_X1Y9_to_NH),
    .from_NI(Tile_X1Y9_to_NI),
    .from_EA(Tile_X0Y8_to_EA),
    .from_EB(Tile_X0Y8_to_EB),
    .from_EC(Tile_X0Y8_to_EC),
    .from_ED(Tile_X0Y8_to_ED),
    .from_EF(Tile_X0Y8_to_EF),
    .from_EG(Tile_X0Y8_to_EG),
    .from_EH(Tile_X0Y8_to_EH),
    .from_EI(Tile_X0Y8_to_EI),
    .from_SA(Tile_X1Y7_to_SA),
    .from_SB(Tile_X1Y7_to_SB),
    .from_SC(Tile_X1Y7_to_SC),
    .from_SD(Tile_X1Y7_to_SD),
    .from_SF(Tile_X1Y7_to_SF),
    .from_SG(Tile_X1Y7_to_SG),
    .from_SH(Tile_X1Y7_to_SH),
    .from_SI(Tile_X1Y7_to_SI),
    .from_WA(Tile_X2Y8_to_WA),
    .from_WB(Tile_X2Y8_to_WB),
    .from_WC(Tile_X2Y8_to_WC),
    .from_WD(Tile_X2Y8_to_WD),
    .from_WF(Tile_X2Y8_to_WF),
    .from_WG(Tile_X2Y8_to_WG),
    .from_WH(Tile_X2Y8_to_WH),
    .from_WI(Tile_X2Y8_to_WI),
    .to_EA(Tile_X1Y8_to_EA),
    .to_EB(Tile_X1Y8_to_EB),
    .to_EC(Tile_X1Y8_to_EC),
    .to_ED(Tile_X1Y8_to_ED),
    .to_EF(Tile_X1Y8_to_EF),
    .to_EG(Tile_X1Y8_to_EG),
    .to_EH(Tile_X1Y8_to_EH),
    .to_EI(Tile_X1Y8_to_EI),
    .to_WA(Tile_X1Y8_to_WA),
    .to_WB(Tile_X1Y8_to_WB),
    .to_WC(Tile_X1Y8_to_WC),
    .to_WD(Tile_X1Y8_to_WD),
    .to_WF(Tile_X1Y8_to_WF),
    .to_WG(Tile_X1Y8_to_WG),
    .to_WH(Tile_X1Y8_to_WH),
    .to_WI(Tile_X1Y8_to_WI),
    .to_NA(Tile_X1Y8_to_NA),
    .to_NB(Tile_X1Y8_to_NB),
    .to_NC(Tile_X1Y8_to_NC),
    .to_ND(Tile_X1Y8_to_ND),
    .to_NF(Tile_X1Y8_to_NF),
    .to_NG(Tile_X1Y8_to_NG),
    .to_NH(Tile_X1Y8_to_NH),
    .to_NI(Tile_X1Y8_to_NI),
    .to_SA(Tile_X1Y8_to_SA),
    .to_SB(Tile_X1Y8_to_SB),
    .to_SC(Tile_X1Y8_to_SC),
    .to_SD(Tile_X1Y8_to_SD),
    .to_SF(Tile_X1Y8_to_SF),
    .to_SG(Tile_X1Y8_to_SG),
    .to_SH(Tile_X1Y8_to_SH),
    .to_SI(Tile_X1Y8_to_SI),
    .F_masked1(Tile_X1Y8_F_masked1),
    .F_masked2(Tile_X1Y8_F_masked2),
    .UserCLK(Tile_X1Y9_UserCLKo),
    .UserCLKo(Tile_X1Y8_UserCLKo),
    .rst(Tile_X1Y9_rsto),
    .rsto(Tile_X1Y8_rsto),
    .FrameData(Tile_X0Y8_FrameData_O),
    .FrameData_O(Tile_X1Y8_FrameData_O),
    .FrameStrobe(Tile_X1Y9_FrameStrobe_O),
    .FrameStrobe_O(Tile_X1Y8_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X2Y8_Emulate_Bitstream)
    )
`endif
    Tile_X2Y8_linear_LMDPL
    (
    .from_NA(Tile_X2Y9_to_NA),
    .from_NB(Tile_X2Y9_to_NB),
    .from_NC(Tile_X2Y9_to_NC),
    .from_ND(Tile_X2Y9_to_ND),
    .from_NF(Tile_X2Y9_to_NF),
    .from_NG(Tile_X2Y9_to_NG),
    .from_NH(Tile_X2Y9_to_NH),
    .from_NI(Tile_X2Y9_to_NI),
    .from_EA(Tile_X1Y8_to_EA),
    .from_EB(Tile_X1Y8_to_EB),
    .from_EC(Tile_X1Y8_to_EC),
    .from_ED(Tile_X1Y8_to_ED),
    .from_EF(Tile_X1Y8_to_EF),
    .from_EG(Tile_X1Y8_to_EG),
    .from_EH(Tile_X1Y8_to_EH),
    .from_EI(Tile_X1Y8_to_EI),
    .from_SA(Tile_X2Y7_to_SA),
    .from_SB(Tile_X2Y7_to_SB),
    .from_SC(Tile_X2Y7_to_SC),
    .from_SD(Tile_X2Y7_to_SD),
    .from_SF(Tile_X2Y7_to_SF),
    .from_SG(Tile_X2Y7_to_SG),
    .from_SH(Tile_X2Y7_to_SH),
    .from_SI(Tile_X2Y7_to_SI),
    .from_WA(Tile_X3Y8_to_WA),
    .from_WB(Tile_X3Y8_to_WB),
    .from_WC(Tile_X3Y8_to_WC),
    .from_WD(Tile_X3Y8_to_WD),
    .from_WF(Tile_X3Y8_to_WF),
    .from_WG(Tile_X3Y8_to_WG),
    .from_WH(Tile_X3Y8_to_WH),
    .from_WI(Tile_X3Y8_to_WI),
    .to_EA(Tile_X2Y8_to_EA),
    .to_EB(Tile_X2Y8_to_EB),
    .to_EC(Tile_X2Y8_to_EC),
    .to_ED(Tile_X2Y8_to_ED),
    .to_EF(Tile_X2Y8_to_EF),
    .to_EG(Tile_X2Y8_to_EG),
    .to_EH(Tile_X2Y8_to_EH),
    .to_EI(Tile_X2Y8_to_EI),
    .to_WA(Tile_X2Y8_to_WA),
    .to_WB(Tile_X2Y8_to_WB),
    .to_WC(Tile_X2Y8_to_WC),
    .to_WD(Tile_X2Y8_to_WD),
    .to_WF(Tile_X2Y8_to_WF),
    .to_WG(Tile_X2Y8_to_WG),
    .to_WH(Tile_X2Y8_to_WH),
    .to_WI(Tile_X2Y8_to_WI),
    .to_NA(Tile_X2Y8_to_NA),
    .to_NB(Tile_X2Y8_to_NB),
    .to_NC(Tile_X2Y8_to_NC),
    .to_ND(Tile_X2Y8_to_ND),
    .to_NF(Tile_X2Y8_to_NF),
    .to_NG(Tile_X2Y8_to_NG),
    .to_NH(Tile_X2Y8_to_NH),
    .to_NI(Tile_X2Y8_to_NI),
    .to_SA(Tile_X2Y8_to_SA),
    .to_SB(Tile_X2Y8_to_SB),
    .to_SC(Tile_X2Y8_to_SC),
    .to_SD(Tile_X2Y8_to_SD),
    .to_SF(Tile_X2Y8_to_SF),
    .to_SG(Tile_X2Y8_to_SG),
    .to_SH(Tile_X2Y8_to_SH),
    .to_SI(Tile_X2Y8_to_SI),
    .F_masked1(Tile_X2Y8_F_masked1),
    .F_masked2(Tile_X2Y8_F_masked2),
    .UserCLK(Tile_X2Y9_UserCLKo),
    .UserCLKo(Tile_X2Y8_UserCLKo),
    .rst(Tile_X2Y9_rsto),
    .rsto(Tile_X2Y8_rsto),
    .FrameData(Tile_X1Y8_FrameData_O),
    .FrameData_O(Tile_X2Y8_FrameData_O),
    .FrameStrobe(Tile_X2Y9_FrameStrobe_O),
    .FrameStrobe_O(Tile_X2Y8_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
nonlinear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X3Y8_Emulate_Bitstream)
    )
`endif
    Tile_X3Y8_nonlinear_LMDPL
    (
    .from_NA(Tile_X3Y9_to_NA),
    .from_NB(Tile_X3Y9_to_NB),
    .from_NC(Tile_X3Y9_to_NC),
    .from_ND(Tile_X3Y9_to_ND),
    .from_NF(Tile_X3Y9_to_NF),
    .from_NG(Tile_X3Y9_to_NG),
    .from_NH(Tile_X3Y9_to_NH),
    .from_NI(Tile_X3Y9_to_NI),
    .from_EA(Tile_X2Y8_to_EA),
    .from_EB(Tile_X2Y8_to_EB),
    .from_EC(Tile_X2Y8_to_EC),
    .from_ED(Tile_X2Y8_to_ED),
    .from_EF(Tile_X2Y8_to_EF),
    .from_EG(Tile_X2Y8_to_EG),
    .from_EH(Tile_X2Y8_to_EH),
    .from_EI(Tile_X2Y8_to_EI),
    .from_SA(Tile_X3Y7_to_SA),
    .from_SB(Tile_X3Y7_to_SB),
    .from_SC(Tile_X3Y7_to_SC),
    .from_SD(Tile_X3Y7_to_SD),
    .from_SF(Tile_X3Y7_to_SF),
    .from_SG(Tile_X3Y7_to_SG),
    .from_SH(Tile_X3Y7_to_SH),
    .from_SI(Tile_X3Y7_to_SI),
    .from_WA(Tile_X4Y8_to_WA),
    .from_WB(Tile_X4Y8_to_WB),
    .from_WC(Tile_X4Y8_to_WC),
    .from_WD(Tile_X4Y8_to_WD),
    .from_WF(Tile_X4Y8_to_WF),
    .from_WG(Tile_X4Y8_to_WG),
    .from_WH(Tile_X4Y8_to_WH),
    .from_WI(Tile_X4Y8_to_WI),
    .to_EA(Tile_X3Y8_to_EA),
    .to_EB(Tile_X3Y8_to_EB),
    .to_EC(Tile_X3Y8_to_EC),
    .to_ED(Tile_X3Y8_to_ED),
    .to_EF(Tile_X3Y8_to_EF),
    .to_EG(Tile_X3Y8_to_EG),
    .to_EH(Tile_X3Y8_to_EH),
    .to_EI(Tile_X3Y8_to_EI),
    .to_WA(Tile_X3Y8_to_WA),
    .to_WB(Tile_X3Y8_to_WB),
    .to_WC(Tile_X3Y8_to_WC),
    .to_WD(Tile_X3Y8_to_WD),
    .to_WF(Tile_X3Y8_to_WF),
    .to_WG(Tile_X3Y8_to_WG),
    .to_WH(Tile_X3Y8_to_WH),
    .to_WI(Tile_X3Y8_to_WI),
    .to_NA(Tile_X3Y8_to_NA),
    .to_NB(Tile_X3Y8_to_NB),
    .to_NC(Tile_X3Y8_to_NC),
    .to_ND(Tile_X3Y8_to_ND),
    .to_NF(Tile_X3Y8_to_NF),
    .to_NG(Tile_X3Y8_to_NG),
    .to_NH(Tile_X3Y8_to_NH),
    .to_NI(Tile_X3Y8_to_NI),
    .to_SA(Tile_X3Y8_to_SA),
    .to_SB(Tile_X3Y8_to_SB),
    .to_SC(Tile_X3Y8_to_SC),
    .to_SD(Tile_X3Y8_to_SD),
    .to_SF(Tile_X3Y8_to_SF),
    .to_SG(Tile_X3Y8_to_SG),
    .to_SH(Tile_X3Y8_to_SH),
    .to_SI(Tile_X3Y8_to_SI),
    .R_t(Tile_X3Y8_R_t),
    .R_f(Tile_X3Y8_R_f),
    .F_masked1(Tile_X3Y8_F_masked1),
    .F_masked2(Tile_X3Y8_F_masked2),
    .UserCLK(Tile_X3Y9_UserCLKo),
    .UserCLKo(Tile_X3Y8_UserCLKo),
    .rst(Tile_X3Y9_rsto),
    .rsto(Tile_X3Y8_rsto),
    .FrameData(Tile_X2Y8_FrameData_O),
    .FrameData_O(Tile_X3Y8_FrameData_O),
    .FrameStrobe(Tile_X3Y9_FrameStrobe_O),
    .FrameStrobe_O(Tile_X3Y8_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X4Y8_Emulate_Bitstream)
    )
`endif
    Tile_X4Y8_linear_LMDPL
    (
    .from_NA(Tile_X4Y9_to_NA),
    .from_NB(Tile_X4Y9_to_NB),
    .from_NC(Tile_X4Y9_to_NC),
    .from_ND(Tile_X4Y9_to_ND),
    .from_NF(Tile_X4Y9_to_NF),
    .from_NG(Tile_X4Y9_to_NG),
    .from_NH(Tile_X4Y9_to_NH),
    .from_NI(Tile_X4Y9_to_NI),
    .from_EA(Tile_X3Y8_to_EA),
    .from_EB(Tile_X3Y8_to_EB),
    .from_EC(Tile_X3Y8_to_EC),
    .from_ED(Tile_X3Y8_to_ED),
    .from_EF(Tile_X3Y8_to_EF),
    .from_EG(Tile_X3Y8_to_EG),
    .from_EH(Tile_X3Y8_to_EH),
    .from_EI(Tile_X3Y8_to_EI),
    .from_SA(Tile_X4Y7_to_SA),
    .from_SB(Tile_X4Y7_to_SB),
    .from_SC(Tile_X4Y7_to_SC),
    .from_SD(Tile_X4Y7_to_SD),
    .from_SF(Tile_X4Y7_to_SF),
    .from_SG(Tile_X4Y7_to_SG),
    .from_SH(Tile_X4Y7_to_SH),
    .from_SI(Tile_X4Y7_to_SI),
    .from_WA(Tile_X5Y8_to_WA),
    .from_WB(Tile_X5Y8_to_WB),
    .from_WC(Tile_X5Y8_to_WC),
    .from_WD(Tile_X5Y8_to_WD),
    .from_WF(Tile_X5Y8_to_WF),
    .from_WG(Tile_X5Y8_to_WG),
    .from_WH(Tile_X5Y8_to_WH),
    .from_WI(Tile_X5Y8_to_WI),
    .to_EA(Tile_X4Y8_to_EA),
    .to_EB(Tile_X4Y8_to_EB),
    .to_EC(Tile_X4Y8_to_EC),
    .to_ED(Tile_X4Y8_to_ED),
    .to_EF(Tile_X4Y8_to_EF),
    .to_EG(Tile_X4Y8_to_EG),
    .to_EH(Tile_X4Y8_to_EH),
    .to_EI(Tile_X4Y8_to_EI),
    .to_WA(Tile_X4Y8_to_WA),
    .to_WB(Tile_X4Y8_to_WB),
    .to_WC(Tile_X4Y8_to_WC),
    .to_WD(Tile_X4Y8_to_WD),
    .to_WF(Tile_X4Y8_to_WF),
    .to_WG(Tile_X4Y8_to_WG),
    .to_WH(Tile_X4Y8_to_WH),
    .to_WI(Tile_X4Y8_to_WI),
    .to_NA(Tile_X4Y8_to_NA),
    .to_NB(Tile_X4Y8_to_NB),
    .to_NC(Tile_X4Y8_to_NC),
    .to_ND(Tile_X4Y8_to_ND),
    .to_NF(Tile_X4Y8_to_NF),
    .to_NG(Tile_X4Y8_to_NG),
    .to_NH(Tile_X4Y8_to_NH),
    .to_NI(Tile_X4Y8_to_NI),
    .to_SA(Tile_X4Y8_to_SA),
    .to_SB(Tile_X4Y8_to_SB),
    .to_SC(Tile_X4Y8_to_SC),
    .to_SD(Tile_X4Y8_to_SD),
    .to_SF(Tile_X4Y8_to_SF),
    .to_SG(Tile_X4Y8_to_SG),
    .to_SH(Tile_X4Y8_to_SH),
    .to_SI(Tile_X4Y8_to_SI),
    .F_masked1(Tile_X4Y8_F_masked1),
    .F_masked2(Tile_X4Y8_F_masked2),
    .UserCLK(Tile_X4Y9_UserCLKo),
    .UserCLKo(Tile_X4Y8_UserCLKo),
    .rst(Tile_X4Y9_rsto),
    .rsto(Tile_X4Y8_rsto),
    .FrameData(Tile_X3Y8_FrameData_O),
    .FrameData_O(Tile_X4Y8_FrameData_O),
    .FrameStrobe(Tile_X4Y9_FrameStrobe_O),
    .FrameStrobe_O(Tile_X4Y8_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X5Y8_Emulate_Bitstream)
    )
`endif
    Tile_X5Y8_linear_LMDPL
    (
    .from_NA(Tile_X5Y9_to_NA),
    .from_NB(Tile_X5Y9_to_NB),
    .from_NC(Tile_X5Y9_to_NC),
    .from_ND(Tile_X5Y9_to_ND),
    .from_NF(Tile_X5Y9_to_NF),
    .from_NG(Tile_X5Y9_to_NG),
    .from_NH(Tile_X5Y9_to_NH),
    .from_NI(Tile_X5Y9_to_NI),
    .from_EA(Tile_X4Y8_to_EA),
    .from_EB(Tile_X4Y8_to_EB),
    .from_EC(Tile_X4Y8_to_EC),
    .from_ED(Tile_X4Y8_to_ED),
    .from_EF(Tile_X4Y8_to_EF),
    .from_EG(Tile_X4Y8_to_EG),
    .from_EH(Tile_X4Y8_to_EH),
    .from_EI(Tile_X4Y8_to_EI),
    .from_SA(Tile_X5Y7_to_SA),
    .from_SB(Tile_X5Y7_to_SB),
    .from_SC(Tile_X5Y7_to_SC),
    .from_SD(Tile_X5Y7_to_SD),
    .from_SF(Tile_X5Y7_to_SF),
    .from_SG(Tile_X5Y7_to_SG),
    .from_SH(Tile_X5Y7_to_SH),
    .from_SI(Tile_X5Y7_to_SI),
    .from_WA(Tile_X6Y8_to_WA),
    .from_WB(Tile_X6Y8_to_WB),
    .from_WC(Tile_X6Y8_to_WC),
    .from_WD(Tile_X6Y8_to_WD),
    .from_WF(Tile_X6Y8_to_WF),
    .from_WG(Tile_X6Y8_to_WG),
    .from_WH(Tile_X6Y8_to_WH),
    .from_WI(Tile_X6Y8_to_WI),
    .to_EA(Tile_X5Y8_to_EA),
    .to_EB(Tile_X5Y8_to_EB),
    .to_EC(Tile_X5Y8_to_EC),
    .to_ED(Tile_X5Y8_to_ED),
    .to_EF(Tile_X5Y8_to_EF),
    .to_EG(Tile_X5Y8_to_EG),
    .to_EH(Tile_X5Y8_to_EH),
    .to_EI(Tile_X5Y8_to_EI),
    .to_WA(Tile_X5Y8_to_WA),
    .to_WB(Tile_X5Y8_to_WB),
    .to_WC(Tile_X5Y8_to_WC),
    .to_WD(Tile_X5Y8_to_WD),
    .to_WF(Tile_X5Y8_to_WF),
    .to_WG(Tile_X5Y8_to_WG),
    .to_WH(Tile_X5Y8_to_WH),
    .to_WI(Tile_X5Y8_to_WI),
    .to_NA(Tile_X5Y8_to_NA),
    .to_NB(Tile_X5Y8_to_NB),
    .to_NC(Tile_X5Y8_to_NC),
    .to_ND(Tile_X5Y8_to_ND),
    .to_NF(Tile_X5Y8_to_NF),
    .to_NG(Tile_X5Y8_to_NG),
    .to_NH(Tile_X5Y8_to_NH),
    .to_NI(Tile_X5Y8_to_NI),
    .to_SA(Tile_X5Y8_to_SA),
    .to_SB(Tile_X5Y8_to_SB),
    .to_SC(Tile_X5Y8_to_SC),
    .to_SD(Tile_X5Y8_to_SD),
    .to_SF(Tile_X5Y8_to_SF),
    .to_SG(Tile_X5Y8_to_SG),
    .to_SH(Tile_X5Y8_to_SH),
    .to_SI(Tile_X5Y8_to_SI),
    .F_masked1(Tile_X5Y8_F_masked1),
    .F_masked2(Tile_X5Y8_F_masked2),
    .UserCLK(Tile_X5Y9_UserCLKo),
    .UserCLKo(Tile_X5Y8_UserCLKo),
    .rst(Tile_X5Y9_rsto),
    .rsto(Tile_X5Y8_rsto),
    .FrameData(Tile_X4Y8_FrameData_O),
    .FrameData_O(Tile_X5Y8_FrameData_O),
    .FrameStrobe(Tile_X5Y9_FrameStrobe_O),
    .FrameStrobe_O(Tile_X5Y8_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
nonlinear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X6Y8_Emulate_Bitstream)
    )
`endif
    Tile_X6Y8_nonlinear_LMDPL
    (
    .from_NA(Tile_X6Y9_to_NA),
    .from_NB(Tile_X6Y9_to_NB),
    .from_NC(Tile_X6Y9_to_NC),
    .from_ND(Tile_X6Y9_to_ND),
    .from_NF(Tile_X6Y9_to_NF),
    .from_NG(Tile_X6Y9_to_NG),
    .from_NH(Tile_X6Y9_to_NH),
    .from_NI(Tile_X6Y9_to_NI),
    .from_EA(Tile_X5Y8_to_EA),
    .from_EB(Tile_X5Y8_to_EB),
    .from_EC(Tile_X5Y8_to_EC),
    .from_ED(Tile_X5Y8_to_ED),
    .from_EF(Tile_X5Y8_to_EF),
    .from_EG(Tile_X5Y8_to_EG),
    .from_EH(Tile_X5Y8_to_EH),
    .from_EI(Tile_X5Y8_to_EI),
    .from_SA(Tile_X6Y7_to_SA),
    .from_SB(Tile_X6Y7_to_SB),
    .from_SC(Tile_X6Y7_to_SC),
    .from_SD(Tile_X6Y7_to_SD),
    .from_SF(Tile_X6Y7_to_SF),
    .from_SG(Tile_X6Y7_to_SG),
    .from_SH(Tile_X6Y7_to_SH),
    .from_SI(Tile_X6Y7_to_SI),
    .from_WA(Tile_X7Y8_to_WA),
    .from_WB(Tile_X7Y8_to_WB),
    .from_WC(Tile_X7Y8_to_WC),
    .from_WD(Tile_X7Y8_to_WD),
    .from_WF(Tile_X7Y8_to_WF),
    .from_WG(Tile_X7Y8_to_WG),
    .from_WH(Tile_X7Y8_to_WH),
    .from_WI(Tile_X7Y8_to_WI),
    .to_EA(Tile_X6Y8_to_EA),
    .to_EB(Tile_X6Y8_to_EB),
    .to_EC(Tile_X6Y8_to_EC),
    .to_ED(Tile_X6Y8_to_ED),
    .to_EF(Tile_X6Y8_to_EF),
    .to_EG(Tile_X6Y8_to_EG),
    .to_EH(Tile_X6Y8_to_EH),
    .to_EI(Tile_X6Y8_to_EI),
    .to_WA(Tile_X6Y8_to_WA),
    .to_WB(Tile_X6Y8_to_WB),
    .to_WC(Tile_X6Y8_to_WC),
    .to_WD(Tile_X6Y8_to_WD),
    .to_WF(Tile_X6Y8_to_WF),
    .to_WG(Tile_X6Y8_to_WG),
    .to_WH(Tile_X6Y8_to_WH),
    .to_WI(Tile_X6Y8_to_WI),
    .to_NA(Tile_X6Y8_to_NA),
    .to_NB(Tile_X6Y8_to_NB),
    .to_NC(Tile_X6Y8_to_NC),
    .to_ND(Tile_X6Y8_to_ND),
    .to_NF(Tile_X6Y8_to_NF),
    .to_NG(Tile_X6Y8_to_NG),
    .to_NH(Tile_X6Y8_to_NH),
    .to_NI(Tile_X6Y8_to_NI),
    .to_SA(Tile_X6Y8_to_SA),
    .to_SB(Tile_X6Y8_to_SB),
    .to_SC(Tile_X6Y8_to_SC),
    .to_SD(Tile_X6Y8_to_SD),
    .to_SF(Tile_X6Y8_to_SF),
    .to_SG(Tile_X6Y8_to_SG),
    .to_SH(Tile_X6Y8_to_SH),
    .to_SI(Tile_X6Y8_to_SI),
    .R_t(Tile_X6Y8_R_t),
    .R_f(Tile_X6Y8_R_f),
    .F_masked1(Tile_X6Y8_F_masked1),
    .F_masked2(Tile_X6Y8_F_masked2),
    .UserCLK(Tile_X6Y9_UserCLKo),
    .UserCLKo(Tile_X6Y8_UserCLKo),
    .rst(Tile_X6Y9_rsto),
    .rsto(Tile_X6Y8_rsto),
    .FrameData(Tile_X5Y8_FrameData_O),
    .FrameData_O(Tile_X6Y8_FrameData_O),
    .FrameStrobe(Tile_X6Y9_FrameStrobe_O),
    .FrameStrobe_O(Tile_X6Y8_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X7Y8_Emulate_Bitstream)
    )
`endif
    Tile_X7Y8_linear_LMDPL
    (
    .from_NA(Tile_X7Y9_to_NA),
    .from_NB(Tile_X7Y9_to_NB),
    .from_NC(Tile_X7Y9_to_NC),
    .from_ND(Tile_X7Y9_to_ND),
    .from_NF(Tile_X7Y9_to_NF),
    .from_NG(Tile_X7Y9_to_NG),
    .from_NH(Tile_X7Y9_to_NH),
    .from_NI(Tile_X7Y9_to_NI),
    .from_EA(Tile_X6Y8_to_EA),
    .from_EB(Tile_X6Y8_to_EB),
    .from_EC(Tile_X6Y8_to_EC),
    .from_ED(Tile_X6Y8_to_ED),
    .from_EF(Tile_X6Y8_to_EF),
    .from_EG(Tile_X6Y8_to_EG),
    .from_EH(Tile_X6Y8_to_EH),
    .from_EI(Tile_X6Y8_to_EI),
    .from_SA(Tile_X7Y7_to_SA),
    .from_SB(Tile_X7Y7_to_SB),
    .from_SC(Tile_X7Y7_to_SC),
    .from_SD(Tile_X7Y7_to_SD),
    .from_SF(Tile_X7Y7_to_SF),
    .from_SG(Tile_X7Y7_to_SG),
    .from_SH(Tile_X7Y7_to_SH),
    .from_SI(Tile_X7Y7_to_SI),
    .from_WA(Tile_X8Y8_to_WA),
    .from_WB(Tile_X8Y8_to_WB),
    .from_WC(Tile_X8Y8_to_WC),
    .from_WD(Tile_X8Y8_to_WD),
    .from_WF(Tile_X8Y8_to_WF),
    .from_WG(Tile_X8Y8_to_WG),
    .from_WH(Tile_X8Y8_to_WH),
    .from_WI(Tile_X8Y8_to_WI),
    .to_EA(Tile_X7Y8_to_EA),
    .to_EB(Tile_X7Y8_to_EB),
    .to_EC(Tile_X7Y8_to_EC),
    .to_ED(Tile_X7Y8_to_ED),
    .to_EF(Tile_X7Y8_to_EF),
    .to_EG(Tile_X7Y8_to_EG),
    .to_EH(Tile_X7Y8_to_EH),
    .to_EI(Tile_X7Y8_to_EI),
    .to_WA(Tile_X7Y8_to_WA),
    .to_WB(Tile_X7Y8_to_WB),
    .to_WC(Tile_X7Y8_to_WC),
    .to_WD(Tile_X7Y8_to_WD),
    .to_WF(Tile_X7Y8_to_WF),
    .to_WG(Tile_X7Y8_to_WG),
    .to_WH(Tile_X7Y8_to_WH),
    .to_WI(Tile_X7Y8_to_WI),
    .to_NA(Tile_X7Y8_to_NA),
    .to_NB(Tile_X7Y8_to_NB),
    .to_NC(Tile_X7Y8_to_NC),
    .to_ND(Tile_X7Y8_to_ND),
    .to_NF(Tile_X7Y8_to_NF),
    .to_NG(Tile_X7Y8_to_NG),
    .to_NH(Tile_X7Y8_to_NH),
    .to_NI(Tile_X7Y8_to_NI),
    .to_SA(Tile_X7Y8_to_SA),
    .to_SB(Tile_X7Y8_to_SB),
    .to_SC(Tile_X7Y8_to_SC),
    .to_SD(Tile_X7Y8_to_SD),
    .to_SF(Tile_X7Y8_to_SF),
    .to_SG(Tile_X7Y8_to_SG),
    .to_SH(Tile_X7Y8_to_SH),
    .to_SI(Tile_X7Y8_to_SI),
    .F_masked1(Tile_X7Y8_F_masked1),
    .F_masked2(Tile_X7Y8_F_masked2),
    .UserCLK(Tile_X7Y9_UserCLKo),
    .UserCLKo(Tile_X7Y8_UserCLKo),
    .rst(Tile_X7Y9_rsto),
    .rsto(Tile_X7Y8_rsto),
    .FrameData(Tile_X6Y8_FrameData_O),
    .FrameData_O(Tile_X7Y8_FrameData_O),
    .FrameStrobe(Tile_X7Y9_FrameStrobe_O),
    .FrameStrobe_O(Tile_X7Y8_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
ctrl_to_sec
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X8Y8_Emulate_Bitstream)
    )
`endif
    Tile_X8Y8_ctrl_to_sec
    (
    .from_NA(Tile_X8Y9_to_NA),
    .from_NB(Tile_X8Y9_to_NB),
    .from_NC(Tile_X8Y9_to_NC),
    .from_ND(Tile_X8Y9_to_ND),
    .from_NF(Tile_X8Y9_to_NF),
    .from_NG(Tile_X8Y9_to_NG),
    .from_NH(Tile_X8Y9_to_NH),
    .from_NI(Tile_X8Y9_to_NI),
    .from_EA(Tile_X7Y8_to_EA),
    .from_EB(Tile_X7Y8_to_EB),
    .from_EC(Tile_X7Y8_to_EC),
    .from_ED(Tile_X7Y8_to_ED),
    .from_EF(Tile_X7Y8_to_EF),
    .from_EG(Tile_X7Y8_to_EG),
    .from_EH(Tile_X7Y8_to_EH),
    .from_EI(Tile_X7Y8_to_EI),
    .from_SA(Tile_X8Y7_to_SA),
    .from_SB(Tile_X8Y7_to_SB),
    .from_SC(Tile_X8Y7_to_SC),
    .from_SD(Tile_X8Y7_to_SD),
    .from_SF(Tile_X8Y7_to_SF),
    .from_SG(Tile_X8Y7_to_SG),
    .from_SH(Tile_X8Y7_to_SH),
    .from_SI(Tile_X8Y7_to_SI),
    .from_WA_1s(Tile_X9Y8_to_WA_1s),
    .from_WB_1s(Tile_X9Y8_to_WB_1s),
    .from_WC_1s(Tile_X9Y8_to_WC_1s),
    .from_WD_1s(Tile_X9Y8_to_WD_1s),
    .from_WF_1s(Tile_X9Y8_to_WF_1s),
    .from_WG_1s(Tile_X9Y8_to_WG_1s),
    .from_WH_1s(Tile_X9Y8_to_WH_1s),
    .from_WI_1s(Tile_X9Y8_to_WI_1s),
    .to_WA(Tile_X8Y8_to_WA),
    .to_WB(Tile_X8Y8_to_WB),
    .to_WC(Tile_X8Y8_to_WC),
    .to_WD(Tile_X8Y8_to_WD),
    .to_WF(Tile_X8Y8_to_WF),
    .to_WG(Tile_X8Y8_to_WG),
    .to_WH(Tile_X8Y8_to_WH),
    .to_WI(Tile_X8Y8_to_WI),
    .to_NA(Tile_X8Y8_to_NA),
    .to_NB(Tile_X8Y8_to_NB),
    .to_NC(Tile_X8Y8_to_NC),
    .to_ND(Tile_X8Y8_to_ND),
    .to_NF(Tile_X8Y8_to_NF),
    .to_NG(Tile_X8Y8_to_NG),
    .to_NH(Tile_X8Y8_to_NH),
    .to_NI(Tile_X8Y8_to_NI),
    .to_SA(Tile_X8Y8_to_SA),
    .to_SB(Tile_X8Y8_to_SB),
    .to_SC(Tile_X8Y8_to_SC),
    .to_SD(Tile_X8Y8_to_SD),
    .to_SF(Tile_X8Y8_to_SF),
    .to_SG(Tile_X8Y8_to_SG),
    .to_SH(Tile_X8Y8_to_SH),
    .to_SI(Tile_X8Y8_to_SI),
    .UserCLK(Tile_X8Y9_UserCLKo),
    .UserCLKo(Tile_X8Y8_UserCLKo),
    .rst(Tile_X8Y9_rsto),
    .rsto(Tile_X8Y8_rsto),
    .FrameData(Tile_X7Y8_FrameData_O),
    .FrameData_O(Tile_X8Y8_FrameData_O),
    .FrameStrobe(Tile_X8Y9_FrameStrobe_O),
    .FrameStrobe_O(Tile_X8Y8_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
combined_WDDL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X9Y8_Emulate_Bitstream)
    )
`endif
    Tile_X9Y8_combined_WDDL
    (
    .from_NA_1s(Tile_X9Y9_to_NA_1s),
    .from_NB_1s(Tile_X9Y9_to_NB_1s),
    .from_NC_1s(Tile_X9Y9_to_NC_1s),
    .from_ND_1s(Tile_X9Y9_to_ND_1s),
    .from_NF_1s(Tile_X9Y9_to_NF_1s),
    .from_NG_1s(Tile_X9Y9_to_NG_1s),
    .from_NH_1s(Tile_X9Y9_to_NH_1s),
    .from_NI_1s(Tile_X9Y9_to_NI_1s),
    .from_SA_1s(Tile_X9Y7_to_SA_1s),
    .from_SB_1s(Tile_X9Y7_to_SB_1s),
    .from_SC_1s(Tile_X9Y7_to_SC_1s),
    .from_SD_1s(Tile_X9Y7_to_SD_1s),
    .from_SF_1s(Tile_X9Y7_to_SF_1s),
    .from_SG_1s(Tile_X9Y7_to_SG_1s),
    .from_SH_1s(Tile_X9Y7_to_SH_1s),
    .from_SI_1s(Tile_X9Y7_to_SI_1s),
    .from_WA_1s(Tile_X10Y8_to_WA_1s),
    .from_WB_1s(Tile_X10Y8_to_WB_1s),
    .from_WC_1s(Tile_X10Y8_to_WC_1s),
    .from_WD_1s(Tile_X10Y8_to_WD_1s),
    .from_WF_1s(Tile_X10Y8_to_WF_1s),
    .from_WG_1s(Tile_X10Y8_to_WG_1s),
    .from_WH_1s(Tile_X10Y8_to_WH_1s),
    .from_WI_1s(Tile_X10Y8_to_WI_1s),
    .to_EA_1s(Tile_X9Y8_to_EA_1s),
    .to_EB_1s(Tile_X9Y8_to_EB_1s),
    .to_EC_1s(Tile_X9Y8_to_EC_1s),
    .to_ED_1s(Tile_X9Y8_to_ED_1s),
    .to_EF_1s(Tile_X9Y8_to_EF_1s),
    .to_EG_1s(Tile_X9Y8_to_EG_1s),
    .to_EH_1s(Tile_X9Y8_to_EH_1s),
    .to_EI_1s(Tile_X9Y8_to_EI_1s),
    .to_WA_1s(Tile_X9Y8_to_WA_1s),
    .to_WB_1s(Tile_X9Y8_to_WB_1s),
    .to_WC_1s(Tile_X9Y8_to_WC_1s),
    .to_WD_1s(Tile_X9Y8_to_WD_1s),
    .to_WF_1s(Tile_X9Y8_to_WF_1s),
    .to_WG_1s(Tile_X9Y8_to_WG_1s),
    .to_WH_1s(Tile_X9Y8_to_WH_1s),
    .to_WI_1s(Tile_X9Y8_to_WI_1s),
    .to_NA_1s(Tile_X9Y8_to_NA_1s),
    .to_NB_1s(Tile_X9Y8_to_NB_1s),
    .to_NC_1s(Tile_X9Y8_to_NC_1s),
    .to_ND_1s(Tile_X9Y8_to_ND_1s),
    .to_NF_1s(Tile_X9Y8_to_NF_1s),
    .to_NG_1s(Tile_X9Y8_to_NG_1s),
    .to_NH_1s(Tile_X9Y8_to_NH_1s),
    .to_NI_1s(Tile_X9Y8_to_NI_1s),
    .to_SA_1s(Tile_X9Y8_to_SA_1s),
    .to_SB_1s(Tile_X9Y8_to_SB_1s),
    .to_SC_1s(Tile_X9Y8_to_SC_1s),
    .to_SD_1s(Tile_X9Y8_to_SD_1s),
    .to_SF_1s(Tile_X9Y8_to_SF_1s),
    .to_SG_1s(Tile_X9Y8_to_SG_1s),
    .to_SH_1s(Tile_X9Y8_to_SH_1s),
    .to_SI_1s(Tile_X9Y8_to_SI_1s),
    .F_ctrl(Tile_X9Y8_F_ctrl),
    .UserCLK(Tile_X9Y9_UserCLKo),
    .UserCLKo(Tile_X9Y8_UserCLKo),
    .rst(Tile_X9Y9_rsto),
    .rsto(Tile_X9Y8_rsto),
    .FrameData(Tile_X8Y8_FrameData_O),
    .FrameData_O(Tile_X9Y8_FrameData_O),
    .FrameStrobe(Tile_X9Y9_FrameStrobe_O),
    .FrameStrobe_O(Tile_X9Y8_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
ctrl_IO
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X10Y8_Emulate_Bitstream)
    )
`endif
    Tile_X10Y8_ctrl_IO
    (
    .from_EA_1s(Tile_X9Y8_to_EA_1s),
    .from_EB_1s(Tile_X9Y8_to_EB_1s),
    .from_EC_1s(Tile_X9Y8_to_EC_1s),
    .from_ED_1s(Tile_X9Y8_to_ED_1s),
    .from_EF_1s(Tile_X9Y8_to_EF_1s),
    .from_EG_1s(Tile_X9Y8_to_EG_1s),
    .from_EH_1s(Tile_X9Y8_to_EH_1s),
    .from_EI_1s(Tile_X9Y8_to_EI_1s),
    .to_WA_1s(Tile_X10Y8_to_WA_1s),
    .to_WB_1s(Tile_X10Y8_to_WB_1s),
    .to_WC_1s(Tile_X10Y8_to_WC_1s),
    .to_WD_1s(Tile_X10Y8_to_WD_1s),
    .to_WF_1s(Tile_X10Y8_to_WF_1s),
    .to_WG_1s(Tile_X10Y8_to_WG_1s),
    .to_WH_1s(Tile_X10Y8_to_WH_1s),
    .to_WI_1s(Tile_X10Y8_to_WI_1s),
    .A_O_top_0_t(Tile_X10Y8_A_O_top_0_t),
    .A_O_top_0_f(Tile_X10Y8_A_O_top_0_f),
    .A_prech2(Tile_X10Y8_A_prech2),
    .A_DR_fault(Tile_X10Y8_A_DR_fault),
    .A_I_top_0_t(Tile_X10Y8_A_I_top_0_t),
    .A_I_top_0_f(Tile_X10Y8_A_I_top_0_f),
    .A_T_top(Tile_X10Y8_A_T_top),
    .A_F_ctrl(Tile_X10Y8_A_F_ctrl),
    .UserCLK(Tile_X10Y9_UserCLKo),
    .UserCLKo(Tile_X10Y8_UserCLKo),
    .rst(Tile_X10Y9_rsto),
    .rsto(Tile_X10Y8_rsto),
    .FrameData(Tile_X9Y8_FrameData_O),
    .FrameData_O(Tile_X10Y8_FrameData_O),
    .FrameStrobe(Tile_X10Y9_FrameStrobe_O),
    .FrameStrobe_O(Tile_X10Y8_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
W_IO_custom
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X0Y9_Emulate_Bitstream)
    )
`endif
    Tile_X0Y9_W_IO_custom
    (
    .from_NA(Tile_X0Y10_to_NA),
    .from_NB(Tile_X0Y10_to_NB),
    .from_NC(Tile_X0Y10_to_NC),
    .from_ND(Tile_X0Y10_to_ND),
    .from_NF(Tile_X0Y10_to_NF),
    .from_NG(Tile_X0Y10_to_NG),
    .from_NH(Tile_X0Y10_to_NH),
    .from_NI(Tile_X0Y10_to_NI),
    .from_SA(Tile_X0Y8_to_SA),
    .from_SB(Tile_X0Y8_to_SB),
    .from_SC(Tile_X0Y8_to_SC),
    .from_SD(Tile_X0Y8_to_SD),
    .from_SF(Tile_X0Y8_to_SF),
    .from_SG(Tile_X0Y8_to_SG),
    .from_SH(Tile_X0Y8_to_SH),
    .from_SI(Tile_X0Y8_to_SI),
    .from_WA(Tile_X1Y9_to_WA),
    .from_WB(Tile_X1Y9_to_WB),
    .from_WC(Tile_X1Y9_to_WC),
    .from_WD(Tile_X1Y9_to_WD),
    .from_WF(Tile_X1Y9_to_WF),
    .from_WG(Tile_X1Y9_to_WG),
    .from_WH(Tile_X1Y9_to_WH),
    .from_WI(Tile_X1Y9_to_WI),
    .to_EA(Tile_X0Y9_to_EA),
    .to_EB(Tile_X0Y9_to_EB),
    .to_EC(Tile_X0Y9_to_EC),
    .to_ED(Tile_X0Y9_to_ED),
    .to_EF(Tile_X0Y9_to_EF),
    .to_EG(Tile_X0Y9_to_EG),
    .to_EH(Tile_X0Y9_to_EH),
    .to_EI(Tile_X0Y9_to_EI),
    .to_NA(Tile_X0Y9_to_NA),
    .to_NB(Tile_X0Y9_to_NB),
    .to_NC(Tile_X0Y9_to_NC),
    .to_ND(Tile_X0Y9_to_ND),
    .to_NF(Tile_X0Y9_to_NF),
    .to_NG(Tile_X0Y9_to_NG),
    .to_NH(Tile_X0Y9_to_NH),
    .to_NI(Tile_X0Y9_to_NI),
    .to_SA(Tile_X0Y9_to_SA),
    .to_SB(Tile_X0Y9_to_SB),
    .to_SC(Tile_X0Y9_to_SC),
    .to_SD(Tile_X0Y9_to_SD),
    .to_SF(Tile_X0Y9_to_SF),
    .to_SG(Tile_X0Y9_to_SG),
    .to_SH(Tile_X0Y9_to_SH),
    .to_SI(Tile_X0Y9_to_SI),
    .A_O_top_0_t(Tile_X0Y9_A_O_top_0_t),
    .A_O_top_0_f(Tile_X0Y9_A_O_top_0_f),
    .A_O_top_1_t(Tile_X0Y9_A_O_top_1_t),
    .A_O_top_1_f(Tile_X0Y9_A_O_top_1_f),
    .A_prech1(Tile_X0Y9_A_prech1),
    .A_prech2(Tile_X0Y9_A_prech2),
    .A_DR_fault(Tile_X0Y9_A_DR_fault),
    .A_I_top_0_t(Tile_X0Y9_A_I_top_0_t),
    .A_I_top_0_f(Tile_X0Y9_A_I_top_0_f),
    .A_I_top_1_t(Tile_X0Y9_A_I_top_1_t),
    .A_I_top_1_f(Tile_X0Y9_A_I_top_1_f),
    .A_T_top(Tile_X0Y9_A_T_top),
    .A_F_masked1(Tile_X0Y9_A_F_masked1),
    .A_F_masked2(Tile_X0Y9_A_F_masked2),
    .A_config_C_bit0(Tile_X0Y9_A_config_C_bit0),
    .A_config_C_bit1(Tile_X0Y9_A_config_C_bit1),
    .A_config_C_bit2(Tile_X0Y9_A_config_C_bit2),
    .A_config_C_bit3(Tile_X0Y9_A_config_C_bit3),
    .B_config_C_bit0(Tile_X0Y9_B_config_C_bit0),
    .B_config_C_bit1(Tile_X0Y9_B_config_C_bit1),
    .B_config_C_bit2(Tile_X0Y9_B_config_C_bit2),
    .B_config_C_bit3(Tile_X0Y9_B_config_C_bit3),
    .UserCLK(Tile_X0Y10_UserCLKo),
    .UserCLKo(Tile_X0Y9_UserCLKo),
    .rst(Tile_X0Y10_rsto),
    .rsto(Tile_X0Y9_rsto),
    .FrameData(Tile_Y9_FrameData),
    .FrameData_O(Tile_X0Y9_FrameData_O),
    .FrameStrobe(Tile_X0Y10_FrameStrobe_O),
    .FrameStrobe_O(Tile_X0Y9_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X1Y9_Emulate_Bitstream)
    )
`endif
    Tile_X1Y9_linear_LMDPL
    (
    .from_NA(Tile_X1Y10_to_NA),
    .from_NB(Tile_X1Y10_to_NB),
    .from_NC(Tile_X1Y10_to_NC),
    .from_ND(Tile_X1Y10_to_ND),
    .from_NF(Tile_X1Y10_to_NF),
    .from_NG(Tile_X1Y10_to_NG),
    .from_NH(Tile_X1Y10_to_NH),
    .from_NI(Tile_X1Y10_to_NI),
    .from_EA(Tile_X0Y9_to_EA),
    .from_EB(Tile_X0Y9_to_EB),
    .from_EC(Tile_X0Y9_to_EC),
    .from_ED(Tile_X0Y9_to_ED),
    .from_EF(Tile_X0Y9_to_EF),
    .from_EG(Tile_X0Y9_to_EG),
    .from_EH(Tile_X0Y9_to_EH),
    .from_EI(Tile_X0Y9_to_EI),
    .from_SA(Tile_X1Y8_to_SA),
    .from_SB(Tile_X1Y8_to_SB),
    .from_SC(Tile_X1Y8_to_SC),
    .from_SD(Tile_X1Y8_to_SD),
    .from_SF(Tile_X1Y8_to_SF),
    .from_SG(Tile_X1Y8_to_SG),
    .from_SH(Tile_X1Y8_to_SH),
    .from_SI(Tile_X1Y8_to_SI),
    .from_WA(Tile_X2Y9_to_WA),
    .from_WB(Tile_X2Y9_to_WB),
    .from_WC(Tile_X2Y9_to_WC),
    .from_WD(Tile_X2Y9_to_WD),
    .from_WF(Tile_X2Y9_to_WF),
    .from_WG(Tile_X2Y9_to_WG),
    .from_WH(Tile_X2Y9_to_WH),
    .from_WI(Tile_X2Y9_to_WI),
    .to_EA(Tile_X1Y9_to_EA),
    .to_EB(Tile_X1Y9_to_EB),
    .to_EC(Tile_X1Y9_to_EC),
    .to_ED(Tile_X1Y9_to_ED),
    .to_EF(Tile_X1Y9_to_EF),
    .to_EG(Tile_X1Y9_to_EG),
    .to_EH(Tile_X1Y9_to_EH),
    .to_EI(Tile_X1Y9_to_EI),
    .to_WA(Tile_X1Y9_to_WA),
    .to_WB(Tile_X1Y9_to_WB),
    .to_WC(Tile_X1Y9_to_WC),
    .to_WD(Tile_X1Y9_to_WD),
    .to_WF(Tile_X1Y9_to_WF),
    .to_WG(Tile_X1Y9_to_WG),
    .to_WH(Tile_X1Y9_to_WH),
    .to_WI(Tile_X1Y9_to_WI),
    .to_NA(Tile_X1Y9_to_NA),
    .to_NB(Tile_X1Y9_to_NB),
    .to_NC(Tile_X1Y9_to_NC),
    .to_ND(Tile_X1Y9_to_ND),
    .to_NF(Tile_X1Y9_to_NF),
    .to_NG(Tile_X1Y9_to_NG),
    .to_NH(Tile_X1Y9_to_NH),
    .to_NI(Tile_X1Y9_to_NI),
    .to_SA(Tile_X1Y9_to_SA),
    .to_SB(Tile_X1Y9_to_SB),
    .to_SC(Tile_X1Y9_to_SC),
    .to_SD(Tile_X1Y9_to_SD),
    .to_SF(Tile_X1Y9_to_SF),
    .to_SG(Tile_X1Y9_to_SG),
    .to_SH(Tile_X1Y9_to_SH),
    .to_SI(Tile_X1Y9_to_SI),
    .F_masked1(Tile_X1Y9_F_masked1),
    .F_masked2(Tile_X1Y9_F_masked2),
    .UserCLK(Tile_X1Y10_UserCLKo),
    .UserCLKo(Tile_X1Y9_UserCLKo),
    .rst(Tile_X1Y10_rsto),
    .rsto(Tile_X1Y9_rsto),
    .FrameData(Tile_X0Y9_FrameData_O),
    .FrameData_O(Tile_X1Y9_FrameData_O),
    .FrameStrobe(Tile_X1Y10_FrameStrobe_O),
    .FrameStrobe_O(Tile_X1Y9_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X2Y9_Emulate_Bitstream)
    )
`endif
    Tile_X2Y9_linear_LMDPL
    (
    .from_NA(Tile_X2Y10_to_NA),
    .from_NB(Tile_X2Y10_to_NB),
    .from_NC(Tile_X2Y10_to_NC),
    .from_ND(Tile_X2Y10_to_ND),
    .from_NF(Tile_X2Y10_to_NF),
    .from_NG(Tile_X2Y10_to_NG),
    .from_NH(Tile_X2Y10_to_NH),
    .from_NI(Tile_X2Y10_to_NI),
    .from_EA(Tile_X1Y9_to_EA),
    .from_EB(Tile_X1Y9_to_EB),
    .from_EC(Tile_X1Y9_to_EC),
    .from_ED(Tile_X1Y9_to_ED),
    .from_EF(Tile_X1Y9_to_EF),
    .from_EG(Tile_X1Y9_to_EG),
    .from_EH(Tile_X1Y9_to_EH),
    .from_EI(Tile_X1Y9_to_EI),
    .from_SA(Tile_X2Y8_to_SA),
    .from_SB(Tile_X2Y8_to_SB),
    .from_SC(Tile_X2Y8_to_SC),
    .from_SD(Tile_X2Y8_to_SD),
    .from_SF(Tile_X2Y8_to_SF),
    .from_SG(Tile_X2Y8_to_SG),
    .from_SH(Tile_X2Y8_to_SH),
    .from_SI(Tile_X2Y8_to_SI),
    .from_WA(Tile_X3Y9_to_WA),
    .from_WB(Tile_X3Y9_to_WB),
    .from_WC(Tile_X3Y9_to_WC),
    .from_WD(Tile_X3Y9_to_WD),
    .from_WF(Tile_X3Y9_to_WF),
    .from_WG(Tile_X3Y9_to_WG),
    .from_WH(Tile_X3Y9_to_WH),
    .from_WI(Tile_X3Y9_to_WI),
    .to_EA(Tile_X2Y9_to_EA),
    .to_EB(Tile_X2Y9_to_EB),
    .to_EC(Tile_X2Y9_to_EC),
    .to_ED(Tile_X2Y9_to_ED),
    .to_EF(Tile_X2Y9_to_EF),
    .to_EG(Tile_X2Y9_to_EG),
    .to_EH(Tile_X2Y9_to_EH),
    .to_EI(Tile_X2Y9_to_EI),
    .to_WA(Tile_X2Y9_to_WA),
    .to_WB(Tile_X2Y9_to_WB),
    .to_WC(Tile_X2Y9_to_WC),
    .to_WD(Tile_X2Y9_to_WD),
    .to_WF(Tile_X2Y9_to_WF),
    .to_WG(Tile_X2Y9_to_WG),
    .to_WH(Tile_X2Y9_to_WH),
    .to_WI(Tile_X2Y9_to_WI),
    .to_NA(Tile_X2Y9_to_NA),
    .to_NB(Tile_X2Y9_to_NB),
    .to_NC(Tile_X2Y9_to_NC),
    .to_ND(Tile_X2Y9_to_ND),
    .to_NF(Tile_X2Y9_to_NF),
    .to_NG(Tile_X2Y9_to_NG),
    .to_NH(Tile_X2Y9_to_NH),
    .to_NI(Tile_X2Y9_to_NI),
    .to_SA(Tile_X2Y9_to_SA),
    .to_SB(Tile_X2Y9_to_SB),
    .to_SC(Tile_X2Y9_to_SC),
    .to_SD(Tile_X2Y9_to_SD),
    .to_SF(Tile_X2Y9_to_SF),
    .to_SG(Tile_X2Y9_to_SG),
    .to_SH(Tile_X2Y9_to_SH),
    .to_SI(Tile_X2Y9_to_SI),
    .F_masked1(Tile_X2Y9_F_masked1),
    .F_masked2(Tile_X2Y9_F_masked2),
    .UserCLK(Tile_X2Y10_UserCLKo),
    .UserCLKo(Tile_X2Y9_UserCLKo),
    .rst(Tile_X2Y10_rsto),
    .rsto(Tile_X2Y9_rsto),
    .FrameData(Tile_X1Y9_FrameData_O),
    .FrameData_O(Tile_X2Y9_FrameData_O),
    .FrameStrobe(Tile_X2Y10_FrameStrobe_O),
    .FrameStrobe_O(Tile_X2Y9_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
nonlinear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X3Y9_Emulate_Bitstream)
    )
`endif
    Tile_X3Y9_nonlinear_LMDPL
    (
    .from_NA(Tile_X3Y10_to_NA),
    .from_NB(Tile_X3Y10_to_NB),
    .from_NC(Tile_X3Y10_to_NC),
    .from_ND(Tile_X3Y10_to_ND),
    .from_NF(Tile_X3Y10_to_NF),
    .from_NG(Tile_X3Y10_to_NG),
    .from_NH(Tile_X3Y10_to_NH),
    .from_NI(Tile_X3Y10_to_NI),
    .from_EA(Tile_X2Y9_to_EA),
    .from_EB(Tile_X2Y9_to_EB),
    .from_EC(Tile_X2Y9_to_EC),
    .from_ED(Tile_X2Y9_to_ED),
    .from_EF(Tile_X2Y9_to_EF),
    .from_EG(Tile_X2Y9_to_EG),
    .from_EH(Tile_X2Y9_to_EH),
    .from_EI(Tile_X2Y9_to_EI),
    .from_SA(Tile_X3Y8_to_SA),
    .from_SB(Tile_X3Y8_to_SB),
    .from_SC(Tile_X3Y8_to_SC),
    .from_SD(Tile_X3Y8_to_SD),
    .from_SF(Tile_X3Y8_to_SF),
    .from_SG(Tile_X3Y8_to_SG),
    .from_SH(Tile_X3Y8_to_SH),
    .from_SI(Tile_X3Y8_to_SI),
    .from_WA(Tile_X4Y9_to_WA),
    .from_WB(Tile_X4Y9_to_WB),
    .from_WC(Tile_X4Y9_to_WC),
    .from_WD(Tile_X4Y9_to_WD),
    .from_WF(Tile_X4Y9_to_WF),
    .from_WG(Tile_X4Y9_to_WG),
    .from_WH(Tile_X4Y9_to_WH),
    .from_WI(Tile_X4Y9_to_WI),
    .to_EA(Tile_X3Y9_to_EA),
    .to_EB(Tile_X3Y9_to_EB),
    .to_EC(Tile_X3Y9_to_EC),
    .to_ED(Tile_X3Y9_to_ED),
    .to_EF(Tile_X3Y9_to_EF),
    .to_EG(Tile_X3Y9_to_EG),
    .to_EH(Tile_X3Y9_to_EH),
    .to_EI(Tile_X3Y9_to_EI),
    .to_WA(Tile_X3Y9_to_WA),
    .to_WB(Tile_X3Y9_to_WB),
    .to_WC(Tile_X3Y9_to_WC),
    .to_WD(Tile_X3Y9_to_WD),
    .to_WF(Tile_X3Y9_to_WF),
    .to_WG(Tile_X3Y9_to_WG),
    .to_WH(Tile_X3Y9_to_WH),
    .to_WI(Tile_X3Y9_to_WI),
    .to_NA(Tile_X3Y9_to_NA),
    .to_NB(Tile_X3Y9_to_NB),
    .to_NC(Tile_X3Y9_to_NC),
    .to_ND(Tile_X3Y9_to_ND),
    .to_NF(Tile_X3Y9_to_NF),
    .to_NG(Tile_X3Y9_to_NG),
    .to_NH(Tile_X3Y9_to_NH),
    .to_NI(Tile_X3Y9_to_NI),
    .to_SA(Tile_X3Y9_to_SA),
    .to_SB(Tile_X3Y9_to_SB),
    .to_SC(Tile_X3Y9_to_SC),
    .to_SD(Tile_X3Y9_to_SD),
    .to_SF(Tile_X3Y9_to_SF),
    .to_SG(Tile_X3Y9_to_SG),
    .to_SH(Tile_X3Y9_to_SH),
    .to_SI(Tile_X3Y9_to_SI),
    .R_t(Tile_X3Y9_R_t),
    .R_f(Tile_X3Y9_R_f),
    .F_masked1(Tile_X3Y9_F_masked1),
    .F_masked2(Tile_X3Y9_F_masked2),
    .UserCLK(Tile_X3Y10_UserCLKo),
    .UserCLKo(Tile_X3Y9_UserCLKo),
    .rst(Tile_X3Y10_rsto),
    .rsto(Tile_X3Y9_rsto),
    .FrameData(Tile_X2Y9_FrameData_O),
    .FrameData_O(Tile_X3Y9_FrameData_O),
    .FrameStrobe(Tile_X3Y10_FrameStrobe_O),
    .FrameStrobe_O(Tile_X3Y9_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X4Y9_Emulate_Bitstream)
    )
`endif
    Tile_X4Y9_linear_LMDPL
    (
    .from_NA(Tile_X4Y10_to_NA),
    .from_NB(Tile_X4Y10_to_NB),
    .from_NC(Tile_X4Y10_to_NC),
    .from_ND(Tile_X4Y10_to_ND),
    .from_NF(Tile_X4Y10_to_NF),
    .from_NG(Tile_X4Y10_to_NG),
    .from_NH(Tile_X4Y10_to_NH),
    .from_NI(Tile_X4Y10_to_NI),
    .from_EA(Tile_X3Y9_to_EA),
    .from_EB(Tile_X3Y9_to_EB),
    .from_EC(Tile_X3Y9_to_EC),
    .from_ED(Tile_X3Y9_to_ED),
    .from_EF(Tile_X3Y9_to_EF),
    .from_EG(Tile_X3Y9_to_EG),
    .from_EH(Tile_X3Y9_to_EH),
    .from_EI(Tile_X3Y9_to_EI),
    .from_SA(Tile_X4Y8_to_SA),
    .from_SB(Tile_X4Y8_to_SB),
    .from_SC(Tile_X4Y8_to_SC),
    .from_SD(Tile_X4Y8_to_SD),
    .from_SF(Tile_X4Y8_to_SF),
    .from_SG(Tile_X4Y8_to_SG),
    .from_SH(Tile_X4Y8_to_SH),
    .from_SI(Tile_X4Y8_to_SI),
    .from_WA(Tile_X5Y9_to_WA),
    .from_WB(Tile_X5Y9_to_WB),
    .from_WC(Tile_X5Y9_to_WC),
    .from_WD(Tile_X5Y9_to_WD),
    .from_WF(Tile_X5Y9_to_WF),
    .from_WG(Tile_X5Y9_to_WG),
    .from_WH(Tile_X5Y9_to_WH),
    .from_WI(Tile_X5Y9_to_WI),
    .to_EA(Tile_X4Y9_to_EA),
    .to_EB(Tile_X4Y9_to_EB),
    .to_EC(Tile_X4Y9_to_EC),
    .to_ED(Tile_X4Y9_to_ED),
    .to_EF(Tile_X4Y9_to_EF),
    .to_EG(Tile_X4Y9_to_EG),
    .to_EH(Tile_X4Y9_to_EH),
    .to_EI(Tile_X4Y9_to_EI),
    .to_WA(Tile_X4Y9_to_WA),
    .to_WB(Tile_X4Y9_to_WB),
    .to_WC(Tile_X4Y9_to_WC),
    .to_WD(Tile_X4Y9_to_WD),
    .to_WF(Tile_X4Y9_to_WF),
    .to_WG(Tile_X4Y9_to_WG),
    .to_WH(Tile_X4Y9_to_WH),
    .to_WI(Tile_X4Y9_to_WI),
    .to_NA(Tile_X4Y9_to_NA),
    .to_NB(Tile_X4Y9_to_NB),
    .to_NC(Tile_X4Y9_to_NC),
    .to_ND(Tile_X4Y9_to_ND),
    .to_NF(Tile_X4Y9_to_NF),
    .to_NG(Tile_X4Y9_to_NG),
    .to_NH(Tile_X4Y9_to_NH),
    .to_NI(Tile_X4Y9_to_NI),
    .to_SA(Tile_X4Y9_to_SA),
    .to_SB(Tile_X4Y9_to_SB),
    .to_SC(Tile_X4Y9_to_SC),
    .to_SD(Tile_X4Y9_to_SD),
    .to_SF(Tile_X4Y9_to_SF),
    .to_SG(Tile_X4Y9_to_SG),
    .to_SH(Tile_X4Y9_to_SH),
    .to_SI(Tile_X4Y9_to_SI),
    .F_masked1(Tile_X4Y9_F_masked1),
    .F_masked2(Tile_X4Y9_F_masked2),
    .UserCLK(Tile_X4Y10_UserCLKo),
    .UserCLKo(Tile_X4Y9_UserCLKo),
    .rst(Tile_X4Y10_rsto),
    .rsto(Tile_X4Y9_rsto),
    .FrameData(Tile_X3Y9_FrameData_O),
    .FrameData_O(Tile_X4Y9_FrameData_O),
    .FrameStrobe(Tile_X4Y10_FrameStrobe_O),
    .FrameStrobe_O(Tile_X4Y9_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X5Y9_Emulate_Bitstream)
    )
`endif
    Tile_X5Y9_linear_LMDPL
    (
    .from_NA(Tile_X5Y10_to_NA),
    .from_NB(Tile_X5Y10_to_NB),
    .from_NC(Tile_X5Y10_to_NC),
    .from_ND(Tile_X5Y10_to_ND),
    .from_NF(Tile_X5Y10_to_NF),
    .from_NG(Tile_X5Y10_to_NG),
    .from_NH(Tile_X5Y10_to_NH),
    .from_NI(Tile_X5Y10_to_NI),
    .from_EA(Tile_X4Y9_to_EA),
    .from_EB(Tile_X4Y9_to_EB),
    .from_EC(Tile_X4Y9_to_EC),
    .from_ED(Tile_X4Y9_to_ED),
    .from_EF(Tile_X4Y9_to_EF),
    .from_EG(Tile_X4Y9_to_EG),
    .from_EH(Tile_X4Y9_to_EH),
    .from_EI(Tile_X4Y9_to_EI),
    .from_SA(Tile_X5Y8_to_SA),
    .from_SB(Tile_X5Y8_to_SB),
    .from_SC(Tile_X5Y8_to_SC),
    .from_SD(Tile_X5Y8_to_SD),
    .from_SF(Tile_X5Y8_to_SF),
    .from_SG(Tile_X5Y8_to_SG),
    .from_SH(Tile_X5Y8_to_SH),
    .from_SI(Tile_X5Y8_to_SI),
    .from_WA(Tile_X6Y9_to_WA),
    .from_WB(Tile_X6Y9_to_WB),
    .from_WC(Tile_X6Y9_to_WC),
    .from_WD(Tile_X6Y9_to_WD),
    .from_WF(Tile_X6Y9_to_WF),
    .from_WG(Tile_X6Y9_to_WG),
    .from_WH(Tile_X6Y9_to_WH),
    .from_WI(Tile_X6Y9_to_WI),
    .to_EA(Tile_X5Y9_to_EA),
    .to_EB(Tile_X5Y9_to_EB),
    .to_EC(Tile_X5Y9_to_EC),
    .to_ED(Tile_X5Y9_to_ED),
    .to_EF(Tile_X5Y9_to_EF),
    .to_EG(Tile_X5Y9_to_EG),
    .to_EH(Tile_X5Y9_to_EH),
    .to_EI(Tile_X5Y9_to_EI),
    .to_WA(Tile_X5Y9_to_WA),
    .to_WB(Tile_X5Y9_to_WB),
    .to_WC(Tile_X5Y9_to_WC),
    .to_WD(Tile_X5Y9_to_WD),
    .to_WF(Tile_X5Y9_to_WF),
    .to_WG(Tile_X5Y9_to_WG),
    .to_WH(Tile_X5Y9_to_WH),
    .to_WI(Tile_X5Y9_to_WI),
    .to_NA(Tile_X5Y9_to_NA),
    .to_NB(Tile_X5Y9_to_NB),
    .to_NC(Tile_X5Y9_to_NC),
    .to_ND(Tile_X5Y9_to_ND),
    .to_NF(Tile_X5Y9_to_NF),
    .to_NG(Tile_X5Y9_to_NG),
    .to_NH(Tile_X5Y9_to_NH),
    .to_NI(Tile_X5Y9_to_NI),
    .to_SA(Tile_X5Y9_to_SA),
    .to_SB(Tile_X5Y9_to_SB),
    .to_SC(Tile_X5Y9_to_SC),
    .to_SD(Tile_X5Y9_to_SD),
    .to_SF(Tile_X5Y9_to_SF),
    .to_SG(Tile_X5Y9_to_SG),
    .to_SH(Tile_X5Y9_to_SH),
    .to_SI(Tile_X5Y9_to_SI),
    .F_masked1(Tile_X5Y9_F_masked1),
    .F_masked2(Tile_X5Y9_F_masked2),
    .UserCLK(Tile_X5Y10_UserCLKo),
    .UserCLKo(Tile_X5Y9_UserCLKo),
    .rst(Tile_X5Y10_rsto),
    .rsto(Tile_X5Y9_rsto),
    .FrameData(Tile_X4Y9_FrameData_O),
    .FrameData_O(Tile_X5Y9_FrameData_O),
    .FrameStrobe(Tile_X5Y10_FrameStrobe_O),
    .FrameStrobe_O(Tile_X5Y9_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
nonlinear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X6Y9_Emulate_Bitstream)
    )
`endif
    Tile_X6Y9_nonlinear_LMDPL
    (
    .from_NA(Tile_X6Y10_to_NA),
    .from_NB(Tile_X6Y10_to_NB),
    .from_NC(Tile_X6Y10_to_NC),
    .from_ND(Tile_X6Y10_to_ND),
    .from_NF(Tile_X6Y10_to_NF),
    .from_NG(Tile_X6Y10_to_NG),
    .from_NH(Tile_X6Y10_to_NH),
    .from_NI(Tile_X6Y10_to_NI),
    .from_EA(Tile_X5Y9_to_EA),
    .from_EB(Tile_X5Y9_to_EB),
    .from_EC(Tile_X5Y9_to_EC),
    .from_ED(Tile_X5Y9_to_ED),
    .from_EF(Tile_X5Y9_to_EF),
    .from_EG(Tile_X5Y9_to_EG),
    .from_EH(Tile_X5Y9_to_EH),
    .from_EI(Tile_X5Y9_to_EI),
    .from_SA(Tile_X6Y8_to_SA),
    .from_SB(Tile_X6Y8_to_SB),
    .from_SC(Tile_X6Y8_to_SC),
    .from_SD(Tile_X6Y8_to_SD),
    .from_SF(Tile_X6Y8_to_SF),
    .from_SG(Tile_X6Y8_to_SG),
    .from_SH(Tile_X6Y8_to_SH),
    .from_SI(Tile_X6Y8_to_SI),
    .from_WA(Tile_X7Y9_to_WA),
    .from_WB(Tile_X7Y9_to_WB),
    .from_WC(Tile_X7Y9_to_WC),
    .from_WD(Tile_X7Y9_to_WD),
    .from_WF(Tile_X7Y9_to_WF),
    .from_WG(Tile_X7Y9_to_WG),
    .from_WH(Tile_X7Y9_to_WH),
    .from_WI(Tile_X7Y9_to_WI),
    .to_EA(Tile_X6Y9_to_EA),
    .to_EB(Tile_X6Y9_to_EB),
    .to_EC(Tile_X6Y9_to_EC),
    .to_ED(Tile_X6Y9_to_ED),
    .to_EF(Tile_X6Y9_to_EF),
    .to_EG(Tile_X6Y9_to_EG),
    .to_EH(Tile_X6Y9_to_EH),
    .to_EI(Tile_X6Y9_to_EI),
    .to_WA(Tile_X6Y9_to_WA),
    .to_WB(Tile_X6Y9_to_WB),
    .to_WC(Tile_X6Y9_to_WC),
    .to_WD(Tile_X6Y9_to_WD),
    .to_WF(Tile_X6Y9_to_WF),
    .to_WG(Tile_X6Y9_to_WG),
    .to_WH(Tile_X6Y9_to_WH),
    .to_WI(Tile_X6Y9_to_WI),
    .to_NA(Tile_X6Y9_to_NA),
    .to_NB(Tile_X6Y9_to_NB),
    .to_NC(Tile_X6Y9_to_NC),
    .to_ND(Tile_X6Y9_to_ND),
    .to_NF(Tile_X6Y9_to_NF),
    .to_NG(Tile_X6Y9_to_NG),
    .to_NH(Tile_X6Y9_to_NH),
    .to_NI(Tile_X6Y9_to_NI),
    .to_SA(Tile_X6Y9_to_SA),
    .to_SB(Tile_X6Y9_to_SB),
    .to_SC(Tile_X6Y9_to_SC),
    .to_SD(Tile_X6Y9_to_SD),
    .to_SF(Tile_X6Y9_to_SF),
    .to_SG(Tile_X6Y9_to_SG),
    .to_SH(Tile_X6Y9_to_SH),
    .to_SI(Tile_X6Y9_to_SI),
    .R_t(Tile_X6Y9_R_t),
    .R_f(Tile_X6Y9_R_f),
    .F_masked1(Tile_X6Y9_F_masked1),
    .F_masked2(Tile_X6Y9_F_masked2),
    .UserCLK(Tile_X6Y10_UserCLKo),
    .UserCLKo(Tile_X6Y9_UserCLKo),
    .rst(Tile_X6Y10_rsto),
    .rsto(Tile_X6Y9_rsto),
    .FrameData(Tile_X5Y9_FrameData_O),
    .FrameData_O(Tile_X6Y9_FrameData_O),
    .FrameStrobe(Tile_X6Y10_FrameStrobe_O),
    .FrameStrobe_O(Tile_X6Y9_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X7Y9_Emulate_Bitstream)
    )
`endif
    Tile_X7Y9_linear_LMDPL
    (
    .from_NA(Tile_X7Y10_to_NA),
    .from_NB(Tile_X7Y10_to_NB),
    .from_NC(Tile_X7Y10_to_NC),
    .from_ND(Tile_X7Y10_to_ND),
    .from_NF(Tile_X7Y10_to_NF),
    .from_NG(Tile_X7Y10_to_NG),
    .from_NH(Tile_X7Y10_to_NH),
    .from_NI(Tile_X7Y10_to_NI),
    .from_EA(Tile_X6Y9_to_EA),
    .from_EB(Tile_X6Y9_to_EB),
    .from_EC(Tile_X6Y9_to_EC),
    .from_ED(Tile_X6Y9_to_ED),
    .from_EF(Tile_X6Y9_to_EF),
    .from_EG(Tile_X6Y9_to_EG),
    .from_EH(Tile_X6Y9_to_EH),
    .from_EI(Tile_X6Y9_to_EI),
    .from_SA(Tile_X7Y8_to_SA),
    .from_SB(Tile_X7Y8_to_SB),
    .from_SC(Tile_X7Y8_to_SC),
    .from_SD(Tile_X7Y8_to_SD),
    .from_SF(Tile_X7Y8_to_SF),
    .from_SG(Tile_X7Y8_to_SG),
    .from_SH(Tile_X7Y8_to_SH),
    .from_SI(Tile_X7Y8_to_SI),
    .from_WA(Tile_X8Y9_to_WA),
    .from_WB(Tile_X8Y9_to_WB),
    .from_WC(Tile_X8Y9_to_WC),
    .from_WD(Tile_X8Y9_to_WD),
    .from_WF(Tile_X8Y9_to_WF),
    .from_WG(Tile_X8Y9_to_WG),
    .from_WH(Tile_X8Y9_to_WH),
    .from_WI(Tile_X8Y9_to_WI),
    .to_EA(Tile_X7Y9_to_EA),
    .to_EB(Tile_X7Y9_to_EB),
    .to_EC(Tile_X7Y9_to_EC),
    .to_ED(Tile_X7Y9_to_ED),
    .to_EF(Tile_X7Y9_to_EF),
    .to_EG(Tile_X7Y9_to_EG),
    .to_EH(Tile_X7Y9_to_EH),
    .to_EI(Tile_X7Y9_to_EI),
    .to_WA(Tile_X7Y9_to_WA),
    .to_WB(Tile_X7Y9_to_WB),
    .to_WC(Tile_X7Y9_to_WC),
    .to_WD(Tile_X7Y9_to_WD),
    .to_WF(Tile_X7Y9_to_WF),
    .to_WG(Tile_X7Y9_to_WG),
    .to_WH(Tile_X7Y9_to_WH),
    .to_WI(Tile_X7Y9_to_WI),
    .to_NA(Tile_X7Y9_to_NA),
    .to_NB(Tile_X7Y9_to_NB),
    .to_NC(Tile_X7Y9_to_NC),
    .to_ND(Tile_X7Y9_to_ND),
    .to_NF(Tile_X7Y9_to_NF),
    .to_NG(Tile_X7Y9_to_NG),
    .to_NH(Tile_X7Y9_to_NH),
    .to_NI(Tile_X7Y9_to_NI),
    .to_SA(Tile_X7Y9_to_SA),
    .to_SB(Tile_X7Y9_to_SB),
    .to_SC(Tile_X7Y9_to_SC),
    .to_SD(Tile_X7Y9_to_SD),
    .to_SF(Tile_X7Y9_to_SF),
    .to_SG(Tile_X7Y9_to_SG),
    .to_SH(Tile_X7Y9_to_SH),
    .to_SI(Tile_X7Y9_to_SI),
    .F_masked1(Tile_X7Y9_F_masked1),
    .F_masked2(Tile_X7Y9_F_masked2),
    .UserCLK(Tile_X7Y10_UserCLKo),
    .UserCLKo(Tile_X7Y9_UserCLKo),
    .rst(Tile_X7Y10_rsto),
    .rsto(Tile_X7Y9_rsto),
    .FrameData(Tile_X6Y9_FrameData_O),
    .FrameData_O(Tile_X7Y9_FrameData_O),
    .FrameStrobe(Tile_X7Y10_FrameStrobe_O),
    .FrameStrobe_O(Tile_X7Y9_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
ctrl_to_sec
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X8Y9_Emulate_Bitstream)
    )
`endif
    Tile_X8Y9_ctrl_to_sec
    (
    .from_NA(Tile_X8Y10_to_NA),
    .from_NB(Tile_X8Y10_to_NB),
    .from_NC(Tile_X8Y10_to_NC),
    .from_ND(Tile_X8Y10_to_ND),
    .from_NF(Tile_X8Y10_to_NF),
    .from_NG(Tile_X8Y10_to_NG),
    .from_NH(Tile_X8Y10_to_NH),
    .from_NI(Tile_X8Y10_to_NI),
    .from_EA(Tile_X7Y9_to_EA),
    .from_EB(Tile_X7Y9_to_EB),
    .from_EC(Tile_X7Y9_to_EC),
    .from_ED(Tile_X7Y9_to_ED),
    .from_EF(Tile_X7Y9_to_EF),
    .from_EG(Tile_X7Y9_to_EG),
    .from_EH(Tile_X7Y9_to_EH),
    .from_EI(Tile_X7Y9_to_EI),
    .from_SA(Tile_X8Y8_to_SA),
    .from_SB(Tile_X8Y8_to_SB),
    .from_SC(Tile_X8Y8_to_SC),
    .from_SD(Tile_X8Y8_to_SD),
    .from_SF(Tile_X8Y8_to_SF),
    .from_SG(Tile_X8Y8_to_SG),
    .from_SH(Tile_X8Y8_to_SH),
    .from_SI(Tile_X8Y8_to_SI),
    .from_WA_1s(Tile_X9Y9_to_WA_1s),
    .from_WB_1s(Tile_X9Y9_to_WB_1s),
    .from_WC_1s(Tile_X9Y9_to_WC_1s),
    .from_WD_1s(Tile_X9Y9_to_WD_1s),
    .from_WF_1s(Tile_X9Y9_to_WF_1s),
    .from_WG_1s(Tile_X9Y9_to_WG_1s),
    .from_WH_1s(Tile_X9Y9_to_WH_1s),
    .from_WI_1s(Tile_X9Y9_to_WI_1s),
    .to_WA(Tile_X8Y9_to_WA),
    .to_WB(Tile_X8Y9_to_WB),
    .to_WC(Tile_X8Y9_to_WC),
    .to_WD(Tile_X8Y9_to_WD),
    .to_WF(Tile_X8Y9_to_WF),
    .to_WG(Tile_X8Y9_to_WG),
    .to_WH(Tile_X8Y9_to_WH),
    .to_WI(Tile_X8Y9_to_WI),
    .to_NA(Tile_X8Y9_to_NA),
    .to_NB(Tile_X8Y9_to_NB),
    .to_NC(Tile_X8Y9_to_NC),
    .to_ND(Tile_X8Y9_to_ND),
    .to_NF(Tile_X8Y9_to_NF),
    .to_NG(Tile_X8Y9_to_NG),
    .to_NH(Tile_X8Y9_to_NH),
    .to_NI(Tile_X8Y9_to_NI),
    .to_SA(Tile_X8Y9_to_SA),
    .to_SB(Tile_X8Y9_to_SB),
    .to_SC(Tile_X8Y9_to_SC),
    .to_SD(Tile_X8Y9_to_SD),
    .to_SF(Tile_X8Y9_to_SF),
    .to_SG(Tile_X8Y9_to_SG),
    .to_SH(Tile_X8Y9_to_SH),
    .to_SI(Tile_X8Y9_to_SI),
    .UserCLK(Tile_X8Y10_UserCLKo),
    .UserCLKo(Tile_X8Y9_UserCLKo),
    .rst(Tile_X8Y10_rsto),
    .rsto(Tile_X8Y9_rsto),
    .FrameData(Tile_X7Y9_FrameData_O),
    .FrameData_O(Tile_X8Y9_FrameData_O),
    .FrameStrobe(Tile_X8Y10_FrameStrobe_O),
    .FrameStrobe_O(Tile_X8Y9_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
combined_WDDL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X9Y9_Emulate_Bitstream)
    )
`endif
    Tile_X9Y9_combined_WDDL
    (
    .from_NA_1s(Tile_X9Y10_to_NA_1s),
    .from_NB_1s(Tile_X9Y10_to_NB_1s),
    .from_NC_1s(Tile_X9Y10_to_NC_1s),
    .from_ND_1s(Tile_X9Y10_to_ND_1s),
    .from_NF_1s(Tile_X9Y10_to_NF_1s),
    .from_NG_1s(Tile_X9Y10_to_NG_1s),
    .from_NH_1s(Tile_X9Y10_to_NH_1s),
    .from_NI_1s(Tile_X9Y10_to_NI_1s),
    .from_SA_1s(Tile_X9Y8_to_SA_1s),
    .from_SB_1s(Tile_X9Y8_to_SB_1s),
    .from_SC_1s(Tile_X9Y8_to_SC_1s),
    .from_SD_1s(Tile_X9Y8_to_SD_1s),
    .from_SF_1s(Tile_X9Y8_to_SF_1s),
    .from_SG_1s(Tile_X9Y8_to_SG_1s),
    .from_SH_1s(Tile_X9Y8_to_SH_1s),
    .from_SI_1s(Tile_X9Y8_to_SI_1s),
    .from_WA_1s(Tile_X10Y9_to_WA_1s),
    .from_WB_1s(Tile_X10Y9_to_WB_1s),
    .from_WC_1s(Tile_X10Y9_to_WC_1s),
    .from_WD_1s(Tile_X10Y9_to_WD_1s),
    .from_WF_1s(Tile_X10Y9_to_WF_1s),
    .from_WG_1s(Tile_X10Y9_to_WG_1s),
    .from_WH_1s(Tile_X10Y9_to_WH_1s),
    .from_WI_1s(Tile_X10Y9_to_WI_1s),
    .to_EA_1s(Tile_X9Y9_to_EA_1s),
    .to_EB_1s(Tile_X9Y9_to_EB_1s),
    .to_EC_1s(Tile_X9Y9_to_EC_1s),
    .to_ED_1s(Tile_X9Y9_to_ED_1s),
    .to_EF_1s(Tile_X9Y9_to_EF_1s),
    .to_EG_1s(Tile_X9Y9_to_EG_1s),
    .to_EH_1s(Tile_X9Y9_to_EH_1s),
    .to_EI_1s(Tile_X9Y9_to_EI_1s),
    .to_WA_1s(Tile_X9Y9_to_WA_1s),
    .to_WB_1s(Tile_X9Y9_to_WB_1s),
    .to_WC_1s(Tile_X9Y9_to_WC_1s),
    .to_WD_1s(Tile_X9Y9_to_WD_1s),
    .to_WF_1s(Tile_X9Y9_to_WF_1s),
    .to_WG_1s(Tile_X9Y9_to_WG_1s),
    .to_WH_1s(Tile_X9Y9_to_WH_1s),
    .to_WI_1s(Tile_X9Y9_to_WI_1s),
    .to_NA_1s(Tile_X9Y9_to_NA_1s),
    .to_NB_1s(Tile_X9Y9_to_NB_1s),
    .to_NC_1s(Tile_X9Y9_to_NC_1s),
    .to_ND_1s(Tile_X9Y9_to_ND_1s),
    .to_NF_1s(Tile_X9Y9_to_NF_1s),
    .to_NG_1s(Tile_X9Y9_to_NG_1s),
    .to_NH_1s(Tile_X9Y9_to_NH_1s),
    .to_NI_1s(Tile_X9Y9_to_NI_1s),
    .to_SA_1s(Tile_X9Y9_to_SA_1s),
    .to_SB_1s(Tile_X9Y9_to_SB_1s),
    .to_SC_1s(Tile_X9Y9_to_SC_1s),
    .to_SD_1s(Tile_X9Y9_to_SD_1s),
    .to_SF_1s(Tile_X9Y9_to_SF_1s),
    .to_SG_1s(Tile_X9Y9_to_SG_1s),
    .to_SH_1s(Tile_X9Y9_to_SH_1s),
    .to_SI_1s(Tile_X9Y9_to_SI_1s),
    .F_ctrl(Tile_X9Y9_F_ctrl),
    .UserCLK(Tile_X9Y10_UserCLKo),
    .UserCLKo(Tile_X9Y9_UserCLKo),
    .rst(Tile_X9Y10_rsto),
    .rsto(Tile_X9Y9_rsto),
    .FrameData(Tile_X8Y9_FrameData_O),
    .FrameData_O(Tile_X9Y9_FrameData_O),
    .FrameStrobe(Tile_X9Y10_FrameStrobe_O),
    .FrameStrobe_O(Tile_X9Y9_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
ctrl_IO
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X10Y9_Emulate_Bitstream)
    )
`endif
    Tile_X10Y9_ctrl_IO
    (
    .from_EA_1s(Tile_X9Y9_to_EA_1s),
    .from_EB_1s(Tile_X9Y9_to_EB_1s),
    .from_EC_1s(Tile_X9Y9_to_EC_1s),
    .from_ED_1s(Tile_X9Y9_to_ED_1s),
    .from_EF_1s(Tile_X9Y9_to_EF_1s),
    .from_EG_1s(Tile_X9Y9_to_EG_1s),
    .from_EH_1s(Tile_X9Y9_to_EH_1s),
    .from_EI_1s(Tile_X9Y9_to_EI_1s),
    .to_WA_1s(Tile_X10Y9_to_WA_1s),
    .to_WB_1s(Tile_X10Y9_to_WB_1s),
    .to_WC_1s(Tile_X10Y9_to_WC_1s),
    .to_WD_1s(Tile_X10Y9_to_WD_1s),
    .to_WF_1s(Tile_X10Y9_to_WF_1s),
    .to_WG_1s(Tile_X10Y9_to_WG_1s),
    .to_WH_1s(Tile_X10Y9_to_WH_1s),
    .to_WI_1s(Tile_X10Y9_to_WI_1s),
    .A_O_top_0_t(Tile_X10Y9_A_O_top_0_t),
    .A_O_top_0_f(Tile_X10Y9_A_O_top_0_f),
    .A_prech2(Tile_X10Y9_A_prech2),
    .A_DR_fault(Tile_X10Y9_A_DR_fault),
    .A_I_top_0_t(Tile_X10Y9_A_I_top_0_t),
    .A_I_top_0_f(Tile_X10Y9_A_I_top_0_f),
    .A_T_top(Tile_X10Y9_A_T_top),
    .A_F_ctrl(Tile_X10Y9_A_F_ctrl),
    .UserCLK(Tile_X10Y10_UserCLKo),
    .UserCLKo(Tile_X10Y9_UserCLKo),
    .rst(Tile_X10Y10_rsto),
    .rsto(Tile_X10Y9_rsto),
    .FrameData(Tile_X9Y9_FrameData_O),
    .FrameData_O(Tile_X10Y9_FrameData_O),
    .FrameStrobe(Tile_X10Y10_FrameStrobe_O),
    .FrameStrobe_O(Tile_X10Y9_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
W_IO_custom
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X0Y10_Emulate_Bitstream)
    )
`endif
    Tile_X0Y10_W_IO_custom
    (
    .from_NA(Tile_X0Y11_to_NA),
    .from_NB(Tile_X0Y11_to_NB),
    .from_NC(Tile_X0Y11_to_NC),
    .from_ND(Tile_X0Y11_to_ND),
    .from_NF(Tile_X0Y11_to_NF),
    .from_NG(Tile_X0Y11_to_NG),
    .from_NH(Tile_X0Y11_to_NH),
    .from_NI(Tile_X0Y11_to_NI),
    .from_SA(Tile_X0Y9_to_SA),
    .from_SB(Tile_X0Y9_to_SB),
    .from_SC(Tile_X0Y9_to_SC),
    .from_SD(Tile_X0Y9_to_SD),
    .from_SF(Tile_X0Y9_to_SF),
    .from_SG(Tile_X0Y9_to_SG),
    .from_SH(Tile_X0Y9_to_SH),
    .from_SI(Tile_X0Y9_to_SI),
    .from_WA(Tile_X1Y10_to_WA),
    .from_WB(Tile_X1Y10_to_WB),
    .from_WC(Tile_X1Y10_to_WC),
    .from_WD(Tile_X1Y10_to_WD),
    .from_WF(Tile_X1Y10_to_WF),
    .from_WG(Tile_X1Y10_to_WG),
    .from_WH(Tile_X1Y10_to_WH),
    .from_WI(Tile_X1Y10_to_WI),
    .to_EA(Tile_X0Y10_to_EA),
    .to_EB(Tile_X0Y10_to_EB),
    .to_EC(Tile_X0Y10_to_EC),
    .to_ED(Tile_X0Y10_to_ED),
    .to_EF(Tile_X0Y10_to_EF),
    .to_EG(Tile_X0Y10_to_EG),
    .to_EH(Tile_X0Y10_to_EH),
    .to_EI(Tile_X0Y10_to_EI),
    .to_NA(Tile_X0Y10_to_NA),
    .to_NB(Tile_X0Y10_to_NB),
    .to_NC(Tile_X0Y10_to_NC),
    .to_ND(Tile_X0Y10_to_ND),
    .to_NF(Tile_X0Y10_to_NF),
    .to_NG(Tile_X0Y10_to_NG),
    .to_NH(Tile_X0Y10_to_NH),
    .to_NI(Tile_X0Y10_to_NI),
    .to_SA(Tile_X0Y10_to_SA),
    .to_SB(Tile_X0Y10_to_SB),
    .to_SC(Tile_X0Y10_to_SC),
    .to_SD(Tile_X0Y10_to_SD),
    .to_SF(Tile_X0Y10_to_SF),
    .to_SG(Tile_X0Y10_to_SG),
    .to_SH(Tile_X0Y10_to_SH),
    .to_SI(Tile_X0Y10_to_SI),
    .A_O_top_0_t(Tile_X0Y10_A_O_top_0_t),
    .A_O_top_0_f(Tile_X0Y10_A_O_top_0_f),
    .A_O_top_1_t(Tile_X0Y10_A_O_top_1_t),
    .A_O_top_1_f(Tile_X0Y10_A_O_top_1_f),
    .A_prech1(Tile_X0Y10_A_prech1),
    .A_prech2(Tile_X0Y10_A_prech2),
    .A_DR_fault(Tile_X0Y10_A_DR_fault),
    .A_I_top_0_t(Tile_X0Y10_A_I_top_0_t),
    .A_I_top_0_f(Tile_X0Y10_A_I_top_0_f),
    .A_I_top_1_t(Tile_X0Y10_A_I_top_1_t),
    .A_I_top_1_f(Tile_X0Y10_A_I_top_1_f),
    .A_T_top(Tile_X0Y10_A_T_top),
    .A_F_masked1(Tile_X0Y10_A_F_masked1),
    .A_F_masked2(Tile_X0Y10_A_F_masked2),
    .A_config_C_bit0(Tile_X0Y10_A_config_C_bit0),
    .A_config_C_bit1(Tile_X0Y10_A_config_C_bit1),
    .A_config_C_bit2(Tile_X0Y10_A_config_C_bit2),
    .A_config_C_bit3(Tile_X0Y10_A_config_C_bit3),
    .B_config_C_bit0(Tile_X0Y10_B_config_C_bit0),
    .B_config_C_bit1(Tile_X0Y10_B_config_C_bit1),
    .B_config_C_bit2(Tile_X0Y10_B_config_C_bit2),
    .B_config_C_bit3(Tile_X0Y10_B_config_C_bit3),
    .UserCLK(Tile_X0Y11_UserCLKo),
    .UserCLKo(Tile_X0Y10_UserCLKo),
    .rst(Tile_X0Y11_rsto),
    .rsto(Tile_X0Y10_rsto),
    .FrameData(Tile_Y10_FrameData),
    .FrameData_O(Tile_X0Y10_FrameData_O),
    .FrameStrobe(Tile_X0Y11_FrameStrobe_O),
    .FrameStrobe_O(Tile_X0Y10_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X1Y10_Emulate_Bitstream)
    )
`endif
    Tile_X1Y10_linear_LMDPL
    (
    .from_NA(Tile_X1Y11_to_NA),
    .from_NB(Tile_X1Y11_to_NB),
    .from_NC(Tile_X1Y11_to_NC),
    .from_ND(Tile_X1Y11_to_ND),
    .from_NF(Tile_X1Y11_to_NF),
    .from_NG(Tile_X1Y11_to_NG),
    .from_NH(Tile_X1Y11_to_NH),
    .from_NI(Tile_X1Y11_to_NI),
    .from_EA(Tile_X0Y10_to_EA),
    .from_EB(Tile_X0Y10_to_EB),
    .from_EC(Tile_X0Y10_to_EC),
    .from_ED(Tile_X0Y10_to_ED),
    .from_EF(Tile_X0Y10_to_EF),
    .from_EG(Tile_X0Y10_to_EG),
    .from_EH(Tile_X0Y10_to_EH),
    .from_EI(Tile_X0Y10_to_EI),
    .from_SA(Tile_X1Y9_to_SA),
    .from_SB(Tile_X1Y9_to_SB),
    .from_SC(Tile_X1Y9_to_SC),
    .from_SD(Tile_X1Y9_to_SD),
    .from_SF(Tile_X1Y9_to_SF),
    .from_SG(Tile_X1Y9_to_SG),
    .from_SH(Tile_X1Y9_to_SH),
    .from_SI(Tile_X1Y9_to_SI),
    .from_WA(Tile_X2Y10_to_WA),
    .from_WB(Tile_X2Y10_to_WB),
    .from_WC(Tile_X2Y10_to_WC),
    .from_WD(Tile_X2Y10_to_WD),
    .from_WF(Tile_X2Y10_to_WF),
    .from_WG(Tile_X2Y10_to_WG),
    .from_WH(Tile_X2Y10_to_WH),
    .from_WI(Tile_X2Y10_to_WI),
    .to_EA(Tile_X1Y10_to_EA),
    .to_EB(Tile_X1Y10_to_EB),
    .to_EC(Tile_X1Y10_to_EC),
    .to_ED(Tile_X1Y10_to_ED),
    .to_EF(Tile_X1Y10_to_EF),
    .to_EG(Tile_X1Y10_to_EG),
    .to_EH(Tile_X1Y10_to_EH),
    .to_EI(Tile_X1Y10_to_EI),
    .to_WA(Tile_X1Y10_to_WA),
    .to_WB(Tile_X1Y10_to_WB),
    .to_WC(Tile_X1Y10_to_WC),
    .to_WD(Tile_X1Y10_to_WD),
    .to_WF(Tile_X1Y10_to_WF),
    .to_WG(Tile_X1Y10_to_WG),
    .to_WH(Tile_X1Y10_to_WH),
    .to_WI(Tile_X1Y10_to_WI),
    .to_NA(Tile_X1Y10_to_NA),
    .to_NB(Tile_X1Y10_to_NB),
    .to_NC(Tile_X1Y10_to_NC),
    .to_ND(Tile_X1Y10_to_ND),
    .to_NF(Tile_X1Y10_to_NF),
    .to_NG(Tile_X1Y10_to_NG),
    .to_NH(Tile_X1Y10_to_NH),
    .to_NI(Tile_X1Y10_to_NI),
    .to_SA(Tile_X1Y10_to_SA),
    .to_SB(Tile_X1Y10_to_SB),
    .to_SC(Tile_X1Y10_to_SC),
    .to_SD(Tile_X1Y10_to_SD),
    .to_SF(Tile_X1Y10_to_SF),
    .to_SG(Tile_X1Y10_to_SG),
    .to_SH(Tile_X1Y10_to_SH),
    .to_SI(Tile_X1Y10_to_SI),
    .F_masked1(Tile_X1Y10_F_masked1),
    .F_masked2(Tile_X1Y10_F_masked2),
    .UserCLK(Tile_X1Y11_UserCLKo),
    .UserCLKo(Tile_X1Y10_UserCLKo),
    .rst(Tile_X1Y11_rsto),
    .rsto(Tile_X1Y10_rsto),
    .FrameData(Tile_X0Y10_FrameData_O),
    .FrameData_O(Tile_X1Y10_FrameData_O),
    .FrameStrobe(Tile_X1Y11_FrameStrobe_O),
    .FrameStrobe_O(Tile_X1Y10_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X2Y10_Emulate_Bitstream)
    )
`endif
    Tile_X2Y10_linear_LMDPL
    (
    .from_NA(Tile_X2Y11_to_NA),
    .from_NB(Tile_X2Y11_to_NB),
    .from_NC(Tile_X2Y11_to_NC),
    .from_ND(Tile_X2Y11_to_ND),
    .from_NF(Tile_X2Y11_to_NF),
    .from_NG(Tile_X2Y11_to_NG),
    .from_NH(Tile_X2Y11_to_NH),
    .from_NI(Tile_X2Y11_to_NI),
    .from_EA(Tile_X1Y10_to_EA),
    .from_EB(Tile_X1Y10_to_EB),
    .from_EC(Tile_X1Y10_to_EC),
    .from_ED(Tile_X1Y10_to_ED),
    .from_EF(Tile_X1Y10_to_EF),
    .from_EG(Tile_X1Y10_to_EG),
    .from_EH(Tile_X1Y10_to_EH),
    .from_EI(Tile_X1Y10_to_EI),
    .from_SA(Tile_X2Y9_to_SA),
    .from_SB(Tile_X2Y9_to_SB),
    .from_SC(Tile_X2Y9_to_SC),
    .from_SD(Tile_X2Y9_to_SD),
    .from_SF(Tile_X2Y9_to_SF),
    .from_SG(Tile_X2Y9_to_SG),
    .from_SH(Tile_X2Y9_to_SH),
    .from_SI(Tile_X2Y9_to_SI),
    .from_WA(Tile_X3Y10_to_WA),
    .from_WB(Tile_X3Y10_to_WB),
    .from_WC(Tile_X3Y10_to_WC),
    .from_WD(Tile_X3Y10_to_WD),
    .from_WF(Tile_X3Y10_to_WF),
    .from_WG(Tile_X3Y10_to_WG),
    .from_WH(Tile_X3Y10_to_WH),
    .from_WI(Tile_X3Y10_to_WI),
    .to_EA(Tile_X2Y10_to_EA),
    .to_EB(Tile_X2Y10_to_EB),
    .to_EC(Tile_X2Y10_to_EC),
    .to_ED(Tile_X2Y10_to_ED),
    .to_EF(Tile_X2Y10_to_EF),
    .to_EG(Tile_X2Y10_to_EG),
    .to_EH(Tile_X2Y10_to_EH),
    .to_EI(Tile_X2Y10_to_EI),
    .to_WA(Tile_X2Y10_to_WA),
    .to_WB(Tile_X2Y10_to_WB),
    .to_WC(Tile_X2Y10_to_WC),
    .to_WD(Tile_X2Y10_to_WD),
    .to_WF(Tile_X2Y10_to_WF),
    .to_WG(Tile_X2Y10_to_WG),
    .to_WH(Tile_X2Y10_to_WH),
    .to_WI(Tile_X2Y10_to_WI),
    .to_NA(Tile_X2Y10_to_NA),
    .to_NB(Tile_X2Y10_to_NB),
    .to_NC(Tile_X2Y10_to_NC),
    .to_ND(Tile_X2Y10_to_ND),
    .to_NF(Tile_X2Y10_to_NF),
    .to_NG(Tile_X2Y10_to_NG),
    .to_NH(Tile_X2Y10_to_NH),
    .to_NI(Tile_X2Y10_to_NI),
    .to_SA(Tile_X2Y10_to_SA),
    .to_SB(Tile_X2Y10_to_SB),
    .to_SC(Tile_X2Y10_to_SC),
    .to_SD(Tile_X2Y10_to_SD),
    .to_SF(Tile_X2Y10_to_SF),
    .to_SG(Tile_X2Y10_to_SG),
    .to_SH(Tile_X2Y10_to_SH),
    .to_SI(Tile_X2Y10_to_SI),
    .F_masked1(Tile_X2Y10_F_masked1),
    .F_masked2(Tile_X2Y10_F_masked2),
    .UserCLK(Tile_X2Y11_UserCLKo),
    .UserCLKo(Tile_X2Y10_UserCLKo),
    .rst(Tile_X2Y11_rsto),
    .rsto(Tile_X2Y10_rsto),
    .FrameData(Tile_X1Y10_FrameData_O),
    .FrameData_O(Tile_X2Y10_FrameData_O),
    .FrameStrobe(Tile_X2Y11_FrameStrobe_O),
    .FrameStrobe_O(Tile_X2Y10_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
nonlinear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X3Y10_Emulate_Bitstream)
    )
`endif
    Tile_X3Y10_nonlinear_LMDPL
    (
    .from_NA(Tile_X3Y11_to_NA),
    .from_NB(Tile_X3Y11_to_NB),
    .from_NC(Tile_X3Y11_to_NC),
    .from_ND(Tile_X3Y11_to_ND),
    .from_NF(Tile_X3Y11_to_NF),
    .from_NG(Tile_X3Y11_to_NG),
    .from_NH(Tile_X3Y11_to_NH),
    .from_NI(Tile_X3Y11_to_NI),
    .from_EA(Tile_X2Y10_to_EA),
    .from_EB(Tile_X2Y10_to_EB),
    .from_EC(Tile_X2Y10_to_EC),
    .from_ED(Tile_X2Y10_to_ED),
    .from_EF(Tile_X2Y10_to_EF),
    .from_EG(Tile_X2Y10_to_EG),
    .from_EH(Tile_X2Y10_to_EH),
    .from_EI(Tile_X2Y10_to_EI),
    .from_SA(Tile_X3Y9_to_SA),
    .from_SB(Tile_X3Y9_to_SB),
    .from_SC(Tile_X3Y9_to_SC),
    .from_SD(Tile_X3Y9_to_SD),
    .from_SF(Tile_X3Y9_to_SF),
    .from_SG(Tile_X3Y9_to_SG),
    .from_SH(Tile_X3Y9_to_SH),
    .from_SI(Tile_X3Y9_to_SI),
    .from_WA(Tile_X4Y10_to_WA),
    .from_WB(Tile_X4Y10_to_WB),
    .from_WC(Tile_X4Y10_to_WC),
    .from_WD(Tile_X4Y10_to_WD),
    .from_WF(Tile_X4Y10_to_WF),
    .from_WG(Tile_X4Y10_to_WG),
    .from_WH(Tile_X4Y10_to_WH),
    .from_WI(Tile_X4Y10_to_WI),
    .to_EA(Tile_X3Y10_to_EA),
    .to_EB(Tile_X3Y10_to_EB),
    .to_EC(Tile_X3Y10_to_EC),
    .to_ED(Tile_X3Y10_to_ED),
    .to_EF(Tile_X3Y10_to_EF),
    .to_EG(Tile_X3Y10_to_EG),
    .to_EH(Tile_X3Y10_to_EH),
    .to_EI(Tile_X3Y10_to_EI),
    .to_WA(Tile_X3Y10_to_WA),
    .to_WB(Tile_X3Y10_to_WB),
    .to_WC(Tile_X3Y10_to_WC),
    .to_WD(Tile_X3Y10_to_WD),
    .to_WF(Tile_X3Y10_to_WF),
    .to_WG(Tile_X3Y10_to_WG),
    .to_WH(Tile_X3Y10_to_WH),
    .to_WI(Tile_X3Y10_to_WI),
    .to_NA(Tile_X3Y10_to_NA),
    .to_NB(Tile_X3Y10_to_NB),
    .to_NC(Tile_X3Y10_to_NC),
    .to_ND(Tile_X3Y10_to_ND),
    .to_NF(Tile_X3Y10_to_NF),
    .to_NG(Tile_X3Y10_to_NG),
    .to_NH(Tile_X3Y10_to_NH),
    .to_NI(Tile_X3Y10_to_NI),
    .to_SA(Tile_X3Y10_to_SA),
    .to_SB(Tile_X3Y10_to_SB),
    .to_SC(Tile_X3Y10_to_SC),
    .to_SD(Tile_X3Y10_to_SD),
    .to_SF(Tile_X3Y10_to_SF),
    .to_SG(Tile_X3Y10_to_SG),
    .to_SH(Tile_X3Y10_to_SH),
    .to_SI(Tile_X3Y10_to_SI),
    .R_t(Tile_X3Y10_R_t),
    .R_f(Tile_X3Y10_R_f),
    .F_masked1(Tile_X3Y10_F_masked1),
    .F_masked2(Tile_X3Y10_F_masked2),
    .UserCLK(Tile_X3Y11_UserCLKo),
    .UserCLKo(Tile_X3Y10_UserCLKo),
    .rst(Tile_X3Y11_rsto),
    .rsto(Tile_X3Y10_rsto),
    .FrameData(Tile_X2Y10_FrameData_O),
    .FrameData_O(Tile_X3Y10_FrameData_O),
    .FrameStrobe(Tile_X3Y11_FrameStrobe_O),
    .FrameStrobe_O(Tile_X3Y10_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X4Y10_Emulate_Bitstream)
    )
`endif
    Tile_X4Y10_linear_LMDPL
    (
    .from_NA(Tile_X4Y11_to_NA),
    .from_NB(Tile_X4Y11_to_NB),
    .from_NC(Tile_X4Y11_to_NC),
    .from_ND(Tile_X4Y11_to_ND),
    .from_NF(Tile_X4Y11_to_NF),
    .from_NG(Tile_X4Y11_to_NG),
    .from_NH(Tile_X4Y11_to_NH),
    .from_NI(Tile_X4Y11_to_NI),
    .from_EA(Tile_X3Y10_to_EA),
    .from_EB(Tile_X3Y10_to_EB),
    .from_EC(Tile_X3Y10_to_EC),
    .from_ED(Tile_X3Y10_to_ED),
    .from_EF(Tile_X3Y10_to_EF),
    .from_EG(Tile_X3Y10_to_EG),
    .from_EH(Tile_X3Y10_to_EH),
    .from_EI(Tile_X3Y10_to_EI),
    .from_SA(Tile_X4Y9_to_SA),
    .from_SB(Tile_X4Y9_to_SB),
    .from_SC(Tile_X4Y9_to_SC),
    .from_SD(Tile_X4Y9_to_SD),
    .from_SF(Tile_X4Y9_to_SF),
    .from_SG(Tile_X4Y9_to_SG),
    .from_SH(Tile_X4Y9_to_SH),
    .from_SI(Tile_X4Y9_to_SI),
    .from_WA(Tile_X5Y10_to_WA),
    .from_WB(Tile_X5Y10_to_WB),
    .from_WC(Tile_X5Y10_to_WC),
    .from_WD(Tile_X5Y10_to_WD),
    .from_WF(Tile_X5Y10_to_WF),
    .from_WG(Tile_X5Y10_to_WG),
    .from_WH(Tile_X5Y10_to_WH),
    .from_WI(Tile_X5Y10_to_WI),
    .to_EA(Tile_X4Y10_to_EA),
    .to_EB(Tile_X4Y10_to_EB),
    .to_EC(Tile_X4Y10_to_EC),
    .to_ED(Tile_X4Y10_to_ED),
    .to_EF(Tile_X4Y10_to_EF),
    .to_EG(Tile_X4Y10_to_EG),
    .to_EH(Tile_X4Y10_to_EH),
    .to_EI(Tile_X4Y10_to_EI),
    .to_WA(Tile_X4Y10_to_WA),
    .to_WB(Tile_X4Y10_to_WB),
    .to_WC(Tile_X4Y10_to_WC),
    .to_WD(Tile_X4Y10_to_WD),
    .to_WF(Tile_X4Y10_to_WF),
    .to_WG(Tile_X4Y10_to_WG),
    .to_WH(Tile_X4Y10_to_WH),
    .to_WI(Tile_X4Y10_to_WI),
    .to_NA(Tile_X4Y10_to_NA),
    .to_NB(Tile_X4Y10_to_NB),
    .to_NC(Tile_X4Y10_to_NC),
    .to_ND(Tile_X4Y10_to_ND),
    .to_NF(Tile_X4Y10_to_NF),
    .to_NG(Tile_X4Y10_to_NG),
    .to_NH(Tile_X4Y10_to_NH),
    .to_NI(Tile_X4Y10_to_NI),
    .to_SA(Tile_X4Y10_to_SA),
    .to_SB(Tile_X4Y10_to_SB),
    .to_SC(Tile_X4Y10_to_SC),
    .to_SD(Tile_X4Y10_to_SD),
    .to_SF(Tile_X4Y10_to_SF),
    .to_SG(Tile_X4Y10_to_SG),
    .to_SH(Tile_X4Y10_to_SH),
    .to_SI(Tile_X4Y10_to_SI),
    .F_masked1(Tile_X4Y10_F_masked1),
    .F_masked2(Tile_X4Y10_F_masked2),
    .UserCLK(Tile_X4Y11_UserCLKo),
    .UserCLKo(Tile_X4Y10_UserCLKo),
    .rst(Tile_X4Y11_rsto),
    .rsto(Tile_X4Y10_rsto),
    .FrameData(Tile_X3Y10_FrameData_O),
    .FrameData_O(Tile_X4Y10_FrameData_O),
    .FrameStrobe(Tile_X4Y11_FrameStrobe_O),
    .FrameStrobe_O(Tile_X4Y10_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X5Y10_Emulate_Bitstream)
    )
`endif
    Tile_X5Y10_linear_LMDPL
    (
    .from_NA(Tile_X5Y11_to_NA),
    .from_NB(Tile_X5Y11_to_NB),
    .from_NC(Tile_X5Y11_to_NC),
    .from_ND(Tile_X5Y11_to_ND),
    .from_NF(Tile_X5Y11_to_NF),
    .from_NG(Tile_X5Y11_to_NG),
    .from_NH(Tile_X5Y11_to_NH),
    .from_NI(Tile_X5Y11_to_NI),
    .from_EA(Tile_X4Y10_to_EA),
    .from_EB(Tile_X4Y10_to_EB),
    .from_EC(Tile_X4Y10_to_EC),
    .from_ED(Tile_X4Y10_to_ED),
    .from_EF(Tile_X4Y10_to_EF),
    .from_EG(Tile_X4Y10_to_EG),
    .from_EH(Tile_X4Y10_to_EH),
    .from_EI(Tile_X4Y10_to_EI),
    .from_SA(Tile_X5Y9_to_SA),
    .from_SB(Tile_X5Y9_to_SB),
    .from_SC(Tile_X5Y9_to_SC),
    .from_SD(Tile_X5Y9_to_SD),
    .from_SF(Tile_X5Y9_to_SF),
    .from_SG(Tile_X5Y9_to_SG),
    .from_SH(Tile_X5Y9_to_SH),
    .from_SI(Tile_X5Y9_to_SI),
    .from_WA(Tile_X6Y10_to_WA),
    .from_WB(Tile_X6Y10_to_WB),
    .from_WC(Tile_X6Y10_to_WC),
    .from_WD(Tile_X6Y10_to_WD),
    .from_WF(Tile_X6Y10_to_WF),
    .from_WG(Tile_X6Y10_to_WG),
    .from_WH(Tile_X6Y10_to_WH),
    .from_WI(Tile_X6Y10_to_WI),
    .to_EA(Tile_X5Y10_to_EA),
    .to_EB(Tile_X5Y10_to_EB),
    .to_EC(Tile_X5Y10_to_EC),
    .to_ED(Tile_X5Y10_to_ED),
    .to_EF(Tile_X5Y10_to_EF),
    .to_EG(Tile_X5Y10_to_EG),
    .to_EH(Tile_X5Y10_to_EH),
    .to_EI(Tile_X5Y10_to_EI),
    .to_WA(Tile_X5Y10_to_WA),
    .to_WB(Tile_X5Y10_to_WB),
    .to_WC(Tile_X5Y10_to_WC),
    .to_WD(Tile_X5Y10_to_WD),
    .to_WF(Tile_X5Y10_to_WF),
    .to_WG(Tile_X5Y10_to_WG),
    .to_WH(Tile_X5Y10_to_WH),
    .to_WI(Tile_X5Y10_to_WI),
    .to_NA(Tile_X5Y10_to_NA),
    .to_NB(Tile_X5Y10_to_NB),
    .to_NC(Tile_X5Y10_to_NC),
    .to_ND(Tile_X5Y10_to_ND),
    .to_NF(Tile_X5Y10_to_NF),
    .to_NG(Tile_X5Y10_to_NG),
    .to_NH(Tile_X5Y10_to_NH),
    .to_NI(Tile_X5Y10_to_NI),
    .to_SA(Tile_X5Y10_to_SA),
    .to_SB(Tile_X5Y10_to_SB),
    .to_SC(Tile_X5Y10_to_SC),
    .to_SD(Tile_X5Y10_to_SD),
    .to_SF(Tile_X5Y10_to_SF),
    .to_SG(Tile_X5Y10_to_SG),
    .to_SH(Tile_X5Y10_to_SH),
    .to_SI(Tile_X5Y10_to_SI),
    .F_masked1(Tile_X5Y10_F_masked1),
    .F_masked2(Tile_X5Y10_F_masked2),
    .UserCLK(Tile_X5Y11_UserCLKo),
    .UserCLKo(Tile_X5Y10_UserCLKo),
    .rst(Tile_X5Y11_rsto),
    .rsto(Tile_X5Y10_rsto),
    .FrameData(Tile_X4Y10_FrameData_O),
    .FrameData_O(Tile_X5Y10_FrameData_O),
    .FrameStrobe(Tile_X5Y11_FrameStrobe_O),
    .FrameStrobe_O(Tile_X5Y10_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
nonlinear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X6Y10_Emulate_Bitstream)
    )
`endif
    Tile_X6Y10_nonlinear_LMDPL
    (
    .from_NA(Tile_X6Y11_to_NA),
    .from_NB(Tile_X6Y11_to_NB),
    .from_NC(Tile_X6Y11_to_NC),
    .from_ND(Tile_X6Y11_to_ND),
    .from_NF(Tile_X6Y11_to_NF),
    .from_NG(Tile_X6Y11_to_NG),
    .from_NH(Tile_X6Y11_to_NH),
    .from_NI(Tile_X6Y11_to_NI),
    .from_EA(Tile_X5Y10_to_EA),
    .from_EB(Tile_X5Y10_to_EB),
    .from_EC(Tile_X5Y10_to_EC),
    .from_ED(Tile_X5Y10_to_ED),
    .from_EF(Tile_X5Y10_to_EF),
    .from_EG(Tile_X5Y10_to_EG),
    .from_EH(Tile_X5Y10_to_EH),
    .from_EI(Tile_X5Y10_to_EI),
    .from_SA(Tile_X6Y9_to_SA),
    .from_SB(Tile_X6Y9_to_SB),
    .from_SC(Tile_X6Y9_to_SC),
    .from_SD(Tile_X6Y9_to_SD),
    .from_SF(Tile_X6Y9_to_SF),
    .from_SG(Tile_X6Y9_to_SG),
    .from_SH(Tile_X6Y9_to_SH),
    .from_SI(Tile_X6Y9_to_SI),
    .from_WA(Tile_X7Y10_to_WA),
    .from_WB(Tile_X7Y10_to_WB),
    .from_WC(Tile_X7Y10_to_WC),
    .from_WD(Tile_X7Y10_to_WD),
    .from_WF(Tile_X7Y10_to_WF),
    .from_WG(Tile_X7Y10_to_WG),
    .from_WH(Tile_X7Y10_to_WH),
    .from_WI(Tile_X7Y10_to_WI),
    .to_EA(Tile_X6Y10_to_EA),
    .to_EB(Tile_X6Y10_to_EB),
    .to_EC(Tile_X6Y10_to_EC),
    .to_ED(Tile_X6Y10_to_ED),
    .to_EF(Tile_X6Y10_to_EF),
    .to_EG(Tile_X6Y10_to_EG),
    .to_EH(Tile_X6Y10_to_EH),
    .to_EI(Tile_X6Y10_to_EI),
    .to_WA(Tile_X6Y10_to_WA),
    .to_WB(Tile_X6Y10_to_WB),
    .to_WC(Tile_X6Y10_to_WC),
    .to_WD(Tile_X6Y10_to_WD),
    .to_WF(Tile_X6Y10_to_WF),
    .to_WG(Tile_X6Y10_to_WG),
    .to_WH(Tile_X6Y10_to_WH),
    .to_WI(Tile_X6Y10_to_WI),
    .to_NA(Tile_X6Y10_to_NA),
    .to_NB(Tile_X6Y10_to_NB),
    .to_NC(Tile_X6Y10_to_NC),
    .to_ND(Tile_X6Y10_to_ND),
    .to_NF(Tile_X6Y10_to_NF),
    .to_NG(Tile_X6Y10_to_NG),
    .to_NH(Tile_X6Y10_to_NH),
    .to_NI(Tile_X6Y10_to_NI),
    .to_SA(Tile_X6Y10_to_SA),
    .to_SB(Tile_X6Y10_to_SB),
    .to_SC(Tile_X6Y10_to_SC),
    .to_SD(Tile_X6Y10_to_SD),
    .to_SF(Tile_X6Y10_to_SF),
    .to_SG(Tile_X6Y10_to_SG),
    .to_SH(Tile_X6Y10_to_SH),
    .to_SI(Tile_X6Y10_to_SI),
    .R_t(Tile_X6Y10_R_t),
    .R_f(Tile_X6Y10_R_f),
    .F_masked1(Tile_X6Y10_F_masked1),
    .F_masked2(Tile_X6Y10_F_masked2),
    .UserCLK(Tile_X6Y11_UserCLKo),
    .UserCLKo(Tile_X6Y10_UserCLKo),
    .rst(Tile_X6Y11_rsto),
    .rsto(Tile_X6Y10_rsto),
    .FrameData(Tile_X5Y10_FrameData_O),
    .FrameData_O(Tile_X6Y10_FrameData_O),
    .FrameStrobe(Tile_X6Y11_FrameStrobe_O),
    .FrameStrobe_O(Tile_X6Y10_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X7Y10_Emulate_Bitstream)
    )
`endif
    Tile_X7Y10_linear_LMDPL
    (
    .from_NA(Tile_X7Y11_to_NA),
    .from_NB(Tile_X7Y11_to_NB),
    .from_NC(Tile_X7Y11_to_NC),
    .from_ND(Tile_X7Y11_to_ND),
    .from_NF(Tile_X7Y11_to_NF),
    .from_NG(Tile_X7Y11_to_NG),
    .from_NH(Tile_X7Y11_to_NH),
    .from_NI(Tile_X7Y11_to_NI),
    .from_EA(Tile_X6Y10_to_EA),
    .from_EB(Tile_X6Y10_to_EB),
    .from_EC(Tile_X6Y10_to_EC),
    .from_ED(Tile_X6Y10_to_ED),
    .from_EF(Tile_X6Y10_to_EF),
    .from_EG(Tile_X6Y10_to_EG),
    .from_EH(Tile_X6Y10_to_EH),
    .from_EI(Tile_X6Y10_to_EI),
    .from_SA(Tile_X7Y9_to_SA),
    .from_SB(Tile_X7Y9_to_SB),
    .from_SC(Tile_X7Y9_to_SC),
    .from_SD(Tile_X7Y9_to_SD),
    .from_SF(Tile_X7Y9_to_SF),
    .from_SG(Tile_X7Y9_to_SG),
    .from_SH(Tile_X7Y9_to_SH),
    .from_SI(Tile_X7Y9_to_SI),
    .from_WA(Tile_X8Y10_to_WA),
    .from_WB(Tile_X8Y10_to_WB),
    .from_WC(Tile_X8Y10_to_WC),
    .from_WD(Tile_X8Y10_to_WD),
    .from_WF(Tile_X8Y10_to_WF),
    .from_WG(Tile_X8Y10_to_WG),
    .from_WH(Tile_X8Y10_to_WH),
    .from_WI(Tile_X8Y10_to_WI),
    .to_EA(Tile_X7Y10_to_EA),
    .to_EB(Tile_X7Y10_to_EB),
    .to_EC(Tile_X7Y10_to_EC),
    .to_ED(Tile_X7Y10_to_ED),
    .to_EF(Tile_X7Y10_to_EF),
    .to_EG(Tile_X7Y10_to_EG),
    .to_EH(Tile_X7Y10_to_EH),
    .to_EI(Tile_X7Y10_to_EI),
    .to_WA(Tile_X7Y10_to_WA),
    .to_WB(Tile_X7Y10_to_WB),
    .to_WC(Tile_X7Y10_to_WC),
    .to_WD(Tile_X7Y10_to_WD),
    .to_WF(Tile_X7Y10_to_WF),
    .to_WG(Tile_X7Y10_to_WG),
    .to_WH(Tile_X7Y10_to_WH),
    .to_WI(Tile_X7Y10_to_WI),
    .to_NA(Tile_X7Y10_to_NA),
    .to_NB(Tile_X7Y10_to_NB),
    .to_NC(Tile_X7Y10_to_NC),
    .to_ND(Tile_X7Y10_to_ND),
    .to_NF(Tile_X7Y10_to_NF),
    .to_NG(Tile_X7Y10_to_NG),
    .to_NH(Tile_X7Y10_to_NH),
    .to_NI(Tile_X7Y10_to_NI),
    .to_SA(Tile_X7Y10_to_SA),
    .to_SB(Tile_X7Y10_to_SB),
    .to_SC(Tile_X7Y10_to_SC),
    .to_SD(Tile_X7Y10_to_SD),
    .to_SF(Tile_X7Y10_to_SF),
    .to_SG(Tile_X7Y10_to_SG),
    .to_SH(Tile_X7Y10_to_SH),
    .to_SI(Tile_X7Y10_to_SI),
    .F_masked1(Tile_X7Y10_F_masked1),
    .F_masked2(Tile_X7Y10_F_masked2),
    .UserCLK(Tile_X7Y11_UserCLKo),
    .UserCLKo(Tile_X7Y10_UserCLKo),
    .rst(Tile_X7Y11_rsto),
    .rsto(Tile_X7Y10_rsto),
    .FrameData(Tile_X6Y10_FrameData_O),
    .FrameData_O(Tile_X7Y10_FrameData_O),
    .FrameStrobe(Tile_X7Y11_FrameStrobe_O),
    .FrameStrobe_O(Tile_X7Y10_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
ctrl_to_sec
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X8Y10_Emulate_Bitstream)
    )
`endif
    Tile_X8Y10_ctrl_to_sec
    (
    .from_NA(Tile_X8Y11_to_NA),
    .from_NB(Tile_X8Y11_to_NB),
    .from_NC(Tile_X8Y11_to_NC),
    .from_ND(Tile_X8Y11_to_ND),
    .from_NF(Tile_X8Y11_to_NF),
    .from_NG(Tile_X8Y11_to_NG),
    .from_NH(Tile_X8Y11_to_NH),
    .from_NI(Tile_X8Y11_to_NI),
    .from_EA(Tile_X7Y10_to_EA),
    .from_EB(Tile_X7Y10_to_EB),
    .from_EC(Tile_X7Y10_to_EC),
    .from_ED(Tile_X7Y10_to_ED),
    .from_EF(Tile_X7Y10_to_EF),
    .from_EG(Tile_X7Y10_to_EG),
    .from_EH(Tile_X7Y10_to_EH),
    .from_EI(Tile_X7Y10_to_EI),
    .from_SA(Tile_X8Y9_to_SA),
    .from_SB(Tile_X8Y9_to_SB),
    .from_SC(Tile_X8Y9_to_SC),
    .from_SD(Tile_X8Y9_to_SD),
    .from_SF(Tile_X8Y9_to_SF),
    .from_SG(Tile_X8Y9_to_SG),
    .from_SH(Tile_X8Y9_to_SH),
    .from_SI(Tile_X8Y9_to_SI),
    .from_WA_1s(Tile_X9Y10_to_WA_1s),
    .from_WB_1s(Tile_X9Y10_to_WB_1s),
    .from_WC_1s(Tile_X9Y10_to_WC_1s),
    .from_WD_1s(Tile_X9Y10_to_WD_1s),
    .from_WF_1s(Tile_X9Y10_to_WF_1s),
    .from_WG_1s(Tile_X9Y10_to_WG_1s),
    .from_WH_1s(Tile_X9Y10_to_WH_1s),
    .from_WI_1s(Tile_X9Y10_to_WI_1s),
    .to_WA(Tile_X8Y10_to_WA),
    .to_WB(Tile_X8Y10_to_WB),
    .to_WC(Tile_X8Y10_to_WC),
    .to_WD(Tile_X8Y10_to_WD),
    .to_WF(Tile_X8Y10_to_WF),
    .to_WG(Tile_X8Y10_to_WG),
    .to_WH(Tile_X8Y10_to_WH),
    .to_WI(Tile_X8Y10_to_WI),
    .to_NA(Tile_X8Y10_to_NA),
    .to_NB(Tile_X8Y10_to_NB),
    .to_NC(Tile_X8Y10_to_NC),
    .to_ND(Tile_X8Y10_to_ND),
    .to_NF(Tile_X8Y10_to_NF),
    .to_NG(Tile_X8Y10_to_NG),
    .to_NH(Tile_X8Y10_to_NH),
    .to_NI(Tile_X8Y10_to_NI),
    .to_SA(Tile_X8Y10_to_SA),
    .to_SB(Tile_X8Y10_to_SB),
    .to_SC(Tile_X8Y10_to_SC),
    .to_SD(Tile_X8Y10_to_SD),
    .to_SF(Tile_X8Y10_to_SF),
    .to_SG(Tile_X8Y10_to_SG),
    .to_SH(Tile_X8Y10_to_SH),
    .to_SI(Tile_X8Y10_to_SI),
    .UserCLK(Tile_X8Y11_UserCLKo),
    .UserCLKo(Tile_X8Y10_UserCLKo),
    .rst(Tile_X8Y11_rsto),
    .rsto(Tile_X8Y10_rsto),
    .FrameData(Tile_X7Y10_FrameData_O),
    .FrameData_O(Tile_X8Y10_FrameData_O),
    .FrameStrobe(Tile_X8Y11_FrameStrobe_O),
    .FrameStrobe_O(Tile_X8Y10_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
combined_WDDL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X9Y10_Emulate_Bitstream)
    )
`endif
    Tile_X9Y10_combined_WDDL
    (
    .from_NA_1s(Tile_X9Y11_to_NA_1s),
    .from_NB_1s(Tile_X9Y11_to_NB_1s),
    .from_NC_1s(Tile_X9Y11_to_NC_1s),
    .from_ND_1s(Tile_X9Y11_to_ND_1s),
    .from_NF_1s(Tile_X9Y11_to_NF_1s),
    .from_NG_1s(Tile_X9Y11_to_NG_1s),
    .from_NH_1s(Tile_X9Y11_to_NH_1s),
    .from_NI_1s(Tile_X9Y11_to_NI_1s),
    .from_SA_1s(Tile_X9Y9_to_SA_1s),
    .from_SB_1s(Tile_X9Y9_to_SB_1s),
    .from_SC_1s(Tile_X9Y9_to_SC_1s),
    .from_SD_1s(Tile_X9Y9_to_SD_1s),
    .from_SF_1s(Tile_X9Y9_to_SF_1s),
    .from_SG_1s(Tile_X9Y9_to_SG_1s),
    .from_SH_1s(Tile_X9Y9_to_SH_1s),
    .from_SI_1s(Tile_X9Y9_to_SI_1s),
    .from_WA_1s(Tile_X10Y10_to_WA_1s),
    .from_WB_1s(Tile_X10Y10_to_WB_1s),
    .from_WC_1s(Tile_X10Y10_to_WC_1s),
    .from_WD_1s(Tile_X10Y10_to_WD_1s),
    .from_WF_1s(Tile_X10Y10_to_WF_1s),
    .from_WG_1s(Tile_X10Y10_to_WG_1s),
    .from_WH_1s(Tile_X10Y10_to_WH_1s),
    .from_WI_1s(Tile_X10Y10_to_WI_1s),
    .to_EA_1s(Tile_X9Y10_to_EA_1s),
    .to_EB_1s(Tile_X9Y10_to_EB_1s),
    .to_EC_1s(Tile_X9Y10_to_EC_1s),
    .to_ED_1s(Tile_X9Y10_to_ED_1s),
    .to_EF_1s(Tile_X9Y10_to_EF_1s),
    .to_EG_1s(Tile_X9Y10_to_EG_1s),
    .to_EH_1s(Tile_X9Y10_to_EH_1s),
    .to_EI_1s(Tile_X9Y10_to_EI_1s),
    .to_WA_1s(Tile_X9Y10_to_WA_1s),
    .to_WB_1s(Tile_X9Y10_to_WB_1s),
    .to_WC_1s(Tile_X9Y10_to_WC_1s),
    .to_WD_1s(Tile_X9Y10_to_WD_1s),
    .to_WF_1s(Tile_X9Y10_to_WF_1s),
    .to_WG_1s(Tile_X9Y10_to_WG_1s),
    .to_WH_1s(Tile_X9Y10_to_WH_1s),
    .to_WI_1s(Tile_X9Y10_to_WI_1s),
    .to_NA_1s(Tile_X9Y10_to_NA_1s),
    .to_NB_1s(Tile_X9Y10_to_NB_1s),
    .to_NC_1s(Tile_X9Y10_to_NC_1s),
    .to_ND_1s(Tile_X9Y10_to_ND_1s),
    .to_NF_1s(Tile_X9Y10_to_NF_1s),
    .to_NG_1s(Tile_X9Y10_to_NG_1s),
    .to_NH_1s(Tile_X9Y10_to_NH_1s),
    .to_NI_1s(Tile_X9Y10_to_NI_1s),
    .to_SA_1s(Tile_X9Y10_to_SA_1s),
    .to_SB_1s(Tile_X9Y10_to_SB_1s),
    .to_SC_1s(Tile_X9Y10_to_SC_1s),
    .to_SD_1s(Tile_X9Y10_to_SD_1s),
    .to_SF_1s(Tile_X9Y10_to_SF_1s),
    .to_SG_1s(Tile_X9Y10_to_SG_1s),
    .to_SH_1s(Tile_X9Y10_to_SH_1s),
    .to_SI_1s(Tile_X9Y10_to_SI_1s),
    .F_ctrl(Tile_X9Y10_F_ctrl),
    .UserCLK(Tile_X9Y11_UserCLKo),
    .UserCLKo(Tile_X9Y10_UserCLKo),
    .rst(Tile_X9Y11_rsto),
    .rsto(Tile_X9Y10_rsto),
    .FrameData(Tile_X8Y10_FrameData_O),
    .FrameData_O(Tile_X9Y10_FrameData_O),
    .FrameStrobe(Tile_X9Y11_FrameStrobe_O),
    .FrameStrobe_O(Tile_X9Y10_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
ctrl_IO
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X10Y10_Emulate_Bitstream)
    )
`endif
    Tile_X10Y10_ctrl_IO
    (
    .from_EA_1s(Tile_X9Y10_to_EA_1s),
    .from_EB_1s(Tile_X9Y10_to_EB_1s),
    .from_EC_1s(Tile_X9Y10_to_EC_1s),
    .from_ED_1s(Tile_X9Y10_to_ED_1s),
    .from_EF_1s(Tile_X9Y10_to_EF_1s),
    .from_EG_1s(Tile_X9Y10_to_EG_1s),
    .from_EH_1s(Tile_X9Y10_to_EH_1s),
    .from_EI_1s(Tile_X9Y10_to_EI_1s),
    .to_WA_1s(Tile_X10Y10_to_WA_1s),
    .to_WB_1s(Tile_X10Y10_to_WB_1s),
    .to_WC_1s(Tile_X10Y10_to_WC_1s),
    .to_WD_1s(Tile_X10Y10_to_WD_1s),
    .to_WF_1s(Tile_X10Y10_to_WF_1s),
    .to_WG_1s(Tile_X10Y10_to_WG_1s),
    .to_WH_1s(Tile_X10Y10_to_WH_1s),
    .to_WI_1s(Tile_X10Y10_to_WI_1s),
    .A_O_top_0_t(Tile_X10Y10_A_O_top_0_t),
    .A_O_top_0_f(Tile_X10Y10_A_O_top_0_f),
    .A_prech2(Tile_X10Y10_A_prech2),
    .A_DR_fault(Tile_X10Y10_A_DR_fault),
    .A_I_top_0_t(Tile_X10Y10_A_I_top_0_t),
    .A_I_top_0_f(Tile_X10Y10_A_I_top_0_f),
    .A_T_top(Tile_X10Y10_A_T_top),
    .A_F_ctrl(Tile_X10Y10_A_F_ctrl),
    .UserCLK(Tile_X10Y11_UserCLKo),
    .UserCLKo(Tile_X10Y10_UserCLKo),
    .rst(Tile_X10Y11_rsto),
    .rsto(Tile_X10Y10_rsto),
    .FrameData(Tile_X9Y10_FrameData_O),
    .FrameData_O(Tile_X10Y10_FrameData_O),
    .FrameStrobe(Tile_X10Y11_FrameStrobe_O),
    .FrameStrobe_O(Tile_X10Y10_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
W_IO_custom
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X0Y11_Emulate_Bitstream)
    )
`endif
    Tile_X0Y11_W_IO_custom
    (
    .from_NA(Tile_X0Y12_to_NA),
    .from_NB(Tile_X0Y12_to_NB),
    .from_NC(Tile_X0Y12_to_NC),
    .from_ND(Tile_X0Y12_to_ND),
    .from_NF(Tile_X0Y12_to_NF),
    .from_NG(Tile_X0Y12_to_NG),
    .from_NH(Tile_X0Y12_to_NH),
    .from_NI(Tile_X0Y12_to_NI),
    .from_SA(Tile_X0Y10_to_SA),
    .from_SB(Tile_X0Y10_to_SB),
    .from_SC(Tile_X0Y10_to_SC),
    .from_SD(Tile_X0Y10_to_SD),
    .from_SF(Tile_X0Y10_to_SF),
    .from_SG(Tile_X0Y10_to_SG),
    .from_SH(Tile_X0Y10_to_SH),
    .from_SI(Tile_X0Y10_to_SI),
    .from_WA(Tile_X1Y11_to_WA),
    .from_WB(Tile_X1Y11_to_WB),
    .from_WC(Tile_X1Y11_to_WC),
    .from_WD(Tile_X1Y11_to_WD),
    .from_WF(Tile_X1Y11_to_WF),
    .from_WG(Tile_X1Y11_to_WG),
    .from_WH(Tile_X1Y11_to_WH),
    .from_WI(Tile_X1Y11_to_WI),
    .to_EA(Tile_X0Y11_to_EA),
    .to_EB(Tile_X0Y11_to_EB),
    .to_EC(Tile_X0Y11_to_EC),
    .to_ED(Tile_X0Y11_to_ED),
    .to_EF(Tile_X0Y11_to_EF),
    .to_EG(Tile_X0Y11_to_EG),
    .to_EH(Tile_X0Y11_to_EH),
    .to_EI(Tile_X0Y11_to_EI),
    .to_NA(Tile_X0Y11_to_NA),
    .to_NB(Tile_X0Y11_to_NB),
    .to_NC(Tile_X0Y11_to_NC),
    .to_ND(Tile_X0Y11_to_ND),
    .to_NF(Tile_X0Y11_to_NF),
    .to_NG(Tile_X0Y11_to_NG),
    .to_NH(Tile_X0Y11_to_NH),
    .to_NI(Tile_X0Y11_to_NI),
    .to_SA(Tile_X0Y11_to_SA),
    .to_SB(Tile_X0Y11_to_SB),
    .to_SC(Tile_X0Y11_to_SC),
    .to_SD(Tile_X0Y11_to_SD),
    .to_SF(Tile_X0Y11_to_SF),
    .to_SG(Tile_X0Y11_to_SG),
    .to_SH(Tile_X0Y11_to_SH),
    .to_SI(Tile_X0Y11_to_SI),
    .A_O_top_0_t(Tile_X0Y11_A_O_top_0_t),
    .A_O_top_0_f(Tile_X0Y11_A_O_top_0_f),
    .A_O_top_1_t(Tile_X0Y11_A_O_top_1_t),
    .A_O_top_1_f(Tile_X0Y11_A_O_top_1_f),
    .A_prech1(Tile_X0Y11_A_prech1),
    .A_prech2(Tile_X0Y11_A_prech2),
    .A_DR_fault(Tile_X0Y11_A_DR_fault),
    .A_I_top_0_t(Tile_X0Y11_A_I_top_0_t),
    .A_I_top_0_f(Tile_X0Y11_A_I_top_0_f),
    .A_I_top_1_t(Tile_X0Y11_A_I_top_1_t),
    .A_I_top_1_f(Tile_X0Y11_A_I_top_1_f),
    .A_T_top(Tile_X0Y11_A_T_top),
    .A_F_masked1(Tile_X0Y11_A_F_masked1),
    .A_F_masked2(Tile_X0Y11_A_F_masked2),
    .A_config_C_bit0(Tile_X0Y11_A_config_C_bit0),
    .A_config_C_bit1(Tile_X0Y11_A_config_C_bit1),
    .A_config_C_bit2(Tile_X0Y11_A_config_C_bit2),
    .A_config_C_bit3(Tile_X0Y11_A_config_C_bit3),
    .B_config_C_bit0(Tile_X0Y11_B_config_C_bit0),
    .B_config_C_bit1(Tile_X0Y11_B_config_C_bit1),
    .B_config_C_bit2(Tile_X0Y11_B_config_C_bit2),
    .B_config_C_bit3(Tile_X0Y11_B_config_C_bit3),
    .UserCLK(Tile_X0Y12_UserCLKo),
    .UserCLKo(Tile_X0Y11_UserCLKo),
    .rst(Tile_X0Y12_rsto),
    .rsto(Tile_X0Y11_rsto),
    .FrameData(Tile_Y11_FrameData),
    .FrameData_O(Tile_X0Y11_FrameData_O),
    .FrameStrobe(Tile_X0Y12_FrameStrobe_O),
    .FrameStrobe_O(Tile_X0Y11_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X1Y11_Emulate_Bitstream)
    )
`endif
    Tile_X1Y11_linear_LMDPL
    (
    .from_NA(Tile_X1Y12_to_NA),
    .from_NB(Tile_X1Y12_to_NB),
    .from_NC(Tile_X1Y12_to_NC),
    .from_ND(Tile_X1Y12_to_ND),
    .from_NF(Tile_X1Y12_to_NF),
    .from_NG(Tile_X1Y12_to_NG),
    .from_NH(Tile_X1Y12_to_NH),
    .from_NI(Tile_X1Y12_to_NI),
    .from_EA(Tile_X0Y11_to_EA),
    .from_EB(Tile_X0Y11_to_EB),
    .from_EC(Tile_X0Y11_to_EC),
    .from_ED(Tile_X0Y11_to_ED),
    .from_EF(Tile_X0Y11_to_EF),
    .from_EG(Tile_X0Y11_to_EG),
    .from_EH(Tile_X0Y11_to_EH),
    .from_EI(Tile_X0Y11_to_EI),
    .from_SA(Tile_X1Y10_to_SA),
    .from_SB(Tile_X1Y10_to_SB),
    .from_SC(Tile_X1Y10_to_SC),
    .from_SD(Tile_X1Y10_to_SD),
    .from_SF(Tile_X1Y10_to_SF),
    .from_SG(Tile_X1Y10_to_SG),
    .from_SH(Tile_X1Y10_to_SH),
    .from_SI(Tile_X1Y10_to_SI),
    .from_WA(Tile_X2Y11_to_WA),
    .from_WB(Tile_X2Y11_to_WB),
    .from_WC(Tile_X2Y11_to_WC),
    .from_WD(Tile_X2Y11_to_WD),
    .from_WF(Tile_X2Y11_to_WF),
    .from_WG(Tile_X2Y11_to_WG),
    .from_WH(Tile_X2Y11_to_WH),
    .from_WI(Tile_X2Y11_to_WI),
    .to_EA(Tile_X1Y11_to_EA),
    .to_EB(Tile_X1Y11_to_EB),
    .to_EC(Tile_X1Y11_to_EC),
    .to_ED(Tile_X1Y11_to_ED),
    .to_EF(Tile_X1Y11_to_EF),
    .to_EG(Tile_X1Y11_to_EG),
    .to_EH(Tile_X1Y11_to_EH),
    .to_EI(Tile_X1Y11_to_EI),
    .to_WA(Tile_X1Y11_to_WA),
    .to_WB(Tile_X1Y11_to_WB),
    .to_WC(Tile_X1Y11_to_WC),
    .to_WD(Tile_X1Y11_to_WD),
    .to_WF(Tile_X1Y11_to_WF),
    .to_WG(Tile_X1Y11_to_WG),
    .to_WH(Tile_X1Y11_to_WH),
    .to_WI(Tile_X1Y11_to_WI),
    .to_NA(Tile_X1Y11_to_NA),
    .to_NB(Tile_X1Y11_to_NB),
    .to_NC(Tile_X1Y11_to_NC),
    .to_ND(Tile_X1Y11_to_ND),
    .to_NF(Tile_X1Y11_to_NF),
    .to_NG(Tile_X1Y11_to_NG),
    .to_NH(Tile_X1Y11_to_NH),
    .to_NI(Tile_X1Y11_to_NI),
    .to_SA(Tile_X1Y11_to_SA),
    .to_SB(Tile_X1Y11_to_SB),
    .to_SC(Tile_X1Y11_to_SC),
    .to_SD(Tile_X1Y11_to_SD),
    .to_SF(Tile_X1Y11_to_SF),
    .to_SG(Tile_X1Y11_to_SG),
    .to_SH(Tile_X1Y11_to_SH),
    .to_SI(Tile_X1Y11_to_SI),
    .F_masked1(Tile_X1Y11_F_masked1),
    .F_masked2(Tile_X1Y11_F_masked2),
    .UserCLK(Tile_X1Y12_UserCLKo),
    .UserCLKo(Tile_X1Y11_UserCLKo),
    .rst(Tile_X1Y12_rsto),
    .rsto(Tile_X1Y11_rsto),
    .FrameData(Tile_X0Y11_FrameData_O),
    .FrameData_O(Tile_X1Y11_FrameData_O),
    .FrameStrobe(Tile_X1Y12_FrameStrobe_O),
    .FrameStrobe_O(Tile_X1Y11_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X2Y11_Emulate_Bitstream)
    )
`endif
    Tile_X2Y11_linear_LMDPL
    (
    .from_NA(Tile_X2Y12_to_NA),
    .from_NB(Tile_X2Y12_to_NB),
    .from_NC(Tile_X2Y12_to_NC),
    .from_ND(Tile_X2Y12_to_ND),
    .from_NF(Tile_X2Y12_to_NF),
    .from_NG(Tile_X2Y12_to_NG),
    .from_NH(Tile_X2Y12_to_NH),
    .from_NI(Tile_X2Y12_to_NI),
    .from_EA(Tile_X1Y11_to_EA),
    .from_EB(Tile_X1Y11_to_EB),
    .from_EC(Tile_X1Y11_to_EC),
    .from_ED(Tile_X1Y11_to_ED),
    .from_EF(Tile_X1Y11_to_EF),
    .from_EG(Tile_X1Y11_to_EG),
    .from_EH(Tile_X1Y11_to_EH),
    .from_EI(Tile_X1Y11_to_EI),
    .from_SA(Tile_X2Y10_to_SA),
    .from_SB(Tile_X2Y10_to_SB),
    .from_SC(Tile_X2Y10_to_SC),
    .from_SD(Tile_X2Y10_to_SD),
    .from_SF(Tile_X2Y10_to_SF),
    .from_SG(Tile_X2Y10_to_SG),
    .from_SH(Tile_X2Y10_to_SH),
    .from_SI(Tile_X2Y10_to_SI),
    .from_WA(Tile_X3Y11_to_WA),
    .from_WB(Tile_X3Y11_to_WB),
    .from_WC(Tile_X3Y11_to_WC),
    .from_WD(Tile_X3Y11_to_WD),
    .from_WF(Tile_X3Y11_to_WF),
    .from_WG(Tile_X3Y11_to_WG),
    .from_WH(Tile_X3Y11_to_WH),
    .from_WI(Tile_X3Y11_to_WI),
    .to_EA(Tile_X2Y11_to_EA),
    .to_EB(Tile_X2Y11_to_EB),
    .to_EC(Tile_X2Y11_to_EC),
    .to_ED(Tile_X2Y11_to_ED),
    .to_EF(Tile_X2Y11_to_EF),
    .to_EG(Tile_X2Y11_to_EG),
    .to_EH(Tile_X2Y11_to_EH),
    .to_EI(Tile_X2Y11_to_EI),
    .to_WA(Tile_X2Y11_to_WA),
    .to_WB(Tile_X2Y11_to_WB),
    .to_WC(Tile_X2Y11_to_WC),
    .to_WD(Tile_X2Y11_to_WD),
    .to_WF(Tile_X2Y11_to_WF),
    .to_WG(Tile_X2Y11_to_WG),
    .to_WH(Tile_X2Y11_to_WH),
    .to_WI(Tile_X2Y11_to_WI),
    .to_NA(Tile_X2Y11_to_NA),
    .to_NB(Tile_X2Y11_to_NB),
    .to_NC(Tile_X2Y11_to_NC),
    .to_ND(Tile_X2Y11_to_ND),
    .to_NF(Tile_X2Y11_to_NF),
    .to_NG(Tile_X2Y11_to_NG),
    .to_NH(Tile_X2Y11_to_NH),
    .to_NI(Tile_X2Y11_to_NI),
    .to_SA(Tile_X2Y11_to_SA),
    .to_SB(Tile_X2Y11_to_SB),
    .to_SC(Tile_X2Y11_to_SC),
    .to_SD(Tile_X2Y11_to_SD),
    .to_SF(Tile_X2Y11_to_SF),
    .to_SG(Tile_X2Y11_to_SG),
    .to_SH(Tile_X2Y11_to_SH),
    .to_SI(Tile_X2Y11_to_SI),
    .F_masked1(Tile_X2Y11_F_masked1),
    .F_masked2(Tile_X2Y11_F_masked2),
    .UserCLK(Tile_X2Y12_UserCLKo),
    .UserCLKo(Tile_X2Y11_UserCLKo),
    .rst(Tile_X2Y12_rsto),
    .rsto(Tile_X2Y11_rsto),
    .FrameData(Tile_X1Y11_FrameData_O),
    .FrameData_O(Tile_X2Y11_FrameData_O),
    .FrameStrobe(Tile_X2Y12_FrameStrobe_O),
    .FrameStrobe_O(Tile_X2Y11_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
nonlinear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X3Y11_Emulate_Bitstream)
    )
`endif
    Tile_X3Y11_nonlinear_LMDPL
    (
    .from_NA(Tile_X3Y12_to_NA),
    .from_NB(Tile_X3Y12_to_NB),
    .from_NC(Tile_X3Y12_to_NC),
    .from_ND(Tile_X3Y12_to_ND),
    .from_NF(Tile_X3Y12_to_NF),
    .from_NG(Tile_X3Y12_to_NG),
    .from_NH(Tile_X3Y12_to_NH),
    .from_NI(Tile_X3Y12_to_NI),
    .from_EA(Tile_X2Y11_to_EA),
    .from_EB(Tile_X2Y11_to_EB),
    .from_EC(Tile_X2Y11_to_EC),
    .from_ED(Tile_X2Y11_to_ED),
    .from_EF(Tile_X2Y11_to_EF),
    .from_EG(Tile_X2Y11_to_EG),
    .from_EH(Tile_X2Y11_to_EH),
    .from_EI(Tile_X2Y11_to_EI),
    .from_SA(Tile_X3Y10_to_SA),
    .from_SB(Tile_X3Y10_to_SB),
    .from_SC(Tile_X3Y10_to_SC),
    .from_SD(Tile_X3Y10_to_SD),
    .from_SF(Tile_X3Y10_to_SF),
    .from_SG(Tile_X3Y10_to_SG),
    .from_SH(Tile_X3Y10_to_SH),
    .from_SI(Tile_X3Y10_to_SI),
    .from_WA(Tile_X4Y11_to_WA),
    .from_WB(Tile_X4Y11_to_WB),
    .from_WC(Tile_X4Y11_to_WC),
    .from_WD(Tile_X4Y11_to_WD),
    .from_WF(Tile_X4Y11_to_WF),
    .from_WG(Tile_X4Y11_to_WG),
    .from_WH(Tile_X4Y11_to_WH),
    .from_WI(Tile_X4Y11_to_WI),
    .to_EA(Tile_X3Y11_to_EA),
    .to_EB(Tile_X3Y11_to_EB),
    .to_EC(Tile_X3Y11_to_EC),
    .to_ED(Tile_X3Y11_to_ED),
    .to_EF(Tile_X3Y11_to_EF),
    .to_EG(Tile_X3Y11_to_EG),
    .to_EH(Tile_X3Y11_to_EH),
    .to_EI(Tile_X3Y11_to_EI),
    .to_WA(Tile_X3Y11_to_WA),
    .to_WB(Tile_X3Y11_to_WB),
    .to_WC(Tile_X3Y11_to_WC),
    .to_WD(Tile_X3Y11_to_WD),
    .to_WF(Tile_X3Y11_to_WF),
    .to_WG(Tile_X3Y11_to_WG),
    .to_WH(Tile_X3Y11_to_WH),
    .to_WI(Tile_X3Y11_to_WI),
    .to_NA(Tile_X3Y11_to_NA),
    .to_NB(Tile_X3Y11_to_NB),
    .to_NC(Tile_X3Y11_to_NC),
    .to_ND(Tile_X3Y11_to_ND),
    .to_NF(Tile_X3Y11_to_NF),
    .to_NG(Tile_X3Y11_to_NG),
    .to_NH(Tile_X3Y11_to_NH),
    .to_NI(Tile_X3Y11_to_NI),
    .to_SA(Tile_X3Y11_to_SA),
    .to_SB(Tile_X3Y11_to_SB),
    .to_SC(Tile_X3Y11_to_SC),
    .to_SD(Tile_X3Y11_to_SD),
    .to_SF(Tile_X3Y11_to_SF),
    .to_SG(Tile_X3Y11_to_SG),
    .to_SH(Tile_X3Y11_to_SH),
    .to_SI(Tile_X3Y11_to_SI),
    .R_t(Tile_X3Y11_R_t),
    .R_f(Tile_X3Y11_R_f),
    .F_masked1(Tile_X3Y11_F_masked1),
    .F_masked2(Tile_X3Y11_F_masked2),
    .UserCLK(Tile_X3Y12_UserCLKo),
    .UserCLKo(Tile_X3Y11_UserCLKo),
    .rst(Tile_X3Y12_rsto),
    .rsto(Tile_X3Y11_rsto),
    .FrameData(Tile_X2Y11_FrameData_O),
    .FrameData_O(Tile_X3Y11_FrameData_O),
    .FrameStrobe(Tile_X3Y12_FrameStrobe_O),
    .FrameStrobe_O(Tile_X3Y11_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X4Y11_Emulate_Bitstream)
    )
`endif
    Tile_X4Y11_linear_LMDPL
    (
    .from_NA(Tile_X4Y12_to_NA),
    .from_NB(Tile_X4Y12_to_NB),
    .from_NC(Tile_X4Y12_to_NC),
    .from_ND(Tile_X4Y12_to_ND),
    .from_NF(Tile_X4Y12_to_NF),
    .from_NG(Tile_X4Y12_to_NG),
    .from_NH(Tile_X4Y12_to_NH),
    .from_NI(Tile_X4Y12_to_NI),
    .from_EA(Tile_X3Y11_to_EA),
    .from_EB(Tile_X3Y11_to_EB),
    .from_EC(Tile_X3Y11_to_EC),
    .from_ED(Tile_X3Y11_to_ED),
    .from_EF(Tile_X3Y11_to_EF),
    .from_EG(Tile_X3Y11_to_EG),
    .from_EH(Tile_X3Y11_to_EH),
    .from_EI(Tile_X3Y11_to_EI),
    .from_SA(Tile_X4Y10_to_SA),
    .from_SB(Tile_X4Y10_to_SB),
    .from_SC(Tile_X4Y10_to_SC),
    .from_SD(Tile_X4Y10_to_SD),
    .from_SF(Tile_X4Y10_to_SF),
    .from_SG(Tile_X4Y10_to_SG),
    .from_SH(Tile_X4Y10_to_SH),
    .from_SI(Tile_X4Y10_to_SI),
    .from_WA(Tile_X5Y11_to_WA),
    .from_WB(Tile_X5Y11_to_WB),
    .from_WC(Tile_X5Y11_to_WC),
    .from_WD(Tile_X5Y11_to_WD),
    .from_WF(Tile_X5Y11_to_WF),
    .from_WG(Tile_X5Y11_to_WG),
    .from_WH(Tile_X5Y11_to_WH),
    .from_WI(Tile_X5Y11_to_WI),
    .to_EA(Tile_X4Y11_to_EA),
    .to_EB(Tile_X4Y11_to_EB),
    .to_EC(Tile_X4Y11_to_EC),
    .to_ED(Tile_X4Y11_to_ED),
    .to_EF(Tile_X4Y11_to_EF),
    .to_EG(Tile_X4Y11_to_EG),
    .to_EH(Tile_X4Y11_to_EH),
    .to_EI(Tile_X4Y11_to_EI),
    .to_WA(Tile_X4Y11_to_WA),
    .to_WB(Tile_X4Y11_to_WB),
    .to_WC(Tile_X4Y11_to_WC),
    .to_WD(Tile_X4Y11_to_WD),
    .to_WF(Tile_X4Y11_to_WF),
    .to_WG(Tile_X4Y11_to_WG),
    .to_WH(Tile_X4Y11_to_WH),
    .to_WI(Tile_X4Y11_to_WI),
    .to_NA(Tile_X4Y11_to_NA),
    .to_NB(Tile_X4Y11_to_NB),
    .to_NC(Tile_X4Y11_to_NC),
    .to_ND(Tile_X4Y11_to_ND),
    .to_NF(Tile_X4Y11_to_NF),
    .to_NG(Tile_X4Y11_to_NG),
    .to_NH(Tile_X4Y11_to_NH),
    .to_NI(Tile_X4Y11_to_NI),
    .to_SA(Tile_X4Y11_to_SA),
    .to_SB(Tile_X4Y11_to_SB),
    .to_SC(Tile_X4Y11_to_SC),
    .to_SD(Tile_X4Y11_to_SD),
    .to_SF(Tile_X4Y11_to_SF),
    .to_SG(Tile_X4Y11_to_SG),
    .to_SH(Tile_X4Y11_to_SH),
    .to_SI(Tile_X4Y11_to_SI),
    .F_masked1(Tile_X4Y11_F_masked1),
    .F_masked2(Tile_X4Y11_F_masked2),
    .UserCLK(Tile_X4Y12_UserCLKo),
    .UserCLKo(Tile_X4Y11_UserCLKo),
    .rst(Tile_X4Y12_rsto),
    .rsto(Tile_X4Y11_rsto),
    .FrameData(Tile_X3Y11_FrameData_O),
    .FrameData_O(Tile_X4Y11_FrameData_O),
    .FrameStrobe(Tile_X4Y12_FrameStrobe_O),
    .FrameStrobe_O(Tile_X4Y11_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X5Y11_Emulate_Bitstream)
    )
`endif
    Tile_X5Y11_linear_LMDPL
    (
    .from_NA(Tile_X5Y12_to_NA),
    .from_NB(Tile_X5Y12_to_NB),
    .from_NC(Tile_X5Y12_to_NC),
    .from_ND(Tile_X5Y12_to_ND),
    .from_NF(Tile_X5Y12_to_NF),
    .from_NG(Tile_X5Y12_to_NG),
    .from_NH(Tile_X5Y12_to_NH),
    .from_NI(Tile_X5Y12_to_NI),
    .from_EA(Tile_X4Y11_to_EA),
    .from_EB(Tile_X4Y11_to_EB),
    .from_EC(Tile_X4Y11_to_EC),
    .from_ED(Tile_X4Y11_to_ED),
    .from_EF(Tile_X4Y11_to_EF),
    .from_EG(Tile_X4Y11_to_EG),
    .from_EH(Tile_X4Y11_to_EH),
    .from_EI(Tile_X4Y11_to_EI),
    .from_SA(Tile_X5Y10_to_SA),
    .from_SB(Tile_X5Y10_to_SB),
    .from_SC(Tile_X5Y10_to_SC),
    .from_SD(Tile_X5Y10_to_SD),
    .from_SF(Tile_X5Y10_to_SF),
    .from_SG(Tile_X5Y10_to_SG),
    .from_SH(Tile_X5Y10_to_SH),
    .from_SI(Tile_X5Y10_to_SI),
    .from_WA(Tile_X6Y11_to_WA),
    .from_WB(Tile_X6Y11_to_WB),
    .from_WC(Tile_X6Y11_to_WC),
    .from_WD(Tile_X6Y11_to_WD),
    .from_WF(Tile_X6Y11_to_WF),
    .from_WG(Tile_X6Y11_to_WG),
    .from_WH(Tile_X6Y11_to_WH),
    .from_WI(Tile_X6Y11_to_WI),
    .to_EA(Tile_X5Y11_to_EA),
    .to_EB(Tile_X5Y11_to_EB),
    .to_EC(Tile_X5Y11_to_EC),
    .to_ED(Tile_X5Y11_to_ED),
    .to_EF(Tile_X5Y11_to_EF),
    .to_EG(Tile_X5Y11_to_EG),
    .to_EH(Tile_X5Y11_to_EH),
    .to_EI(Tile_X5Y11_to_EI),
    .to_WA(Tile_X5Y11_to_WA),
    .to_WB(Tile_X5Y11_to_WB),
    .to_WC(Tile_X5Y11_to_WC),
    .to_WD(Tile_X5Y11_to_WD),
    .to_WF(Tile_X5Y11_to_WF),
    .to_WG(Tile_X5Y11_to_WG),
    .to_WH(Tile_X5Y11_to_WH),
    .to_WI(Tile_X5Y11_to_WI),
    .to_NA(Tile_X5Y11_to_NA),
    .to_NB(Tile_X5Y11_to_NB),
    .to_NC(Tile_X5Y11_to_NC),
    .to_ND(Tile_X5Y11_to_ND),
    .to_NF(Tile_X5Y11_to_NF),
    .to_NG(Tile_X5Y11_to_NG),
    .to_NH(Tile_X5Y11_to_NH),
    .to_NI(Tile_X5Y11_to_NI),
    .to_SA(Tile_X5Y11_to_SA),
    .to_SB(Tile_X5Y11_to_SB),
    .to_SC(Tile_X5Y11_to_SC),
    .to_SD(Tile_X5Y11_to_SD),
    .to_SF(Tile_X5Y11_to_SF),
    .to_SG(Tile_X5Y11_to_SG),
    .to_SH(Tile_X5Y11_to_SH),
    .to_SI(Tile_X5Y11_to_SI),
    .F_masked1(Tile_X5Y11_F_masked1),
    .F_masked2(Tile_X5Y11_F_masked2),
    .UserCLK(Tile_X5Y12_UserCLKo),
    .UserCLKo(Tile_X5Y11_UserCLKo),
    .rst(Tile_X5Y12_rsto),
    .rsto(Tile_X5Y11_rsto),
    .FrameData(Tile_X4Y11_FrameData_O),
    .FrameData_O(Tile_X5Y11_FrameData_O),
    .FrameStrobe(Tile_X5Y12_FrameStrobe_O),
    .FrameStrobe_O(Tile_X5Y11_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
nonlinear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X6Y11_Emulate_Bitstream)
    )
`endif
    Tile_X6Y11_nonlinear_LMDPL
    (
    .from_NA(Tile_X6Y12_to_NA),
    .from_NB(Tile_X6Y12_to_NB),
    .from_NC(Tile_X6Y12_to_NC),
    .from_ND(Tile_X6Y12_to_ND),
    .from_NF(Tile_X6Y12_to_NF),
    .from_NG(Tile_X6Y12_to_NG),
    .from_NH(Tile_X6Y12_to_NH),
    .from_NI(Tile_X6Y12_to_NI),
    .from_EA(Tile_X5Y11_to_EA),
    .from_EB(Tile_X5Y11_to_EB),
    .from_EC(Tile_X5Y11_to_EC),
    .from_ED(Tile_X5Y11_to_ED),
    .from_EF(Tile_X5Y11_to_EF),
    .from_EG(Tile_X5Y11_to_EG),
    .from_EH(Tile_X5Y11_to_EH),
    .from_EI(Tile_X5Y11_to_EI),
    .from_SA(Tile_X6Y10_to_SA),
    .from_SB(Tile_X6Y10_to_SB),
    .from_SC(Tile_X6Y10_to_SC),
    .from_SD(Tile_X6Y10_to_SD),
    .from_SF(Tile_X6Y10_to_SF),
    .from_SG(Tile_X6Y10_to_SG),
    .from_SH(Tile_X6Y10_to_SH),
    .from_SI(Tile_X6Y10_to_SI),
    .from_WA(Tile_X7Y11_to_WA),
    .from_WB(Tile_X7Y11_to_WB),
    .from_WC(Tile_X7Y11_to_WC),
    .from_WD(Tile_X7Y11_to_WD),
    .from_WF(Tile_X7Y11_to_WF),
    .from_WG(Tile_X7Y11_to_WG),
    .from_WH(Tile_X7Y11_to_WH),
    .from_WI(Tile_X7Y11_to_WI),
    .to_EA(Tile_X6Y11_to_EA),
    .to_EB(Tile_X6Y11_to_EB),
    .to_EC(Tile_X6Y11_to_EC),
    .to_ED(Tile_X6Y11_to_ED),
    .to_EF(Tile_X6Y11_to_EF),
    .to_EG(Tile_X6Y11_to_EG),
    .to_EH(Tile_X6Y11_to_EH),
    .to_EI(Tile_X6Y11_to_EI),
    .to_WA(Tile_X6Y11_to_WA),
    .to_WB(Tile_X6Y11_to_WB),
    .to_WC(Tile_X6Y11_to_WC),
    .to_WD(Tile_X6Y11_to_WD),
    .to_WF(Tile_X6Y11_to_WF),
    .to_WG(Tile_X6Y11_to_WG),
    .to_WH(Tile_X6Y11_to_WH),
    .to_WI(Tile_X6Y11_to_WI),
    .to_NA(Tile_X6Y11_to_NA),
    .to_NB(Tile_X6Y11_to_NB),
    .to_NC(Tile_X6Y11_to_NC),
    .to_ND(Tile_X6Y11_to_ND),
    .to_NF(Tile_X6Y11_to_NF),
    .to_NG(Tile_X6Y11_to_NG),
    .to_NH(Tile_X6Y11_to_NH),
    .to_NI(Tile_X6Y11_to_NI),
    .to_SA(Tile_X6Y11_to_SA),
    .to_SB(Tile_X6Y11_to_SB),
    .to_SC(Tile_X6Y11_to_SC),
    .to_SD(Tile_X6Y11_to_SD),
    .to_SF(Tile_X6Y11_to_SF),
    .to_SG(Tile_X6Y11_to_SG),
    .to_SH(Tile_X6Y11_to_SH),
    .to_SI(Tile_X6Y11_to_SI),
    .R_t(Tile_X6Y11_R_t),
    .R_f(Tile_X6Y11_R_f),
    .F_masked1(Tile_X6Y11_F_masked1),
    .F_masked2(Tile_X6Y11_F_masked2),
    .UserCLK(Tile_X6Y12_UserCLKo),
    .UserCLKo(Tile_X6Y11_UserCLKo),
    .rst(Tile_X6Y12_rsto),
    .rsto(Tile_X6Y11_rsto),
    .FrameData(Tile_X5Y11_FrameData_O),
    .FrameData_O(Tile_X6Y11_FrameData_O),
    .FrameStrobe(Tile_X6Y12_FrameStrobe_O),
    .FrameStrobe_O(Tile_X6Y11_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X7Y11_Emulate_Bitstream)
    )
`endif
    Tile_X7Y11_linear_LMDPL
    (
    .from_NA(Tile_X7Y12_to_NA),
    .from_NB(Tile_X7Y12_to_NB),
    .from_NC(Tile_X7Y12_to_NC),
    .from_ND(Tile_X7Y12_to_ND),
    .from_NF(Tile_X7Y12_to_NF),
    .from_NG(Tile_X7Y12_to_NG),
    .from_NH(Tile_X7Y12_to_NH),
    .from_NI(Tile_X7Y12_to_NI),
    .from_EA(Tile_X6Y11_to_EA),
    .from_EB(Tile_X6Y11_to_EB),
    .from_EC(Tile_X6Y11_to_EC),
    .from_ED(Tile_X6Y11_to_ED),
    .from_EF(Tile_X6Y11_to_EF),
    .from_EG(Tile_X6Y11_to_EG),
    .from_EH(Tile_X6Y11_to_EH),
    .from_EI(Tile_X6Y11_to_EI),
    .from_SA(Tile_X7Y10_to_SA),
    .from_SB(Tile_X7Y10_to_SB),
    .from_SC(Tile_X7Y10_to_SC),
    .from_SD(Tile_X7Y10_to_SD),
    .from_SF(Tile_X7Y10_to_SF),
    .from_SG(Tile_X7Y10_to_SG),
    .from_SH(Tile_X7Y10_to_SH),
    .from_SI(Tile_X7Y10_to_SI),
    .from_WA(Tile_X8Y11_to_WA),
    .from_WB(Tile_X8Y11_to_WB),
    .from_WC(Tile_X8Y11_to_WC),
    .from_WD(Tile_X8Y11_to_WD),
    .from_WF(Tile_X8Y11_to_WF),
    .from_WG(Tile_X8Y11_to_WG),
    .from_WH(Tile_X8Y11_to_WH),
    .from_WI(Tile_X8Y11_to_WI),
    .to_EA(Tile_X7Y11_to_EA),
    .to_EB(Tile_X7Y11_to_EB),
    .to_EC(Tile_X7Y11_to_EC),
    .to_ED(Tile_X7Y11_to_ED),
    .to_EF(Tile_X7Y11_to_EF),
    .to_EG(Tile_X7Y11_to_EG),
    .to_EH(Tile_X7Y11_to_EH),
    .to_EI(Tile_X7Y11_to_EI),
    .to_WA(Tile_X7Y11_to_WA),
    .to_WB(Tile_X7Y11_to_WB),
    .to_WC(Tile_X7Y11_to_WC),
    .to_WD(Tile_X7Y11_to_WD),
    .to_WF(Tile_X7Y11_to_WF),
    .to_WG(Tile_X7Y11_to_WG),
    .to_WH(Tile_X7Y11_to_WH),
    .to_WI(Tile_X7Y11_to_WI),
    .to_NA(Tile_X7Y11_to_NA),
    .to_NB(Tile_X7Y11_to_NB),
    .to_NC(Tile_X7Y11_to_NC),
    .to_ND(Tile_X7Y11_to_ND),
    .to_NF(Tile_X7Y11_to_NF),
    .to_NG(Tile_X7Y11_to_NG),
    .to_NH(Tile_X7Y11_to_NH),
    .to_NI(Tile_X7Y11_to_NI),
    .to_SA(Tile_X7Y11_to_SA),
    .to_SB(Tile_X7Y11_to_SB),
    .to_SC(Tile_X7Y11_to_SC),
    .to_SD(Tile_X7Y11_to_SD),
    .to_SF(Tile_X7Y11_to_SF),
    .to_SG(Tile_X7Y11_to_SG),
    .to_SH(Tile_X7Y11_to_SH),
    .to_SI(Tile_X7Y11_to_SI),
    .F_masked1(Tile_X7Y11_F_masked1),
    .F_masked2(Tile_X7Y11_F_masked2),
    .UserCLK(Tile_X7Y12_UserCLKo),
    .UserCLKo(Tile_X7Y11_UserCLKo),
    .rst(Tile_X7Y12_rsto),
    .rsto(Tile_X7Y11_rsto),
    .FrameData(Tile_X6Y11_FrameData_O),
    .FrameData_O(Tile_X7Y11_FrameData_O),
    .FrameStrobe(Tile_X7Y12_FrameStrobe_O),
    .FrameStrobe_O(Tile_X7Y11_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
ctrl_to_sec
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X8Y11_Emulate_Bitstream)
    )
`endif
    Tile_X8Y11_ctrl_to_sec
    (
    .from_NA(Tile_X8Y12_to_NA),
    .from_NB(Tile_X8Y12_to_NB),
    .from_NC(Tile_X8Y12_to_NC),
    .from_ND(Tile_X8Y12_to_ND),
    .from_NF(Tile_X8Y12_to_NF),
    .from_NG(Tile_X8Y12_to_NG),
    .from_NH(Tile_X8Y12_to_NH),
    .from_NI(Tile_X8Y12_to_NI),
    .from_EA(Tile_X7Y11_to_EA),
    .from_EB(Tile_X7Y11_to_EB),
    .from_EC(Tile_X7Y11_to_EC),
    .from_ED(Tile_X7Y11_to_ED),
    .from_EF(Tile_X7Y11_to_EF),
    .from_EG(Tile_X7Y11_to_EG),
    .from_EH(Tile_X7Y11_to_EH),
    .from_EI(Tile_X7Y11_to_EI),
    .from_SA(Tile_X8Y10_to_SA),
    .from_SB(Tile_X8Y10_to_SB),
    .from_SC(Tile_X8Y10_to_SC),
    .from_SD(Tile_X8Y10_to_SD),
    .from_SF(Tile_X8Y10_to_SF),
    .from_SG(Tile_X8Y10_to_SG),
    .from_SH(Tile_X8Y10_to_SH),
    .from_SI(Tile_X8Y10_to_SI),
    .from_WA_1s(Tile_X9Y11_to_WA_1s),
    .from_WB_1s(Tile_X9Y11_to_WB_1s),
    .from_WC_1s(Tile_X9Y11_to_WC_1s),
    .from_WD_1s(Tile_X9Y11_to_WD_1s),
    .from_WF_1s(Tile_X9Y11_to_WF_1s),
    .from_WG_1s(Tile_X9Y11_to_WG_1s),
    .from_WH_1s(Tile_X9Y11_to_WH_1s),
    .from_WI_1s(Tile_X9Y11_to_WI_1s),
    .to_WA(Tile_X8Y11_to_WA),
    .to_WB(Tile_X8Y11_to_WB),
    .to_WC(Tile_X8Y11_to_WC),
    .to_WD(Tile_X8Y11_to_WD),
    .to_WF(Tile_X8Y11_to_WF),
    .to_WG(Tile_X8Y11_to_WG),
    .to_WH(Tile_X8Y11_to_WH),
    .to_WI(Tile_X8Y11_to_WI),
    .to_NA(Tile_X8Y11_to_NA),
    .to_NB(Tile_X8Y11_to_NB),
    .to_NC(Tile_X8Y11_to_NC),
    .to_ND(Tile_X8Y11_to_ND),
    .to_NF(Tile_X8Y11_to_NF),
    .to_NG(Tile_X8Y11_to_NG),
    .to_NH(Tile_X8Y11_to_NH),
    .to_NI(Tile_X8Y11_to_NI),
    .to_SA(Tile_X8Y11_to_SA),
    .to_SB(Tile_X8Y11_to_SB),
    .to_SC(Tile_X8Y11_to_SC),
    .to_SD(Tile_X8Y11_to_SD),
    .to_SF(Tile_X8Y11_to_SF),
    .to_SG(Tile_X8Y11_to_SG),
    .to_SH(Tile_X8Y11_to_SH),
    .to_SI(Tile_X8Y11_to_SI),
    .UserCLK(Tile_X8Y12_UserCLKo),
    .UserCLKo(Tile_X8Y11_UserCLKo),
    .rst(Tile_X8Y12_rsto),
    .rsto(Tile_X8Y11_rsto),
    .FrameData(Tile_X7Y11_FrameData_O),
    .FrameData_O(Tile_X8Y11_FrameData_O),
    .FrameStrobe(Tile_X8Y12_FrameStrobe_O),
    .FrameStrobe_O(Tile_X8Y11_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
combined_WDDL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X9Y11_Emulate_Bitstream)
    )
`endif
    Tile_X9Y11_combined_WDDL
    (
    .from_NA_1s(Tile_X9Y12_to_NA_1s),
    .from_NB_1s(Tile_X9Y12_to_NB_1s),
    .from_NC_1s(Tile_X9Y12_to_NC_1s),
    .from_ND_1s(Tile_X9Y12_to_ND_1s),
    .from_NF_1s(Tile_X9Y12_to_NF_1s),
    .from_NG_1s(Tile_X9Y12_to_NG_1s),
    .from_NH_1s(Tile_X9Y12_to_NH_1s),
    .from_NI_1s(Tile_X9Y12_to_NI_1s),
    .from_SA_1s(Tile_X9Y10_to_SA_1s),
    .from_SB_1s(Tile_X9Y10_to_SB_1s),
    .from_SC_1s(Tile_X9Y10_to_SC_1s),
    .from_SD_1s(Tile_X9Y10_to_SD_1s),
    .from_SF_1s(Tile_X9Y10_to_SF_1s),
    .from_SG_1s(Tile_X9Y10_to_SG_1s),
    .from_SH_1s(Tile_X9Y10_to_SH_1s),
    .from_SI_1s(Tile_X9Y10_to_SI_1s),
    .from_WA_1s(Tile_X10Y11_to_WA_1s),
    .from_WB_1s(Tile_X10Y11_to_WB_1s),
    .from_WC_1s(Tile_X10Y11_to_WC_1s),
    .from_WD_1s(Tile_X10Y11_to_WD_1s),
    .from_WF_1s(Tile_X10Y11_to_WF_1s),
    .from_WG_1s(Tile_X10Y11_to_WG_1s),
    .from_WH_1s(Tile_X10Y11_to_WH_1s),
    .from_WI_1s(Tile_X10Y11_to_WI_1s),
    .to_EA_1s(Tile_X9Y11_to_EA_1s),
    .to_EB_1s(Tile_X9Y11_to_EB_1s),
    .to_EC_1s(Tile_X9Y11_to_EC_1s),
    .to_ED_1s(Tile_X9Y11_to_ED_1s),
    .to_EF_1s(Tile_X9Y11_to_EF_1s),
    .to_EG_1s(Tile_X9Y11_to_EG_1s),
    .to_EH_1s(Tile_X9Y11_to_EH_1s),
    .to_EI_1s(Tile_X9Y11_to_EI_1s),
    .to_WA_1s(Tile_X9Y11_to_WA_1s),
    .to_WB_1s(Tile_X9Y11_to_WB_1s),
    .to_WC_1s(Tile_X9Y11_to_WC_1s),
    .to_WD_1s(Tile_X9Y11_to_WD_1s),
    .to_WF_1s(Tile_X9Y11_to_WF_1s),
    .to_WG_1s(Tile_X9Y11_to_WG_1s),
    .to_WH_1s(Tile_X9Y11_to_WH_1s),
    .to_WI_1s(Tile_X9Y11_to_WI_1s),
    .to_NA_1s(Tile_X9Y11_to_NA_1s),
    .to_NB_1s(Tile_X9Y11_to_NB_1s),
    .to_NC_1s(Tile_X9Y11_to_NC_1s),
    .to_ND_1s(Tile_X9Y11_to_ND_1s),
    .to_NF_1s(Tile_X9Y11_to_NF_1s),
    .to_NG_1s(Tile_X9Y11_to_NG_1s),
    .to_NH_1s(Tile_X9Y11_to_NH_1s),
    .to_NI_1s(Tile_X9Y11_to_NI_1s),
    .to_SA_1s(Tile_X9Y11_to_SA_1s),
    .to_SB_1s(Tile_X9Y11_to_SB_1s),
    .to_SC_1s(Tile_X9Y11_to_SC_1s),
    .to_SD_1s(Tile_X9Y11_to_SD_1s),
    .to_SF_1s(Tile_X9Y11_to_SF_1s),
    .to_SG_1s(Tile_X9Y11_to_SG_1s),
    .to_SH_1s(Tile_X9Y11_to_SH_1s),
    .to_SI_1s(Tile_X9Y11_to_SI_1s),
    .F_ctrl(Tile_X9Y11_F_ctrl),
    .UserCLK(Tile_X9Y12_UserCLKo),
    .UserCLKo(Tile_X9Y11_UserCLKo),
    .rst(Tile_X9Y12_rsto),
    .rsto(Tile_X9Y11_rsto),
    .FrameData(Tile_X8Y11_FrameData_O),
    .FrameData_O(Tile_X9Y11_FrameData_O),
    .FrameStrobe(Tile_X9Y12_FrameStrobe_O),
    .FrameStrobe_O(Tile_X9Y11_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
ctrl_IO
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X10Y11_Emulate_Bitstream)
    )
`endif
    Tile_X10Y11_ctrl_IO
    (
    .from_EA_1s(Tile_X9Y11_to_EA_1s),
    .from_EB_1s(Tile_X9Y11_to_EB_1s),
    .from_EC_1s(Tile_X9Y11_to_EC_1s),
    .from_ED_1s(Tile_X9Y11_to_ED_1s),
    .from_EF_1s(Tile_X9Y11_to_EF_1s),
    .from_EG_1s(Tile_X9Y11_to_EG_1s),
    .from_EH_1s(Tile_X9Y11_to_EH_1s),
    .from_EI_1s(Tile_X9Y11_to_EI_1s),
    .to_WA_1s(Tile_X10Y11_to_WA_1s),
    .to_WB_1s(Tile_X10Y11_to_WB_1s),
    .to_WC_1s(Tile_X10Y11_to_WC_1s),
    .to_WD_1s(Tile_X10Y11_to_WD_1s),
    .to_WF_1s(Tile_X10Y11_to_WF_1s),
    .to_WG_1s(Tile_X10Y11_to_WG_1s),
    .to_WH_1s(Tile_X10Y11_to_WH_1s),
    .to_WI_1s(Tile_X10Y11_to_WI_1s),
    .A_O_top_0_t(Tile_X10Y11_A_O_top_0_t),
    .A_O_top_0_f(Tile_X10Y11_A_O_top_0_f),
    .A_prech2(Tile_X10Y11_A_prech2),
    .A_DR_fault(Tile_X10Y11_A_DR_fault),
    .A_I_top_0_t(Tile_X10Y11_A_I_top_0_t),
    .A_I_top_0_f(Tile_X10Y11_A_I_top_0_f),
    .A_T_top(Tile_X10Y11_A_T_top),
    .A_F_ctrl(Tile_X10Y11_A_F_ctrl),
    .UserCLK(Tile_X10Y12_UserCLKo),
    .UserCLKo(Tile_X10Y11_UserCLKo),
    .rst(Tile_X10Y12_rsto),
    .rsto(Tile_X10Y11_rsto),
    .FrameData(Tile_X9Y11_FrameData_O),
    .FrameData_O(Tile_X10Y11_FrameData_O),
    .FrameStrobe(Tile_X10Y12_FrameStrobe_O),
    .FrameStrobe_O(Tile_X10Y11_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
W_IO_custom
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X0Y12_Emulate_Bitstream)
    )
`endif
    Tile_X0Y12_W_IO_custom
    (
    .from_NA(Tile_X0Y13_to_NA),
    .from_NB(Tile_X0Y13_to_NB),
    .from_NC(Tile_X0Y13_to_NC),
    .from_ND(Tile_X0Y13_to_ND),
    .from_NF(Tile_X0Y13_to_NF),
    .from_NG(Tile_X0Y13_to_NG),
    .from_NH(Tile_X0Y13_to_NH),
    .from_NI(Tile_X0Y13_to_NI),
    .from_SA(Tile_X0Y11_to_SA),
    .from_SB(Tile_X0Y11_to_SB),
    .from_SC(Tile_X0Y11_to_SC),
    .from_SD(Tile_X0Y11_to_SD),
    .from_SF(Tile_X0Y11_to_SF),
    .from_SG(Tile_X0Y11_to_SG),
    .from_SH(Tile_X0Y11_to_SH),
    .from_SI(Tile_X0Y11_to_SI),
    .from_WA(Tile_X1Y12_to_WA),
    .from_WB(Tile_X1Y12_to_WB),
    .from_WC(Tile_X1Y12_to_WC),
    .from_WD(Tile_X1Y12_to_WD),
    .from_WF(Tile_X1Y12_to_WF),
    .from_WG(Tile_X1Y12_to_WG),
    .from_WH(Tile_X1Y12_to_WH),
    .from_WI(Tile_X1Y12_to_WI),
    .to_EA(Tile_X0Y12_to_EA),
    .to_EB(Tile_X0Y12_to_EB),
    .to_EC(Tile_X0Y12_to_EC),
    .to_ED(Tile_X0Y12_to_ED),
    .to_EF(Tile_X0Y12_to_EF),
    .to_EG(Tile_X0Y12_to_EG),
    .to_EH(Tile_X0Y12_to_EH),
    .to_EI(Tile_X0Y12_to_EI),
    .to_NA(Tile_X0Y12_to_NA),
    .to_NB(Tile_X0Y12_to_NB),
    .to_NC(Tile_X0Y12_to_NC),
    .to_ND(Tile_X0Y12_to_ND),
    .to_NF(Tile_X0Y12_to_NF),
    .to_NG(Tile_X0Y12_to_NG),
    .to_NH(Tile_X0Y12_to_NH),
    .to_NI(Tile_X0Y12_to_NI),
    .to_SA(Tile_X0Y12_to_SA),
    .to_SB(Tile_X0Y12_to_SB),
    .to_SC(Tile_X0Y12_to_SC),
    .to_SD(Tile_X0Y12_to_SD),
    .to_SF(Tile_X0Y12_to_SF),
    .to_SG(Tile_X0Y12_to_SG),
    .to_SH(Tile_X0Y12_to_SH),
    .to_SI(Tile_X0Y12_to_SI),
    .A_O_top_0_t(Tile_X0Y12_A_O_top_0_t),
    .A_O_top_0_f(Tile_X0Y12_A_O_top_0_f),
    .A_O_top_1_t(Tile_X0Y12_A_O_top_1_t),
    .A_O_top_1_f(Tile_X0Y12_A_O_top_1_f),
    .A_prech1(Tile_X0Y12_A_prech1),
    .A_prech2(Tile_X0Y12_A_prech2),
    .A_DR_fault(Tile_X0Y12_A_DR_fault),
    .A_I_top_0_t(Tile_X0Y12_A_I_top_0_t),
    .A_I_top_0_f(Tile_X0Y12_A_I_top_0_f),
    .A_I_top_1_t(Tile_X0Y12_A_I_top_1_t),
    .A_I_top_1_f(Tile_X0Y12_A_I_top_1_f),
    .A_T_top(Tile_X0Y12_A_T_top),
    .A_F_masked1(Tile_X0Y12_A_F_masked1),
    .A_F_masked2(Tile_X0Y12_A_F_masked2),
    .A_config_C_bit0(Tile_X0Y12_A_config_C_bit0),
    .A_config_C_bit1(Tile_X0Y12_A_config_C_bit1),
    .A_config_C_bit2(Tile_X0Y12_A_config_C_bit2),
    .A_config_C_bit3(Tile_X0Y12_A_config_C_bit3),
    .B_config_C_bit0(Tile_X0Y12_B_config_C_bit0),
    .B_config_C_bit1(Tile_X0Y12_B_config_C_bit1),
    .B_config_C_bit2(Tile_X0Y12_B_config_C_bit2),
    .B_config_C_bit3(Tile_X0Y12_B_config_C_bit3),
    .UserCLK(Tile_X0Y13_UserCLKo),
    .UserCLKo(Tile_X0Y12_UserCLKo),
    .rst(Tile_X0Y13_rsto),
    .rsto(Tile_X0Y12_rsto),
    .FrameData(Tile_Y12_FrameData),
    .FrameData_O(Tile_X0Y12_FrameData_O),
    .FrameStrobe(Tile_X0Y13_FrameStrobe_O),
    .FrameStrobe_O(Tile_X0Y12_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X1Y12_Emulate_Bitstream)
    )
`endif
    Tile_X1Y12_linear_LMDPL
    (
    .from_NA(Tile_X1Y13_to_NA),
    .from_NB(Tile_X1Y13_to_NB),
    .from_NC(Tile_X1Y13_to_NC),
    .from_ND(Tile_X1Y13_to_ND),
    .from_NF(Tile_X1Y13_to_NF),
    .from_NG(Tile_X1Y13_to_NG),
    .from_NH(Tile_X1Y13_to_NH),
    .from_NI(Tile_X1Y13_to_NI),
    .from_EA(Tile_X0Y12_to_EA),
    .from_EB(Tile_X0Y12_to_EB),
    .from_EC(Tile_X0Y12_to_EC),
    .from_ED(Tile_X0Y12_to_ED),
    .from_EF(Tile_X0Y12_to_EF),
    .from_EG(Tile_X0Y12_to_EG),
    .from_EH(Tile_X0Y12_to_EH),
    .from_EI(Tile_X0Y12_to_EI),
    .from_SA(Tile_X1Y11_to_SA),
    .from_SB(Tile_X1Y11_to_SB),
    .from_SC(Tile_X1Y11_to_SC),
    .from_SD(Tile_X1Y11_to_SD),
    .from_SF(Tile_X1Y11_to_SF),
    .from_SG(Tile_X1Y11_to_SG),
    .from_SH(Tile_X1Y11_to_SH),
    .from_SI(Tile_X1Y11_to_SI),
    .from_WA(Tile_X2Y12_to_WA),
    .from_WB(Tile_X2Y12_to_WB),
    .from_WC(Tile_X2Y12_to_WC),
    .from_WD(Tile_X2Y12_to_WD),
    .from_WF(Tile_X2Y12_to_WF),
    .from_WG(Tile_X2Y12_to_WG),
    .from_WH(Tile_X2Y12_to_WH),
    .from_WI(Tile_X2Y12_to_WI),
    .to_EA(Tile_X1Y12_to_EA),
    .to_EB(Tile_X1Y12_to_EB),
    .to_EC(Tile_X1Y12_to_EC),
    .to_ED(Tile_X1Y12_to_ED),
    .to_EF(Tile_X1Y12_to_EF),
    .to_EG(Tile_X1Y12_to_EG),
    .to_EH(Tile_X1Y12_to_EH),
    .to_EI(Tile_X1Y12_to_EI),
    .to_WA(Tile_X1Y12_to_WA),
    .to_WB(Tile_X1Y12_to_WB),
    .to_WC(Tile_X1Y12_to_WC),
    .to_WD(Tile_X1Y12_to_WD),
    .to_WF(Tile_X1Y12_to_WF),
    .to_WG(Tile_X1Y12_to_WG),
    .to_WH(Tile_X1Y12_to_WH),
    .to_WI(Tile_X1Y12_to_WI),
    .to_NA(Tile_X1Y12_to_NA),
    .to_NB(Tile_X1Y12_to_NB),
    .to_NC(Tile_X1Y12_to_NC),
    .to_ND(Tile_X1Y12_to_ND),
    .to_NF(Tile_X1Y12_to_NF),
    .to_NG(Tile_X1Y12_to_NG),
    .to_NH(Tile_X1Y12_to_NH),
    .to_NI(Tile_X1Y12_to_NI),
    .to_SA(Tile_X1Y12_to_SA),
    .to_SB(Tile_X1Y12_to_SB),
    .to_SC(Tile_X1Y12_to_SC),
    .to_SD(Tile_X1Y12_to_SD),
    .to_SF(Tile_X1Y12_to_SF),
    .to_SG(Tile_X1Y12_to_SG),
    .to_SH(Tile_X1Y12_to_SH),
    .to_SI(Tile_X1Y12_to_SI),
    .F_masked1(Tile_X1Y12_F_masked1),
    .F_masked2(Tile_X1Y12_F_masked2),
    .UserCLK(Tile_X1Y13_UserCLKo),
    .UserCLKo(Tile_X1Y12_UserCLKo),
    .rst(Tile_X1Y13_rsto),
    .rsto(Tile_X1Y12_rsto),
    .FrameData(Tile_X0Y12_FrameData_O),
    .FrameData_O(Tile_X1Y12_FrameData_O),
    .FrameStrobe(Tile_X1Y13_FrameStrobe_O),
    .FrameStrobe_O(Tile_X1Y12_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X2Y12_Emulate_Bitstream)
    )
`endif
    Tile_X2Y12_linear_LMDPL
    (
    .from_NA(Tile_X2Y13_to_NA),
    .from_NB(Tile_X2Y13_to_NB),
    .from_NC(Tile_X2Y13_to_NC),
    .from_ND(Tile_X2Y13_to_ND),
    .from_NF(Tile_X2Y13_to_NF),
    .from_NG(Tile_X2Y13_to_NG),
    .from_NH(Tile_X2Y13_to_NH),
    .from_NI(Tile_X2Y13_to_NI),
    .from_EA(Tile_X1Y12_to_EA),
    .from_EB(Tile_X1Y12_to_EB),
    .from_EC(Tile_X1Y12_to_EC),
    .from_ED(Tile_X1Y12_to_ED),
    .from_EF(Tile_X1Y12_to_EF),
    .from_EG(Tile_X1Y12_to_EG),
    .from_EH(Tile_X1Y12_to_EH),
    .from_EI(Tile_X1Y12_to_EI),
    .from_SA(Tile_X2Y11_to_SA),
    .from_SB(Tile_X2Y11_to_SB),
    .from_SC(Tile_X2Y11_to_SC),
    .from_SD(Tile_X2Y11_to_SD),
    .from_SF(Tile_X2Y11_to_SF),
    .from_SG(Tile_X2Y11_to_SG),
    .from_SH(Tile_X2Y11_to_SH),
    .from_SI(Tile_X2Y11_to_SI),
    .from_WA(Tile_X3Y12_to_WA),
    .from_WB(Tile_X3Y12_to_WB),
    .from_WC(Tile_X3Y12_to_WC),
    .from_WD(Tile_X3Y12_to_WD),
    .from_WF(Tile_X3Y12_to_WF),
    .from_WG(Tile_X3Y12_to_WG),
    .from_WH(Tile_X3Y12_to_WH),
    .from_WI(Tile_X3Y12_to_WI),
    .to_EA(Tile_X2Y12_to_EA),
    .to_EB(Tile_X2Y12_to_EB),
    .to_EC(Tile_X2Y12_to_EC),
    .to_ED(Tile_X2Y12_to_ED),
    .to_EF(Tile_X2Y12_to_EF),
    .to_EG(Tile_X2Y12_to_EG),
    .to_EH(Tile_X2Y12_to_EH),
    .to_EI(Tile_X2Y12_to_EI),
    .to_WA(Tile_X2Y12_to_WA),
    .to_WB(Tile_X2Y12_to_WB),
    .to_WC(Tile_X2Y12_to_WC),
    .to_WD(Tile_X2Y12_to_WD),
    .to_WF(Tile_X2Y12_to_WF),
    .to_WG(Tile_X2Y12_to_WG),
    .to_WH(Tile_X2Y12_to_WH),
    .to_WI(Tile_X2Y12_to_WI),
    .to_NA(Tile_X2Y12_to_NA),
    .to_NB(Tile_X2Y12_to_NB),
    .to_NC(Tile_X2Y12_to_NC),
    .to_ND(Tile_X2Y12_to_ND),
    .to_NF(Tile_X2Y12_to_NF),
    .to_NG(Tile_X2Y12_to_NG),
    .to_NH(Tile_X2Y12_to_NH),
    .to_NI(Tile_X2Y12_to_NI),
    .to_SA(Tile_X2Y12_to_SA),
    .to_SB(Tile_X2Y12_to_SB),
    .to_SC(Tile_X2Y12_to_SC),
    .to_SD(Tile_X2Y12_to_SD),
    .to_SF(Tile_X2Y12_to_SF),
    .to_SG(Tile_X2Y12_to_SG),
    .to_SH(Tile_X2Y12_to_SH),
    .to_SI(Tile_X2Y12_to_SI),
    .F_masked1(Tile_X2Y12_F_masked1),
    .F_masked2(Tile_X2Y12_F_masked2),
    .UserCLK(Tile_X2Y13_UserCLKo),
    .UserCLKo(Tile_X2Y12_UserCLKo),
    .rst(Tile_X2Y13_rsto),
    .rsto(Tile_X2Y12_rsto),
    .FrameData(Tile_X1Y12_FrameData_O),
    .FrameData_O(Tile_X2Y12_FrameData_O),
    .FrameStrobe(Tile_X2Y13_FrameStrobe_O),
    .FrameStrobe_O(Tile_X2Y12_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
nonlinear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X3Y12_Emulate_Bitstream)
    )
`endif
    Tile_X3Y12_nonlinear_LMDPL
    (
    .from_NA(Tile_X3Y13_to_NA),
    .from_NB(Tile_X3Y13_to_NB),
    .from_NC(Tile_X3Y13_to_NC),
    .from_ND(Tile_X3Y13_to_ND),
    .from_NF(Tile_X3Y13_to_NF),
    .from_NG(Tile_X3Y13_to_NG),
    .from_NH(Tile_X3Y13_to_NH),
    .from_NI(Tile_X3Y13_to_NI),
    .from_EA(Tile_X2Y12_to_EA),
    .from_EB(Tile_X2Y12_to_EB),
    .from_EC(Tile_X2Y12_to_EC),
    .from_ED(Tile_X2Y12_to_ED),
    .from_EF(Tile_X2Y12_to_EF),
    .from_EG(Tile_X2Y12_to_EG),
    .from_EH(Tile_X2Y12_to_EH),
    .from_EI(Tile_X2Y12_to_EI),
    .from_SA(Tile_X3Y11_to_SA),
    .from_SB(Tile_X3Y11_to_SB),
    .from_SC(Tile_X3Y11_to_SC),
    .from_SD(Tile_X3Y11_to_SD),
    .from_SF(Tile_X3Y11_to_SF),
    .from_SG(Tile_X3Y11_to_SG),
    .from_SH(Tile_X3Y11_to_SH),
    .from_SI(Tile_X3Y11_to_SI),
    .from_WA(Tile_X4Y12_to_WA),
    .from_WB(Tile_X4Y12_to_WB),
    .from_WC(Tile_X4Y12_to_WC),
    .from_WD(Tile_X4Y12_to_WD),
    .from_WF(Tile_X4Y12_to_WF),
    .from_WG(Tile_X4Y12_to_WG),
    .from_WH(Tile_X4Y12_to_WH),
    .from_WI(Tile_X4Y12_to_WI),
    .to_EA(Tile_X3Y12_to_EA),
    .to_EB(Tile_X3Y12_to_EB),
    .to_EC(Tile_X3Y12_to_EC),
    .to_ED(Tile_X3Y12_to_ED),
    .to_EF(Tile_X3Y12_to_EF),
    .to_EG(Tile_X3Y12_to_EG),
    .to_EH(Tile_X3Y12_to_EH),
    .to_EI(Tile_X3Y12_to_EI),
    .to_WA(Tile_X3Y12_to_WA),
    .to_WB(Tile_X3Y12_to_WB),
    .to_WC(Tile_X3Y12_to_WC),
    .to_WD(Tile_X3Y12_to_WD),
    .to_WF(Tile_X3Y12_to_WF),
    .to_WG(Tile_X3Y12_to_WG),
    .to_WH(Tile_X3Y12_to_WH),
    .to_WI(Tile_X3Y12_to_WI),
    .to_NA(Tile_X3Y12_to_NA),
    .to_NB(Tile_X3Y12_to_NB),
    .to_NC(Tile_X3Y12_to_NC),
    .to_ND(Tile_X3Y12_to_ND),
    .to_NF(Tile_X3Y12_to_NF),
    .to_NG(Tile_X3Y12_to_NG),
    .to_NH(Tile_X3Y12_to_NH),
    .to_NI(Tile_X3Y12_to_NI),
    .to_SA(Tile_X3Y12_to_SA),
    .to_SB(Tile_X3Y12_to_SB),
    .to_SC(Tile_X3Y12_to_SC),
    .to_SD(Tile_X3Y12_to_SD),
    .to_SF(Tile_X3Y12_to_SF),
    .to_SG(Tile_X3Y12_to_SG),
    .to_SH(Tile_X3Y12_to_SH),
    .to_SI(Tile_X3Y12_to_SI),
    .R_t(Tile_X3Y12_R_t),
    .R_f(Tile_X3Y12_R_f),
    .F_masked1(Tile_X3Y12_F_masked1),
    .F_masked2(Tile_X3Y12_F_masked2),
    .UserCLK(Tile_X3Y13_UserCLKo),
    .UserCLKo(Tile_X3Y12_UserCLKo),
    .rst(Tile_X3Y13_rsto),
    .rsto(Tile_X3Y12_rsto),
    .FrameData(Tile_X2Y12_FrameData_O),
    .FrameData_O(Tile_X3Y12_FrameData_O),
    .FrameStrobe(Tile_X3Y13_FrameStrobe_O),
    .FrameStrobe_O(Tile_X3Y12_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X4Y12_Emulate_Bitstream)
    )
`endif
    Tile_X4Y12_linear_LMDPL
    (
    .from_NA(Tile_X4Y13_to_NA),
    .from_NB(Tile_X4Y13_to_NB),
    .from_NC(Tile_X4Y13_to_NC),
    .from_ND(Tile_X4Y13_to_ND),
    .from_NF(Tile_X4Y13_to_NF),
    .from_NG(Tile_X4Y13_to_NG),
    .from_NH(Tile_X4Y13_to_NH),
    .from_NI(Tile_X4Y13_to_NI),
    .from_EA(Tile_X3Y12_to_EA),
    .from_EB(Tile_X3Y12_to_EB),
    .from_EC(Tile_X3Y12_to_EC),
    .from_ED(Tile_X3Y12_to_ED),
    .from_EF(Tile_X3Y12_to_EF),
    .from_EG(Tile_X3Y12_to_EG),
    .from_EH(Tile_X3Y12_to_EH),
    .from_EI(Tile_X3Y12_to_EI),
    .from_SA(Tile_X4Y11_to_SA),
    .from_SB(Tile_X4Y11_to_SB),
    .from_SC(Tile_X4Y11_to_SC),
    .from_SD(Tile_X4Y11_to_SD),
    .from_SF(Tile_X4Y11_to_SF),
    .from_SG(Tile_X4Y11_to_SG),
    .from_SH(Tile_X4Y11_to_SH),
    .from_SI(Tile_X4Y11_to_SI),
    .from_WA(Tile_X5Y12_to_WA),
    .from_WB(Tile_X5Y12_to_WB),
    .from_WC(Tile_X5Y12_to_WC),
    .from_WD(Tile_X5Y12_to_WD),
    .from_WF(Tile_X5Y12_to_WF),
    .from_WG(Tile_X5Y12_to_WG),
    .from_WH(Tile_X5Y12_to_WH),
    .from_WI(Tile_X5Y12_to_WI),
    .to_EA(Tile_X4Y12_to_EA),
    .to_EB(Tile_X4Y12_to_EB),
    .to_EC(Tile_X4Y12_to_EC),
    .to_ED(Tile_X4Y12_to_ED),
    .to_EF(Tile_X4Y12_to_EF),
    .to_EG(Tile_X4Y12_to_EG),
    .to_EH(Tile_X4Y12_to_EH),
    .to_EI(Tile_X4Y12_to_EI),
    .to_WA(Tile_X4Y12_to_WA),
    .to_WB(Tile_X4Y12_to_WB),
    .to_WC(Tile_X4Y12_to_WC),
    .to_WD(Tile_X4Y12_to_WD),
    .to_WF(Tile_X4Y12_to_WF),
    .to_WG(Tile_X4Y12_to_WG),
    .to_WH(Tile_X4Y12_to_WH),
    .to_WI(Tile_X4Y12_to_WI),
    .to_NA(Tile_X4Y12_to_NA),
    .to_NB(Tile_X4Y12_to_NB),
    .to_NC(Tile_X4Y12_to_NC),
    .to_ND(Tile_X4Y12_to_ND),
    .to_NF(Tile_X4Y12_to_NF),
    .to_NG(Tile_X4Y12_to_NG),
    .to_NH(Tile_X4Y12_to_NH),
    .to_NI(Tile_X4Y12_to_NI),
    .to_SA(Tile_X4Y12_to_SA),
    .to_SB(Tile_X4Y12_to_SB),
    .to_SC(Tile_X4Y12_to_SC),
    .to_SD(Tile_X4Y12_to_SD),
    .to_SF(Tile_X4Y12_to_SF),
    .to_SG(Tile_X4Y12_to_SG),
    .to_SH(Tile_X4Y12_to_SH),
    .to_SI(Tile_X4Y12_to_SI),
    .F_masked1(Tile_X4Y12_F_masked1),
    .F_masked2(Tile_X4Y12_F_masked2),
    .UserCLK(Tile_X4Y13_UserCLKo),
    .UserCLKo(Tile_X4Y12_UserCLKo),
    .rst(Tile_X4Y13_rsto),
    .rsto(Tile_X4Y12_rsto),
    .FrameData(Tile_X3Y12_FrameData_O),
    .FrameData_O(Tile_X4Y12_FrameData_O),
    .FrameStrobe(Tile_X4Y13_FrameStrobe_O),
    .FrameStrobe_O(Tile_X4Y12_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X5Y12_Emulate_Bitstream)
    )
`endif
    Tile_X5Y12_linear_LMDPL
    (
    .from_NA(Tile_X5Y13_to_NA),
    .from_NB(Tile_X5Y13_to_NB),
    .from_NC(Tile_X5Y13_to_NC),
    .from_ND(Tile_X5Y13_to_ND),
    .from_NF(Tile_X5Y13_to_NF),
    .from_NG(Tile_X5Y13_to_NG),
    .from_NH(Tile_X5Y13_to_NH),
    .from_NI(Tile_X5Y13_to_NI),
    .from_EA(Tile_X4Y12_to_EA),
    .from_EB(Tile_X4Y12_to_EB),
    .from_EC(Tile_X4Y12_to_EC),
    .from_ED(Tile_X4Y12_to_ED),
    .from_EF(Tile_X4Y12_to_EF),
    .from_EG(Tile_X4Y12_to_EG),
    .from_EH(Tile_X4Y12_to_EH),
    .from_EI(Tile_X4Y12_to_EI),
    .from_SA(Tile_X5Y11_to_SA),
    .from_SB(Tile_X5Y11_to_SB),
    .from_SC(Tile_X5Y11_to_SC),
    .from_SD(Tile_X5Y11_to_SD),
    .from_SF(Tile_X5Y11_to_SF),
    .from_SG(Tile_X5Y11_to_SG),
    .from_SH(Tile_X5Y11_to_SH),
    .from_SI(Tile_X5Y11_to_SI),
    .from_WA(Tile_X6Y12_to_WA),
    .from_WB(Tile_X6Y12_to_WB),
    .from_WC(Tile_X6Y12_to_WC),
    .from_WD(Tile_X6Y12_to_WD),
    .from_WF(Tile_X6Y12_to_WF),
    .from_WG(Tile_X6Y12_to_WG),
    .from_WH(Tile_X6Y12_to_WH),
    .from_WI(Tile_X6Y12_to_WI),
    .to_EA(Tile_X5Y12_to_EA),
    .to_EB(Tile_X5Y12_to_EB),
    .to_EC(Tile_X5Y12_to_EC),
    .to_ED(Tile_X5Y12_to_ED),
    .to_EF(Tile_X5Y12_to_EF),
    .to_EG(Tile_X5Y12_to_EG),
    .to_EH(Tile_X5Y12_to_EH),
    .to_EI(Tile_X5Y12_to_EI),
    .to_WA(Tile_X5Y12_to_WA),
    .to_WB(Tile_X5Y12_to_WB),
    .to_WC(Tile_X5Y12_to_WC),
    .to_WD(Tile_X5Y12_to_WD),
    .to_WF(Tile_X5Y12_to_WF),
    .to_WG(Tile_X5Y12_to_WG),
    .to_WH(Tile_X5Y12_to_WH),
    .to_WI(Tile_X5Y12_to_WI),
    .to_NA(Tile_X5Y12_to_NA),
    .to_NB(Tile_X5Y12_to_NB),
    .to_NC(Tile_X5Y12_to_NC),
    .to_ND(Tile_X5Y12_to_ND),
    .to_NF(Tile_X5Y12_to_NF),
    .to_NG(Tile_X5Y12_to_NG),
    .to_NH(Tile_X5Y12_to_NH),
    .to_NI(Tile_X5Y12_to_NI),
    .to_SA(Tile_X5Y12_to_SA),
    .to_SB(Tile_X5Y12_to_SB),
    .to_SC(Tile_X5Y12_to_SC),
    .to_SD(Tile_X5Y12_to_SD),
    .to_SF(Tile_X5Y12_to_SF),
    .to_SG(Tile_X5Y12_to_SG),
    .to_SH(Tile_X5Y12_to_SH),
    .to_SI(Tile_X5Y12_to_SI),
    .F_masked1(Tile_X5Y12_F_masked1),
    .F_masked2(Tile_X5Y12_F_masked2),
    .UserCLK(Tile_X5Y13_UserCLKo),
    .UserCLKo(Tile_X5Y12_UserCLKo),
    .rst(Tile_X5Y13_rsto),
    .rsto(Tile_X5Y12_rsto),
    .FrameData(Tile_X4Y12_FrameData_O),
    .FrameData_O(Tile_X5Y12_FrameData_O),
    .FrameStrobe(Tile_X5Y13_FrameStrobe_O),
    .FrameStrobe_O(Tile_X5Y12_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
nonlinear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X6Y12_Emulate_Bitstream)
    )
`endif
    Tile_X6Y12_nonlinear_LMDPL
    (
    .from_NA(Tile_X6Y13_to_NA),
    .from_NB(Tile_X6Y13_to_NB),
    .from_NC(Tile_X6Y13_to_NC),
    .from_ND(Tile_X6Y13_to_ND),
    .from_NF(Tile_X6Y13_to_NF),
    .from_NG(Tile_X6Y13_to_NG),
    .from_NH(Tile_X6Y13_to_NH),
    .from_NI(Tile_X6Y13_to_NI),
    .from_EA(Tile_X5Y12_to_EA),
    .from_EB(Tile_X5Y12_to_EB),
    .from_EC(Tile_X5Y12_to_EC),
    .from_ED(Tile_X5Y12_to_ED),
    .from_EF(Tile_X5Y12_to_EF),
    .from_EG(Tile_X5Y12_to_EG),
    .from_EH(Tile_X5Y12_to_EH),
    .from_EI(Tile_X5Y12_to_EI),
    .from_SA(Tile_X6Y11_to_SA),
    .from_SB(Tile_X6Y11_to_SB),
    .from_SC(Tile_X6Y11_to_SC),
    .from_SD(Tile_X6Y11_to_SD),
    .from_SF(Tile_X6Y11_to_SF),
    .from_SG(Tile_X6Y11_to_SG),
    .from_SH(Tile_X6Y11_to_SH),
    .from_SI(Tile_X6Y11_to_SI),
    .from_WA(Tile_X7Y12_to_WA),
    .from_WB(Tile_X7Y12_to_WB),
    .from_WC(Tile_X7Y12_to_WC),
    .from_WD(Tile_X7Y12_to_WD),
    .from_WF(Tile_X7Y12_to_WF),
    .from_WG(Tile_X7Y12_to_WG),
    .from_WH(Tile_X7Y12_to_WH),
    .from_WI(Tile_X7Y12_to_WI),
    .to_EA(Tile_X6Y12_to_EA),
    .to_EB(Tile_X6Y12_to_EB),
    .to_EC(Tile_X6Y12_to_EC),
    .to_ED(Tile_X6Y12_to_ED),
    .to_EF(Tile_X6Y12_to_EF),
    .to_EG(Tile_X6Y12_to_EG),
    .to_EH(Tile_X6Y12_to_EH),
    .to_EI(Tile_X6Y12_to_EI),
    .to_WA(Tile_X6Y12_to_WA),
    .to_WB(Tile_X6Y12_to_WB),
    .to_WC(Tile_X6Y12_to_WC),
    .to_WD(Tile_X6Y12_to_WD),
    .to_WF(Tile_X6Y12_to_WF),
    .to_WG(Tile_X6Y12_to_WG),
    .to_WH(Tile_X6Y12_to_WH),
    .to_WI(Tile_X6Y12_to_WI),
    .to_NA(Tile_X6Y12_to_NA),
    .to_NB(Tile_X6Y12_to_NB),
    .to_NC(Tile_X6Y12_to_NC),
    .to_ND(Tile_X6Y12_to_ND),
    .to_NF(Tile_X6Y12_to_NF),
    .to_NG(Tile_X6Y12_to_NG),
    .to_NH(Tile_X6Y12_to_NH),
    .to_NI(Tile_X6Y12_to_NI),
    .to_SA(Tile_X6Y12_to_SA),
    .to_SB(Tile_X6Y12_to_SB),
    .to_SC(Tile_X6Y12_to_SC),
    .to_SD(Tile_X6Y12_to_SD),
    .to_SF(Tile_X6Y12_to_SF),
    .to_SG(Tile_X6Y12_to_SG),
    .to_SH(Tile_X6Y12_to_SH),
    .to_SI(Tile_X6Y12_to_SI),
    .R_t(Tile_X6Y12_R_t),
    .R_f(Tile_X6Y12_R_f),
    .F_masked1(Tile_X6Y12_F_masked1),
    .F_masked2(Tile_X6Y12_F_masked2),
    .UserCLK(Tile_X6Y13_UserCLKo),
    .UserCLKo(Tile_X6Y12_UserCLKo),
    .rst(Tile_X6Y13_rsto),
    .rsto(Tile_X6Y12_rsto),
    .FrameData(Tile_X5Y12_FrameData_O),
    .FrameData_O(Tile_X6Y12_FrameData_O),
    .FrameStrobe(Tile_X6Y13_FrameStrobe_O),
    .FrameStrobe_O(Tile_X6Y12_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X7Y12_Emulate_Bitstream)
    )
`endif
    Tile_X7Y12_linear_LMDPL
    (
    .from_NA(Tile_X7Y13_to_NA),
    .from_NB(Tile_X7Y13_to_NB),
    .from_NC(Tile_X7Y13_to_NC),
    .from_ND(Tile_X7Y13_to_ND),
    .from_NF(Tile_X7Y13_to_NF),
    .from_NG(Tile_X7Y13_to_NG),
    .from_NH(Tile_X7Y13_to_NH),
    .from_NI(Tile_X7Y13_to_NI),
    .from_EA(Tile_X6Y12_to_EA),
    .from_EB(Tile_X6Y12_to_EB),
    .from_EC(Tile_X6Y12_to_EC),
    .from_ED(Tile_X6Y12_to_ED),
    .from_EF(Tile_X6Y12_to_EF),
    .from_EG(Tile_X6Y12_to_EG),
    .from_EH(Tile_X6Y12_to_EH),
    .from_EI(Tile_X6Y12_to_EI),
    .from_SA(Tile_X7Y11_to_SA),
    .from_SB(Tile_X7Y11_to_SB),
    .from_SC(Tile_X7Y11_to_SC),
    .from_SD(Tile_X7Y11_to_SD),
    .from_SF(Tile_X7Y11_to_SF),
    .from_SG(Tile_X7Y11_to_SG),
    .from_SH(Tile_X7Y11_to_SH),
    .from_SI(Tile_X7Y11_to_SI),
    .from_WA(Tile_X8Y12_to_WA),
    .from_WB(Tile_X8Y12_to_WB),
    .from_WC(Tile_X8Y12_to_WC),
    .from_WD(Tile_X8Y12_to_WD),
    .from_WF(Tile_X8Y12_to_WF),
    .from_WG(Tile_X8Y12_to_WG),
    .from_WH(Tile_X8Y12_to_WH),
    .from_WI(Tile_X8Y12_to_WI),
    .to_EA(Tile_X7Y12_to_EA),
    .to_EB(Tile_X7Y12_to_EB),
    .to_EC(Tile_X7Y12_to_EC),
    .to_ED(Tile_X7Y12_to_ED),
    .to_EF(Tile_X7Y12_to_EF),
    .to_EG(Tile_X7Y12_to_EG),
    .to_EH(Tile_X7Y12_to_EH),
    .to_EI(Tile_X7Y12_to_EI),
    .to_WA(Tile_X7Y12_to_WA),
    .to_WB(Tile_X7Y12_to_WB),
    .to_WC(Tile_X7Y12_to_WC),
    .to_WD(Tile_X7Y12_to_WD),
    .to_WF(Tile_X7Y12_to_WF),
    .to_WG(Tile_X7Y12_to_WG),
    .to_WH(Tile_X7Y12_to_WH),
    .to_WI(Tile_X7Y12_to_WI),
    .to_NA(Tile_X7Y12_to_NA),
    .to_NB(Tile_X7Y12_to_NB),
    .to_NC(Tile_X7Y12_to_NC),
    .to_ND(Tile_X7Y12_to_ND),
    .to_NF(Tile_X7Y12_to_NF),
    .to_NG(Tile_X7Y12_to_NG),
    .to_NH(Tile_X7Y12_to_NH),
    .to_NI(Tile_X7Y12_to_NI),
    .to_SA(Tile_X7Y12_to_SA),
    .to_SB(Tile_X7Y12_to_SB),
    .to_SC(Tile_X7Y12_to_SC),
    .to_SD(Tile_X7Y12_to_SD),
    .to_SF(Tile_X7Y12_to_SF),
    .to_SG(Tile_X7Y12_to_SG),
    .to_SH(Tile_X7Y12_to_SH),
    .to_SI(Tile_X7Y12_to_SI),
    .F_masked1(Tile_X7Y12_F_masked1),
    .F_masked2(Tile_X7Y12_F_masked2),
    .UserCLK(Tile_X7Y13_UserCLKo),
    .UserCLKo(Tile_X7Y12_UserCLKo),
    .rst(Tile_X7Y13_rsto),
    .rsto(Tile_X7Y12_rsto),
    .FrameData(Tile_X6Y12_FrameData_O),
    .FrameData_O(Tile_X7Y12_FrameData_O),
    .FrameStrobe(Tile_X7Y13_FrameStrobe_O),
    .FrameStrobe_O(Tile_X7Y12_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
ctrl_to_sec
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X8Y12_Emulate_Bitstream)
    )
`endif
    Tile_X8Y12_ctrl_to_sec
    (
    .from_NA(Tile_X8Y13_to_NA),
    .from_NB(Tile_X8Y13_to_NB),
    .from_NC(Tile_X8Y13_to_NC),
    .from_ND(Tile_X8Y13_to_ND),
    .from_NF(Tile_X8Y13_to_NF),
    .from_NG(Tile_X8Y13_to_NG),
    .from_NH(Tile_X8Y13_to_NH),
    .from_NI(Tile_X8Y13_to_NI),
    .from_EA(Tile_X7Y12_to_EA),
    .from_EB(Tile_X7Y12_to_EB),
    .from_EC(Tile_X7Y12_to_EC),
    .from_ED(Tile_X7Y12_to_ED),
    .from_EF(Tile_X7Y12_to_EF),
    .from_EG(Tile_X7Y12_to_EG),
    .from_EH(Tile_X7Y12_to_EH),
    .from_EI(Tile_X7Y12_to_EI),
    .from_SA(Tile_X8Y11_to_SA),
    .from_SB(Tile_X8Y11_to_SB),
    .from_SC(Tile_X8Y11_to_SC),
    .from_SD(Tile_X8Y11_to_SD),
    .from_SF(Tile_X8Y11_to_SF),
    .from_SG(Tile_X8Y11_to_SG),
    .from_SH(Tile_X8Y11_to_SH),
    .from_SI(Tile_X8Y11_to_SI),
    .from_WA_1s(Tile_X9Y12_to_WA_1s),
    .from_WB_1s(Tile_X9Y12_to_WB_1s),
    .from_WC_1s(Tile_X9Y12_to_WC_1s),
    .from_WD_1s(Tile_X9Y12_to_WD_1s),
    .from_WF_1s(Tile_X9Y12_to_WF_1s),
    .from_WG_1s(Tile_X9Y12_to_WG_1s),
    .from_WH_1s(Tile_X9Y12_to_WH_1s),
    .from_WI_1s(Tile_X9Y12_to_WI_1s),
    .to_WA(Tile_X8Y12_to_WA),
    .to_WB(Tile_X8Y12_to_WB),
    .to_WC(Tile_X8Y12_to_WC),
    .to_WD(Tile_X8Y12_to_WD),
    .to_WF(Tile_X8Y12_to_WF),
    .to_WG(Tile_X8Y12_to_WG),
    .to_WH(Tile_X8Y12_to_WH),
    .to_WI(Tile_X8Y12_to_WI),
    .to_NA(Tile_X8Y12_to_NA),
    .to_NB(Tile_X8Y12_to_NB),
    .to_NC(Tile_X8Y12_to_NC),
    .to_ND(Tile_X8Y12_to_ND),
    .to_NF(Tile_X8Y12_to_NF),
    .to_NG(Tile_X8Y12_to_NG),
    .to_NH(Tile_X8Y12_to_NH),
    .to_NI(Tile_X8Y12_to_NI),
    .to_SA(Tile_X8Y12_to_SA),
    .to_SB(Tile_X8Y12_to_SB),
    .to_SC(Tile_X8Y12_to_SC),
    .to_SD(Tile_X8Y12_to_SD),
    .to_SF(Tile_X8Y12_to_SF),
    .to_SG(Tile_X8Y12_to_SG),
    .to_SH(Tile_X8Y12_to_SH),
    .to_SI(Tile_X8Y12_to_SI),
    .UserCLK(Tile_X8Y13_UserCLKo),
    .UserCLKo(Tile_X8Y12_UserCLKo),
    .rst(Tile_X8Y13_rsto),
    .rsto(Tile_X8Y12_rsto),
    .FrameData(Tile_X7Y12_FrameData_O),
    .FrameData_O(Tile_X8Y12_FrameData_O),
    .FrameStrobe(Tile_X8Y13_FrameStrobe_O),
    .FrameStrobe_O(Tile_X8Y12_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
combined_WDDL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X9Y12_Emulate_Bitstream)
    )
`endif
    Tile_X9Y12_combined_WDDL
    (
    .from_NA_1s(Tile_X9Y13_to_NA_1s),
    .from_NB_1s(Tile_X9Y13_to_NB_1s),
    .from_NC_1s(Tile_X9Y13_to_NC_1s),
    .from_ND_1s(Tile_X9Y13_to_ND_1s),
    .from_NF_1s(Tile_X9Y13_to_NF_1s),
    .from_NG_1s(Tile_X9Y13_to_NG_1s),
    .from_NH_1s(Tile_X9Y13_to_NH_1s),
    .from_NI_1s(Tile_X9Y13_to_NI_1s),
    .from_SA_1s(Tile_X9Y11_to_SA_1s),
    .from_SB_1s(Tile_X9Y11_to_SB_1s),
    .from_SC_1s(Tile_X9Y11_to_SC_1s),
    .from_SD_1s(Tile_X9Y11_to_SD_1s),
    .from_SF_1s(Tile_X9Y11_to_SF_1s),
    .from_SG_1s(Tile_X9Y11_to_SG_1s),
    .from_SH_1s(Tile_X9Y11_to_SH_1s),
    .from_SI_1s(Tile_X9Y11_to_SI_1s),
    .from_WA_1s(Tile_X10Y12_to_WA_1s),
    .from_WB_1s(Tile_X10Y12_to_WB_1s),
    .from_WC_1s(Tile_X10Y12_to_WC_1s),
    .from_WD_1s(Tile_X10Y12_to_WD_1s),
    .from_WF_1s(Tile_X10Y12_to_WF_1s),
    .from_WG_1s(Tile_X10Y12_to_WG_1s),
    .from_WH_1s(Tile_X10Y12_to_WH_1s),
    .from_WI_1s(Tile_X10Y12_to_WI_1s),
    .to_EA_1s(Tile_X9Y12_to_EA_1s),
    .to_EB_1s(Tile_X9Y12_to_EB_1s),
    .to_EC_1s(Tile_X9Y12_to_EC_1s),
    .to_ED_1s(Tile_X9Y12_to_ED_1s),
    .to_EF_1s(Tile_X9Y12_to_EF_1s),
    .to_EG_1s(Tile_X9Y12_to_EG_1s),
    .to_EH_1s(Tile_X9Y12_to_EH_1s),
    .to_EI_1s(Tile_X9Y12_to_EI_1s),
    .to_WA_1s(Tile_X9Y12_to_WA_1s),
    .to_WB_1s(Tile_X9Y12_to_WB_1s),
    .to_WC_1s(Tile_X9Y12_to_WC_1s),
    .to_WD_1s(Tile_X9Y12_to_WD_1s),
    .to_WF_1s(Tile_X9Y12_to_WF_1s),
    .to_WG_1s(Tile_X9Y12_to_WG_1s),
    .to_WH_1s(Tile_X9Y12_to_WH_1s),
    .to_WI_1s(Tile_X9Y12_to_WI_1s),
    .to_NA_1s(Tile_X9Y12_to_NA_1s),
    .to_NB_1s(Tile_X9Y12_to_NB_1s),
    .to_NC_1s(Tile_X9Y12_to_NC_1s),
    .to_ND_1s(Tile_X9Y12_to_ND_1s),
    .to_NF_1s(Tile_X9Y12_to_NF_1s),
    .to_NG_1s(Tile_X9Y12_to_NG_1s),
    .to_NH_1s(Tile_X9Y12_to_NH_1s),
    .to_NI_1s(Tile_X9Y12_to_NI_1s),
    .to_SA_1s(Tile_X9Y12_to_SA_1s),
    .to_SB_1s(Tile_X9Y12_to_SB_1s),
    .to_SC_1s(Tile_X9Y12_to_SC_1s),
    .to_SD_1s(Tile_X9Y12_to_SD_1s),
    .to_SF_1s(Tile_X9Y12_to_SF_1s),
    .to_SG_1s(Tile_X9Y12_to_SG_1s),
    .to_SH_1s(Tile_X9Y12_to_SH_1s),
    .to_SI_1s(Tile_X9Y12_to_SI_1s),
    .F_ctrl(Tile_X9Y12_F_ctrl),
    .UserCLK(Tile_X9Y13_UserCLKo),
    .UserCLKo(Tile_X9Y12_UserCLKo),
    .rst(Tile_X9Y13_rsto),
    .rsto(Tile_X9Y12_rsto),
    .FrameData(Tile_X8Y12_FrameData_O),
    .FrameData_O(Tile_X9Y12_FrameData_O),
    .FrameStrobe(Tile_X9Y13_FrameStrobe_O),
    .FrameStrobe_O(Tile_X9Y12_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
ctrl_IO
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X10Y12_Emulate_Bitstream)
    )
`endif
    Tile_X10Y12_ctrl_IO
    (
    .from_EA_1s(Tile_X9Y12_to_EA_1s),
    .from_EB_1s(Tile_X9Y12_to_EB_1s),
    .from_EC_1s(Tile_X9Y12_to_EC_1s),
    .from_ED_1s(Tile_X9Y12_to_ED_1s),
    .from_EF_1s(Tile_X9Y12_to_EF_1s),
    .from_EG_1s(Tile_X9Y12_to_EG_1s),
    .from_EH_1s(Tile_X9Y12_to_EH_1s),
    .from_EI_1s(Tile_X9Y12_to_EI_1s),
    .to_WA_1s(Tile_X10Y12_to_WA_1s),
    .to_WB_1s(Tile_X10Y12_to_WB_1s),
    .to_WC_1s(Tile_X10Y12_to_WC_1s),
    .to_WD_1s(Tile_X10Y12_to_WD_1s),
    .to_WF_1s(Tile_X10Y12_to_WF_1s),
    .to_WG_1s(Tile_X10Y12_to_WG_1s),
    .to_WH_1s(Tile_X10Y12_to_WH_1s),
    .to_WI_1s(Tile_X10Y12_to_WI_1s),
    .A_O_top_0_t(Tile_X10Y12_A_O_top_0_t),
    .A_O_top_0_f(Tile_X10Y12_A_O_top_0_f),
    .A_prech2(Tile_X10Y12_A_prech2),
    .A_DR_fault(Tile_X10Y12_A_DR_fault),
    .A_I_top_0_t(Tile_X10Y12_A_I_top_0_t),
    .A_I_top_0_f(Tile_X10Y12_A_I_top_0_f),
    .A_T_top(Tile_X10Y12_A_T_top),
    .A_F_ctrl(Tile_X10Y12_A_F_ctrl),
    .UserCLK(Tile_X10Y13_UserCLKo),
    .UserCLKo(Tile_X10Y12_UserCLKo),
    .rst(Tile_X10Y13_rsto),
    .rsto(Tile_X10Y12_rsto),
    .FrameData(Tile_X9Y12_FrameData_O),
    .FrameData_O(Tile_X10Y12_FrameData_O),
    .FrameStrobe(Tile_X10Y13_FrameStrobe_O),
    .FrameStrobe_O(Tile_X10Y12_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
W_IO_custom
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X0Y13_Emulate_Bitstream)
    )
`endif
    Tile_X0Y13_W_IO_custom
    (
    .from_NA(Tile_X0Y14_to_NA),
    .from_NB(Tile_X0Y14_to_NB),
    .from_NC(Tile_X0Y14_to_NC),
    .from_ND(Tile_X0Y14_to_ND),
    .from_NF(Tile_X0Y14_to_NF),
    .from_NG(Tile_X0Y14_to_NG),
    .from_NH(Tile_X0Y14_to_NH),
    .from_NI(Tile_X0Y14_to_NI),
    .from_SA(Tile_X0Y12_to_SA),
    .from_SB(Tile_X0Y12_to_SB),
    .from_SC(Tile_X0Y12_to_SC),
    .from_SD(Tile_X0Y12_to_SD),
    .from_SF(Tile_X0Y12_to_SF),
    .from_SG(Tile_X0Y12_to_SG),
    .from_SH(Tile_X0Y12_to_SH),
    .from_SI(Tile_X0Y12_to_SI),
    .from_WA(Tile_X1Y13_to_WA),
    .from_WB(Tile_X1Y13_to_WB),
    .from_WC(Tile_X1Y13_to_WC),
    .from_WD(Tile_X1Y13_to_WD),
    .from_WF(Tile_X1Y13_to_WF),
    .from_WG(Tile_X1Y13_to_WG),
    .from_WH(Tile_X1Y13_to_WH),
    .from_WI(Tile_X1Y13_to_WI),
    .to_EA(Tile_X0Y13_to_EA),
    .to_EB(Tile_X0Y13_to_EB),
    .to_EC(Tile_X0Y13_to_EC),
    .to_ED(Tile_X0Y13_to_ED),
    .to_EF(Tile_X0Y13_to_EF),
    .to_EG(Tile_X0Y13_to_EG),
    .to_EH(Tile_X0Y13_to_EH),
    .to_EI(Tile_X0Y13_to_EI),
    .to_NA(Tile_X0Y13_to_NA),
    .to_NB(Tile_X0Y13_to_NB),
    .to_NC(Tile_X0Y13_to_NC),
    .to_ND(Tile_X0Y13_to_ND),
    .to_NF(Tile_X0Y13_to_NF),
    .to_NG(Tile_X0Y13_to_NG),
    .to_NH(Tile_X0Y13_to_NH),
    .to_NI(Tile_X0Y13_to_NI),
    .to_SA(Tile_X0Y13_to_SA),
    .to_SB(Tile_X0Y13_to_SB),
    .to_SC(Tile_X0Y13_to_SC),
    .to_SD(Tile_X0Y13_to_SD),
    .to_SF(Tile_X0Y13_to_SF),
    .to_SG(Tile_X0Y13_to_SG),
    .to_SH(Tile_X0Y13_to_SH),
    .to_SI(Tile_X0Y13_to_SI),
    .A_O_top_0_t(Tile_X0Y13_A_O_top_0_t),
    .A_O_top_0_f(Tile_X0Y13_A_O_top_0_f),
    .A_O_top_1_t(Tile_X0Y13_A_O_top_1_t),
    .A_O_top_1_f(Tile_X0Y13_A_O_top_1_f),
    .A_prech1(Tile_X0Y13_A_prech1),
    .A_prech2(Tile_X0Y13_A_prech2),
    .A_DR_fault(Tile_X0Y13_A_DR_fault),
    .A_I_top_0_t(Tile_X0Y13_A_I_top_0_t),
    .A_I_top_0_f(Tile_X0Y13_A_I_top_0_f),
    .A_I_top_1_t(Tile_X0Y13_A_I_top_1_t),
    .A_I_top_1_f(Tile_X0Y13_A_I_top_1_f),
    .A_T_top(Tile_X0Y13_A_T_top),
    .A_F_masked1(Tile_X0Y13_A_F_masked1),
    .A_F_masked2(Tile_X0Y13_A_F_masked2),
    .A_config_C_bit0(Tile_X0Y13_A_config_C_bit0),
    .A_config_C_bit1(Tile_X0Y13_A_config_C_bit1),
    .A_config_C_bit2(Tile_X0Y13_A_config_C_bit2),
    .A_config_C_bit3(Tile_X0Y13_A_config_C_bit3),
    .B_config_C_bit0(Tile_X0Y13_B_config_C_bit0),
    .B_config_C_bit1(Tile_X0Y13_B_config_C_bit1),
    .B_config_C_bit2(Tile_X0Y13_B_config_C_bit2),
    .B_config_C_bit3(Tile_X0Y13_B_config_C_bit3),
    .UserCLK(Tile_X0Y14_UserCLKo),
    .UserCLKo(Tile_X0Y13_UserCLKo),
    .rst(Tile_X0Y14_rsto),
    .rsto(Tile_X0Y13_rsto),
    .FrameData(Tile_Y13_FrameData),
    .FrameData_O(Tile_X0Y13_FrameData_O),
    .FrameStrobe(Tile_X0Y14_FrameStrobe_O),
    .FrameStrobe_O(Tile_X0Y13_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X1Y13_Emulate_Bitstream)
    )
`endif
    Tile_X1Y13_linear_LMDPL
    (
    .from_NA(Tile_X1Y14_to_NA),
    .from_NB(Tile_X1Y14_to_NB),
    .from_NC(Tile_X1Y14_to_NC),
    .from_ND(Tile_X1Y14_to_ND),
    .from_NF(Tile_X1Y14_to_NF),
    .from_NG(Tile_X1Y14_to_NG),
    .from_NH(Tile_X1Y14_to_NH),
    .from_NI(Tile_X1Y14_to_NI),
    .from_EA(Tile_X0Y13_to_EA),
    .from_EB(Tile_X0Y13_to_EB),
    .from_EC(Tile_X0Y13_to_EC),
    .from_ED(Tile_X0Y13_to_ED),
    .from_EF(Tile_X0Y13_to_EF),
    .from_EG(Tile_X0Y13_to_EG),
    .from_EH(Tile_X0Y13_to_EH),
    .from_EI(Tile_X0Y13_to_EI),
    .from_SA(Tile_X1Y12_to_SA),
    .from_SB(Tile_X1Y12_to_SB),
    .from_SC(Tile_X1Y12_to_SC),
    .from_SD(Tile_X1Y12_to_SD),
    .from_SF(Tile_X1Y12_to_SF),
    .from_SG(Tile_X1Y12_to_SG),
    .from_SH(Tile_X1Y12_to_SH),
    .from_SI(Tile_X1Y12_to_SI),
    .from_WA(Tile_X2Y13_to_WA),
    .from_WB(Tile_X2Y13_to_WB),
    .from_WC(Tile_X2Y13_to_WC),
    .from_WD(Tile_X2Y13_to_WD),
    .from_WF(Tile_X2Y13_to_WF),
    .from_WG(Tile_X2Y13_to_WG),
    .from_WH(Tile_X2Y13_to_WH),
    .from_WI(Tile_X2Y13_to_WI),
    .to_EA(Tile_X1Y13_to_EA),
    .to_EB(Tile_X1Y13_to_EB),
    .to_EC(Tile_X1Y13_to_EC),
    .to_ED(Tile_X1Y13_to_ED),
    .to_EF(Tile_X1Y13_to_EF),
    .to_EG(Tile_X1Y13_to_EG),
    .to_EH(Tile_X1Y13_to_EH),
    .to_EI(Tile_X1Y13_to_EI),
    .to_WA(Tile_X1Y13_to_WA),
    .to_WB(Tile_X1Y13_to_WB),
    .to_WC(Tile_X1Y13_to_WC),
    .to_WD(Tile_X1Y13_to_WD),
    .to_WF(Tile_X1Y13_to_WF),
    .to_WG(Tile_X1Y13_to_WG),
    .to_WH(Tile_X1Y13_to_WH),
    .to_WI(Tile_X1Y13_to_WI),
    .to_NA(Tile_X1Y13_to_NA),
    .to_NB(Tile_X1Y13_to_NB),
    .to_NC(Tile_X1Y13_to_NC),
    .to_ND(Tile_X1Y13_to_ND),
    .to_NF(Tile_X1Y13_to_NF),
    .to_NG(Tile_X1Y13_to_NG),
    .to_NH(Tile_X1Y13_to_NH),
    .to_NI(Tile_X1Y13_to_NI),
    .to_SA(Tile_X1Y13_to_SA),
    .to_SB(Tile_X1Y13_to_SB),
    .to_SC(Tile_X1Y13_to_SC),
    .to_SD(Tile_X1Y13_to_SD),
    .to_SF(Tile_X1Y13_to_SF),
    .to_SG(Tile_X1Y13_to_SG),
    .to_SH(Tile_X1Y13_to_SH),
    .to_SI(Tile_X1Y13_to_SI),
    .F_masked1(Tile_X1Y13_F_masked1),
    .F_masked2(Tile_X1Y13_F_masked2),
    .UserCLK(Tile_X1Y14_UserCLKo),
    .UserCLKo(Tile_X1Y13_UserCLKo),
    .rst(Tile_X1Y14_rsto),
    .rsto(Tile_X1Y13_rsto),
    .FrameData(Tile_X0Y13_FrameData_O),
    .FrameData_O(Tile_X1Y13_FrameData_O),
    .FrameStrobe(Tile_X1Y14_FrameStrobe_O),
    .FrameStrobe_O(Tile_X1Y13_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X2Y13_Emulate_Bitstream)
    )
`endif
    Tile_X2Y13_linear_LMDPL
    (
    .from_NA(Tile_X2Y14_to_NA),
    .from_NB(Tile_X2Y14_to_NB),
    .from_NC(Tile_X2Y14_to_NC),
    .from_ND(Tile_X2Y14_to_ND),
    .from_NF(Tile_X2Y14_to_NF),
    .from_NG(Tile_X2Y14_to_NG),
    .from_NH(Tile_X2Y14_to_NH),
    .from_NI(Tile_X2Y14_to_NI),
    .from_EA(Tile_X1Y13_to_EA),
    .from_EB(Tile_X1Y13_to_EB),
    .from_EC(Tile_X1Y13_to_EC),
    .from_ED(Tile_X1Y13_to_ED),
    .from_EF(Tile_X1Y13_to_EF),
    .from_EG(Tile_X1Y13_to_EG),
    .from_EH(Tile_X1Y13_to_EH),
    .from_EI(Tile_X1Y13_to_EI),
    .from_SA(Tile_X2Y12_to_SA),
    .from_SB(Tile_X2Y12_to_SB),
    .from_SC(Tile_X2Y12_to_SC),
    .from_SD(Tile_X2Y12_to_SD),
    .from_SF(Tile_X2Y12_to_SF),
    .from_SG(Tile_X2Y12_to_SG),
    .from_SH(Tile_X2Y12_to_SH),
    .from_SI(Tile_X2Y12_to_SI),
    .from_WA(Tile_X3Y13_to_WA),
    .from_WB(Tile_X3Y13_to_WB),
    .from_WC(Tile_X3Y13_to_WC),
    .from_WD(Tile_X3Y13_to_WD),
    .from_WF(Tile_X3Y13_to_WF),
    .from_WG(Tile_X3Y13_to_WG),
    .from_WH(Tile_X3Y13_to_WH),
    .from_WI(Tile_X3Y13_to_WI),
    .to_EA(Tile_X2Y13_to_EA),
    .to_EB(Tile_X2Y13_to_EB),
    .to_EC(Tile_X2Y13_to_EC),
    .to_ED(Tile_X2Y13_to_ED),
    .to_EF(Tile_X2Y13_to_EF),
    .to_EG(Tile_X2Y13_to_EG),
    .to_EH(Tile_X2Y13_to_EH),
    .to_EI(Tile_X2Y13_to_EI),
    .to_WA(Tile_X2Y13_to_WA),
    .to_WB(Tile_X2Y13_to_WB),
    .to_WC(Tile_X2Y13_to_WC),
    .to_WD(Tile_X2Y13_to_WD),
    .to_WF(Tile_X2Y13_to_WF),
    .to_WG(Tile_X2Y13_to_WG),
    .to_WH(Tile_X2Y13_to_WH),
    .to_WI(Tile_X2Y13_to_WI),
    .to_NA(Tile_X2Y13_to_NA),
    .to_NB(Tile_X2Y13_to_NB),
    .to_NC(Tile_X2Y13_to_NC),
    .to_ND(Tile_X2Y13_to_ND),
    .to_NF(Tile_X2Y13_to_NF),
    .to_NG(Tile_X2Y13_to_NG),
    .to_NH(Tile_X2Y13_to_NH),
    .to_NI(Tile_X2Y13_to_NI),
    .to_SA(Tile_X2Y13_to_SA),
    .to_SB(Tile_X2Y13_to_SB),
    .to_SC(Tile_X2Y13_to_SC),
    .to_SD(Tile_X2Y13_to_SD),
    .to_SF(Tile_X2Y13_to_SF),
    .to_SG(Tile_X2Y13_to_SG),
    .to_SH(Tile_X2Y13_to_SH),
    .to_SI(Tile_X2Y13_to_SI),
    .F_masked1(Tile_X2Y13_F_masked1),
    .F_masked2(Tile_X2Y13_F_masked2),
    .UserCLK(Tile_X2Y14_UserCLKo),
    .UserCLKo(Tile_X2Y13_UserCLKo),
    .rst(Tile_X2Y14_rsto),
    .rsto(Tile_X2Y13_rsto),
    .FrameData(Tile_X1Y13_FrameData_O),
    .FrameData_O(Tile_X2Y13_FrameData_O),
    .FrameStrobe(Tile_X2Y14_FrameStrobe_O),
    .FrameStrobe_O(Tile_X2Y13_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
nonlinear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X3Y13_Emulate_Bitstream)
    )
`endif
    Tile_X3Y13_nonlinear_LMDPL
    (
    .from_NA(Tile_X3Y14_to_NA),
    .from_NB(Tile_X3Y14_to_NB),
    .from_NC(Tile_X3Y14_to_NC),
    .from_ND(Tile_X3Y14_to_ND),
    .from_NF(Tile_X3Y14_to_NF),
    .from_NG(Tile_X3Y14_to_NG),
    .from_NH(Tile_X3Y14_to_NH),
    .from_NI(Tile_X3Y14_to_NI),
    .from_EA(Tile_X2Y13_to_EA),
    .from_EB(Tile_X2Y13_to_EB),
    .from_EC(Tile_X2Y13_to_EC),
    .from_ED(Tile_X2Y13_to_ED),
    .from_EF(Tile_X2Y13_to_EF),
    .from_EG(Tile_X2Y13_to_EG),
    .from_EH(Tile_X2Y13_to_EH),
    .from_EI(Tile_X2Y13_to_EI),
    .from_SA(Tile_X3Y12_to_SA),
    .from_SB(Tile_X3Y12_to_SB),
    .from_SC(Tile_X3Y12_to_SC),
    .from_SD(Tile_X3Y12_to_SD),
    .from_SF(Tile_X3Y12_to_SF),
    .from_SG(Tile_X3Y12_to_SG),
    .from_SH(Tile_X3Y12_to_SH),
    .from_SI(Tile_X3Y12_to_SI),
    .from_WA(Tile_X4Y13_to_WA),
    .from_WB(Tile_X4Y13_to_WB),
    .from_WC(Tile_X4Y13_to_WC),
    .from_WD(Tile_X4Y13_to_WD),
    .from_WF(Tile_X4Y13_to_WF),
    .from_WG(Tile_X4Y13_to_WG),
    .from_WH(Tile_X4Y13_to_WH),
    .from_WI(Tile_X4Y13_to_WI),
    .to_EA(Tile_X3Y13_to_EA),
    .to_EB(Tile_X3Y13_to_EB),
    .to_EC(Tile_X3Y13_to_EC),
    .to_ED(Tile_X3Y13_to_ED),
    .to_EF(Tile_X3Y13_to_EF),
    .to_EG(Tile_X3Y13_to_EG),
    .to_EH(Tile_X3Y13_to_EH),
    .to_EI(Tile_X3Y13_to_EI),
    .to_WA(Tile_X3Y13_to_WA),
    .to_WB(Tile_X3Y13_to_WB),
    .to_WC(Tile_X3Y13_to_WC),
    .to_WD(Tile_X3Y13_to_WD),
    .to_WF(Tile_X3Y13_to_WF),
    .to_WG(Tile_X3Y13_to_WG),
    .to_WH(Tile_X3Y13_to_WH),
    .to_WI(Tile_X3Y13_to_WI),
    .to_NA(Tile_X3Y13_to_NA),
    .to_NB(Tile_X3Y13_to_NB),
    .to_NC(Tile_X3Y13_to_NC),
    .to_ND(Tile_X3Y13_to_ND),
    .to_NF(Tile_X3Y13_to_NF),
    .to_NG(Tile_X3Y13_to_NG),
    .to_NH(Tile_X3Y13_to_NH),
    .to_NI(Tile_X3Y13_to_NI),
    .to_SA(Tile_X3Y13_to_SA),
    .to_SB(Tile_X3Y13_to_SB),
    .to_SC(Tile_X3Y13_to_SC),
    .to_SD(Tile_X3Y13_to_SD),
    .to_SF(Tile_X3Y13_to_SF),
    .to_SG(Tile_X3Y13_to_SG),
    .to_SH(Tile_X3Y13_to_SH),
    .to_SI(Tile_X3Y13_to_SI),
    .R_t(Tile_X3Y13_R_t),
    .R_f(Tile_X3Y13_R_f),
    .F_masked1(Tile_X3Y13_F_masked1),
    .F_masked2(Tile_X3Y13_F_masked2),
    .UserCLK(Tile_X3Y14_UserCLKo),
    .UserCLKo(Tile_X3Y13_UserCLKo),
    .rst(Tile_X3Y14_rsto),
    .rsto(Tile_X3Y13_rsto),
    .FrameData(Tile_X2Y13_FrameData_O),
    .FrameData_O(Tile_X3Y13_FrameData_O),
    .FrameStrobe(Tile_X3Y14_FrameStrobe_O),
    .FrameStrobe_O(Tile_X3Y13_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X4Y13_Emulate_Bitstream)
    )
`endif
    Tile_X4Y13_linear_LMDPL
    (
    .from_NA(Tile_X4Y14_to_NA),
    .from_NB(Tile_X4Y14_to_NB),
    .from_NC(Tile_X4Y14_to_NC),
    .from_ND(Tile_X4Y14_to_ND),
    .from_NF(Tile_X4Y14_to_NF),
    .from_NG(Tile_X4Y14_to_NG),
    .from_NH(Tile_X4Y14_to_NH),
    .from_NI(Tile_X4Y14_to_NI),
    .from_EA(Tile_X3Y13_to_EA),
    .from_EB(Tile_X3Y13_to_EB),
    .from_EC(Tile_X3Y13_to_EC),
    .from_ED(Tile_X3Y13_to_ED),
    .from_EF(Tile_X3Y13_to_EF),
    .from_EG(Tile_X3Y13_to_EG),
    .from_EH(Tile_X3Y13_to_EH),
    .from_EI(Tile_X3Y13_to_EI),
    .from_SA(Tile_X4Y12_to_SA),
    .from_SB(Tile_X4Y12_to_SB),
    .from_SC(Tile_X4Y12_to_SC),
    .from_SD(Tile_X4Y12_to_SD),
    .from_SF(Tile_X4Y12_to_SF),
    .from_SG(Tile_X4Y12_to_SG),
    .from_SH(Tile_X4Y12_to_SH),
    .from_SI(Tile_X4Y12_to_SI),
    .from_WA(Tile_X5Y13_to_WA),
    .from_WB(Tile_X5Y13_to_WB),
    .from_WC(Tile_X5Y13_to_WC),
    .from_WD(Tile_X5Y13_to_WD),
    .from_WF(Tile_X5Y13_to_WF),
    .from_WG(Tile_X5Y13_to_WG),
    .from_WH(Tile_X5Y13_to_WH),
    .from_WI(Tile_X5Y13_to_WI),
    .to_EA(Tile_X4Y13_to_EA),
    .to_EB(Tile_X4Y13_to_EB),
    .to_EC(Tile_X4Y13_to_EC),
    .to_ED(Tile_X4Y13_to_ED),
    .to_EF(Tile_X4Y13_to_EF),
    .to_EG(Tile_X4Y13_to_EG),
    .to_EH(Tile_X4Y13_to_EH),
    .to_EI(Tile_X4Y13_to_EI),
    .to_WA(Tile_X4Y13_to_WA),
    .to_WB(Tile_X4Y13_to_WB),
    .to_WC(Tile_X4Y13_to_WC),
    .to_WD(Tile_X4Y13_to_WD),
    .to_WF(Tile_X4Y13_to_WF),
    .to_WG(Tile_X4Y13_to_WG),
    .to_WH(Tile_X4Y13_to_WH),
    .to_WI(Tile_X4Y13_to_WI),
    .to_NA(Tile_X4Y13_to_NA),
    .to_NB(Tile_X4Y13_to_NB),
    .to_NC(Tile_X4Y13_to_NC),
    .to_ND(Tile_X4Y13_to_ND),
    .to_NF(Tile_X4Y13_to_NF),
    .to_NG(Tile_X4Y13_to_NG),
    .to_NH(Tile_X4Y13_to_NH),
    .to_NI(Tile_X4Y13_to_NI),
    .to_SA(Tile_X4Y13_to_SA),
    .to_SB(Tile_X4Y13_to_SB),
    .to_SC(Tile_X4Y13_to_SC),
    .to_SD(Tile_X4Y13_to_SD),
    .to_SF(Tile_X4Y13_to_SF),
    .to_SG(Tile_X4Y13_to_SG),
    .to_SH(Tile_X4Y13_to_SH),
    .to_SI(Tile_X4Y13_to_SI),
    .F_masked1(Tile_X4Y13_F_masked1),
    .F_masked2(Tile_X4Y13_F_masked2),
    .UserCLK(Tile_X4Y14_UserCLKo),
    .UserCLKo(Tile_X4Y13_UserCLKo),
    .rst(Tile_X4Y14_rsto),
    .rsto(Tile_X4Y13_rsto),
    .FrameData(Tile_X3Y13_FrameData_O),
    .FrameData_O(Tile_X4Y13_FrameData_O),
    .FrameStrobe(Tile_X4Y14_FrameStrobe_O),
    .FrameStrobe_O(Tile_X4Y13_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X5Y13_Emulate_Bitstream)
    )
`endif
    Tile_X5Y13_linear_LMDPL
    (
    .from_NA(Tile_X5Y14_to_NA),
    .from_NB(Tile_X5Y14_to_NB),
    .from_NC(Tile_X5Y14_to_NC),
    .from_ND(Tile_X5Y14_to_ND),
    .from_NF(Tile_X5Y14_to_NF),
    .from_NG(Tile_X5Y14_to_NG),
    .from_NH(Tile_X5Y14_to_NH),
    .from_NI(Tile_X5Y14_to_NI),
    .from_EA(Tile_X4Y13_to_EA),
    .from_EB(Tile_X4Y13_to_EB),
    .from_EC(Tile_X4Y13_to_EC),
    .from_ED(Tile_X4Y13_to_ED),
    .from_EF(Tile_X4Y13_to_EF),
    .from_EG(Tile_X4Y13_to_EG),
    .from_EH(Tile_X4Y13_to_EH),
    .from_EI(Tile_X4Y13_to_EI),
    .from_SA(Tile_X5Y12_to_SA),
    .from_SB(Tile_X5Y12_to_SB),
    .from_SC(Tile_X5Y12_to_SC),
    .from_SD(Tile_X5Y12_to_SD),
    .from_SF(Tile_X5Y12_to_SF),
    .from_SG(Tile_X5Y12_to_SG),
    .from_SH(Tile_X5Y12_to_SH),
    .from_SI(Tile_X5Y12_to_SI),
    .from_WA(Tile_X6Y13_to_WA),
    .from_WB(Tile_X6Y13_to_WB),
    .from_WC(Tile_X6Y13_to_WC),
    .from_WD(Tile_X6Y13_to_WD),
    .from_WF(Tile_X6Y13_to_WF),
    .from_WG(Tile_X6Y13_to_WG),
    .from_WH(Tile_X6Y13_to_WH),
    .from_WI(Tile_X6Y13_to_WI),
    .to_EA(Tile_X5Y13_to_EA),
    .to_EB(Tile_X5Y13_to_EB),
    .to_EC(Tile_X5Y13_to_EC),
    .to_ED(Tile_X5Y13_to_ED),
    .to_EF(Tile_X5Y13_to_EF),
    .to_EG(Tile_X5Y13_to_EG),
    .to_EH(Tile_X5Y13_to_EH),
    .to_EI(Tile_X5Y13_to_EI),
    .to_WA(Tile_X5Y13_to_WA),
    .to_WB(Tile_X5Y13_to_WB),
    .to_WC(Tile_X5Y13_to_WC),
    .to_WD(Tile_X5Y13_to_WD),
    .to_WF(Tile_X5Y13_to_WF),
    .to_WG(Tile_X5Y13_to_WG),
    .to_WH(Tile_X5Y13_to_WH),
    .to_WI(Tile_X5Y13_to_WI),
    .to_NA(Tile_X5Y13_to_NA),
    .to_NB(Tile_X5Y13_to_NB),
    .to_NC(Tile_X5Y13_to_NC),
    .to_ND(Tile_X5Y13_to_ND),
    .to_NF(Tile_X5Y13_to_NF),
    .to_NG(Tile_X5Y13_to_NG),
    .to_NH(Tile_X5Y13_to_NH),
    .to_NI(Tile_X5Y13_to_NI),
    .to_SA(Tile_X5Y13_to_SA),
    .to_SB(Tile_X5Y13_to_SB),
    .to_SC(Tile_X5Y13_to_SC),
    .to_SD(Tile_X5Y13_to_SD),
    .to_SF(Tile_X5Y13_to_SF),
    .to_SG(Tile_X5Y13_to_SG),
    .to_SH(Tile_X5Y13_to_SH),
    .to_SI(Tile_X5Y13_to_SI),
    .F_masked1(Tile_X5Y13_F_masked1),
    .F_masked2(Tile_X5Y13_F_masked2),
    .UserCLK(Tile_X5Y14_UserCLKo),
    .UserCLKo(Tile_X5Y13_UserCLKo),
    .rst(Tile_X5Y14_rsto),
    .rsto(Tile_X5Y13_rsto),
    .FrameData(Tile_X4Y13_FrameData_O),
    .FrameData_O(Tile_X5Y13_FrameData_O),
    .FrameStrobe(Tile_X5Y14_FrameStrobe_O),
    .FrameStrobe_O(Tile_X5Y13_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
nonlinear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X6Y13_Emulate_Bitstream)
    )
`endif
    Tile_X6Y13_nonlinear_LMDPL
    (
    .from_NA(Tile_X6Y14_to_NA),
    .from_NB(Tile_X6Y14_to_NB),
    .from_NC(Tile_X6Y14_to_NC),
    .from_ND(Tile_X6Y14_to_ND),
    .from_NF(Tile_X6Y14_to_NF),
    .from_NG(Tile_X6Y14_to_NG),
    .from_NH(Tile_X6Y14_to_NH),
    .from_NI(Tile_X6Y14_to_NI),
    .from_EA(Tile_X5Y13_to_EA),
    .from_EB(Tile_X5Y13_to_EB),
    .from_EC(Tile_X5Y13_to_EC),
    .from_ED(Tile_X5Y13_to_ED),
    .from_EF(Tile_X5Y13_to_EF),
    .from_EG(Tile_X5Y13_to_EG),
    .from_EH(Tile_X5Y13_to_EH),
    .from_EI(Tile_X5Y13_to_EI),
    .from_SA(Tile_X6Y12_to_SA),
    .from_SB(Tile_X6Y12_to_SB),
    .from_SC(Tile_X6Y12_to_SC),
    .from_SD(Tile_X6Y12_to_SD),
    .from_SF(Tile_X6Y12_to_SF),
    .from_SG(Tile_X6Y12_to_SG),
    .from_SH(Tile_X6Y12_to_SH),
    .from_SI(Tile_X6Y12_to_SI),
    .from_WA(Tile_X7Y13_to_WA),
    .from_WB(Tile_X7Y13_to_WB),
    .from_WC(Tile_X7Y13_to_WC),
    .from_WD(Tile_X7Y13_to_WD),
    .from_WF(Tile_X7Y13_to_WF),
    .from_WG(Tile_X7Y13_to_WG),
    .from_WH(Tile_X7Y13_to_WH),
    .from_WI(Tile_X7Y13_to_WI),
    .to_EA(Tile_X6Y13_to_EA),
    .to_EB(Tile_X6Y13_to_EB),
    .to_EC(Tile_X6Y13_to_EC),
    .to_ED(Tile_X6Y13_to_ED),
    .to_EF(Tile_X6Y13_to_EF),
    .to_EG(Tile_X6Y13_to_EG),
    .to_EH(Tile_X6Y13_to_EH),
    .to_EI(Tile_X6Y13_to_EI),
    .to_WA(Tile_X6Y13_to_WA),
    .to_WB(Tile_X6Y13_to_WB),
    .to_WC(Tile_X6Y13_to_WC),
    .to_WD(Tile_X6Y13_to_WD),
    .to_WF(Tile_X6Y13_to_WF),
    .to_WG(Tile_X6Y13_to_WG),
    .to_WH(Tile_X6Y13_to_WH),
    .to_WI(Tile_X6Y13_to_WI),
    .to_NA(Tile_X6Y13_to_NA),
    .to_NB(Tile_X6Y13_to_NB),
    .to_NC(Tile_X6Y13_to_NC),
    .to_ND(Tile_X6Y13_to_ND),
    .to_NF(Tile_X6Y13_to_NF),
    .to_NG(Tile_X6Y13_to_NG),
    .to_NH(Tile_X6Y13_to_NH),
    .to_NI(Tile_X6Y13_to_NI),
    .to_SA(Tile_X6Y13_to_SA),
    .to_SB(Tile_X6Y13_to_SB),
    .to_SC(Tile_X6Y13_to_SC),
    .to_SD(Tile_X6Y13_to_SD),
    .to_SF(Tile_X6Y13_to_SF),
    .to_SG(Tile_X6Y13_to_SG),
    .to_SH(Tile_X6Y13_to_SH),
    .to_SI(Tile_X6Y13_to_SI),
    .R_t(Tile_X6Y13_R_t),
    .R_f(Tile_X6Y13_R_f),
    .F_masked1(Tile_X6Y13_F_masked1),
    .F_masked2(Tile_X6Y13_F_masked2),
    .UserCLK(Tile_X6Y14_UserCLKo),
    .UserCLKo(Tile_X6Y13_UserCLKo),
    .rst(Tile_X6Y14_rsto),
    .rsto(Tile_X6Y13_rsto),
    .FrameData(Tile_X5Y13_FrameData_O),
    .FrameData_O(Tile_X6Y13_FrameData_O),
    .FrameStrobe(Tile_X6Y14_FrameStrobe_O),
    .FrameStrobe_O(Tile_X6Y13_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X7Y13_Emulate_Bitstream)
    )
`endif
    Tile_X7Y13_linear_LMDPL
    (
    .from_NA(Tile_X7Y14_to_NA),
    .from_NB(Tile_X7Y14_to_NB),
    .from_NC(Tile_X7Y14_to_NC),
    .from_ND(Tile_X7Y14_to_ND),
    .from_NF(Tile_X7Y14_to_NF),
    .from_NG(Tile_X7Y14_to_NG),
    .from_NH(Tile_X7Y14_to_NH),
    .from_NI(Tile_X7Y14_to_NI),
    .from_EA(Tile_X6Y13_to_EA),
    .from_EB(Tile_X6Y13_to_EB),
    .from_EC(Tile_X6Y13_to_EC),
    .from_ED(Tile_X6Y13_to_ED),
    .from_EF(Tile_X6Y13_to_EF),
    .from_EG(Tile_X6Y13_to_EG),
    .from_EH(Tile_X6Y13_to_EH),
    .from_EI(Tile_X6Y13_to_EI),
    .from_SA(Tile_X7Y12_to_SA),
    .from_SB(Tile_X7Y12_to_SB),
    .from_SC(Tile_X7Y12_to_SC),
    .from_SD(Tile_X7Y12_to_SD),
    .from_SF(Tile_X7Y12_to_SF),
    .from_SG(Tile_X7Y12_to_SG),
    .from_SH(Tile_X7Y12_to_SH),
    .from_SI(Tile_X7Y12_to_SI),
    .from_WA(Tile_X8Y13_to_WA),
    .from_WB(Tile_X8Y13_to_WB),
    .from_WC(Tile_X8Y13_to_WC),
    .from_WD(Tile_X8Y13_to_WD),
    .from_WF(Tile_X8Y13_to_WF),
    .from_WG(Tile_X8Y13_to_WG),
    .from_WH(Tile_X8Y13_to_WH),
    .from_WI(Tile_X8Y13_to_WI),
    .to_EA(Tile_X7Y13_to_EA),
    .to_EB(Tile_X7Y13_to_EB),
    .to_EC(Tile_X7Y13_to_EC),
    .to_ED(Tile_X7Y13_to_ED),
    .to_EF(Tile_X7Y13_to_EF),
    .to_EG(Tile_X7Y13_to_EG),
    .to_EH(Tile_X7Y13_to_EH),
    .to_EI(Tile_X7Y13_to_EI),
    .to_WA(Tile_X7Y13_to_WA),
    .to_WB(Tile_X7Y13_to_WB),
    .to_WC(Tile_X7Y13_to_WC),
    .to_WD(Tile_X7Y13_to_WD),
    .to_WF(Tile_X7Y13_to_WF),
    .to_WG(Tile_X7Y13_to_WG),
    .to_WH(Tile_X7Y13_to_WH),
    .to_WI(Tile_X7Y13_to_WI),
    .to_NA(Tile_X7Y13_to_NA),
    .to_NB(Tile_X7Y13_to_NB),
    .to_NC(Tile_X7Y13_to_NC),
    .to_ND(Tile_X7Y13_to_ND),
    .to_NF(Tile_X7Y13_to_NF),
    .to_NG(Tile_X7Y13_to_NG),
    .to_NH(Tile_X7Y13_to_NH),
    .to_NI(Tile_X7Y13_to_NI),
    .to_SA(Tile_X7Y13_to_SA),
    .to_SB(Tile_X7Y13_to_SB),
    .to_SC(Tile_X7Y13_to_SC),
    .to_SD(Tile_X7Y13_to_SD),
    .to_SF(Tile_X7Y13_to_SF),
    .to_SG(Tile_X7Y13_to_SG),
    .to_SH(Tile_X7Y13_to_SH),
    .to_SI(Tile_X7Y13_to_SI),
    .F_masked1(Tile_X7Y13_F_masked1),
    .F_masked2(Tile_X7Y13_F_masked2),
    .UserCLK(Tile_X7Y14_UserCLKo),
    .UserCLKo(Tile_X7Y13_UserCLKo),
    .rst(Tile_X7Y14_rsto),
    .rsto(Tile_X7Y13_rsto),
    .FrameData(Tile_X6Y13_FrameData_O),
    .FrameData_O(Tile_X7Y13_FrameData_O),
    .FrameStrobe(Tile_X7Y14_FrameStrobe_O),
    .FrameStrobe_O(Tile_X7Y13_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
ctrl_to_sec
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X8Y13_Emulate_Bitstream)
    )
`endif
    Tile_X8Y13_ctrl_to_sec
    (
    .from_NA(Tile_X8Y14_to_NA),
    .from_NB(Tile_X8Y14_to_NB),
    .from_NC(Tile_X8Y14_to_NC),
    .from_ND(Tile_X8Y14_to_ND),
    .from_NF(Tile_X8Y14_to_NF),
    .from_NG(Tile_X8Y14_to_NG),
    .from_NH(Tile_X8Y14_to_NH),
    .from_NI(Tile_X8Y14_to_NI),
    .from_EA(Tile_X7Y13_to_EA),
    .from_EB(Tile_X7Y13_to_EB),
    .from_EC(Tile_X7Y13_to_EC),
    .from_ED(Tile_X7Y13_to_ED),
    .from_EF(Tile_X7Y13_to_EF),
    .from_EG(Tile_X7Y13_to_EG),
    .from_EH(Tile_X7Y13_to_EH),
    .from_EI(Tile_X7Y13_to_EI),
    .from_SA(Tile_X8Y12_to_SA),
    .from_SB(Tile_X8Y12_to_SB),
    .from_SC(Tile_X8Y12_to_SC),
    .from_SD(Tile_X8Y12_to_SD),
    .from_SF(Tile_X8Y12_to_SF),
    .from_SG(Tile_X8Y12_to_SG),
    .from_SH(Tile_X8Y12_to_SH),
    .from_SI(Tile_X8Y12_to_SI),
    .from_WA_1s(Tile_X9Y13_to_WA_1s),
    .from_WB_1s(Tile_X9Y13_to_WB_1s),
    .from_WC_1s(Tile_X9Y13_to_WC_1s),
    .from_WD_1s(Tile_X9Y13_to_WD_1s),
    .from_WF_1s(Tile_X9Y13_to_WF_1s),
    .from_WG_1s(Tile_X9Y13_to_WG_1s),
    .from_WH_1s(Tile_X9Y13_to_WH_1s),
    .from_WI_1s(Tile_X9Y13_to_WI_1s),
    .to_WA(Tile_X8Y13_to_WA),
    .to_WB(Tile_X8Y13_to_WB),
    .to_WC(Tile_X8Y13_to_WC),
    .to_WD(Tile_X8Y13_to_WD),
    .to_WF(Tile_X8Y13_to_WF),
    .to_WG(Tile_X8Y13_to_WG),
    .to_WH(Tile_X8Y13_to_WH),
    .to_WI(Tile_X8Y13_to_WI),
    .to_NA(Tile_X8Y13_to_NA),
    .to_NB(Tile_X8Y13_to_NB),
    .to_NC(Tile_X8Y13_to_NC),
    .to_ND(Tile_X8Y13_to_ND),
    .to_NF(Tile_X8Y13_to_NF),
    .to_NG(Tile_X8Y13_to_NG),
    .to_NH(Tile_X8Y13_to_NH),
    .to_NI(Tile_X8Y13_to_NI),
    .to_SA(Tile_X8Y13_to_SA),
    .to_SB(Tile_X8Y13_to_SB),
    .to_SC(Tile_X8Y13_to_SC),
    .to_SD(Tile_X8Y13_to_SD),
    .to_SF(Tile_X8Y13_to_SF),
    .to_SG(Tile_X8Y13_to_SG),
    .to_SH(Tile_X8Y13_to_SH),
    .to_SI(Tile_X8Y13_to_SI),
    .UserCLK(Tile_X8Y14_UserCLKo),
    .UserCLKo(Tile_X8Y13_UserCLKo),
    .rst(Tile_X8Y14_rsto),
    .rsto(Tile_X8Y13_rsto),
    .FrameData(Tile_X7Y13_FrameData_O),
    .FrameData_O(Tile_X8Y13_FrameData_O),
    .FrameStrobe(Tile_X8Y14_FrameStrobe_O),
    .FrameStrobe_O(Tile_X8Y13_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
combined_WDDL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X9Y13_Emulate_Bitstream)
    )
`endif
    Tile_X9Y13_combined_WDDL
    (
    .from_NA_1s(Tile_X9Y14_to_NA_1s),
    .from_NB_1s(Tile_X9Y14_to_NB_1s),
    .from_NC_1s(Tile_X9Y14_to_NC_1s),
    .from_ND_1s(Tile_X9Y14_to_ND_1s),
    .from_NF_1s(Tile_X9Y14_to_NF_1s),
    .from_NG_1s(Tile_X9Y14_to_NG_1s),
    .from_NH_1s(Tile_X9Y14_to_NH_1s),
    .from_NI_1s(Tile_X9Y14_to_NI_1s),
    .from_SA_1s(Tile_X9Y12_to_SA_1s),
    .from_SB_1s(Tile_X9Y12_to_SB_1s),
    .from_SC_1s(Tile_X9Y12_to_SC_1s),
    .from_SD_1s(Tile_X9Y12_to_SD_1s),
    .from_SF_1s(Tile_X9Y12_to_SF_1s),
    .from_SG_1s(Tile_X9Y12_to_SG_1s),
    .from_SH_1s(Tile_X9Y12_to_SH_1s),
    .from_SI_1s(Tile_X9Y12_to_SI_1s),
    .from_WA_1s(Tile_X10Y13_to_WA_1s),
    .from_WB_1s(Tile_X10Y13_to_WB_1s),
    .from_WC_1s(Tile_X10Y13_to_WC_1s),
    .from_WD_1s(Tile_X10Y13_to_WD_1s),
    .from_WF_1s(Tile_X10Y13_to_WF_1s),
    .from_WG_1s(Tile_X10Y13_to_WG_1s),
    .from_WH_1s(Tile_X10Y13_to_WH_1s),
    .from_WI_1s(Tile_X10Y13_to_WI_1s),
    .to_EA_1s(Tile_X9Y13_to_EA_1s),
    .to_EB_1s(Tile_X9Y13_to_EB_1s),
    .to_EC_1s(Tile_X9Y13_to_EC_1s),
    .to_ED_1s(Tile_X9Y13_to_ED_1s),
    .to_EF_1s(Tile_X9Y13_to_EF_1s),
    .to_EG_1s(Tile_X9Y13_to_EG_1s),
    .to_EH_1s(Tile_X9Y13_to_EH_1s),
    .to_EI_1s(Tile_X9Y13_to_EI_1s),
    .to_WA_1s(Tile_X9Y13_to_WA_1s),
    .to_WB_1s(Tile_X9Y13_to_WB_1s),
    .to_WC_1s(Tile_X9Y13_to_WC_1s),
    .to_WD_1s(Tile_X9Y13_to_WD_1s),
    .to_WF_1s(Tile_X9Y13_to_WF_1s),
    .to_WG_1s(Tile_X9Y13_to_WG_1s),
    .to_WH_1s(Tile_X9Y13_to_WH_1s),
    .to_WI_1s(Tile_X9Y13_to_WI_1s),
    .to_NA_1s(Tile_X9Y13_to_NA_1s),
    .to_NB_1s(Tile_X9Y13_to_NB_1s),
    .to_NC_1s(Tile_X9Y13_to_NC_1s),
    .to_ND_1s(Tile_X9Y13_to_ND_1s),
    .to_NF_1s(Tile_X9Y13_to_NF_1s),
    .to_NG_1s(Tile_X9Y13_to_NG_1s),
    .to_NH_1s(Tile_X9Y13_to_NH_1s),
    .to_NI_1s(Tile_X9Y13_to_NI_1s),
    .to_SA_1s(Tile_X9Y13_to_SA_1s),
    .to_SB_1s(Tile_X9Y13_to_SB_1s),
    .to_SC_1s(Tile_X9Y13_to_SC_1s),
    .to_SD_1s(Tile_X9Y13_to_SD_1s),
    .to_SF_1s(Tile_X9Y13_to_SF_1s),
    .to_SG_1s(Tile_X9Y13_to_SG_1s),
    .to_SH_1s(Tile_X9Y13_to_SH_1s),
    .to_SI_1s(Tile_X9Y13_to_SI_1s),
    .F_ctrl(Tile_X9Y13_F_ctrl),
    .UserCLK(Tile_X9Y14_UserCLKo),
    .UserCLKo(Tile_X9Y13_UserCLKo),
    .rst(Tile_X9Y14_rsto),
    .rsto(Tile_X9Y13_rsto),
    .FrameData(Tile_X8Y13_FrameData_O),
    .FrameData_O(Tile_X9Y13_FrameData_O),
    .FrameStrobe(Tile_X9Y14_FrameStrobe_O),
    .FrameStrobe_O(Tile_X9Y13_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
ctrl_IO
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X10Y13_Emulate_Bitstream)
    )
`endif
    Tile_X10Y13_ctrl_IO
    (
    .from_EA_1s(Tile_X9Y13_to_EA_1s),
    .from_EB_1s(Tile_X9Y13_to_EB_1s),
    .from_EC_1s(Tile_X9Y13_to_EC_1s),
    .from_ED_1s(Tile_X9Y13_to_ED_1s),
    .from_EF_1s(Tile_X9Y13_to_EF_1s),
    .from_EG_1s(Tile_X9Y13_to_EG_1s),
    .from_EH_1s(Tile_X9Y13_to_EH_1s),
    .from_EI_1s(Tile_X9Y13_to_EI_1s),
    .to_WA_1s(Tile_X10Y13_to_WA_1s),
    .to_WB_1s(Tile_X10Y13_to_WB_1s),
    .to_WC_1s(Tile_X10Y13_to_WC_1s),
    .to_WD_1s(Tile_X10Y13_to_WD_1s),
    .to_WF_1s(Tile_X10Y13_to_WF_1s),
    .to_WG_1s(Tile_X10Y13_to_WG_1s),
    .to_WH_1s(Tile_X10Y13_to_WH_1s),
    .to_WI_1s(Tile_X10Y13_to_WI_1s),
    .A_O_top_0_t(Tile_X10Y13_A_O_top_0_t),
    .A_O_top_0_f(Tile_X10Y13_A_O_top_0_f),
    .A_prech2(Tile_X10Y13_A_prech2),
    .A_DR_fault(Tile_X10Y13_A_DR_fault),
    .A_I_top_0_t(Tile_X10Y13_A_I_top_0_t),
    .A_I_top_0_f(Tile_X10Y13_A_I_top_0_f),
    .A_T_top(Tile_X10Y13_A_T_top),
    .A_F_ctrl(Tile_X10Y13_A_F_ctrl),
    .UserCLK(Tile_X10Y14_UserCLKo),
    .UserCLKo(Tile_X10Y13_UserCLKo),
    .rst(Tile_X10Y14_rsto),
    .rsto(Tile_X10Y13_rsto),
    .FrameData(Tile_X9Y13_FrameData_O),
    .FrameData_O(Tile_X10Y13_FrameData_O),
    .FrameStrobe(Tile_X10Y14_FrameStrobe_O),
    .FrameStrobe_O(Tile_X10Y13_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
W_IO_custom
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X0Y14_Emulate_Bitstream)
    )
`endif
    Tile_X0Y14_W_IO_custom
    (
    .from_NA(Tile_X0Y15_to_NA),
    .from_NB(Tile_X0Y15_to_NB),
    .from_NC(Tile_X0Y15_to_NC),
    .from_ND(Tile_X0Y15_to_ND),
    .from_NF(Tile_X0Y15_to_NF),
    .from_NG(Tile_X0Y15_to_NG),
    .from_NH(Tile_X0Y15_to_NH),
    .from_NI(Tile_X0Y15_to_NI),
    .from_SA(Tile_X0Y13_to_SA),
    .from_SB(Tile_X0Y13_to_SB),
    .from_SC(Tile_X0Y13_to_SC),
    .from_SD(Tile_X0Y13_to_SD),
    .from_SF(Tile_X0Y13_to_SF),
    .from_SG(Tile_X0Y13_to_SG),
    .from_SH(Tile_X0Y13_to_SH),
    .from_SI(Tile_X0Y13_to_SI),
    .from_WA(Tile_X1Y14_to_WA),
    .from_WB(Tile_X1Y14_to_WB),
    .from_WC(Tile_X1Y14_to_WC),
    .from_WD(Tile_X1Y14_to_WD),
    .from_WF(Tile_X1Y14_to_WF),
    .from_WG(Tile_X1Y14_to_WG),
    .from_WH(Tile_X1Y14_to_WH),
    .from_WI(Tile_X1Y14_to_WI),
    .to_EA(Tile_X0Y14_to_EA),
    .to_EB(Tile_X0Y14_to_EB),
    .to_EC(Tile_X0Y14_to_EC),
    .to_ED(Tile_X0Y14_to_ED),
    .to_EF(Tile_X0Y14_to_EF),
    .to_EG(Tile_X0Y14_to_EG),
    .to_EH(Tile_X0Y14_to_EH),
    .to_EI(Tile_X0Y14_to_EI),
    .to_NA(Tile_X0Y14_to_NA),
    .to_NB(Tile_X0Y14_to_NB),
    .to_NC(Tile_X0Y14_to_NC),
    .to_ND(Tile_X0Y14_to_ND),
    .to_NF(Tile_X0Y14_to_NF),
    .to_NG(Tile_X0Y14_to_NG),
    .to_NH(Tile_X0Y14_to_NH),
    .to_NI(Tile_X0Y14_to_NI),
    .to_SA(Tile_X0Y14_to_SA),
    .to_SB(Tile_X0Y14_to_SB),
    .to_SC(Tile_X0Y14_to_SC),
    .to_SD(Tile_X0Y14_to_SD),
    .to_SF(Tile_X0Y14_to_SF),
    .to_SG(Tile_X0Y14_to_SG),
    .to_SH(Tile_X0Y14_to_SH),
    .to_SI(Tile_X0Y14_to_SI),
    .A_O_top_0_t(Tile_X0Y14_A_O_top_0_t),
    .A_O_top_0_f(Tile_X0Y14_A_O_top_0_f),
    .A_O_top_1_t(Tile_X0Y14_A_O_top_1_t),
    .A_O_top_1_f(Tile_X0Y14_A_O_top_1_f),
    .A_prech1(Tile_X0Y14_A_prech1),
    .A_prech2(Tile_X0Y14_A_prech2),
    .A_DR_fault(Tile_X0Y14_A_DR_fault),
    .A_I_top_0_t(Tile_X0Y14_A_I_top_0_t),
    .A_I_top_0_f(Tile_X0Y14_A_I_top_0_f),
    .A_I_top_1_t(Tile_X0Y14_A_I_top_1_t),
    .A_I_top_1_f(Tile_X0Y14_A_I_top_1_f),
    .A_T_top(Tile_X0Y14_A_T_top),
    .A_F_masked1(Tile_X0Y14_A_F_masked1),
    .A_F_masked2(Tile_X0Y14_A_F_masked2),
    .A_config_C_bit0(Tile_X0Y14_A_config_C_bit0),
    .A_config_C_bit1(Tile_X0Y14_A_config_C_bit1),
    .A_config_C_bit2(Tile_X0Y14_A_config_C_bit2),
    .A_config_C_bit3(Tile_X0Y14_A_config_C_bit3),
    .B_config_C_bit0(Tile_X0Y14_B_config_C_bit0),
    .B_config_C_bit1(Tile_X0Y14_B_config_C_bit1),
    .B_config_C_bit2(Tile_X0Y14_B_config_C_bit2),
    .B_config_C_bit3(Tile_X0Y14_B_config_C_bit3),
    .UserCLK(Tile_X0Y15_UserCLKo),
    .UserCLKo(Tile_X0Y14_UserCLKo),
    .rst(Tile_X0Y15_rsto),
    .rsto(Tile_X0Y14_rsto),
    .FrameData(Tile_Y14_FrameData),
    .FrameData_O(Tile_X0Y14_FrameData_O),
    .FrameStrobe(Tile_X0Y15_FrameStrobe_O),
    .FrameStrobe_O(Tile_X0Y14_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X1Y14_Emulate_Bitstream)
    )
`endif
    Tile_X1Y14_linear_LMDPL
    (
    .from_NA(Tile_X1Y15_to_NA),
    .from_NB(Tile_X1Y15_to_NB),
    .from_NC(Tile_X1Y15_to_NC),
    .from_ND(Tile_X1Y15_to_ND),
    .from_NF(Tile_X1Y15_to_NF),
    .from_NG(Tile_X1Y15_to_NG),
    .from_NH(Tile_X1Y15_to_NH),
    .from_NI(Tile_X1Y15_to_NI),
    .from_EA(Tile_X0Y14_to_EA),
    .from_EB(Tile_X0Y14_to_EB),
    .from_EC(Tile_X0Y14_to_EC),
    .from_ED(Tile_X0Y14_to_ED),
    .from_EF(Tile_X0Y14_to_EF),
    .from_EG(Tile_X0Y14_to_EG),
    .from_EH(Tile_X0Y14_to_EH),
    .from_EI(Tile_X0Y14_to_EI),
    .from_SA(Tile_X1Y13_to_SA),
    .from_SB(Tile_X1Y13_to_SB),
    .from_SC(Tile_X1Y13_to_SC),
    .from_SD(Tile_X1Y13_to_SD),
    .from_SF(Tile_X1Y13_to_SF),
    .from_SG(Tile_X1Y13_to_SG),
    .from_SH(Tile_X1Y13_to_SH),
    .from_SI(Tile_X1Y13_to_SI),
    .from_WA(Tile_X2Y14_to_WA),
    .from_WB(Tile_X2Y14_to_WB),
    .from_WC(Tile_X2Y14_to_WC),
    .from_WD(Tile_X2Y14_to_WD),
    .from_WF(Tile_X2Y14_to_WF),
    .from_WG(Tile_X2Y14_to_WG),
    .from_WH(Tile_X2Y14_to_WH),
    .from_WI(Tile_X2Y14_to_WI),
    .to_EA(Tile_X1Y14_to_EA),
    .to_EB(Tile_X1Y14_to_EB),
    .to_EC(Tile_X1Y14_to_EC),
    .to_ED(Tile_X1Y14_to_ED),
    .to_EF(Tile_X1Y14_to_EF),
    .to_EG(Tile_X1Y14_to_EG),
    .to_EH(Tile_X1Y14_to_EH),
    .to_EI(Tile_X1Y14_to_EI),
    .to_WA(Tile_X1Y14_to_WA),
    .to_WB(Tile_X1Y14_to_WB),
    .to_WC(Tile_X1Y14_to_WC),
    .to_WD(Tile_X1Y14_to_WD),
    .to_WF(Tile_X1Y14_to_WF),
    .to_WG(Tile_X1Y14_to_WG),
    .to_WH(Tile_X1Y14_to_WH),
    .to_WI(Tile_X1Y14_to_WI),
    .to_NA(Tile_X1Y14_to_NA),
    .to_NB(Tile_X1Y14_to_NB),
    .to_NC(Tile_X1Y14_to_NC),
    .to_ND(Tile_X1Y14_to_ND),
    .to_NF(Tile_X1Y14_to_NF),
    .to_NG(Tile_X1Y14_to_NG),
    .to_NH(Tile_X1Y14_to_NH),
    .to_NI(Tile_X1Y14_to_NI),
    .to_SA(Tile_X1Y14_to_SA),
    .to_SB(Tile_X1Y14_to_SB),
    .to_SC(Tile_X1Y14_to_SC),
    .to_SD(Tile_X1Y14_to_SD),
    .to_SF(Tile_X1Y14_to_SF),
    .to_SG(Tile_X1Y14_to_SG),
    .to_SH(Tile_X1Y14_to_SH),
    .to_SI(Tile_X1Y14_to_SI),
    .F_masked1(Tile_X1Y14_F_masked1),
    .F_masked2(Tile_X1Y14_F_masked2),
    .UserCLK(Tile_X1Y15_UserCLKo),
    .UserCLKo(Tile_X1Y14_UserCLKo),
    .rst(Tile_X1Y15_rsto),
    .rsto(Tile_X1Y14_rsto),
    .FrameData(Tile_X0Y14_FrameData_O),
    .FrameData_O(Tile_X1Y14_FrameData_O),
    .FrameStrobe(Tile_X1Y15_FrameStrobe_O),
    .FrameStrobe_O(Tile_X1Y14_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X2Y14_Emulate_Bitstream)
    )
`endif
    Tile_X2Y14_linear_LMDPL
    (
    .from_NA(Tile_X2Y15_to_NA),
    .from_NB(Tile_X2Y15_to_NB),
    .from_NC(Tile_X2Y15_to_NC),
    .from_ND(Tile_X2Y15_to_ND),
    .from_NF(Tile_X2Y15_to_NF),
    .from_NG(Tile_X2Y15_to_NG),
    .from_NH(Tile_X2Y15_to_NH),
    .from_NI(Tile_X2Y15_to_NI),
    .from_EA(Tile_X1Y14_to_EA),
    .from_EB(Tile_X1Y14_to_EB),
    .from_EC(Tile_X1Y14_to_EC),
    .from_ED(Tile_X1Y14_to_ED),
    .from_EF(Tile_X1Y14_to_EF),
    .from_EG(Tile_X1Y14_to_EG),
    .from_EH(Tile_X1Y14_to_EH),
    .from_EI(Tile_X1Y14_to_EI),
    .from_SA(Tile_X2Y13_to_SA),
    .from_SB(Tile_X2Y13_to_SB),
    .from_SC(Tile_X2Y13_to_SC),
    .from_SD(Tile_X2Y13_to_SD),
    .from_SF(Tile_X2Y13_to_SF),
    .from_SG(Tile_X2Y13_to_SG),
    .from_SH(Tile_X2Y13_to_SH),
    .from_SI(Tile_X2Y13_to_SI),
    .from_WA(Tile_X3Y14_to_WA),
    .from_WB(Tile_X3Y14_to_WB),
    .from_WC(Tile_X3Y14_to_WC),
    .from_WD(Tile_X3Y14_to_WD),
    .from_WF(Tile_X3Y14_to_WF),
    .from_WG(Tile_X3Y14_to_WG),
    .from_WH(Tile_X3Y14_to_WH),
    .from_WI(Tile_X3Y14_to_WI),
    .to_EA(Tile_X2Y14_to_EA),
    .to_EB(Tile_X2Y14_to_EB),
    .to_EC(Tile_X2Y14_to_EC),
    .to_ED(Tile_X2Y14_to_ED),
    .to_EF(Tile_X2Y14_to_EF),
    .to_EG(Tile_X2Y14_to_EG),
    .to_EH(Tile_X2Y14_to_EH),
    .to_EI(Tile_X2Y14_to_EI),
    .to_WA(Tile_X2Y14_to_WA),
    .to_WB(Tile_X2Y14_to_WB),
    .to_WC(Tile_X2Y14_to_WC),
    .to_WD(Tile_X2Y14_to_WD),
    .to_WF(Tile_X2Y14_to_WF),
    .to_WG(Tile_X2Y14_to_WG),
    .to_WH(Tile_X2Y14_to_WH),
    .to_WI(Tile_X2Y14_to_WI),
    .to_NA(Tile_X2Y14_to_NA),
    .to_NB(Tile_X2Y14_to_NB),
    .to_NC(Tile_X2Y14_to_NC),
    .to_ND(Tile_X2Y14_to_ND),
    .to_NF(Tile_X2Y14_to_NF),
    .to_NG(Tile_X2Y14_to_NG),
    .to_NH(Tile_X2Y14_to_NH),
    .to_NI(Tile_X2Y14_to_NI),
    .to_SA(Tile_X2Y14_to_SA),
    .to_SB(Tile_X2Y14_to_SB),
    .to_SC(Tile_X2Y14_to_SC),
    .to_SD(Tile_X2Y14_to_SD),
    .to_SF(Tile_X2Y14_to_SF),
    .to_SG(Tile_X2Y14_to_SG),
    .to_SH(Tile_X2Y14_to_SH),
    .to_SI(Tile_X2Y14_to_SI),
    .F_masked1(Tile_X2Y14_F_masked1),
    .F_masked2(Tile_X2Y14_F_masked2),
    .UserCLK(Tile_X2Y15_UserCLKo),
    .UserCLKo(Tile_X2Y14_UserCLKo),
    .rst(Tile_X2Y15_rsto),
    .rsto(Tile_X2Y14_rsto),
    .FrameData(Tile_X1Y14_FrameData_O),
    .FrameData_O(Tile_X2Y14_FrameData_O),
    .FrameStrobe(Tile_X2Y15_FrameStrobe_O),
    .FrameStrobe_O(Tile_X2Y14_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
nonlinear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X3Y14_Emulate_Bitstream)
    )
`endif
    Tile_X3Y14_nonlinear_LMDPL
    (
    .from_NA(Tile_X3Y15_to_NA),
    .from_NB(Tile_X3Y15_to_NB),
    .from_NC(Tile_X3Y15_to_NC),
    .from_ND(Tile_X3Y15_to_ND),
    .from_NF(Tile_X3Y15_to_NF),
    .from_NG(Tile_X3Y15_to_NG),
    .from_NH(Tile_X3Y15_to_NH),
    .from_NI(Tile_X3Y15_to_NI),
    .from_EA(Tile_X2Y14_to_EA),
    .from_EB(Tile_X2Y14_to_EB),
    .from_EC(Tile_X2Y14_to_EC),
    .from_ED(Tile_X2Y14_to_ED),
    .from_EF(Tile_X2Y14_to_EF),
    .from_EG(Tile_X2Y14_to_EG),
    .from_EH(Tile_X2Y14_to_EH),
    .from_EI(Tile_X2Y14_to_EI),
    .from_SA(Tile_X3Y13_to_SA),
    .from_SB(Tile_X3Y13_to_SB),
    .from_SC(Tile_X3Y13_to_SC),
    .from_SD(Tile_X3Y13_to_SD),
    .from_SF(Tile_X3Y13_to_SF),
    .from_SG(Tile_X3Y13_to_SG),
    .from_SH(Tile_X3Y13_to_SH),
    .from_SI(Tile_X3Y13_to_SI),
    .from_WA(Tile_X4Y14_to_WA),
    .from_WB(Tile_X4Y14_to_WB),
    .from_WC(Tile_X4Y14_to_WC),
    .from_WD(Tile_X4Y14_to_WD),
    .from_WF(Tile_X4Y14_to_WF),
    .from_WG(Tile_X4Y14_to_WG),
    .from_WH(Tile_X4Y14_to_WH),
    .from_WI(Tile_X4Y14_to_WI),
    .to_EA(Tile_X3Y14_to_EA),
    .to_EB(Tile_X3Y14_to_EB),
    .to_EC(Tile_X3Y14_to_EC),
    .to_ED(Tile_X3Y14_to_ED),
    .to_EF(Tile_X3Y14_to_EF),
    .to_EG(Tile_X3Y14_to_EG),
    .to_EH(Tile_X3Y14_to_EH),
    .to_EI(Tile_X3Y14_to_EI),
    .to_WA(Tile_X3Y14_to_WA),
    .to_WB(Tile_X3Y14_to_WB),
    .to_WC(Tile_X3Y14_to_WC),
    .to_WD(Tile_X3Y14_to_WD),
    .to_WF(Tile_X3Y14_to_WF),
    .to_WG(Tile_X3Y14_to_WG),
    .to_WH(Tile_X3Y14_to_WH),
    .to_WI(Tile_X3Y14_to_WI),
    .to_NA(Tile_X3Y14_to_NA),
    .to_NB(Tile_X3Y14_to_NB),
    .to_NC(Tile_X3Y14_to_NC),
    .to_ND(Tile_X3Y14_to_ND),
    .to_NF(Tile_X3Y14_to_NF),
    .to_NG(Tile_X3Y14_to_NG),
    .to_NH(Tile_X3Y14_to_NH),
    .to_NI(Tile_X3Y14_to_NI),
    .to_SA(Tile_X3Y14_to_SA),
    .to_SB(Tile_X3Y14_to_SB),
    .to_SC(Tile_X3Y14_to_SC),
    .to_SD(Tile_X3Y14_to_SD),
    .to_SF(Tile_X3Y14_to_SF),
    .to_SG(Tile_X3Y14_to_SG),
    .to_SH(Tile_X3Y14_to_SH),
    .to_SI(Tile_X3Y14_to_SI),
    .R_t(Tile_X3Y14_R_t),
    .R_f(Tile_X3Y14_R_f),
    .F_masked1(Tile_X3Y14_F_masked1),
    .F_masked2(Tile_X3Y14_F_masked2),
    .UserCLK(Tile_X3Y15_UserCLKo),
    .UserCLKo(Tile_X3Y14_UserCLKo),
    .rst(Tile_X3Y15_rsto),
    .rsto(Tile_X3Y14_rsto),
    .FrameData(Tile_X2Y14_FrameData_O),
    .FrameData_O(Tile_X3Y14_FrameData_O),
    .FrameStrobe(Tile_X3Y15_FrameStrobe_O),
    .FrameStrobe_O(Tile_X3Y14_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X4Y14_Emulate_Bitstream)
    )
`endif
    Tile_X4Y14_linear_LMDPL
    (
    .from_NA(Tile_X4Y15_to_NA),
    .from_NB(Tile_X4Y15_to_NB),
    .from_NC(Tile_X4Y15_to_NC),
    .from_ND(Tile_X4Y15_to_ND),
    .from_NF(Tile_X4Y15_to_NF),
    .from_NG(Tile_X4Y15_to_NG),
    .from_NH(Tile_X4Y15_to_NH),
    .from_NI(Tile_X4Y15_to_NI),
    .from_EA(Tile_X3Y14_to_EA),
    .from_EB(Tile_X3Y14_to_EB),
    .from_EC(Tile_X3Y14_to_EC),
    .from_ED(Tile_X3Y14_to_ED),
    .from_EF(Tile_X3Y14_to_EF),
    .from_EG(Tile_X3Y14_to_EG),
    .from_EH(Tile_X3Y14_to_EH),
    .from_EI(Tile_X3Y14_to_EI),
    .from_SA(Tile_X4Y13_to_SA),
    .from_SB(Tile_X4Y13_to_SB),
    .from_SC(Tile_X4Y13_to_SC),
    .from_SD(Tile_X4Y13_to_SD),
    .from_SF(Tile_X4Y13_to_SF),
    .from_SG(Tile_X4Y13_to_SG),
    .from_SH(Tile_X4Y13_to_SH),
    .from_SI(Tile_X4Y13_to_SI),
    .from_WA(Tile_X5Y14_to_WA),
    .from_WB(Tile_X5Y14_to_WB),
    .from_WC(Tile_X5Y14_to_WC),
    .from_WD(Tile_X5Y14_to_WD),
    .from_WF(Tile_X5Y14_to_WF),
    .from_WG(Tile_X5Y14_to_WG),
    .from_WH(Tile_X5Y14_to_WH),
    .from_WI(Tile_X5Y14_to_WI),
    .to_EA(Tile_X4Y14_to_EA),
    .to_EB(Tile_X4Y14_to_EB),
    .to_EC(Tile_X4Y14_to_EC),
    .to_ED(Tile_X4Y14_to_ED),
    .to_EF(Tile_X4Y14_to_EF),
    .to_EG(Tile_X4Y14_to_EG),
    .to_EH(Tile_X4Y14_to_EH),
    .to_EI(Tile_X4Y14_to_EI),
    .to_WA(Tile_X4Y14_to_WA),
    .to_WB(Tile_X4Y14_to_WB),
    .to_WC(Tile_X4Y14_to_WC),
    .to_WD(Tile_X4Y14_to_WD),
    .to_WF(Tile_X4Y14_to_WF),
    .to_WG(Tile_X4Y14_to_WG),
    .to_WH(Tile_X4Y14_to_WH),
    .to_WI(Tile_X4Y14_to_WI),
    .to_NA(Tile_X4Y14_to_NA),
    .to_NB(Tile_X4Y14_to_NB),
    .to_NC(Tile_X4Y14_to_NC),
    .to_ND(Tile_X4Y14_to_ND),
    .to_NF(Tile_X4Y14_to_NF),
    .to_NG(Tile_X4Y14_to_NG),
    .to_NH(Tile_X4Y14_to_NH),
    .to_NI(Tile_X4Y14_to_NI),
    .to_SA(Tile_X4Y14_to_SA),
    .to_SB(Tile_X4Y14_to_SB),
    .to_SC(Tile_X4Y14_to_SC),
    .to_SD(Tile_X4Y14_to_SD),
    .to_SF(Tile_X4Y14_to_SF),
    .to_SG(Tile_X4Y14_to_SG),
    .to_SH(Tile_X4Y14_to_SH),
    .to_SI(Tile_X4Y14_to_SI),
    .F_masked1(Tile_X4Y14_F_masked1),
    .F_masked2(Tile_X4Y14_F_masked2),
    .UserCLK(Tile_X4Y15_UserCLKo),
    .UserCLKo(Tile_X4Y14_UserCLKo),
    .rst(Tile_X4Y15_rsto),
    .rsto(Tile_X4Y14_rsto),
    .FrameData(Tile_X3Y14_FrameData_O),
    .FrameData_O(Tile_X4Y14_FrameData_O),
    .FrameStrobe(Tile_X4Y15_FrameStrobe_O),
    .FrameStrobe_O(Tile_X4Y14_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X5Y14_Emulate_Bitstream)
    )
`endif
    Tile_X5Y14_linear_LMDPL
    (
    .from_NA(Tile_X5Y15_to_NA),
    .from_NB(Tile_X5Y15_to_NB),
    .from_NC(Tile_X5Y15_to_NC),
    .from_ND(Tile_X5Y15_to_ND),
    .from_NF(Tile_X5Y15_to_NF),
    .from_NG(Tile_X5Y15_to_NG),
    .from_NH(Tile_X5Y15_to_NH),
    .from_NI(Tile_X5Y15_to_NI),
    .from_EA(Tile_X4Y14_to_EA),
    .from_EB(Tile_X4Y14_to_EB),
    .from_EC(Tile_X4Y14_to_EC),
    .from_ED(Tile_X4Y14_to_ED),
    .from_EF(Tile_X4Y14_to_EF),
    .from_EG(Tile_X4Y14_to_EG),
    .from_EH(Tile_X4Y14_to_EH),
    .from_EI(Tile_X4Y14_to_EI),
    .from_SA(Tile_X5Y13_to_SA),
    .from_SB(Tile_X5Y13_to_SB),
    .from_SC(Tile_X5Y13_to_SC),
    .from_SD(Tile_X5Y13_to_SD),
    .from_SF(Tile_X5Y13_to_SF),
    .from_SG(Tile_X5Y13_to_SG),
    .from_SH(Tile_X5Y13_to_SH),
    .from_SI(Tile_X5Y13_to_SI),
    .from_WA(Tile_X6Y14_to_WA),
    .from_WB(Tile_X6Y14_to_WB),
    .from_WC(Tile_X6Y14_to_WC),
    .from_WD(Tile_X6Y14_to_WD),
    .from_WF(Tile_X6Y14_to_WF),
    .from_WG(Tile_X6Y14_to_WG),
    .from_WH(Tile_X6Y14_to_WH),
    .from_WI(Tile_X6Y14_to_WI),
    .to_EA(Tile_X5Y14_to_EA),
    .to_EB(Tile_X5Y14_to_EB),
    .to_EC(Tile_X5Y14_to_EC),
    .to_ED(Tile_X5Y14_to_ED),
    .to_EF(Tile_X5Y14_to_EF),
    .to_EG(Tile_X5Y14_to_EG),
    .to_EH(Tile_X5Y14_to_EH),
    .to_EI(Tile_X5Y14_to_EI),
    .to_WA(Tile_X5Y14_to_WA),
    .to_WB(Tile_X5Y14_to_WB),
    .to_WC(Tile_X5Y14_to_WC),
    .to_WD(Tile_X5Y14_to_WD),
    .to_WF(Tile_X5Y14_to_WF),
    .to_WG(Tile_X5Y14_to_WG),
    .to_WH(Tile_X5Y14_to_WH),
    .to_WI(Tile_X5Y14_to_WI),
    .to_NA(Tile_X5Y14_to_NA),
    .to_NB(Tile_X5Y14_to_NB),
    .to_NC(Tile_X5Y14_to_NC),
    .to_ND(Tile_X5Y14_to_ND),
    .to_NF(Tile_X5Y14_to_NF),
    .to_NG(Tile_X5Y14_to_NG),
    .to_NH(Tile_X5Y14_to_NH),
    .to_NI(Tile_X5Y14_to_NI),
    .to_SA(Tile_X5Y14_to_SA),
    .to_SB(Tile_X5Y14_to_SB),
    .to_SC(Tile_X5Y14_to_SC),
    .to_SD(Tile_X5Y14_to_SD),
    .to_SF(Tile_X5Y14_to_SF),
    .to_SG(Tile_X5Y14_to_SG),
    .to_SH(Tile_X5Y14_to_SH),
    .to_SI(Tile_X5Y14_to_SI),
    .F_masked1(Tile_X5Y14_F_masked1),
    .F_masked2(Tile_X5Y14_F_masked2),
    .UserCLK(Tile_X5Y15_UserCLKo),
    .UserCLKo(Tile_X5Y14_UserCLKo),
    .rst(Tile_X5Y15_rsto),
    .rsto(Tile_X5Y14_rsto),
    .FrameData(Tile_X4Y14_FrameData_O),
    .FrameData_O(Tile_X5Y14_FrameData_O),
    .FrameStrobe(Tile_X5Y15_FrameStrobe_O),
    .FrameStrobe_O(Tile_X5Y14_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
nonlinear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X6Y14_Emulate_Bitstream)
    )
`endif
    Tile_X6Y14_nonlinear_LMDPL
    (
    .from_NA(Tile_X6Y15_to_NA),
    .from_NB(Tile_X6Y15_to_NB),
    .from_NC(Tile_X6Y15_to_NC),
    .from_ND(Tile_X6Y15_to_ND),
    .from_NF(Tile_X6Y15_to_NF),
    .from_NG(Tile_X6Y15_to_NG),
    .from_NH(Tile_X6Y15_to_NH),
    .from_NI(Tile_X6Y15_to_NI),
    .from_EA(Tile_X5Y14_to_EA),
    .from_EB(Tile_X5Y14_to_EB),
    .from_EC(Tile_X5Y14_to_EC),
    .from_ED(Tile_X5Y14_to_ED),
    .from_EF(Tile_X5Y14_to_EF),
    .from_EG(Tile_X5Y14_to_EG),
    .from_EH(Tile_X5Y14_to_EH),
    .from_EI(Tile_X5Y14_to_EI),
    .from_SA(Tile_X6Y13_to_SA),
    .from_SB(Tile_X6Y13_to_SB),
    .from_SC(Tile_X6Y13_to_SC),
    .from_SD(Tile_X6Y13_to_SD),
    .from_SF(Tile_X6Y13_to_SF),
    .from_SG(Tile_X6Y13_to_SG),
    .from_SH(Tile_X6Y13_to_SH),
    .from_SI(Tile_X6Y13_to_SI),
    .from_WA(Tile_X7Y14_to_WA),
    .from_WB(Tile_X7Y14_to_WB),
    .from_WC(Tile_X7Y14_to_WC),
    .from_WD(Tile_X7Y14_to_WD),
    .from_WF(Tile_X7Y14_to_WF),
    .from_WG(Tile_X7Y14_to_WG),
    .from_WH(Tile_X7Y14_to_WH),
    .from_WI(Tile_X7Y14_to_WI),
    .to_EA(Tile_X6Y14_to_EA),
    .to_EB(Tile_X6Y14_to_EB),
    .to_EC(Tile_X6Y14_to_EC),
    .to_ED(Tile_X6Y14_to_ED),
    .to_EF(Tile_X6Y14_to_EF),
    .to_EG(Tile_X6Y14_to_EG),
    .to_EH(Tile_X6Y14_to_EH),
    .to_EI(Tile_X6Y14_to_EI),
    .to_WA(Tile_X6Y14_to_WA),
    .to_WB(Tile_X6Y14_to_WB),
    .to_WC(Tile_X6Y14_to_WC),
    .to_WD(Tile_X6Y14_to_WD),
    .to_WF(Tile_X6Y14_to_WF),
    .to_WG(Tile_X6Y14_to_WG),
    .to_WH(Tile_X6Y14_to_WH),
    .to_WI(Tile_X6Y14_to_WI),
    .to_NA(Tile_X6Y14_to_NA),
    .to_NB(Tile_X6Y14_to_NB),
    .to_NC(Tile_X6Y14_to_NC),
    .to_ND(Tile_X6Y14_to_ND),
    .to_NF(Tile_X6Y14_to_NF),
    .to_NG(Tile_X6Y14_to_NG),
    .to_NH(Tile_X6Y14_to_NH),
    .to_NI(Tile_X6Y14_to_NI),
    .to_SA(Tile_X6Y14_to_SA),
    .to_SB(Tile_X6Y14_to_SB),
    .to_SC(Tile_X6Y14_to_SC),
    .to_SD(Tile_X6Y14_to_SD),
    .to_SF(Tile_X6Y14_to_SF),
    .to_SG(Tile_X6Y14_to_SG),
    .to_SH(Tile_X6Y14_to_SH),
    .to_SI(Tile_X6Y14_to_SI),
    .R_t(Tile_X6Y14_R_t),
    .R_f(Tile_X6Y14_R_f),
    .F_masked1(Tile_X6Y14_F_masked1),
    .F_masked2(Tile_X6Y14_F_masked2),
    .UserCLK(Tile_X6Y15_UserCLKo),
    .UserCLKo(Tile_X6Y14_UserCLKo),
    .rst(Tile_X6Y15_rsto),
    .rsto(Tile_X6Y14_rsto),
    .FrameData(Tile_X5Y14_FrameData_O),
    .FrameData_O(Tile_X6Y14_FrameData_O),
    .FrameStrobe(Tile_X6Y15_FrameStrobe_O),
    .FrameStrobe_O(Tile_X6Y14_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X7Y14_Emulate_Bitstream)
    )
`endif
    Tile_X7Y14_linear_LMDPL
    (
    .from_NA(Tile_X7Y15_to_NA),
    .from_NB(Tile_X7Y15_to_NB),
    .from_NC(Tile_X7Y15_to_NC),
    .from_ND(Tile_X7Y15_to_ND),
    .from_NF(Tile_X7Y15_to_NF),
    .from_NG(Tile_X7Y15_to_NG),
    .from_NH(Tile_X7Y15_to_NH),
    .from_NI(Tile_X7Y15_to_NI),
    .from_EA(Tile_X6Y14_to_EA),
    .from_EB(Tile_X6Y14_to_EB),
    .from_EC(Tile_X6Y14_to_EC),
    .from_ED(Tile_X6Y14_to_ED),
    .from_EF(Tile_X6Y14_to_EF),
    .from_EG(Tile_X6Y14_to_EG),
    .from_EH(Tile_X6Y14_to_EH),
    .from_EI(Tile_X6Y14_to_EI),
    .from_SA(Tile_X7Y13_to_SA),
    .from_SB(Tile_X7Y13_to_SB),
    .from_SC(Tile_X7Y13_to_SC),
    .from_SD(Tile_X7Y13_to_SD),
    .from_SF(Tile_X7Y13_to_SF),
    .from_SG(Tile_X7Y13_to_SG),
    .from_SH(Tile_X7Y13_to_SH),
    .from_SI(Tile_X7Y13_to_SI),
    .from_WA(Tile_X8Y14_to_WA),
    .from_WB(Tile_X8Y14_to_WB),
    .from_WC(Tile_X8Y14_to_WC),
    .from_WD(Tile_X8Y14_to_WD),
    .from_WF(Tile_X8Y14_to_WF),
    .from_WG(Tile_X8Y14_to_WG),
    .from_WH(Tile_X8Y14_to_WH),
    .from_WI(Tile_X8Y14_to_WI),
    .to_EA(Tile_X7Y14_to_EA),
    .to_EB(Tile_X7Y14_to_EB),
    .to_EC(Tile_X7Y14_to_EC),
    .to_ED(Tile_X7Y14_to_ED),
    .to_EF(Tile_X7Y14_to_EF),
    .to_EG(Tile_X7Y14_to_EG),
    .to_EH(Tile_X7Y14_to_EH),
    .to_EI(Tile_X7Y14_to_EI),
    .to_WA(Tile_X7Y14_to_WA),
    .to_WB(Tile_X7Y14_to_WB),
    .to_WC(Tile_X7Y14_to_WC),
    .to_WD(Tile_X7Y14_to_WD),
    .to_WF(Tile_X7Y14_to_WF),
    .to_WG(Tile_X7Y14_to_WG),
    .to_WH(Tile_X7Y14_to_WH),
    .to_WI(Tile_X7Y14_to_WI),
    .to_NA(Tile_X7Y14_to_NA),
    .to_NB(Tile_X7Y14_to_NB),
    .to_NC(Tile_X7Y14_to_NC),
    .to_ND(Tile_X7Y14_to_ND),
    .to_NF(Tile_X7Y14_to_NF),
    .to_NG(Tile_X7Y14_to_NG),
    .to_NH(Tile_X7Y14_to_NH),
    .to_NI(Tile_X7Y14_to_NI),
    .to_SA(Tile_X7Y14_to_SA),
    .to_SB(Tile_X7Y14_to_SB),
    .to_SC(Tile_X7Y14_to_SC),
    .to_SD(Tile_X7Y14_to_SD),
    .to_SF(Tile_X7Y14_to_SF),
    .to_SG(Tile_X7Y14_to_SG),
    .to_SH(Tile_X7Y14_to_SH),
    .to_SI(Tile_X7Y14_to_SI),
    .F_masked1(Tile_X7Y14_F_masked1),
    .F_masked2(Tile_X7Y14_F_masked2),
    .UserCLK(Tile_X7Y15_UserCLKo),
    .UserCLKo(Tile_X7Y14_UserCLKo),
    .rst(Tile_X7Y15_rsto),
    .rsto(Tile_X7Y14_rsto),
    .FrameData(Tile_X6Y14_FrameData_O),
    .FrameData_O(Tile_X7Y14_FrameData_O),
    .FrameStrobe(Tile_X7Y15_FrameStrobe_O),
    .FrameStrobe_O(Tile_X7Y14_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
ctrl_to_sec
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X8Y14_Emulate_Bitstream)
    )
`endif
    Tile_X8Y14_ctrl_to_sec
    (
    .from_NA(Tile_X8Y15_to_NA),
    .from_NB(Tile_X8Y15_to_NB),
    .from_NC(Tile_X8Y15_to_NC),
    .from_ND(Tile_X8Y15_to_ND),
    .from_NF(Tile_X8Y15_to_NF),
    .from_NG(Tile_X8Y15_to_NG),
    .from_NH(Tile_X8Y15_to_NH),
    .from_NI(Tile_X8Y15_to_NI),
    .from_EA(Tile_X7Y14_to_EA),
    .from_EB(Tile_X7Y14_to_EB),
    .from_EC(Tile_X7Y14_to_EC),
    .from_ED(Tile_X7Y14_to_ED),
    .from_EF(Tile_X7Y14_to_EF),
    .from_EG(Tile_X7Y14_to_EG),
    .from_EH(Tile_X7Y14_to_EH),
    .from_EI(Tile_X7Y14_to_EI),
    .from_SA(Tile_X8Y13_to_SA),
    .from_SB(Tile_X8Y13_to_SB),
    .from_SC(Tile_X8Y13_to_SC),
    .from_SD(Tile_X8Y13_to_SD),
    .from_SF(Tile_X8Y13_to_SF),
    .from_SG(Tile_X8Y13_to_SG),
    .from_SH(Tile_X8Y13_to_SH),
    .from_SI(Tile_X8Y13_to_SI),
    .from_WA_1s(Tile_X9Y14_to_WA_1s),
    .from_WB_1s(Tile_X9Y14_to_WB_1s),
    .from_WC_1s(Tile_X9Y14_to_WC_1s),
    .from_WD_1s(Tile_X9Y14_to_WD_1s),
    .from_WF_1s(Tile_X9Y14_to_WF_1s),
    .from_WG_1s(Tile_X9Y14_to_WG_1s),
    .from_WH_1s(Tile_X9Y14_to_WH_1s),
    .from_WI_1s(Tile_X9Y14_to_WI_1s),
    .to_WA(Tile_X8Y14_to_WA),
    .to_WB(Tile_X8Y14_to_WB),
    .to_WC(Tile_X8Y14_to_WC),
    .to_WD(Tile_X8Y14_to_WD),
    .to_WF(Tile_X8Y14_to_WF),
    .to_WG(Tile_X8Y14_to_WG),
    .to_WH(Tile_X8Y14_to_WH),
    .to_WI(Tile_X8Y14_to_WI),
    .to_NA(Tile_X8Y14_to_NA),
    .to_NB(Tile_X8Y14_to_NB),
    .to_NC(Tile_X8Y14_to_NC),
    .to_ND(Tile_X8Y14_to_ND),
    .to_NF(Tile_X8Y14_to_NF),
    .to_NG(Tile_X8Y14_to_NG),
    .to_NH(Tile_X8Y14_to_NH),
    .to_NI(Tile_X8Y14_to_NI),
    .to_SA(Tile_X8Y14_to_SA),
    .to_SB(Tile_X8Y14_to_SB),
    .to_SC(Tile_X8Y14_to_SC),
    .to_SD(Tile_X8Y14_to_SD),
    .to_SF(Tile_X8Y14_to_SF),
    .to_SG(Tile_X8Y14_to_SG),
    .to_SH(Tile_X8Y14_to_SH),
    .to_SI(Tile_X8Y14_to_SI),
    .UserCLK(Tile_X8Y15_UserCLKo),
    .UserCLKo(Tile_X8Y14_UserCLKo),
    .rst(Tile_X8Y15_rsto),
    .rsto(Tile_X8Y14_rsto),
    .FrameData(Tile_X7Y14_FrameData_O),
    .FrameData_O(Tile_X8Y14_FrameData_O),
    .FrameStrobe(Tile_X8Y15_FrameStrobe_O),
    .FrameStrobe_O(Tile_X8Y14_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
combined_WDDL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X9Y14_Emulate_Bitstream)
    )
`endif
    Tile_X9Y14_combined_WDDL
    (
    .from_NA_1s(Tile_X9Y15_to_NA_1s),
    .from_NB_1s(Tile_X9Y15_to_NB_1s),
    .from_NC_1s(Tile_X9Y15_to_NC_1s),
    .from_ND_1s(Tile_X9Y15_to_ND_1s),
    .from_NF_1s(Tile_X9Y15_to_NF_1s),
    .from_NG_1s(Tile_X9Y15_to_NG_1s),
    .from_NH_1s(Tile_X9Y15_to_NH_1s),
    .from_NI_1s(Tile_X9Y15_to_NI_1s),
    .from_SA_1s(Tile_X9Y13_to_SA_1s),
    .from_SB_1s(Tile_X9Y13_to_SB_1s),
    .from_SC_1s(Tile_X9Y13_to_SC_1s),
    .from_SD_1s(Tile_X9Y13_to_SD_1s),
    .from_SF_1s(Tile_X9Y13_to_SF_1s),
    .from_SG_1s(Tile_X9Y13_to_SG_1s),
    .from_SH_1s(Tile_X9Y13_to_SH_1s),
    .from_SI_1s(Tile_X9Y13_to_SI_1s),
    .from_WA_1s(Tile_X10Y14_to_WA_1s),
    .from_WB_1s(Tile_X10Y14_to_WB_1s),
    .from_WC_1s(Tile_X10Y14_to_WC_1s),
    .from_WD_1s(Tile_X10Y14_to_WD_1s),
    .from_WF_1s(Tile_X10Y14_to_WF_1s),
    .from_WG_1s(Tile_X10Y14_to_WG_1s),
    .from_WH_1s(Tile_X10Y14_to_WH_1s),
    .from_WI_1s(Tile_X10Y14_to_WI_1s),
    .to_EA_1s(Tile_X9Y14_to_EA_1s),
    .to_EB_1s(Tile_X9Y14_to_EB_1s),
    .to_EC_1s(Tile_X9Y14_to_EC_1s),
    .to_ED_1s(Tile_X9Y14_to_ED_1s),
    .to_EF_1s(Tile_X9Y14_to_EF_1s),
    .to_EG_1s(Tile_X9Y14_to_EG_1s),
    .to_EH_1s(Tile_X9Y14_to_EH_1s),
    .to_EI_1s(Tile_X9Y14_to_EI_1s),
    .to_WA_1s(Tile_X9Y14_to_WA_1s),
    .to_WB_1s(Tile_X9Y14_to_WB_1s),
    .to_WC_1s(Tile_X9Y14_to_WC_1s),
    .to_WD_1s(Tile_X9Y14_to_WD_1s),
    .to_WF_1s(Tile_X9Y14_to_WF_1s),
    .to_WG_1s(Tile_X9Y14_to_WG_1s),
    .to_WH_1s(Tile_X9Y14_to_WH_1s),
    .to_WI_1s(Tile_X9Y14_to_WI_1s),
    .to_NA_1s(Tile_X9Y14_to_NA_1s),
    .to_NB_1s(Tile_X9Y14_to_NB_1s),
    .to_NC_1s(Tile_X9Y14_to_NC_1s),
    .to_ND_1s(Tile_X9Y14_to_ND_1s),
    .to_NF_1s(Tile_X9Y14_to_NF_1s),
    .to_NG_1s(Tile_X9Y14_to_NG_1s),
    .to_NH_1s(Tile_X9Y14_to_NH_1s),
    .to_NI_1s(Tile_X9Y14_to_NI_1s),
    .to_SA_1s(Tile_X9Y14_to_SA_1s),
    .to_SB_1s(Tile_X9Y14_to_SB_1s),
    .to_SC_1s(Tile_X9Y14_to_SC_1s),
    .to_SD_1s(Tile_X9Y14_to_SD_1s),
    .to_SF_1s(Tile_X9Y14_to_SF_1s),
    .to_SG_1s(Tile_X9Y14_to_SG_1s),
    .to_SH_1s(Tile_X9Y14_to_SH_1s),
    .to_SI_1s(Tile_X9Y14_to_SI_1s),
    .F_ctrl(Tile_X9Y14_F_ctrl),
    .UserCLK(Tile_X9Y15_UserCLKo),
    .UserCLKo(Tile_X9Y14_UserCLKo),
    .rst(Tile_X9Y15_rsto),
    .rsto(Tile_X9Y14_rsto),
    .FrameData(Tile_X8Y14_FrameData_O),
    .FrameData_O(Tile_X9Y14_FrameData_O),
    .FrameStrobe(Tile_X9Y15_FrameStrobe_O),
    .FrameStrobe_O(Tile_X9Y14_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
ctrl_IO
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X10Y14_Emulate_Bitstream)
    )
`endif
    Tile_X10Y14_ctrl_IO
    (
    .from_EA_1s(Tile_X9Y14_to_EA_1s),
    .from_EB_1s(Tile_X9Y14_to_EB_1s),
    .from_EC_1s(Tile_X9Y14_to_EC_1s),
    .from_ED_1s(Tile_X9Y14_to_ED_1s),
    .from_EF_1s(Tile_X9Y14_to_EF_1s),
    .from_EG_1s(Tile_X9Y14_to_EG_1s),
    .from_EH_1s(Tile_X9Y14_to_EH_1s),
    .from_EI_1s(Tile_X9Y14_to_EI_1s),
    .to_WA_1s(Tile_X10Y14_to_WA_1s),
    .to_WB_1s(Tile_X10Y14_to_WB_1s),
    .to_WC_1s(Tile_X10Y14_to_WC_1s),
    .to_WD_1s(Tile_X10Y14_to_WD_1s),
    .to_WF_1s(Tile_X10Y14_to_WF_1s),
    .to_WG_1s(Tile_X10Y14_to_WG_1s),
    .to_WH_1s(Tile_X10Y14_to_WH_1s),
    .to_WI_1s(Tile_X10Y14_to_WI_1s),
    .A_O_top_0_t(Tile_X10Y14_A_O_top_0_t),
    .A_O_top_0_f(Tile_X10Y14_A_O_top_0_f),
    .A_prech2(Tile_X10Y14_A_prech2),
    .A_DR_fault(Tile_X10Y14_A_DR_fault),
    .A_I_top_0_t(Tile_X10Y14_A_I_top_0_t),
    .A_I_top_0_f(Tile_X10Y14_A_I_top_0_f),
    .A_T_top(Tile_X10Y14_A_T_top),
    .A_F_ctrl(Tile_X10Y14_A_F_ctrl),
    .UserCLK(Tile_X10Y15_UserCLKo),
    .UserCLKo(Tile_X10Y14_UserCLKo),
    .rst(Tile_X10Y15_rsto),
    .rsto(Tile_X10Y14_rsto),
    .FrameData(Tile_X9Y14_FrameData_O),
    .FrameData_O(Tile_X10Y14_FrameData_O),
    .FrameStrobe(Tile_X10Y15_FrameStrobe_O),
    .FrameStrobe_O(Tile_X10Y14_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
W_IO_custom
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X0Y15_Emulate_Bitstream)
    )
`endif
    Tile_X0Y15_W_IO_custom
    (
    .from_NA(Tile_X0Y16_to_NA),
    .from_NB(Tile_X0Y16_to_NB),
    .from_NC(Tile_X0Y16_to_NC),
    .from_ND(Tile_X0Y16_to_ND),
    .from_NF(Tile_X0Y16_to_NF),
    .from_NG(Tile_X0Y16_to_NG),
    .from_NH(Tile_X0Y16_to_NH),
    .from_NI(Tile_X0Y16_to_NI),
    .from_SA(Tile_X0Y14_to_SA),
    .from_SB(Tile_X0Y14_to_SB),
    .from_SC(Tile_X0Y14_to_SC),
    .from_SD(Tile_X0Y14_to_SD),
    .from_SF(Tile_X0Y14_to_SF),
    .from_SG(Tile_X0Y14_to_SG),
    .from_SH(Tile_X0Y14_to_SH),
    .from_SI(Tile_X0Y14_to_SI),
    .from_WA(Tile_X1Y15_to_WA),
    .from_WB(Tile_X1Y15_to_WB),
    .from_WC(Tile_X1Y15_to_WC),
    .from_WD(Tile_X1Y15_to_WD),
    .from_WF(Tile_X1Y15_to_WF),
    .from_WG(Tile_X1Y15_to_WG),
    .from_WH(Tile_X1Y15_to_WH),
    .from_WI(Tile_X1Y15_to_WI),
    .to_EA(Tile_X0Y15_to_EA),
    .to_EB(Tile_X0Y15_to_EB),
    .to_EC(Tile_X0Y15_to_EC),
    .to_ED(Tile_X0Y15_to_ED),
    .to_EF(Tile_X0Y15_to_EF),
    .to_EG(Tile_X0Y15_to_EG),
    .to_EH(Tile_X0Y15_to_EH),
    .to_EI(Tile_X0Y15_to_EI),
    .to_NA(Tile_X0Y15_to_NA),
    .to_NB(Tile_X0Y15_to_NB),
    .to_NC(Tile_X0Y15_to_NC),
    .to_ND(Tile_X0Y15_to_ND),
    .to_NF(Tile_X0Y15_to_NF),
    .to_NG(Tile_X0Y15_to_NG),
    .to_NH(Tile_X0Y15_to_NH),
    .to_NI(Tile_X0Y15_to_NI),
    .to_SA(Tile_X0Y15_to_SA),
    .to_SB(Tile_X0Y15_to_SB),
    .to_SC(Tile_X0Y15_to_SC),
    .to_SD(Tile_X0Y15_to_SD),
    .to_SF(Tile_X0Y15_to_SF),
    .to_SG(Tile_X0Y15_to_SG),
    .to_SH(Tile_X0Y15_to_SH),
    .to_SI(Tile_X0Y15_to_SI),
    .A_O_top_0_t(Tile_X0Y15_A_O_top_0_t),
    .A_O_top_0_f(Tile_X0Y15_A_O_top_0_f),
    .A_O_top_1_t(Tile_X0Y15_A_O_top_1_t),
    .A_O_top_1_f(Tile_X0Y15_A_O_top_1_f),
    .A_prech1(Tile_X0Y15_A_prech1),
    .A_prech2(Tile_X0Y15_A_prech2),
    .A_DR_fault(Tile_X0Y15_A_DR_fault),
    .A_I_top_0_t(Tile_X0Y15_A_I_top_0_t),
    .A_I_top_0_f(Tile_X0Y15_A_I_top_0_f),
    .A_I_top_1_t(Tile_X0Y15_A_I_top_1_t),
    .A_I_top_1_f(Tile_X0Y15_A_I_top_1_f),
    .A_T_top(Tile_X0Y15_A_T_top),
    .A_F_masked1(Tile_X0Y15_A_F_masked1),
    .A_F_masked2(Tile_X0Y15_A_F_masked2),
    .A_config_C_bit0(Tile_X0Y15_A_config_C_bit0),
    .A_config_C_bit1(Tile_X0Y15_A_config_C_bit1),
    .A_config_C_bit2(Tile_X0Y15_A_config_C_bit2),
    .A_config_C_bit3(Tile_X0Y15_A_config_C_bit3),
    .B_config_C_bit0(Tile_X0Y15_B_config_C_bit0),
    .B_config_C_bit1(Tile_X0Y15_B_config_C_bit1),
    .B_config_C_bit2(Tile_X0Y15_B_config_C_bit2),
    .B_config_C_bit3(Tile_X0Y15_B_config_C_bit3),
    .UserCLK(Tile_X0Y16_UserCLKo),
    .UserCLKo(Tile_X0Y15_UserCLKo),
    .rst(Tile_X0Y16_rsto),
    .rsto(Tile_X0Y15_rsto),
    .FrameData(Tile_Y15_FrameData),
    .FrameData_O(Tile_X0Y15_FrameData_O),
    .FrameStrobe(Tile_X0Y16_FrameStrobe_O),
    .FrameStrobe_O(Tile_X0Y15_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X1Y15_Emulate_Bitstream)
    )
`endif
    Tile_X1Y15_linear_LMDPL
    (
    .from_NA(Tile_X1Y16_to_NA),
    .from_NB(Tile_X1Y16_to_NB),
    .from_NC(Tile_X1Y16_to_NC),
    .from_ND(Tile_X1Y16_to_ND),
    .from_NF(Tile_X1Y16_to_NF),
    .from_NG(Tile_X1Y16_to_NG),
    .from_NH(Tile_X1Y16_to_NH),
    .from_NI(Tile_X1Y16_to_NI),
    .from_EA(Tile_X0Y15_to_EA),
    .from_EB(Tile_X0Y15_to_EB),
    .from_EC(Tile_X0Y15_to_EC),
    .from_ED(Tile_X0Y15_to_ED),
    .from_EF(Tile_X0Y15_to_EF),
    .from_EG(Tile_X0Y15_to_EG),
    .from_EH(Tile_X0Y15_to_EH),
    .from_EI(Tile_X0Y15_to_EI),
    .from_SA(Tile_X1Y14_to_SA),
    .from_SB(Tile_X1Y14_to_SB),
    .from_SC(Tile_X1Y14_to_SC),
    .from_SD(Tile_X1Y14_to_SD),
    .from_SF(Tile_X1Y14_to_SF),
    .from_SG(Tile_X1Y14_to_SG),
    .from_SH(Tile_X1Y14_to_SH),
    .from_SI(Tile_X1Y14_to_SI),
    .from_WA(Tile_X2Y15_to_WA),
    .from_WB(Tile_X2Y15_to_WB),
    .from_WC(Tile_X2Y15_to_WC),
    .from_WD(Tile_X2Y15_to_WD),
    .from_WF(Tile_X2Y15_to_WF),
    .from_WG(Tile_X2Y15_to_WG),
    .from_WH(Tile_X2Y15_to_WH),
    .from_WI(Tile_X2Y15_to_WI),
    .to_EA(Tile_X1Y15_to_EA),
    .to_EB(Tile_X1Y15_to_EB),
    .to_EC(Tile_X1Y15_to_EC),
    .to_ED(Tile_X1Y15_to_ED),
    .to_EF(Tile_X1Y15_to_EF),
    .to_EG(Tile_X1Y15_to_EG),
    .to_EH(Tile_X1Y15_to_EH),
    .to_EI(Tile_X1Y15_to_EI),
    .to_WA(Tile_X1Y15_to_WA),
    .to_WB(Tile_X1Y15_to_WB),
    .to_WC(Tile_X1Y15_to_WC),
    .to_WD(Tile_X1Y15_to_WD),
    .to_WF(Tile_X1Y15_to_WF),
    .to_WG(Tile_X1Y15_to_WG),
    .to_WH(Tile_X1Y15_to_WH),
    .to_WI(Tile_X1Y15_to_WI),
    .to_NA(Tile_X1Y15_to_NA),
    .to_NB(Tile_X1Y15_to_NB),
    .to_NC(Tile_X1Y15_to_NC),
    .to_ND(Tile_X1Y15_to_ND),
    .to_NF(Tile_X1Y15_to_NF),
    .to_NG(Tile_X1Y15_to_NG),
    .to_NH(Tile_X1Y15_to_NH),
    .to_NI(Tile_X1Y15_to_NI),
    .to_SA(Tile_X1Y15_to_SA),
    .to_SB(Tile_X1Y15_to_SB),
    .to_SC(Tile_X1Y15_to_SC),
    .to_SD(Tile_X1Y15_to_SD),
    .to_SF(Tile_X1Y15_to_SF),
    .to_SG(Tile_X1Y15_to_SG),
    .to_SH(Tile_X1Y15_to_SH),
    .to_SI(Tile_X1Y15_to_SI),
    .F_masked1(Tile_X1Y15_F_masked1),
    .F_masked2(Tile_X1Y15_F_masked2),
    .UserCLK(Tile_X1Y16_UserCLKo),
    .UserCLKo(Tile_X1Y15_UserCLKo),
    .rst(Tile_X1Y16_rsto),
    .rsto(Tile_X1Y15_rsto),
    .FrameData(Tile_X0Y15_FrameData_O),
    .FrameData_O(Tile_X1Y15_FrameData_O),
    .FrameStrobe(Tile_X1Y16_FrameStrobe_O),
    .FrameStrobe_O(Tile_X1Y15_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X2Y15_Emulate_Bitstream)
    )
`endif
    Tile_X2Y15_linear_LMDPL
    (
    .from_NA(Tile_X2Y16_to_NA),
    .from_NB(Tile_X2Y16_to_NB),
    .from_NC(Tile_X2Y16_to_NC),
    .from_ND(Tile_X2Y16_to_ND),
    .from_NF(Tile_X2Y16_to_NF),
    .from_NG(Tile_X2Y16_to_NG),
    .from_NH(Tile_X2Y16_to_NH),
    .from_NI(Tile_X2Y16_to_NI),
    .from_EA(Tile_X1Y15_to_EA),
    .from_EB(Tile_X1Y15_to_EB),
    .from_EC(Tile_X1Y15_to_EC),
    .from_ED(Tile_X1Y15_to_ED),
    .from_EF(Tile_X1Y15_to_EF),
    .from_EG(Tile_X1Y15_to_EG),
    .from_EH(Tile_X1Y15_to_EH),
    .from_EI(Tile_X1Y15_to_EI),
    .from_SA(Tile_X2Y14_to_SA),
    .from_SB(Tile_X2Y14_to_SB),
    .from_SC(Tile_X2Y14_to_SC),
    .from_SD(Tile_X2Y14_to_SD),
    .from_SF(Tile_X2Y14_to_SF),
    .from_SG(Tile_X2Y14_to_SG),
    .from_SH(Tile_X2Y14_to_SH),
    .from_SI(Tile_X2Y14_to_SI),
    .from_WA(Tile_X3Y15_to_WA),
    .from_WB(Tile_X3Y15_to_WB),
    .from_WC(Tile_X3Y15_to_WC),
    .from_WD(Tile_X3Y15_to_WD),
    .from_WF(Tile_X3Y15_to_WF),
    .from_WG(Tile_X3Y15_to_WG),
    .from_WH(Tile_X3Y15_to_WH),
    .from_WI(Tile_X3Y15_to_WI),
    .to_EA(Tile_X2Y15_to_EA),
    .to_EB(Tile_X2Y15_to_EB),
    .to_EC(Tile_X2Y15_to_EC),
    .to_ED(Tile_X2Y15_to_ED),
    .to_EF(Tile_X2Y15_to_EF),
    .to_EG(Tile_X2Y15_to_EG),
    .to_EH(Tile_X2Y15_to_EH),
    .to_EI(Tile_X2Y15_to_EI),
    .to_WA(Tile_X2Y15_to_WA),
    .to_WB(Tile_X2Y15_to_WB),
    .to_WC(Tile_X2Y15_to_WC),
    .to_WD(Tile_X2Y15_to_WD),
    .to_WF(Tile_X2Y15_to_WF),
    .to_WG(Tile_X2Y15_to_WG),
    .to_WH(Tile_X2Y15_to_WH),
    .to_WI(Tile_X2Y15_to_WI),
    .to_NA(Tile_X2Y15_to_NA),
    .to_NB(Tile_X2Y15_to_NB),
    .to_NC(Tile_X2Y15_to_NC),
    .to_ND(Tile_X2Y15_to_ND),
    .to_NF(Tile_X2Y15_to_NF),
    .to_NG(Tile_X2Y15_to_NG),
    .to_NH(Tile_X2Y15_to_NH),
    .to_NI(Tile_X2Y15_to_NI),
    .to_SA(Tile_X2Y15_to_SA),
    .to_SB(Tile_X2Y15_to_SB),
    .to_SC(Tile_X2Y15_to_SC),
    .to_SD(Tile_X2Y15_to_SD),
    .to_SF(Tile_X2Y15_to_SF),
    .to_SG(Tile_X2Y15_to_SG),
    .to_SH(Tile_X2Y15_to_SH),
    .to_SI(Tile_X2Y15_to_SI),
    .F_masked1(Tile_X2Y15_F_masked1),
    .F_masked2(Tile_X2Y15_F_masked2),
    .UserCLK(Tile_X2Y16_UserCLKo),
    .UserCLKo(Tile_X2Y15_UserCLKo),
    .rst(Tile_X2Y16_rsto),
    .rsto(Tile_X2Y15_rsto),
    .FrameData(Tile_X1Y15_FrameData_O),
    .FrameData_O(Tile_X2Y15_FrameData_O),
    .FrameStrobe(Tile_X2Y16_FrameStrobe_O),
    .FrameStrobe_O(Tile_X2Y15_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
nonlinear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X3Y15_Emulate_Bitstream)
    )
`endif
    Tile_X3Y15_nonlinear_LMDPL
    (
    .from_NA(Tile_X3Y16_to_NA),
    .from_NB(Tile_X3Y16_to_NB),
    .from_NC(Tile_X3Y16_to_NC),
    .from_ND(Tile_X3Y16_to_ND),
    .from_NF(Tile_X3Y16_to_NF),
    .from_NG(Tile_X3Y16_to_NG),
    .from_NH(Tile_X3Y16_to_NH),
    .from_NI(Tile_X3Y16_to_NI),
    .from_EA(Tile_X2Y15_to_EA),
    .from_EB(Tile_X2Y15_to_EB),
    .from_EC(Tile_X2Y15_to_EC),
    .from_ED(Tile_X2Y15_to_ED),
    .from_EF(Tile_X2Y15_to_EF),
    .from_EG(Tile_X2Y15_to_EG),
    .from_EH(Tile_X2Y15_to_EH),
    .from_EI(Tile_X2Y15_to_EI),
    .from_SA(Tile_X3Y14_to_SA),
    .from_SB(Tile_X3Y14_to_SB),
    .from_SC(Tile_X3Y14_to_SC),
    .from_SD(Tile_X3Y14_to_SD),
    .from_SF(Tile_X3Y14_to_SF),
    .from_SG(Tile_X3Y14_to_SG),
    .from_SH(Tile_X3Y14_to_SH),
    .from_SI(Tile_X3Y14_to_SI),
    .from_WA(Tile_X4Y15_to_WA),
    .from_WB(Tile_X4Y15_to_WB),
    .from_WC(Tile_X4Y15_to_WC),
    .from_WD(Tile_X4Y15_to_WD),
    .from_WF(Tile_X4Y15_to_WF),
    .from_WG(Tile_X4Y15_to_WG),
    .from_WH(Tile_X4Y15_to_WH),
    .from_WI(Tile_X4Y15_to_WI),
    .to_EA(Tile_X3Y15_to_EA),
    .to_EB(Tile_X3Y15_to_EB),
    .to_EC(Tile_X3Y15_to_EC),
    .to_ED(Tile_X3Y15_to_ED),
    .to_EF(Tile_X3Y15_to_EF),
    .to_EG(Tile_X3Y15_to_EG),
    .to_EH(Tile_X3Y15_to_EH),
    .to_EI(Tile_X3Y15_to_EI),
    .to_WA(Tile_X3Y15_to_WA),
    .to_WB(Tile_X3Y15_to_WB),
    .to_WC(Tile_X3Y15_to_WC),
    .to_WD(Tile_X3Y15_to_WD),
    .to_WF(Tile_X3Y15_to_WF),
    .to_WG(Tile_X3Y15_to_WG),
    .to_WH(Tile_X3Y15_to_WH),
    .to_WI(Tile_X3Y15_to_WI),
    .to_NA(Tile_X3Y15_to_NA),
    .to_NB(Tile_X3Y15_to_NB),
    .to_NC(Tile_X3Y15_to_NC),
    .to_ND(Tile_X3Y15_to_ND),
    .to_NF(Tile_X3Y15_to_NF),
    .to_NG(Tile_X3Y15_to_NG),
    .to_NH(Tile_X3Y15_to_NH),
    .to_NI(Tile_X3Y15_to_NI),
    .to_SA(Tile_X3Y15_to_SA),
    .to_SB(Tile_X3Y15_to_SB),
    .to_SC(Tile_X3Y15_to_SC),
    .to_SD(Tile_X3Y15_to_SD),
    .to_SF(Tile_X3Y15_to_SF),
    .to_SG(Tile_X3Y15_to_SG),
    .to_SH(Tile_X3Y15_to_SH),
    .to_SI(Tile_X3Y15_to_SI),
    .R_t(Tile_X3Y15_R_t),
    .R_f(Tile_X3Y15_R_f),
    .F_masked1(Tile_X3Y15_F_masked1),
    .F_masked2(Tile_X3Y15_F_masked2),
    .UserCLK(Tile_X3Y16_UserCLKo),
    .UserCLKo(Tile_X3Y15_UserCLKo),
    .rst(Tile_X3Y16_rsto),
    .rsto(Tile_X3Y15_rsto),
    .FrameData(Tile_X2Y15_FrameData_O),
    .FrameData_O(Tile_X3Y15_FrameData_O),
    .FrameStrobe(Tile_X3Y16_FrameStrobe_O),
    .FrameStrobe_O(Tile_X3Y15_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X4Y15_Emulate_Bitstream)
    )
`endif
    Tile_X4Y15_linear_LMDPL
    (
    .from_NA(Tile_X4Y16_to_NA),
    .from_NB(Tile_X4Y16_to_NB),
    .from_NC(Tile_X4Y16_to_NC),
    .from_ND(Tile_X4Y16_to_ND),
    .from_NF(Tile_X4Y16_to_NF),
    .from_NG(Tile_X4Y16_to_NG),
    .from_NH(Tile_X4Y16_to_NH),
    .from_NI(Tile_X4Y16_to_NI),
    .from_EA(Tile_X3Y15_to_EA),
    .from_EB(Tile_X3Y15_to_EB),
    .from_EC(Tile_X3Y15_to_EC),
    .from_ED(Tile_X3Y15_to_ED),
    .from_EF(Tile_X3Y15_to_EF),
    .from_EG(Tile_X3Y15_to_EG),
    .from_EH(Tile_X3Y15_to_EH),
    .from_EI(Tile_X3Y15_to_EI),
    .from_SA(Tile_X4Y14_to_SA),
    .from_SB(Tile_X4Y14_to_SB),
    .from_SC(Tile_X4Y14_to_SC),
    .from_SD(Tile_X4Y14_to_SD),
    .from_SF(Tile_X4Y14_to_SF),
    .from_SG(Tile_X4Y14_to_SG),
    .from_SH(Tile_X4Y14_to_SH),
    .from_SI(Tile_X4Y14_to_SI),
    .from_WA(Tile_X5Y15_to_WA),
    .from_WB(Tile_X5Y15_to_WB),
    .from_WC(Tile_X5Y15_to_WC),
    .from_WD(Tile_X5Y15_to_WD),
    .from_WF(Tile_X5Y15_to_WF),
    .from_WG(Tile_X5Y15_to_WG),
    .from_WH(Tile_X5Y15_to_WH),
    .from_WI(Tile_X5Y15_to_WI),
    .to_EA(Tile_X4Y15_to_EA),
    .to_EB(Tile_X4Y15_to_EB),
    .to_EC(Tile_X4Y15_to_EC),
    .to_ED(Tile_X4Y15_to_ED),
    .to_EF(Tile_X4Y15_to_EF),
    .to_EG(Tile_X4Y15_to_EG),
    .to_EH(Tile_X4Y15_to_EH),
    .to_EI(Tile_X4Y15_to_EI),
    .to_WA(Tile_X4Y15_to_WA),
    .to_WB(Tile_X4Y15_to_WB),
    .to_WC(Tile_X4Y15_to_WC),
    .to_WD(Tile_X4Y15_to_WD),
    .to_WF(Tile_X4Y15_to_WF),
    .to_WG(Tile_X4Y15_to_WG),
    .to_WH(Tile_X4Y15_to_WH),
    .to_WI(Tile_X4Y15_to_WI),
    .to_NA(Tile_X4Y15_to_NA),
    .to_NB(Tile_X4Y15_to_NB),
    .to_NC(Tile_X4Y15_to_NC),
    .to_ND(Tile_X4Y15_to_ND),
    .to_NF(Tile_X4Y15_to_NF),
    .to_NG(Tile_X4Y15_to_NG),
    .to_NH(Tile_X4Y15_to_NH),
    .to_NI(Tile_X4Y15_to_NI),
    .to_SA(Tile_X4Y15_to_SA),
    .to_SB(Tile_X4Y15_to_SB),
    .to_SC(Tile_X4Y15_to_SC),
    .to_SD(Tile_X4Y15_to_SD),
    .to_SF(Tile_X4Y15_to_SF),
    .to_SG(Tile_X4Y15_to_SG),
    .to_SH(Tile_X4Y15_to_SH),
    .to_SI(Tile_X4Y15_to_SI),
    .F_masked1(Tile_X4Y15_F_masked1),
    .F_masked2(Tile_X4Y15_F_masked2),
    .UserCLK(Tile_X4Y16_UserCLKo),
    .UserCLKo(Tile_X4Y15_UserCLKo),
    .rst(Tile_X4Y16_rsto),
    .rsto(Tile_X4Y15_rsto),
    .FrameData(Tile_X3Y15_FrameData_O),
    .FrameData_O(Tile_X4Y15_FrameData_O),
    .FrameStrobe(Tile_X4Y16_FrameStrobe_O),
    .FrameStrobe_O(Tile_X4Y15_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X5Y15_Emulate_Bitstream)
    )
`endif
    Tile_X5Y15_linear_LMDPL
    (
    .from_NA(Tile_X5Y16_to_NA),
    .from_NB(Tile_X5Y16_to_NB),
    .from_NC(Tile_X5Y16_to_NC),
    .from_ND(Tile_X5Y16_to_ND),
    .from_NF(Tile_X5Y16_to_NF),
    .from_NG(Tile_X5Y16_to_NG),
    .from_NH(Tile_X5Y16_to_NH),
    .from_NI(Tile_X5Y16_to_NI),
    .from_EA(Tile_X4Y15_to_EA),
    .from_EB(Tile_X4Y15_to_EB),
    .from_EC(Tile_X4Y15_to_EC),
    .from_ED(Tile_X4Y15_to_ED),
    .from_EF(Tile_X4Y15_to_EF),
    .from_EG(Tile_X4Y15_to_EG),
    .from_EH(Tile_X4Y15_to_EH),
    .from_EI(Tile_X4Y15_to_EI),
    .from_SA(Tile_X5Y14_to_SA),
    .from_SB(Tile_X5Y14_to_SB),
    .from_SC(Tile_X5Y14_to_SC),
    .from_SD(Tile_X5Y14_to_SD),
    .from_SF(Tile_X5Y14_to_SF),
    .from_SG(Tile_X5Y14_to_SG),
    .from_SH(Tile_X5Y14_to_SH),
    .from_SI(Tile_X5Y14_to_SI),
    .from_WA(Tile_X6Y15_to_WA),
    .from_WB(Tile_X6Y15_to_WB),
    .from_WC(Tile_X6Y15_to_WC),
    .from_WD(Tile_X6Y15_to_WD),
    .from_WF(Tile_X6Y15_to_WF),
    .from_WG(Tile_X6Y15_to_WG),
    .from_WH(Tile_X6Y15_to_WH),
    .from_WI(Tile_X6Y15_to_WI),
    .to_EA(Tile_X5Y15_to_EA),
    .to_EB(Tile_X5Y15_to_EB),
    .to_EC(Tile_X5Y15_to_EC),
    .to_ED(Tile_X5Y15_to_ED),
    .to_EF(Tile_X5Y15_to_EF),
    .to_EG(Tile_X5Y15_to_EG),
    .to_EH(Tile_X5Y15_to_EH),
    .to_EI(Tile_X5Y15_to_EI),
    .to_WA(Tile_X5Y15_to_WA),
    .to_WB(Tile_X5Y15_to_WB),
    .to_WC(Tile_X5Y15_to_WC),
    .to_WD(Tile_X5Y15_to_WD),
    .to_WF(Tile_X5Y15_to_WF),
    .to_WG(Tile_X5Y15_to_WG),
    .to_WH(Tile_X5Y15_to_WH),
    .to_WI(Tile_X5Y15_to_WI),
    .to_NA(Tile_X5Y15_to_NA),
    .to_NB(Tile_X5Y15_to_NB),
    .to_NC(Tile_X5Y15_to_NC),
    .to_ND(Tile_X5Y15_to_ND),
    .to_NF(Tile_X5Y15_to_NF),
    .to_NG(Tile_X5Y15_to_NG),
    .to_NH(Tile_X5Y15_to_NH),
    .to_NI(Tile_X5Y15_to_NI),
    .to_SA(Tile_X5Y15_to_SA),
    .to_SB(Tile_X5Y15_to_SB),
    .to_SC(Tile_X5Y15_to_SC),
    .to_SD(Tile_X5Y15_to_SD),
    .to_SF(Tile_X5Y15_to_SF),
    .to_SG(Tile_X5Y15_to_SG),
    .to_SH(Tile_X5Y15_to_SH),
    .to_SI(Tile_X5Y15_to_SI),
    .F_masked1(Tile_X5Y15_F_masked1),
    .F_masked2(Tile_X5Y15_F_masked2),
    .UserCLK(Tile_X5Y16_UserCLKo),
    .UserCLKo(Tile_X5Y15_UserCLKo),
    .rst(Tile_X5Y16_rsto),
    .rsto(Tile_X5Y15_rsto),
    .FrameData(Tile_X4Y15_FrameData_O),
    .FrameData_O(Tile_X5Y15_FrameData_O),
    .FrameStrobe(Tile_X5Y16_FrameStrobe_O),
    .FrameStrobe_O(Tile_X5Y15_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
nonlinear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X6Y15_Emulate_Bitstream)
    )
`endif
    Tile_X6Y15_nonlinear_LMDPL
    (
    .from_NA(Tile_X6Y16_to_NA),
    .from_NB(Tile_X6Y16_to_NB),
    .from_NC(Tile_X6Y16_to_NC),
    .from_ND(Tile_X6Y16_to_ND),
    .from_NF(Tile_X6Y16_to_NF),
    .from_NG(Tile_X6Y16_to_NG),
    .from_NH(Tile_X6Y16_to_NH),
    .from_NI(Tile_X6Y16_to_NI),
    .from_EA(Tile_X5Y15_to_EA),
    .from_EB(Tile_X5Y15_to_EB),
    .from_EC(Tile_X5Y15_to_EC),
    .from_ED(Tile_X5Y15_to_ED),
    .from_EF(Tile_X5Y15_to_EF),
    .from_EG(Tile_X5Y15_to_EG),
    .from_EH(Tile_X5Y15_to_EH),
    .from_EI(Tile_X5Y15_to_EI),
    .from_SA(Tile_X6Y14_to_SA),
    .from_SB(Tile_X6Y14_to_SB),
    .from_SC(Tile_X6Y14_to_SC),
    .from_SD(Tile_X6Y14_to_SD),
    .from_SF(Tile_X6Y14_to_SF),
    .from_SG(Tile_X6Y14_to_SG),
    .from_SH(Tile_X6Y14_to_SH),
    .from_SI(Tile_X6Y14_to_SI),
    .from_WA(Tile_X7Y15_to_WA),
    .from_WB(Tile_X7Y15_to_WB),
    .from_WC(Tile_X7Y15_to_WC),
    .from_WD(Tile_X7Y15_to_WD),
    .from_WF(Tile_X7Y15_to_WF),
    .from_WG(Tile_X7Y15_to_WG),
    .from_WH(Tile_X7Y15_to_WH),
    .from_WI(Tile_X7Y15_to_WI),
    .to_EA(Tile_X6Y15_to_EA),
    .to_EB(Tile_X6Y15_to_EB),
    .to_EC(Tile_X6Y15_to_EC),
    .to_ED(Tile_X6Y15_to_ED),
    .to_EF(Tile_X6Y15_to_EF),
    .to_EG(Tile_X6Y15_to_EG),
    .to_EH(Tile_X6Y15_to_EH),
    .to_EI(Tile_X6Y15_to_EI),
    .to_WA(Tile_X6Y15_to_WA),
    .to_WB(Tile_X6Y15_to_WB),
    .to_WC(Tile_X6Y15_to_WC),
    .to_WD(Tile_X6Y15_to_WD),
    .to_WF(Tile_X6Y15_to_WF),
    .to_WG(Tile_X6Y15_to_WG),
    .to_WH(Tile_X6Y15_to_WH),
    .to_WI(Tile_X6Y15_to_WI),
    .to_NA(Tile_X6Y15_to_NA),
    .to_NB(Tile_X6Y15_to_NB),
    .to_NC(Tile_X6Y15_to_NC),
    .to_ND(Tile_X6Y15_to_ND),
    .to_NF(Tile_X6Y15_to_NF),
    .to_NG(Tile_X6Y15_to_NG),
    .to_NH(Tile_X6Y15_to_NH),
    .to_NI(Tile_X6Y15_to_NI),
    .to_SA(Tile_X6Y15_to_SA),
    .to_SB(Tile_X6Y15_to_SB),
    .to_SC(Tile_X6Y15_to_SC),
    .to_SD(Tile_X6Y15_to_SD),
    .to_SF(Tile_X6Y15_to_SF),
    .to_SG(Tile_X6Y15_to_SG),
    .to_SH(Tile_X6Y15_to_SH),
    .to_SI(Tile_X6Y15_to_SI),
    .R_t(Tile_X6Y15_R_t),
    .R_f(Tile_X6Y15_R_f),
    .F_masked1(Tile_X6Y15_F_masked1),
    .F_masked2(Tile_X6Y15_F_masked2),
    .UserCLK(Tile_X6Y16_UserCLKo),
    .UserCLKo(Tile_X6Y15_UserCLKo),
    .rst(Tile_X6Y16_rsto),
    .rsto(Tile_X6Y15_rsto),
    .FrameData(Tile_X5Y15_FrameData_O),
    .FrameData_O(Tile_X6Y15_FrameData_O),
    .FrameStrobe(Tile_X6Y16_FrameStrobe_O),
    .FrameStrobe_O(Tile_X6Y15_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X7Y15_Emulate_Bitstream)
    )
`endif
    Tile_X7Y15_linear_LMDPL
    (
    .from_NA(Tile_X7Y16_to_NA),
    .from_NB(Tile_X7Y16_to_NB),
    .from_NC(Tile_X7Y16_to_NC),
    .from_ND(Tile_X7Y16_to_ND),
    .from_NF(Tile_X7Y16_to_NF),
    .from_NG(Tile_X7Y16_to_NG),
    .from_NH(Tile_X7Y16_to_NH),
    .from_NI(Tile_X7Y16_to_NI),
    .from_EA(Tile_X6Y15_to_EA),
    .from_EB(Tile_X6Y15_to_EB),
    .from_EC(Tile_X6Y15_to_EC),
    .from_ED(Tile_X6Y15_to_ED),
    .from_EF(Tile_X6Y15_to_EF),
    .from_EG(Tile_X6Y15_to_EG),
    .from_EH(Tile_X6Y15_to_EH),
    .from_EI(Tile_X6Y15_to_EI),
    .from_SA(Tile_X7Y14_to_SA),
    .from_SB(Tile_X7Y14_to_SB),
    .from_SC(Tile_X7Y14_to_SC),
    .from_SD(Tile_X7Y14_to_SD),
    .from_SF(Tile_X7Y14_to_SF),
    .from_SG(Tile_X7Y14_to_SG),
    .from_SH(Tile_X7Y14_to_SH),
    .from_SI(Tile_X7Y14_to_SI),
    .from_WA(Tile_X8Y15_to_WA),
    .from_WB(Tile_X8Y15_to_WB),
    .from_WC(Tile_X8Y15_to_WC),
    .from_WD(Tile_X8Y15_to_WD),
    .from_WF(Tile_X8Y15_to_WF),
    .from_WG(Tile_X8Y15_to_WG),
    .from_WH(Tile_X8Y15_to_WH),
    .from_WI(Tile_X8Y15_to_WI),
    .to_EA(Tile_X7Y15_to_EA),
    .to_EB(Tile_X7Y15_to_EB),
    .to_EC(Tile_X7Y15_to_EC),
    .to_ED(Tile_X7Y15_to_ED),
    .to_EF(Tile_X7Y15_to_EF),
    .to_EG(Tile_X7Y15_to_EG),
    .to_EH(Tile_X7Y15_to_EH),
    .to_EI(Tile_X7Y15_to_EI),
    .to_WA(Tile_X7Y15_to_WA),
    .to_WB(Tile_X7Y15_to_WB),
    .to_WC(Tile_X7Y15_to_WC),
    .to_WD(Tile_X7Y15_to_WD),
    .to_WF(Tile_X7Y15_to_WF),
    .to_WG(Tile_X7Y15_to_WG),
    .to_WH(Tile_X7Y15_to_WH),
    .to_WI(Tile_X7Y15_to_WI),
    .to_NA(Tile_X7Y15_to_NA),
    .to_NB(Tile_X7Y15_to_NB),
    .to_NC(Tile_X7Y15_to_NC),
    .to_ND(Tile_X7Y15_to_ND),
    .to_NF(Tile_X7Y15_to_NF),
    .to_NG(Tile_X7Y15_to_NG),
    .to_NH(Tile_X7Y15_to_NH),
    .to_NI(Tile_X7Y15_to_NI),
    .to_SA(Tile_X7Y15_to_SA),
    .to_SB(Tile_X7Y15_to_SB),
    .to_SC(Tile_X7Y15_to_SC),
    .to_SD(Tile_X7Y15_to_SD),
    .to_SF(Tile_X7Y15_to_SF),
    .to_SG(Tile_X7Y15_to_SG),
    .to_SH(Tile_X7Y15_to_SH),
    .to_SI(Tile_X7Y15_to_SI),
    .F_masked1(Tile_X7Y15_F_masked1),
    .F_masked2(Tile_X7Y15_F_masked2),
    .UserCLK(Tile_X7Y16_UserCLKo),
    .UserCLKo(Tile_X7Y15_UserCLKo),
    .rst(Tile_X7Y16_rsto),
    .rsto(Tile_X7Y15_rsto),
    .FrameData(Tile_X6Y15_FrameData_O),
    .FrameData_O(Tile_X7Y15_FrameData_O),
    .FrameStrobe(Tile_X7Y16_FrameStrobe_O),
    .FrameStrobe_O(Tile_X7Y15_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
ctrl_to_sec
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X8Y15_Emulate_Bitstream)
    )
`endif
    Tile_X8Y15_ctrl_to_sec
    (
    .from_NA(Tile_X8Y16_to_NA),
    .from_NB(Tile_X8Y16_to_NB),
    .from_NC(Tile_X8Y16_to_NC),
    .from_ND(Tile_X8Y16_to_ND),
    .from_NF(Tile_X8Y16_to_NF),
    .from_NG(Tile_X8Y16_to_NG),
    .from_NH(Tile_X8Y16_to_NH),
    .from_NI(Tile_X8Y16_to_NI),
    .from_EA(Tile_X7Y15_to_EA),
    .from_EB(Tile_X7Y15_to_EB),
    .from_EC(Tile_X7Y15_to_EC),
    .from_ED(Tile_X7Y15_to_ED),
    .from_EF(Tile_X7Y15_to_EF),
    .from_EG(Tile_X7Y15_to_EG),
    .from_EH(Tile_X7Y15_to_EH),
    .from_EI(Tile_X7Y15_to_EI),
    .from_SA(Tile_X8Y14_to_SA),
    .from_SB(Tile_X8Y14_to_SB),
    .from_SC(Tile_X8Y14_to_SC),
    .from_SD(Tile_X8Y14_to_SD),
    .from_SF(Tile_X8Y14_to_SF),
    .from_SG(Tile_X8Y14_to_SG),
    .from_SH(Tile_X8Y14_to_SH),
    .from_SI(Tile_X8Y14_to_SI),
    .from_WA_1s(Tile_X9Y15_to_WA_1s),
    .from_WB_1s(Tile_X9Y15_to_WB_1s),
    .from_WC_1s(Tile_X9Y15_to_WC_1s),
    .from_WD_1s(Tile_X9Y15_to_WD_1s),
    .from_WF_1s(Tile_X9Y15_to_WF_1s),
    .from_WG_1s(Tile_X9Y15_to_WG_1s),
    .from_WH_1s(Tile_X9Y15_to_WH_1s),
    .from_WI_1s(Tile_X9Y15_to_WI_1s),
    .to_WA(Tile_X8Y15_to_WA),
    .to_WB(Tile_X8Y15_to_WB),
    .to_WC(Tile_X8Y15_to_WC),
    .to_WD(Tile_X8Y15_to_WD),
    .to_WF(Tile_X8Y15_to_WF),
    .to_WG(Tile_X8Y15_to_WG),
    .to_WH(Tile_X8Y15_to_WH),
    .to_WI(Tile_X8Y15_to_WI),
    .to_NA(Tile_X8Y15_to_NA),
    .to_NB(Tile_X8Y15_to_NB),
    .to_NC(Tile_X8Y15_to_NC),
    .to_ND(Tile_X8Y15_to_ND),
    .to_NF(Tile_X8Y15_to_NF),
    .to_NG(Tile_X8Y15_to_NG),
    .to_NH(Tile_X8Y15_to_NH),
    .to_NI(Tile_X8Y15_to_NI),
    .to_SA(Tile_X8Y15_to_SA),
    .to_SB(Tile_X8Y15_to_SB),
    .to_SC(Tile_X8Y15_to_SC),
    .to_SD(Tile_X8Y15_to_SD),
    .to_SF(Tile_X8Y15_to_SF),
    .to_SG(Tile_X8Y15_to_SG),
    .to_SH(Tile_X8Y15_to_SH),
    .to_SI(Tile_X8Y15_to_SI),
    .UserCLK(Tile_X8Y16_UserCLKo),
    .UserCLKo(Tile_X8Y15_UserCLKo),
    .rst(Tile_X8Y16_rsto),
    .rsto(Tile_X8Y15_rsto),
    .FrameData(Tile_X7Y15_FrameData_O),
    .FrameData_O(Tile_X8Y15_FrameData_O),
    .FrameStrobe(Tile_X8Y16_FrameStrobe_O),
    .FrameStrobe_O(Tile_X8Y15_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
combined_WDDL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X9Y15_Emulate_Bitstream)
    )
`endif
    Tile_X9Y15_combined_WDDL
    (
    .from_NA_1s(Tile_X9Y16_to_NA_1s),
    .from_NB_1s(Tile_X9Y16_to_NB_1s),
    .from_NC_1s(Tile_X9Y16_to_NC_1s),
    .from_ND_1s(Tile_X9Y16_to_ND_1s),
    .from_NF_1s(Tile_X9Y16_to_NF_1s),
    .from_NG_1s(Tile_X9Y16_to_NG_1s),
    .from_NH_1s(Tile_X9Y16_to_NH_1s),
    .from_NI_1s(Tile_X9Y16_to_NI_1s),
    .from_SA_1s(Tile_X9Y14_to_SA_1s),
    .from_SB_1s(Tile_X9Y14_to_SB_1s),
    .from_SC_1s(Tile_X9Y14_to_SC_1s),
    .from_SD_1s(Tile_X9Y14_to_SD_1s),
    .from_SF_1s(Tile_X9Y14_to_SF_1s),
    .from_SG_1s(Tile_X9Y14_to_SG_1s),
    .from_SH_1s(Tile_X9Y14_to_SH_1s),
    .from_SI_1s(Tile_X9Y14_to_SI_1s),
    .from_WA_1s(Tile_X10Y15_to_WA_1s),
    .from_WB_1s(Tile_X10Y15_to_WB_1s),
    .from_WC_1s(Tile_X10Y15_to_WC_1s),
    .from_WD_1s(Tile_X10Y15_to_WD_1s),
    .from_WF_1s(Tile_X10Y15_to_WF_1s),
    .from_WG_1s(Tile_X10Y15_to_WG_1s),
    .from_WH_1s(Tile_X10Y15_to_WH_1s),
    .from_WI_1s(Tile_X10Y15_to_WI_1s),
    .to_EA_1s(Tile_X9Y15_to_EA_1s),
    .to_EB_1s(Tile_X9Y15_to_EB_1s),
    .to_EC_1s(Tile_X9Y15_to_EC_1s),
    .to_ED_1s(Tile_X9Y15_to_ED_1s),
    .to_EF_1s(Tile_X9Y15_to_EF_1s),
    .to_EG_1s(Tile_X9Y15_to_EG_1s),
    .to_EH_1s(Tile_X9Y15_to_EH_1s),
    .to_EI_1s(Tile_X9Y15_to_EI_1s),
    .to_WA_1s(Tile_X9Y15_to_WA_1s),
    .to_WB_1s(Tile_X9Y15_to_WB_1s),
    .to_WC_1s(Tile_X9Y15_to_WC_1s),
    .to_WD_1s(Tile_X9Y15_to_WD_1s),
    .to_WF_1s(Tile_X9Y15_to_WF_1s),
    .to_WG_1s(Tile_X9Y15_to_WG_1s),
    .to_WH_1s(Tile_X9Y15_to_WH_1s),
    .to_WI_1s(Tile_X9Y15_to_WI_1s),
    .to_NA_1s(Tile_X9Y15_to_NA_1s),
    .to_NB_1s(Tile_X9Y15_to_NB_1s),
    .to_NC_1s(Tile_X9Y15_to_NC_1s),
    .to_ND_1s(Tile_X9Y15_to_ND_1s),
    .to_NF_1s(Tile_X9Y15_to_NF_1s),
    .to_NG_1s(Tile_X9Y15_to_NG_1s),
    .to_NH_1s(Tile_X9Y15_to_NH_1s),
    .to_NI_1s(Tile_X9Y15_to_NI_1s),
    .to_SA_1s(Tile_X9Y15_to_SA_1s),
    .to_SB_1s(Tile_X9Y15_to_SB_1s),
    .to_SC_1s(Tile_X9Y15_to_SC_1s),
    .to_SD_1s(Tile_X9Y15_to_SD_1s),
    .to_SF_1s(Tile_X9Y15_to_SF_1s),
    .to_SG_1s(Tile_X9Y15_to_SG_1s),
    .to_SH_1s(Tile_X9Y15_to_SH_1s),
    .to_SI_1s(Tile_X9Y15_to_SI_1s),
    .F_ctrl(Tile_X9Y15_F_ctrl),
    .UserCLK(Tile_X9Y16_UserCLKo),
    .UserCLKo(Tile_X9Y15_UserCLKo),
    .rst(Tile_X9Y16_rsto),
    .rsto(Tile_X9Y15_rsto),
    .FrameData(Tile_X8Y15_FrameData_O),
    .FrameData_O(Tile_X9Y15_FrameData_O),
    .FrameStrobe(Tile_X9Y16_FrameStrobe_O),
    .FrameStrobe_O(Tile_X9Y15_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
ctrl_IO
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X10Y15_Emulate_Bitstream)
    )
`endif
    Tile_X10Y15_ctrl_IO
    (
    .from_EA_1s(Tile_X9Y15_to_EA_1s),
    .from_EB_1s(Tile_X9Y15_to_EB_1s),
    .from_EC_1s(Tile_X9Y15_to_EC_1s),
    .from_ED_1s(Tile_X9Y15_to_ED_1s),
    .from_EF_1s(Tile_X9Y15_to_EF_1s),
    .from_EG_1s(Tile_X9Y15_to_EG_1s),
    .from_EH_1s(Tile_X9Y15_to_EH_1s),
    .from_EI_1s(Tile_X9Y15_to_EI_1s),
    .to_WA_1s(Tile_X10Y15_to_WA_1s),
    .to_WB_1s(Tile_X10Y15_to_WB_1s),
    .to_WC_1s(Tile_X10Y15_to_WC_1s),
    .to_WD_1s(Tile_X10Y15_to_WD_1s),
    .to_WF_1s(Tile_X10Y15_to_WF_1s),
    .to_WG_1s(Tile_X10Y15_to_WG_1s),
    .to_WH_1s(Tile_X10Y15_to_WH_1s),
    .to_WI_1s(Tile_X10Y15_to_WI_1s),
    .A_O_top_0_t(Tile_X10Y15_A_O_top_0_t),
    .A_O_top_0_f(Tile_X10Y15_A_O_top_0_f),
    .A_prech2(Tile_X10Y15_A_prech2),
    .A_DR_fault(Tile_X10Y15_A_DR_fault),
    .A_I_top_0_t(Tile_X10Y15_A_I_top_0_t),
    .A_I_top_0_f(Tile_X10Y15_A_I_top_0_f),
    .A_T_top(Tile_X10Y15_A_T_top),
    .A_F_ctrl(Tile_X10Y15_A_F_ctrl),
    .UserCLK(Tile_X10Y16_UserCLKo),
    .UserCLKo(Tile_X10Y15_UserCLKo),
    .rst(Tile_X10Y16_rsto),
    .rsto(Tile_X10Y15_rsto),
    .FrameData(Tile_X9Y15_FrameData_O),
    .FrameData_O(Tile_X10Y15_FrameData_O),
    .FrameStrobe(Tile_X10Y16_FrameStrobe_O),
    .FrameStrobe_O(Tile_X10Y15_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
W_IO_custom
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X0Y16_Emulate_Bitstream)
    )
`endif
    Tile_X0Y16_W_IO_custom
    (
    .from_NA(Tile_X0Y17_to_NA),
    .from_NB(Tile_X0Y17_to_NB),
    .from_NC(Tile_X0Y17_to_NC),
    .from_ND(Tile_X0Y17_to_ND),
    .from_NF(Tile_X0Y17_to_NF),
    .from_NG(Tile_X0Y17_to_NG),
    .from_NH(Tile_X0Y17_to_NH),
    .from_NI(Tile_X0Y17_to_NI),
    .from_SA(Tile_X0Y15_to_SA),
    .from_SB(Tile_X0Y15_to_SB),
    .from_SC(Tile_X0Y15_to_SC),
    .from_SD(Tile_X0Y15_to_SD),
    .from_SF(Tile_X0Y15_to_SF),
    .from_SG(Tile_X0Y15_to_SG),
    .from_SH(Tile_X0Y15_to_SH),
    .from_SI(Tile_X0Y15_to_SI),
    .from_WA(Tile_X1Y16_to_WA),
    .from_WB(Tile_X1Y16_to_WB),
    .from_WC(Tile_X1Y16_to_WC),
    .from_WD(Tile_X1Y16_to_WD),
    .from_WF(Tile_X1Y16_to_WF),
    .from_WG(Tile_X1Y16_to_WG),
    .from_WH(Tile_X1Y16_to_WH),
    .from_WI(Tile_X1Y16_to_WI),
    .to_EA(Tile_X0Y16_to_EA),
    .to_EB(Tile_X0Y16_to_EB),
    .to_EC(Tile_X0Y16_to_EC),
    .to_ED(Tile_X0Y16_to_ED),
    .to_EF(Tile_X0Y16_to_EF),
    .to_EG(Tile_X0Y16_to_EG),
    .to_EH(Tile_X0Y16_to_EH),
    .to_EI(Tile_X0Y16_to_EI),
    .to_NA(Tile_X0Y16_to_NA),
    .to_NB(Tile_X0Y16_to_NB),
    .to_NC(Tile_X0Y16_to_NC),
    .to_ND(Tile_X0Y16_to_ND),
    .to_NF(Tile_X0Y16_to_NF),
    .to_NG(Tile_X0Y16_to_NG),
    .to_NH(Tile_X0Y16_to_NH),
    .to_NI(Tile_X0Y16_to_NI),
    .to_SA(Tile_X0Y16_to_SA),
    .to_SB(Tile_X0Y16_to_SB),
    .to_SC(Tile_X0Y16_to_SC),
    .to_SD(Tile_X0Y16_to_SD),
    .to_SF(Tile_X0Y16_to_SF),
    .to_SG(Tile_X0Y16_to_SG),
    .to_SH(Tile_X0Y16_to_SH),
    .to_SI(Tile_X0Y16_to_SI),
    .A_O_top_0_t(Tile_X0Y16_A_O_top_0_t),
    .A_O_top_0_f(Tile_X0Y16_A_O_top_0_f),
    .A_O_top_1_t(Tile_X0Y16_A_O_top_1_t),
    .A_O_top_1_f(Tile_X0Y16_A_O_top_1_f),
    .A_prech1(Tile_X0Y16_A_prech1),
    .A_prech2(Tile_X0Y16_A_prech2),
    .A_DR_fault(Tile_X0Y16_A_DR_fault),
    .A_I_top_0_t(Tile_X0Y16_A_I_top_0_t),
    .A_I_top_0_f(Tile_X0Y16_A_I_top_0_f),
    .A_I_top_1_t(Tile_X0Y16_A_I_top_1_t),
    .A_I_top_1_f(Tile_X0Y16_A_I_top_1_f),
    .A_T_top(Tile_X0Y16_A_T_top),
    .A_F_masked1(Tile_X0Y16_A_F_masked1),
    .A_F_masked2(Tile_X0Y16_A_F_masked2),
    .A_config_C_bit0(Tile_X0Y16_A_config_C_bit0),
    .A_config_C_bit1(Tile_X0Y16_A_config_C_bit1),
    .A_config_C_bit2(Tile_X0Y16_A_config_C_bit2),
    .A_config_C_bit3(Tile_X0Y16_A_config_C_bit3),
    .B_config_C_bit0(Tile_X0Y16_B_config_C_bit0),
    .B_config_C_bit1(Tile_X0Y16_B_config_C_bit1),
    .B_config_C_bit2(Tile_X0Y16_B_config_C_bit2),
    .B_config_C_bit3(Tile_X0Y16_B_config_C_bit3),
    .UserCLK(Tile_X0Y17_UserCLKo),
    .UserCLKo(Tile_X0Y16_UserCLKo),
    .rst(Tile_X0Y17_rsto),
    .rsto(Tile_X0Y16_rsto),
    .FrameData(Tile_Y16_FrameData),
    .FrameData_O(Tile_X0Y16_FrameData_O),
    .FrameStrobe(Tile_X0Y17_FrameStrobe_O),
    .FrameStrobe_O(Tile_X0Y16_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X1Y16_Emulate_Bitstream)
    )
`endif
    Tile_X1Y16_linear_LMDPL
    (
    .from_NA(Tile_X1Y17_to_NA),
    .from_NB(Tile_X1Y17_to_NB),
    .from_NC(Tile_X1Y17_to_NC),
    .from_ND(Tile_X1Y17_to_ND),
    .from_NF(Tile_X1Y17_to_NF),
    .from_NG(Tile_X1Y17_to_NG),
    .from_NH(Tile_X1Y17_to_NH),
    .from_NI(Tile_X1Y17_to_NI),
    .from_EA(Tile_X0Y16_to_EA),
    .from_EB(Tile_X0Y16_to_EB),
    .from_EC(Tile_X0Y16_to_EC),
    .from_ED(Tile_X0Y16_to_ED),
    .from_EF(Tile_X0Y16_to_EF),
    .from_EG(Tile_X0Y16_to_EG),
    .from_EH(Tile_X0Y16_to_EH),
    .from_EI(Tile_X0Y16_to_EI),
    .from_SA(Tile_X1Y15_to_SA),
    .from_SB(Tile_X1Y15_to_SB),
    .from_SC(Tile_X1Y15_to_SC),
    .from_SD(Tile_X1Y15_to_SD),
    .from_SF(Tile_X1Y15_to_SF),
    .from_SG(Tile_X1Y15_to_SG),
    .from_SH(Tile_X1Y15_to_SH),
    .from_SI(Tile_X1Y15_to_SI),
    .from_WA(Tile_X2Y16_to_WA),
    .from_WB(Tile_X2Y16_to_WB),
    .from_WC(Tile_X2Y16_to_WC),
    .from_WD(Tile_X2Y16_to_WD),
    .from_WF(Tile_X2Y16_to_WF),
    .from_WG(Tile_X2Y16_to_WG),
    .from_WH(Tile_X2Y16_to_WH),
    .from_WI(Tile_X2Y16_to_WI),
    .to_EA(Tile_X1Y16_to_EA),
    .to_EB(Tile_X1Y16_to_EB),
    .to_EC(Tile_X1Y16_to_EC),
    .to_ED(Tile_X1Y16_to_ED),
    .to_EF(Tile_X1Y16_to_EF),
    .to_EG(Tile_X1Y16_to_EG),
    .to_EH(Tile_X1Y16_to_EH),
    .to_EI(Tile_X1Y16_to_EI),
    .to_WA(Tile_X1Y16_to_WA),
    .to_WB(Tile_X1Y16_to_WB),
    .to_WC(Tile_X1Y16_to_WC),
    .to_WD(Tile_X1Y16_to_WD),
    .to_WF(Tile_X1Y16_to_WF),
    .to_WG(Tile_X1Y16_to_WG),
    .to_WH(Tile_X1Y16_to_WH),
    .to_WI(Tile_X1Y16_to_WI),
    .to_NA(Tile_X1Y16_to_NA),
    .to_NB(Tile_X1Y16_to_NB),
    .to_NC(Tile_X1Y16_to_NC),
    .to_ND(Tile_X1Y16_to_ND),
    .to_NF(Tile_X1Y16_to_NF),
    .to_NG(Tile_X1Y16_to_NG),
    .to_NH(Tile_X1Y16_to_NH),
    .to_NI(Tile_X1Y16_to_NI),
    .to_SA(Tile_X1Y16_to_SA),
    .to_SB(Tile_X1Y16_to_SB),
    .to_SC(Tile_X1Y16_to_SC),
    .to_SD(Tile_X1Y16_to_SD),
    .to_SF(Tile_X1Y16_to_SF),
    .to_SG(Tile_X1Y16_to_SG),
    .to_SH(Tile_X1Y16_to_SH),
    .to_SI(Tile_X1Y16_to_SI),
    .F_masked1(Tile_X1Y16_F_masked1),
    .F_masked2(Tile_X1Y16_F_masked2),
    .UserCLK(Tile_X1Y17_UserCLKo),
    .UserCLKo(Tile_X1Y16_UserCLKo),
    .rst(Tile_X1Y17_rsto),
    .rsto(Tile_X1Y16_rsto),
    .FrameData(Tile_X0Y16_FrameData_O),
    .FrameData_O(Tile_X1Y16_FrameData_O),
    .FrameStrobe(Tile_X1Y17_FrameStrobe_O),
    .FrameStrobe_O(Tile_X1Y16_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X2Y16_Emulate_Bitstream)
    )
`endif
    Tile_X2Y16_linear_LMDPL
    (
    .from_NA(Tile_X2Y17_to_NA),
    .from_NB(Tile_X2Y17_to_NB),
    .from_NC(Tile_X2Y17_to_NC),
    .from_ND(Tile_X2Y17_to_ND),
    .from_NF(Tile_X2Y17_to_NF),
    .from_NG(Tile_X2Y17_to_NG),
    .from_NH(Tile_X2Y17_to_NH),
    .from_NI(Tile_X2Y17_to_NI),
    .from_EA(Tile_X1Y16_to_EA),
    .from_EB(Tile_X1Y16_to_EB),
    .from_EC(Tile_X1Y16_to_EC),
    .from_ED(Tile_X1Y16_to_ED),
    .from_EF(Tile_X1Y16_to_EF),
    .from_EG(Tile_X1Y16_to_EG),
    .from_EH(Tile_X1Y16_to_EH),
    .from_EI(Tile_X1Y16_to_EI),
    .from_SA(Tile_X2Y15_to_SA),
    .from_SB(Tile_X2Y15_to_SB),
    .from_SC(Tile_X2Y15_to_SC),
    .from_SD(Tile_X2Y15_to_SD),
    .from_SF(Tile_X2Y15_to_SF),
    .from_SG(Tile_X2Y15_to_SG),
    .from_SH(Tile_X2Y15_to_SH),
    .from_SI(Tile_X2Y15_to_SI),
    .from_WA(Tile_X3Y16_to_WA),
    .from_WB(Tile_X3Y16_to_WB),
    .from_WC(Tile_X3Y16_to_WC),
    .from_WD(Tile_X3Y16_to_WD),
    .from_WF(Tile_X3Y16_to_WF),
    .from_WG(Tile_X3Y16_to_WG),
    .from_WH(Tile_X3Y16_to_WH),
    .from_WI(Tile_X3Y16_to_WI),
    .to_EA(Tile_X2Y16_to_EA),
    .to_EB(Tile_X2Y16_to_EB),
    .to_EC(Tile_X2Y16_to_EC),
    .to_ED(Tile_X2Y16_to_ED),
    .to_EF(Tile_X2Y16_to_EF),
    .to_EG(Tile_X2Y16_to_EG),
    .to_EH(Tile_X2Y16_to_EH),
    .to_EI(Tile_X2Y16_to_EI),
    .to_WA(Tile_X2Y16_to_WA),
    .to_WB(Tile_X2Y16_to_WB),
    .to_WC(Tile_X2Y16_to_WC),
    .to_WD(Tile_X2Y16_to_WD),
    .to_WF(Tile_X2Y16_to_WF),
    .to_WG(Tile_X2Y16_to_WG),
    .to_WH(Tile_X2Y16_to_WH),
    .to_WI(Tile_X2Y16_to_WI),
    .to_NA(Tile_X2Y16_to_NA),
    .to_NB(Tile_X2Y16_to_NB),
    .to_NC(Tile_X2Y16_to_NC),
    .to_ND(Tile_X2Y16_to_ND),
    .to_NF(Tile_X2Y16_to_NF),
    .to_NG(Tile_X2Y16_to_NG),
    .to_NH(Tile_X2Y16_to_NH),
    .to_NI(Tile_X2Y16_to_NI),
    .to_SA(Tile_X2Y16_to_SA),
    .to_SB(Tile_X2Y16_to_SB),
    .to_SC(Tile_X2Y16_to_SC),
    .to_SD(Tile_X2Y16_to_SD),
    .to_SF(Tile_X2Y16_to_SF),
    .to_SG(Tile_X2Y16_to_SG),
    .to_SH(Tile_X2Y16_to_SH),
    .to_SI(Tile_X2Y16_to_SI),
    .F_masked1(Tile_X2Y16_F_masked1),
    .F_masked2(Tile_X2Y16_F_masked2),
    .UserCLK(Tile_X2Y17_UserCLKo),
    .UserCLKo(Tile_X2Y16_UserCLKo),
    .rst(Tile_X2Y17_rsto),
    .rsto(Tile_X2Y16_rsto),
    .FrameData(Tile_X1Y16_FrameData_O),
    .FrameData_O(Tile_X2Y16_FrameData_O),
    .FrameStrobe(Tile_X2Y17_FrameStrobe_O),
    .FrameStrobe_O(Tile_X2Y16_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
nonlinear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X3Y16_Emulate_Bitstream)
    )
`endif
    Tile_X3Y16_nonlinear_LMDPL
    (
    .from_NA(Tile_X3Y17_to_NA),
    .from_NB(Tile_X3Y17_to_NB),
    .from_NC(Tile_X3Y17_to_NC),
    .from_ND(Tile_X3Y17_to_ND),
    .from_NF(Tile_X3Y17_to_NF),
    .from_NG(Tile_X3Y17_to_NG),
    .from_NH(Tile_X3Y17_to_NH),
    .from_NI(Tile_X3Y17_to_NI),
    .from_EA(Tile_X2Y16_to_EA),
    .from_EB(Tile_X2Y16_to_EB),
    .from_EC(Tile_X2Y16_to_EC),
    .from_ED(Tile_X2Y16_to_ED),
    .from_EF(Tile_X2Y16_to_EF),
    .from_EG(Tile_X2Y16_to_EG),
    .from_EH(Tile_X2Y16_to_EH),
    .from_EI(Tile_X2Y16_to_EI),
    .from_SA(Tile_X3Y15_to_SA),
    .from_SB(Tile_X3Y15_to_SB),
    .from_SC(Tile_X3Y15_to_SC),
    .from_SD(Tile_X3Y15_to_SD),
    .from_SF(Tile_X3Y15_to_SF),
    .from_SG(Tile_X3Y15_to_SG),
    .from_SH(Tile_X3Y15_to_SH),
    .from_SI(Tile_X3Y15_to_SI),
    .from_WA(Tile_X4Y16_to_WA),
    .from_WB(Tile_X4Y16_to_WB),
    .from_WC(Tile_X4Y16_to_WC),
    .from_WD(Tile_X4Y16_to_WD),
    .from_WF(Tile_X4Y16_to_WF),
    .from_WG(Tile_X4Y16_to_WG),
    .from_WH(Tile_X4Y16_to_WH),
    .from_WI(Tile_X4Y16_to_WI),
    .to_EA(Tile_X3Y16_to_EA),
    .to_EB(Tile_X3Y16_to_EB),
    .to_EC(Tile_X3Y16_to_EC),
    .to_ED(Tile_X3Y16_to_ED),
    .to_EF(Tile_X3Y16_to_EF),
    .to_EG(Tile_X3Y16_to_EG),
    .to_EH(Tile_X3Y16_to_EH),
    .to_EI(Tile_X3Y16_to_EI),
    .to_WA(Tile_X3Y16_to_WA),
    .to_WB(Tile_X3Y16_to_WB),
    .to_WC(Tile_X3Y16_to_WC),
    .to_WD(Tile_X3Y16_to_WD),
    .to_WF(Tile_X3Y16_to_WF),
    .to_WG(Tile_X3Y16_to_WG),
    .to_WH(Tile_X3Y16_to_WH),
    .to_WI(Tile_X3Y16_to_WI),
    .to_NA(Tile_X3Y16_to_NA),
    .to_NB(Tile_X3Y16_to_NB),
    .to_NC(Tile_X3Y16_to_NC),
    .to_ND(Tile_X3Y16_to_ND),
    .to_NF(Tile_X3Y16_to_NF),
    .to_NG(Tile_X3Y16_to_NG),
    .to_NH(Tile_X3Y16_to_NH),
    .to_NI(Tile_X3Y16_to_NI),
    .to_SA(Tile_X3Y16_to_SA),
    .to_SB(Tile_X3Y16_to_SB),
    .to_SC(Tile_X3Y16_to_SC),
    .to_SD(Tile_X3Y16_to_SD),
    .to_SF(Tile_X3Y16_to_SF),
    .to_SG(Tile_X3Y16_to_SG),
    .to_SH(Tile_X3Y16_to_SH),
    .to_SI(Tile_X3Y16_to_SI),
    .R_t(Tile_X3Y16_R_t),
    .R_f(Tile_X3Y16_R_f),
    .F_masked1(Tile_X3Y16_F_masked1),
    .F_masked2(Tile_X3Y16_F_masked2),
    .UserCLK(Tile_X3Y17_UserCLKo),
    .UserCLKo(Tile_X3Y16_UserCLKo),
    .rst(Tile_X3Y17_rsto),
    .rsto(Tile_X3Y16_rsto),
    .FrameData(Tile_X2Y16_FrameData_O),
    .FrameData_O(Tile_X3Y16_FrameData_O),
    .FrameStrobe(Tile_X3Y17_FrameStrobe_O),
    .FrameStrobe_O(Tile_X3Y16_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X4Y16_Emulate_Bitstream)
    )
`endif
    Tile_X4Y16_linear_LMDPL
    (
    .from_NA(Tile_X4Y17_to_NA),
    .from_NB(Tile_X4Y17_to_NB),
    .from_NC(Tile_X4Y17_to_NC),
    .from_ND(Tile_X4Y17_to_ND),
    .from_NF(Tile_X4Y17_to_NF),
    .from_NG(Tile_X4Y17_to_NG),
    .from_NH(Tile_X4Y17_to_NH),
    .from_NI(Tile_X4Y17_to_NI),
    .from_EA(Tile_X3Y16_to_EA),
    .from_EB(Tile_X3Y16_to_EB),
    .from_EC(Tile_X3Y16_to_EC),
    .from_ED(Tile_X3Y16_to_ED),
    .from_EF(Tile_X3Y16_to_EF),
    .from_EG(Tile_X3Y16_to_EG),
    .from_EH(Tile_X3Y16_to_EH),
    .from_EI(Tile_X3Y16_to_EI),
    .from_SA(Tile_X4Y15_to_SA),
    .from_SB(Tile_X4Y15_to_SB),
    .from_SC(Tile_X4Y15_to_SC),
    .from_SD(Tile_X4Y15_to_SD),
    .from_SF(Tile_X4Y15_to_SF),
    .from_SG(Tile_X4Y15_to_SG),
    .from_SH(Tile_X4Y15_to_SH),
    .from_SI(Tile_X4Y15_to_SI),
    .from_WA(Tile_X5Y16_to_WA),
    .from_WB(Tile_X5Y16_to_WB),
    .from_WC(Tile_X5Y16_to_WC),
    .from_WD(Tile_X5Y16_to_WD),
    .from_WF(Tile_X5Y16_to_WF),
    .from_WG(Tile_X5Y16_to_WG),
    .from_WH(Tile_X5Y16_to_WH),
    .from_WI(Tile_X5Y16_to_WI),
    .to_EA(Tile_X4Y16_to_EA),
    .to_EB(Tile_X4Y16_to_EB),
    .to_EC(Tile_X4Y16_to_EC),
    .to_ED(Tile_X4Y16_to_ED),
    .to_EF(Tile_X4Y16_to_EF),
    .to_EG(Tile_X4Y16_to_EG),
    .to_EH(Tile_X4Y16_to_EH),
    .to_EI(Tile_X4Y16_to_EI),
    .to_WA(Tile_X4Y16_to_WA),
    .to_WB(Tile_X4Y16_to_WB),
    .to_WC(Tile_X4Y16_to_WC),
    .to_WD(Tile_X4Y16_to_WD),
    .to_WF(Tile_X4Y16_to_WF),
    .to_WG(Tile_X4Y16_to_WG),
    .to_WH(Tile_X4Y16_to_WH),
    .to_WI(Tile_X4Y16_to_WI),
    .to_NA(Tile_X4Y16_to_NA),
    .to_NB(Tile_X4Y16_to_NB),
    .to_NC(Tile_X4Y16_to_NC),
    .to_ND(Tile_X4Y16_to_ND),
    .to_NF(Tile_X4Y16_to_NF),
    .to_NG(Tile_X4Y16_to_NG),
    .to_NH(Tile_X4Y16_to_NH),
    .to_NI(Tile_X4Y16_to_NI),
    .to_SA(Tile_X4Y16_to_SA),
    .to_SB(Tile_X4Y16_to_SB),
    .to_SC(Tile_X4Y16_to_SC),
    .to_SD(Tile_X4Y16_to_SD),
    .to_SF(Tile_X4Y16_to_SF),
    .to_SG(Tile_X4Y16_to_SG),
    .to_SH(Tile_X4Y16_to_SH),
    .to_SI(Tile_X4Y16_to_SI),
    .F_masked1(Tile_X4Y16_F_masked1),
    .F_masked2(Tile_X4Y16_F_masked2),
    .UserCLK(Tile_X4Y17_UserCLKo),
    .UserCLKo(Tile_X4Y16_UserCLKo),
    .rst(Tile_X4Y17_rsto),
    .rsto(Tile_X4Y16_rsto),
    .FrameData(Tile_X3Y16_FrameData_O),
    .FrameData_O(Tile_X4Y16_FrameData_O),
    .FrameStrobe(Tile_X4Y17_FrameStrobe_O),
    .FrameStrobe_O(Tile_X4Y16_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X5Y16_Emulate_Bitstream)
    )
`endif
    Tile_X5Y16_linear_LMDPL
    (
    .from_NA(Tile_X5Y17_to_NA),
    .from_NB(Tile_X5Y17_to_NB),
    .from_NC(Tile_X5Y17_to_NC),
    .from_ND(Tile_X5Y17_to_ND),
    .from_NF(Tile_X5Y17_to_NF),
    .from_NG(Tile_X5Y17_to_NG),
    .from_NH(Tile_X5Y17_to_NH),
    .from_NI(Tile_X5Y17_to_NI),
    .from_EA(Tile_X4Y16_to_EA),
    .from_EB(Tile_X4Y16_to_EB),
    .from_EC(Tile_X4Y16_to_EC),
    .from_ED(Tile_X4Y16_to_ED),
    .from_EF(Tile_X4Y16_to_EF),
    .from_EG(Tile_X4Y16_to_EG),
    .from_EH(Tile_X4Y16_to_EH),
    .from_EI(Tile_X4Y16_to_EI),
    .from_SA(Tile_X5Y15_to_SA),
    .from_SB(Tile_X5Y15_to_SB),
    .from_SC(Tile_X5Y15_to_SC),
    .from_SD(Tile_X5Y15_to_SD),
    .from_SF(Tile_X5Y15_to_SF),
    .from_SG(Tile_X5Y15_to_SG),
    .from_SH(Tile_X5Y15_to_SH),
    .from_SI(Tile_X5Y15_to_SI),
    .from_WA(Tile_X6Y16_to_WA),
    .from_WB(Tile_X6Y16_to_WB),
    .from_WC(Tile_X6Y16_to_WC),
    .from_WD(Tile_X6Y16_to_WD),
    .from_WF(Tile_X6Y16_to_WF),
    .from_WG(Tile_X6Y16_to_WG),
    .from_WH(Tile_X6Y16_to_WH),
    .from_WI(Tile_X6Y16_to_WI),
    .to_EA(Tile_X5Y16_to_EA),
    .to_EB(Tile_X5Y16_to_EB),
    .to_EC(Tile_X5Y16_to_EC),
    .to_ED(Tile_X5Y16_to_ED),
    .to_EF(Tile_X5Y16_to_EF),
    .to_EG(Tile_X5Y16_to_EG),
    .to_EH(Tile_X5Y16_to_EH),
    .to_EI(Tile_X5Y16_to_EI),
    .to_WA(Tile_X5Y16_to_WA),
    .to_WB(Tile_X5Y16_to_WB),
    .to_WC(Tile_X5Y16_to_WC),
    .to_WD(Tile_X5Y16_to_WD),
    .to_WF(Tile_X5Y16_to_WF),
    .to_WG(Tile_X5Y16_to_WG),
    .to_WH(Tile_X5Y16_to_WH),
    .to_WI(Tile_X5Y16_to_WI),
    .to_NA(Tile_X5Y16_to_NA),
    .to_NB(Tile_X5Y16_to_NB),
    .to_NC(Tile_X5Y16_to_NC),
    .to_ND(Tile_X5Y16_to_ND),
    .to_NF(Tile_X5Y16_to_NF),
    .to_NG(Tile_X5Y16_to_NG),
    .to_NH(Tile_X5Y16_to_NH),
    .to_NI(Tile_X5Y16_to_NI),
    .to_SA(Tile_X5Y16_to_SA),
    .to_SB(Tile_X5Y16_to_SB),
    .to_SC(Tile_X5Y16_to_SC),
    .to_SD(Tile_X5Y16_to_SD),
    .to_SF(Tile_X5Y16_to_SF),
    .to_SG(Tile_X5Y16_to_SG),
    .to_SH(Tile_X5Y16_to_SH),
    .to_SI(Tile_X5Y16_to_SI),
    .F_masked1(Tile_X5Y16_F_masked1),
    .F_masked2(Tile_X5Y16_F_masked2),
    .UserCLK(Tile_X5Y17_UserCLKo),
    .UserCLKo(Tile_X5Y16_UserCLKo),
    .rst(Tile_X5Y17_rsto),
    .rsto(Tile_X5Y16_rsto),
    .FrameData(Tile_X4Y16_FrameData_O),
    .FrameData_O(Tile_X5Y16_FrameData_O),
    .FrameStrobe(Tile_X5Y17_FrameStrobe_O),
    .FrameStrobe_O(Tile_X5Y16_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
nonlinear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X6Y16_Emulate_Bitstream)
    )
`endif
    Tile_X6Y16_nonlinear_LMDPL
    (
    .from_NA(Tile_X6Y17_to_NA),
    .from_NB(Tile_X6Y17_to_NB),
    .from_NC(Tile_X6Y17_to_NC),
    .from_ND(Tile_X6Y17_to_ND),
    .from_NF(Tile_X6Y17_to_NF),
    .from_NG(Tile_X6Y17_to_NG),
    .from_NH(Tile_X6Y17_to_NH),
    .from_NI(Tile_X6Y17_to_NI),
    .from_EA(Tile_X5Y16_to_EA),
    .from_EB(Tile_X5Y16_to_EB),
    .from_EC(Tile_X5Y16_to_EC),
    .from_ED(Tile_X5Y16_to_ED),
    .from_EF(Tile_X5Y16_to_EF),
    .from_EG(Tile_X5Y16_to_EG),
    .from_EH(Tile_X5Y16_to_EH),
    .from_EI(Tile_X5Y16_to_EI),
    .from_SA(Tile_X6Y15_to_SA),
    .from_SB(Tile_X6Y15_to_SB),
    .from_SC(Tile_X6Y15_to_SC),
    .from_SD(Tile_X6Y15_to_SD),
    .from_SF(Tile_X6Y15_to_SF),
    .from_SG(Tile_X6Y15_to_SG),
    .from_SH(Tile_X6Y15_to_SH),
    .from_SI(Tile_X6Y15_to_SI),
    .from_WA(Tile_X7Y16_to_WA),
    .from_WB(Tile_X7Y16_to_WB),
    .from_WC(Tile_X7Y16_to_WC),
    .from_WD(Tile_X7Y16_to_WD),
    .from_WF(Tile_X7Y16_to_WF),
    .from_WG(Tile_X7Y16_to_WG),
    .from_WH(Tile_X7Y16_to_WH),
    .from_WI(Tile_X7Y16_to_WI),
    .to_EA(Tile_X6Y16_to_EA),
    .to_EB(Tile_X6Y16_to_EB),
    .to_EC(Tile_X6Y16_to_EC),
    .to_ED(Tile_X6Y16_to_ED),
    .to_EF(Tile_X6Y16_to_EF),
    .to_EG(Tile_X6Y16_to_EG),
    .to_EH(Tile_X6Y16_to_EH),
    .to_EI(Tile_X6Y16_to_EI),
    .to_WA(Tile_X6Y16_to_WA),
    .to_WB(Tile_X6Y16_to_WB),
    .to_WC(Tile_X6Y16_to_WC),
    .to_WD(Tile_X6Y16_to_WD),
    .to_WF(Tile_X6Y16_to_WF),
    .to_WG(Tile_X6Y16_to_WG),
    .to_WH(Tile_X6Y16_to_WH),
    .to_WI(Tile_X6Y16_to_WI),
    .to_NA(Tile_X6Y16_to_NA),
    .to_NB(Tile_X6Y16_to_NB),
    .to_NC(Tile_X6Y16_to_NC),
    .to_ND(Tile_X6Y16_to_ND),
    .to_NF(Tile_X6Y16_to_NF),
    .to_NG(Tile_X6Y16_to_NG),
    .to_NH(Tile_X6Y16_to_NH),
    .to_NI(Tile_X6Y16_to_NI),
    .to_SA(Tile_X6Y16_to_SA),
    .to_SB(Tile_X6Y16_to_SB),
    .to_SC(Tile_X6Y16_to_SC),
    .to_SD(Tile_X6Y16_to_SD),
    .to_SF(Tile_X6Y16_to_SF),
    .to_SG(Tile_X6Y16_to_SG),
    .to_SH(Tile_X6Y16_to_SH),
    .to_SI(Tile_X6Y16_to_SI),
    .R_t(Tile_X6Y16_R_t),
    .R_f(Tile_X6Y16_R_f),
    .F_masked1(Tile_X6Y16_F_masked1),
    .F_masked2(Tile_X6Y16_F_masked2),
    .UserCLK(Tile_X6Y17_UserCLKo),
    .UserCLKo(Tile_X6Y16_UserCLKo),
    .rst(Tile_X6Y17_rsto),
    .rsto(Tile_X6Y16_rsto),
    .FrameData(Tile_X5Y16_FrameData_O),
    .FrameData_O(Tile_X6Y16_FrameData_O),
    .FrameStrobe(Tile_X6Y17_FrameStrobe_O),
    .FrameStrobe_O(Tile_X6Y16_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X7Y16_Emulate_Bitstream)
    )
`endif
    Tile_X7Y16_linear_LMDPL
    (
    .from_NA(Tile_X7Y17_to_NA),
    .from_NB(Tile_X7Y17_to_NB),
    .from_NC(Tile_X7Y17_to_NC),
    .from_ND(Tile_X7Y17_to_ND),
    .from_NF(Tile_X7Y17_to_NF),
    .from_NG(Tile_X7Y17_to_NG),
    .from_NH(Tile_X7Y17_to_NH),
    .from_NI(Tile_X7Y17_to_NI),
    .from_EA(Tile_X6Y16_to_EA),
    .from_EB(Tile_X6Y16_to_EB),
    .from_EC(Tile_X6Y16_to_EC),
    .from_ED(Tile_X6Y16_to_ED),
    .from_EF(Tile_X6Y16_to_EF),
    .from_EG(Tile_X6Y16_to_EG),
    .from_EH(Tile_X6Y16_to_EH),
    .from_EI(Tile_X6Y16_to_EI),
    .from_SA(Tile_X7Y15_to_SA),
    .from_SB(Tile_X7Y15_to_SB),
    .from_SC(Tile_X7Y15_to_SC),
    .from_SD(Tile_X7Y15_to_SD),
    .from_SF(Tile_X7Y15_to_SF),
    .from_SG(Tile_X7Y15_to_SG),
    .from_SH(Tile_X7Y15_to_SH),
    .from_SI(Tile_X7Y15_to_SI),
    .from_WA(Tile_X8Y16_to_WA),
    .from_WB(Tile_X8Y16_to_WB),
    .from_WC(Tile_X8Y16_to_WC),
    .from_WD(Tile_X8Y16_to_WD),
    .from_WF(Tile_X8Y16_to_WF),
    .from_WG(Tile_X8Y16_to_WG),
    .from_WH(Tile_X8Y16_to_WH),
    .from_WI(Tile_X8Y16_to_WI),
    .to_EA(Tile_X7Y16_to_EA),
    .to_EB(Tile_X7Y16_to_EB),
    .to_EC(Tile_X7Y16_to_EC),
    .to_ED(Tile_X7Y16_to_ED),
    .to_EF(Tile_X7Y16_to_EF),
    .to_EG(Tile_X7Y16_to_EG),
    .to_EH(Tile_X7Y16_to_EH),
    .to_EI(Tile_X7Y16_to_EI),
    .to_WA(Tile_X7Y16_to_WA),
    .to_WB(Tile_X7Y16_to_WB),
    .to_WC(Tile_X7Y16_to_WC),
    .to_WD(Tile_X7Y16_to_WD),
    .to_WF(Tile_X7Y16_to_WF),
    .to_WG(Tile_X7Y16_to_WG),
    .to_WH(Tile_X7Y16_to_WH),
    .to_WI(Tile_X7Y16_to_WI),
    .to_NA(Tile_X7Y16_to_NA),
    .to_NB(Tile_X7Y16_to_NB),
    .to_NC(Tile_X7Y16_to_NC),
    .to_ND(Tile_X7Y16_to_ND),
    .to_NF(Tile_X7Y16_to_NF),
    .to_NG(Tile_X7Y16_to_NG),
    .to_NH(Tile_X7Y16_to_NH),
    .to_NI(Tile_X7Y16_to_NI),
    .to_SA(Tile_X7Y16_to_SA),
    .to_SB(Tile_X7Y16_to_SB),
    .to_SC(Tile_X7Y16_to_SC),
    .to_SD(Tile_X7Y16_to_SD),
    .to_SF(Tile_X7Y16_to_SF),
    .to_SG(Tile_X7Y16_to_SG),
    .to_SH(Tile_X7Y16_to_SH),
    .to_SI(Tile_X7Y16_to_SI),
    .F_masked1(Tile_X7Y16_F_masked1),
    .F_masked2(Tile_X7Y16_F_masked2),
    .UserCLK(Tile_X7Y17_UserCLKo),
    .UserCLKo(Tile_X7Y16_UserCLKo),
    .rst(Tile_X7Y17_rsto),
    .rsto(Tile_X7Y16_rsto),
    .FrameData(Tile_X6Y16_FrameData_O),
    .FrameData_O(Tile_X7Y16_FrameData_O),
    .FrameStrobe(Tile_X7Y17_FrameStrobe_O),
    .FrameStrobe_O(Tile_X7Y16_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
ctrl_to_sec
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X8Y16_Emulate_Bitstream)
    )
`endif
    Tile_X8Y16_ctrl_to_sec
    (
    .from_NA(Tile_X8Y17_to_NA),
    .from_NB(Tile_X8Y17_to_NB),
    .from_NC(Tile_X8Y17_to_NC),
    .from_ND(Tile_X8Y17_to_ND),
    .from_NF(Tile_X8Y17_to_NF),
    .from_NG(Tile_X8Y17_to_NG),
    .from_NH(Tile_X8Y17_to_NH),
    .from_NI(Tile_X8Y17_to_NI),
    .from_EA(Tile_X7Y16_to_EA),
    .from_EB(Tile_X7Y16_to_EB),
    .from_EC(Tile_X7Y16_to_EC),
    .from_ED(Tile_X7Y16_to_ED),
    .from_EF(Tile_X7Y16_to_EF),
    .from_EG(Tile_X7Y16_to_EG),
    .from_EH(Tile_X7Y16_to_EH),
    .from_EI(Tile_X7Y16_to_EI),
    .from_SA(Tile_X8Y15_to_SA),
    .from_SB(Tile_X8Y15_to_SB),
    .from_SC(Tile_X8Y15_to_SC),
    .from_SD(Tile_X8Y15_to_SD),
    .from_SF(Tile_X8Y15_to_SF),
    .from_SG(Tile_X8Y15_to_SG),
    .from_SH(Tile_X8Y15_to_SH),
    .from_SI(Tile_X8Y15_to_SI),
    .from_WA_1s(Tile_X9Y16_to_WA_1s),
    .from_WB_1s(Tile_X9Y16_to_WB_1s),
    .from_WC_1s(Tile_X9Y16_to_WC_1s),
    .from_WD_1s(Tile_X9Y16_to_WD_1s),
    .from_WF_1s(Tile_X9Y16_to_WF_1s),
    .from_WG_1s(Tile_X9Y16_to_WG_1s),
    .from_WH_1s(Tile_X9Y16_to_WH_1s),
    .from_WI_1s(Tile_X9Y16_to_WI_1s),
    .to_WA(Tile_X8Y16_to_WA),
    .to_WB(Tile_X8Y16_to_WB),
    .to_WC(Tile_X8Y16_to_WC),
    .to_WD(Tile_X8Y16_to_WD),
    .to_WF(Tile_X8Y16_to_WF),
    .to_WG(Tile_X8Y16_to_WG),
    .to_WH(Tile_X8Y16_to_WH),
    .to_WI(Tile_X8Y16_to_WI),
    .to_NA(Tile_X8Y16_to_NA),
    .to_NB(Tile_X8Y16_to_NB),
    .to_NC(Tile_X8Y16_to_NC),
    .to_ND(Tile_X8Y16_to_ND),
    .to_NF(Tile_X8Y16_to_NF),
    .to_NG(Tile_X8Y16_to_NG),
    .to_NH(Tile_X8Y16_to_NH),
    .to_NI(Tile_X8Y16_to_NI),
    .to_SA(Tile_X8Y16_to_SA),
    .to_SB(Tile_X8Y16_to_SB),
    .to_SC(Tile_X8Y16_to_SC),
    .to_SD(Tile_X8Y16_to_SD),
    .to_SF(Tile_X8Y16_to_SF),
    .to_SG(Tile_X8Y16_to_SG),
    .to_SH(Tile_X8Y16_to_SH),
    .to_SI(Tile_X8Y16_to_SI),
    .UserCLK(Tile_X8Y17_UserCLKo),
    .UserCLKo(Tile_X8Y16_UserCLKo),
    .rst(Tile_X8Y17_rsto),
    .rsto(Tile_X8Y16_rsto),
    .FrameData(Tile_X7Y16_FrameData_O),
    .FrameData_O(Tile_X8Y16_FrameData_O),
    .FrameStrobe(Tile_X8Y17_FrameStrobe_O),
    .FrameStrobe_O(Tile_X8Y16_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
combined_WDDL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X9Y16_Emulate_Bitstream)
    )
`endif
    Tile_X9Y16_combined_WDDL
    (
    .from_NA_1s(Tile_X9Y17_to_NA_1s),
    .from_NB_1s(Tile_X9Y17_to_NB_1s),
    .from_NC_1s(Tile_X9Y17_to_NC_1s),
    .from_ND_1s(Tile_X9Y17_to_ND_1s),
    .from_NF_1s(Tile_X9Y17_to_NF_1s),
    .from_NG_1s(Tile_X9Y17_to_NG_1s),
    .from_NH_1s(Tile_X9Y17_to_NH_1s),
    .from_NI_1s(Tile_X9Y17_to_NI_1s),
    .from_SA_1s(Tile_X9Y15_to_SA_1s),
    .from_SB_1s(Tile_X9Y15_to_SB_1s),
    .from_SC_1s(Tile_X9Y15_to_SC_1s),
    .from_SD_1s(Tile_X9Y15_to_SD_1s),
    .from_SF_1s(Tile_X9Y15_to_SF_1s),
    .from_SG_1s(Tile_X9Y15_to_SG_1s),
    .from_SH_1s(Tile_X9Y15_to_SH_1s),
    .from_SI_1s(Tile_X9Y15_to_SI_1s),
    .from_WA_1s(Tile_X10Y16_to_WA_1s),
    .from_WB_1s(Tile_X10Y16_to_WB_1s),
    .from_WC_1s(Tile_X10Y16_to_WC_1s),
    .from_WD_1s(Tile_X10Y16_to_WD_1s),
    .from_WF_1s(Tile_X10Y16_to_WF_1s),
    .from_WG_1s(Tile_X10Y16_to_WG_1s),
    .from_WH_1s(Tile_X10Y16_to_WH_1s),
    .from_WI_1s(Tile_X10Y16_to_WI_1s),
    .to_EA_1s(Tile_X9Y16_to_EA_1s),
    .to_EB_1s(Tile_X9Y16_to_EB_1s),
    .to_EC_1s(Tile_X9Y16_to_EC_1s),
    .to_ED_1s(Tile_X9Y16_to_ED_1s),
    .to_EF_1s(Tile_X9Y16_to_EF_1s),
    .to_EG_1s(Tile_X9Y16_to_EG_1s),
    .to_EH_1s(Tile_X9Y16_to_EH_1s),
    .to_EI_1s(Tile_X9Y16_to_EI_1s),
    .to_WA_1s(Tile_X9Y16_to_WA_1s),
    .to_WB_1s(Tile_X9Y16_to_WB_1s),
    .to_WC_1s(Tile_X9Y16_to_WC_1s),
    .to_WD_1s(Tile_X9Y16_to_WD_1s),
    .to_WF_1s(Tile_X9Y16_to_WF_1s),
    .to_WG_1s(Tile_X9Y16_to_WG_1s),
    .to_WH_1s(Tile_X9Y16_to_WH_1s),
    .to_WI_1s(Tile_X9Y16_to_WI_1s),
    .to_NA_1s(Tile_X9Y16_to_NA_1s),
    .to_NB_1s(Tile_X9Y16_to_NB_1s),
    .to_NC_1s(Tile_X9Y16_to_NC_1s),
    .to_ND_1s(Tile_X9Y16_to_ND_1s),
    .to_NF_1s(Tile_X9Y16_to_NF_1s),
    .to_NG_1s(Tile_X9Y16_to_NG_1s),
    .to_NH_1s(Tile_X9Y16_to_NH_1s),
    .to_NI_1s(Tile_X9Y16_to_NI_1s),
    .to_SA_1s(Tile_X9Y16_to_SA_1s),
    .to_SB_1s(Tile_X9Y16_to_SB_1s),
    .to_SC_1s(Tile_X9Y16_to_SC_1s),
    .to_SD_1s(Tile_X9Y16_to_SD_1s),
    .to_SF_1s(Tile_X9Y16_to_SF_1s),
    .to_SG_1s(Tile_X9Y16_to_SG_1s),
    .to_SH_1s(Tile_X9Y16_to_SH_1s),
    .to_SI_1s(Tile_X9Y16_to_SI_1s),
    .F_ctrl(Tile_X9Y16_F_ctrl),
    .UserCLK(Tile_X9Y17_UserCLKo),
    .UserCLKo(Tile_X9Y16_UserCLKo),
    .rst(Tile_X9Y17_rsto),
    .rsto(Tile_X9Y16_rsto),
    .FrameData(Tile_X8Y16_FrameData_O),
    .FrameData_O(Tile_X9Y16_FrameData_O),
    .FrameStrobe(Tile_X9Y17_FrameStrobe_O),
    .FrameStrobe_O(Tile_X9Y16_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
ctrl_IO
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X10Y16_Emulate_Bitstream)
    )
`endif
    Tile_X10Y16_ctrl_IO
    (
    .from_EA_1s(Tile_X9Y16_to_EA_1s),
    .from_EB_1s(Tile_X9Y16_to_EB_1s),
    .from_EC_1s(Tile_X9Y16_to_EC_1s),
    .from_ED_1s(Tile_X9Y16_to_ED_1s),
    .from_EF_1s(Tile_X9Y16_to_EF_1s),
    .from_EG_1s(Tile_X9Y16_to_EG_1s),
    .from_EH_1s(Tile_X9Y16_to_EH_1s),
    .from_EI_1s(Tile_X9Y16_to_EI_1s),
    .to_WA_1s(Tile_X10Y16_to_WA_1s),
    .to_WB_1s(Tile_X10Y16_to_WB_1s),
    .to_WC_1s(Tile_X10Y16_to_WC_1s),
    .to_WD_1s(Tile_X10Y16_to_WD_1s),
    .to_WF_1s(Tile_X10Y16_to_WF_1s),
    .to_WG_1s(Tile_X10Y16_to_WG_1s),
    .to_WH_1s(Tile_X10Y16_to_WH_1s),
    .to_WI_1s(Tile_X10Y16_to_WI_1s),
    .A_O_top_0_t(Tile_X10Y16_A_O_top_0_t),
    .A_O_top_0_f(Tile_X10Y16_A_O_top_0_f),
    .A_prech2(Tile_X10Y16_A_prech2),
    .A_DR_fault(Tile_X10Y16_A_DR_fault),
    .A_I_top_0_t(Tile_X10Y16_A_I_top_0_t),
    .A_I_top_0_f(Tile_X10Y16_A_I_top_0_f),
    .A_T_top(Tile_X10Y16_A_T_top),
    .A_F_ctrl(Tile_X10Y16_A_F_ctrl),
    .UserCLK(Tile_X10Y17_UserCLKo),
    .UserCLKo(Tile_X10Y16_UserCLKo),
    .rst(Tile_X10Y17_rsto),
    .rsto(Tile_X10Y16_rsto),
    .FrameData(Tile_X9Y16_FrameData_O),
    .FrameData_O(Tile_X10Y16_FrameData_O),
    .FrameStrobe(Tile_X10Y17_FrameStrobe_O),
    .FrameStrobe_O(Tile_X10Y16_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
W_IO_custom
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X0Y17_Emulate_Bitstream)
    )
`endif
    Tile_X0Y17_W_IO_custom
    (
    .from_NA(Tile_X0Y18_to_NA),
    .from_NB(Tile_X0Y18_to_NB),
    .from_NC(Tile_X0Y18_to_NC),
    .from_ND(Tile_X0Y18_to_ND),
    .from_NF(Tile_X0Y18_to_NF),
    .from_NG(Tile_X0Y18_to_NG),
    .from_NH(Tile_X0Y18_to_NH),
    .from_NI(Tile_X0Y18_to_NI),
    .from_SA(Tile_X0Y16_to_SA),
    .from_SB(Tile_X0Y16_to_SB),
    .from_SC(Tile_X0Y16_to_SC),
    .from_SD(Tile_X0Y16_to_SD),
    .from_SF(Tile_X0Y16_to_SF),
    .from_SG(Tile_X0Y16_to_SG),
    .from_SH(Tile_X0Y16_to_SH),
    .from_SI(Tile_X0Y16_to_SI),
    .from_WA(Tile_X1Y17_to_WA),
    .from_WB(Tile_X1Y17_to_WB),
    .from_WC(Tile_X1Y17_to_WC),
    .from_WD(Tile_X1Y17_to_WD),
    .from_WF(Tile_X1Y17_to_WF),
    .from_WG(Tile_X1Y17_to_WG),
    .from_WH(Tile_X1Y17_to_WH),
    .from_WI(Tile_X1Y17_to_WI),
    .to_EA(Tile_X0Y17_to_EA),
    .to_EB(Tile_X0Y17_to_EB),
    .to_EC(Tile_X0Y17_to_EC),
    .to_ED(Tile_X0Y17_to_ED),
    .to_EF(Tile_X0Y17_to_EF),
    .to_EG(Tile_X0Y17_to_EG),
    .to_EH(Tile_X0Y17_to_EH),
    .to_EI(Tile_X0Y17_to_EI),
    .to_NA(Tile_X0Y17_to_NA),
    .to_NB(Tile_X0Y17_to_NB),
    .to_NC(Tile_X0Y17_to_NC),
    .to_ND(Tile_X0Y17_to_ND),
    .to_NF(Tile_X0Y17_to_NF),
    .to_NG(Tile_X0Y17_to_NG),
    .to_NH(Tile_X0Y17_to_NH),
    .to_NI(Tile_X0Y17_to_NI),
    .to_SA(Tile_X0Y17_to_SA),
    .to_SB(Tile_X0Y17_to_SB),
    .to_SC(Tile_X0Y17_to_SC),
    .to_SD(Tile_X0Y17_to_SD),
    .to_SF(Tile_X0Y17_to_SF),
    .to_SG(Tile_X0Y17_to_SG),
    .to_SH(Tile_X0Y17_to_SH),
    .to_SI(Tile_X0Y17_to_SI),
    .A_O_top_0_t(Tile_X0Y17_A_O_top_0_t),
    .A_O_top_0_f(Tile_X0Y17_A_O_top_0_f),
    .A_O_top_1_t(Tile_X0Y17_A_O_top_1_t),
    .A_O_top_1_f(Tile_X0Y17_A_O_top_1_f),
    .A_prech1(Tile_X0Y17_A_prech1),
    .A_prech2(Tile_X0Y17_A_prech2),
    .A_DR_fault(Tile_X0Y17_A_DR_fault),
    .A_I_top_0_t(Tile_X0Y17_A_I_top_0_t),
    .A_I_top_0_f(Tile_X0Y17_A_I_top_0_f),
    .A_I_top_1_t(Tile_X0Y17_A_I_top_1_t),
    .A_I_top_1_f(Tile_X0Y17_A_I_top_1_f),
    .A_T_top(Tile_X0Y17_A_T_top),
    .A_F_masked1(Tile_X0Y17_A_F_masked1),
    .A_F_masked2(Tile_X0Y17_A_F_masked2),
    .A_config_C_bit0(Tile_X0Y17_A_config_C_bit0),
    .A_config_C_bit1(Tile_X0Y17_A_config_C_bit1),
    .A_config_C_bit2(Tile_X0Y17_A_config_C_bit2),
    .A_config_C_bit3(Tile_X0Y17_A_config_C_bit3),
    .B_config_C_bit0(Tile_X0Y17_B_config_C_bit0),
    .B_config_C_bit1(Tile_X0Y17_B_config_C_bit1),
    .B_config_C_bit2(Tile_X0Y17_B_config_C_bit2),
    .B_config_C_bit3(Tile_X0Y17_B_config_C_bit3),
    .UserCLK(Tile_X0Y18_UserCLKo),
    .UserCLKo(Tile_X0Y17_UserCLKo),
    .rst(Tile_X0Y18_rsto),
    .rsto(Tile_X0Y17_rsto),
    .FrameData(Tile_Y17_FrameData),
    .FrameData_O(Tile_X0Y17_FrameData_O),
    .FrameStrobe(Tile_X0Y18_FrameStrobe_O),
    .FrameStrobe_O(Tile_X0Y17_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X1Y17_Emulate_Bitstream)
    )
`endif
    Tile_X1Y17_linear_LMDPL
    (
    .from_NA(Tile_X1Y18_to_NA),
    .from_NB(Tile_X1Y18_to_NB),
    .from_NC(Tile_X1Y18_to_NC),
    .from_ND(Tile_X1Y18_to_ND),
    .from_NF(Tile_X1Y18_to_NF),
    .from_NG(Tile_X1Y18_to_NG),
    .from_NH(Tile_X1Y18_to_NH),
    .from_NI(Tile_X1Y18_to_NI),
    .from_EA(Tile_X0Y17_to_EA),
    .from_EB(Tile_X0Y17_to_EB),
    .from_EC(Tile_X0Y17_to_EC),
    .from_ED(Tile_X0Y17_to_ED),
    .from_EF(Tile_X0Y17_to_EF),
    .from_EG(Tile_X0Y17_to_EG),
    .from_EH(Tile_X0Y17_to_EH),
    .from_EI(Tile_X0Y17_to_EI),
    .from_SA(Tile_X1Y16_to_SA),
    .from_SB(Tile_X1Y16_to_SB),
    .from_SC(Tile_X1Y16_to_SC),
    .from_SD(Tile_X1Y16_to_SD),
    .from_SF(Tile_X1Y16_to_SF),
    .from_SG(Tile_X1Y16_to_SG),
    .from_SH(Tile_X1Y16_to_SH),
    .from_SI(Tile_X1Y16_to_SI),
    .from_WA(Tile_X2Y17_to_WA),
    .from_WB(Tile_X2Y17_to_WB),
    .from_WC(Tile_X2Y17_to_WC),
    .from_WD(Tile_X2Y17_to_WD),
    .from_WF(Tile_X2Y17_to_WF),
    .from_WG(Tile_X2Y17_to_WG),
    .from_WH(Tile_X2Y17_to_WH),
    .from_WI(Tile_X2Y17_to_WI),
    .to_EA(Tile_X1Y17_to_EA),
    .to_EB(Tile_X1Y17_to_EB),
    .to_EC(Tile_X1Y17_to_EC),
    .to_ED(Tile_X1Y17_to_ED),
    .to_EF(Tile_X1Y17_to_EF),
    .to_EG(Tile_X1Y17_to_EG),
    .to_EH(Tile_X1Y17_to_EH),
    .to_EI(Tile_X1Y17_to_EI),
    .to_WA(Tile_X1Y17_to_WA),
    .to_WB(Tile_X1Y17_to_WB),
    .to_WC(Tile_X1Y17_to_WC),
    .to_WD(Tile_X1Y17_to_WD),
    .to_WF(Tile_X1Y17_to_WF),
    .to_WG(Tile_X1Y17_to_WG),
    .to_WH(Tile_X1Y17_to_WH),
    .to_WI(Tile_X1Y17_to_WI),
    .to_NA(Tile_X1Y17_to_NA),
    .to_NB(Tile_X1Y17_to_NB),
    .to_NC(Tile_X1Y17_to_NC),
    .to_ND(Tile_X1Y17_to_ND),
    .to_NF(Tile_X1Y17_to_NF),
    .to_NG(Tile_X1Y17_to_NG),
    .to_NH(Tile_X1Y17_to_NH),
    .to_NI(Tile_X1Y17_to_NI),
    .to_SA(Tile_X1Y17_to_SA),
    .to_SB(Tile_X1Y17_to_SB),
    .to_SC(Tile_X1Y17_to_SC),
    .to_SD(Tile_X1Y17_to_SD),
    .to_SF(Tile_X1Y17_to_SF),
    .to_SG(Tile_X1Y17_to_SG),
    .to_SH(Tile_X1Y17_to_SH),
    .to_SI(Tile_X1Y17_to_SI),
    .F_masked1(Tile_X1Y17_F_masked1),
    .F_masked2(Tile_X1Y17_F_masked2),
    .UserCLK(Tile_X1Y18_UserCLKo),
    .UserCLKo(Tile_X1Y17_UserCLKo),
    .rst(Tile_X1Y18_rsto),
    .rsto(Tile_X1Y17_rsto),
    .FrameData(Tile_X0Y17_FrameData_O),
    .FrameData_O(Tile_X1Y17_FrameData_O),
    .FrameStrobe(Tile_X1Y18_FrameStrobe_O),
    .FrameStrobe_O(Tile_X1Y17_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X2Y17_Emulate_Bitstream)
    )
`endif
    Tile_X2Y17_linear_LMDPL
    (
    .from_NA(Tile_X2Y18_to_NA),
    .from_NB(Tile_X2Y18_to_NB),
    .from_NC(Tile_X2Y18_to_NC),
    .from_ND(Tile_X2Y18_to_ND),
    .from_NF(Tile_X2Y18_to_NF),
    .from_NG(Tile_X2Y18_to_NG),
    .from_NH(Tile_X2Y18_to_NH),
    .from_NI(Tile_X2Y18_to_NI),
    .from_EA(Tile_X1Y17_to_EA),
    .from_EB(Tile_X1Y17_to_EB),
    .from_EC(Tile_X1Y17_to_EC),
    .from_ED(Tile_X1Y17_to_ED),
    .from_EF(Tile_X1Y17_to_EF),
    .from_EG(Tile_X1Y17_to_EG),
    .from_EH(Tile_X1Y17_to_EH),
    .from_EI(Tile_X1Y17_to_EI),
    .from_SA(Tile_X2Y16_to_SA),
    .from_SB(Tile_X2Y16_to_SB),
    .from_SC(Tile_X2Y16_to_SC),
    .from_SD(Tile_X2Y16_to_SD),
    .from_SF(Tile_X2Y16_to_SF),
    .from_SG(Tile_X2Y16_to_SG),
    .from_SH(Tile_X2Y16_to_SH),
    .from_SI(Tile_X2Y16_to_SI),
    .from_WA(Tile_X3Y17_to_WA),
    .from_WB(Tile_X3Y17_to_WB),
    .from_WC(Tile_X3Y17_to_WC),
    .from_WD(Tile_X3Y17_to_WD),
    .from_WF(Tile_X3Y17_to_WF),
    .from_WG(Tile_X3Y17_to_WG),
    .from_WH(Tile_X3Y17_to_WH),
    .from_WI(Tile_X3Y17_to_WI),
    .to_EA(Tile_X2Y17_to_EA),
    .to_EB(Tile_X2Y17_to_EB),
    .to_EC(Tile_X2Y17_to_EC),
    .to_ED(Tile_X2Y17_to_ED),
    .to_EF(Tile_X2Y17_to_EF),
    .to_EG(Tile_X2Y17_to_EG),
    .to_EH(Tile_X2Y17_to_EH),
    .to_EI(Tile_X2Y17_to_EI),
    .to_WA(Tile_X2Y17_to_WA),
    .to_WB(Tile_X2Y17_to_WB),
    .to_WC(Tile_X2Y17_to_WC),
    .to_WD(Tile_X2Y17_to_WD),
    .to_WF(Tile_X2Y17_to_WF),
    .to_WG(Tile_X2Y17_to_WG),
    .to_WH(Tile_X2Y17_to_WH),
    .to_WI(Tile_X2Y17_to_WI),
    .to_NA(Tile_X2Y17_to_NA),
    .to_NB(Tile_X2Y17_to_NB),
    .to_NC(Tile_X2Y17_to_NC),
    .to_ND(Tile_X2Y17_to_ND),
    .to_NF(Tile_X2Y17_to_NF),
    .to_NG(Tile_X2Y17_to_NG),
    .to_NH(Tile_X2Y17_to_NH),
    .to_NI(Tile_X2Y17_to_NI),
    .to_SA(Tile_X2Y17_to_SA),
    .to_SB(Tile_X2Y17_to_SB),
    .to_SC(Tile_X2Y17_to_SC),
    .to_SD(Tile_X2Y17_to_SD),
    .to_SF(Tile_X2Y17_to_SF),
    .to_SG(Tile_X2Y17_to_SG),
    .to_SH(Tile_X2Y17_to_SH),
    .to_SI(Tile_X2Y17_to_SI),
    .F_masked1(Tile_X2Y17_F_masked1),
    .F_masked2(Tile_X2Y17_F_masked2),
    .UserCLK(Tile_X2Y18_UserCLKo),
    .UserCLKo(Tile_X2Y17_UserCLKo),
    .rst(Tile_X2Y18_rsto),
    .rsto(Tile_X2Y17_rsto),
    .FrameData(Tile_X1Y17_FrameData_O),
    .FrameData_O(Tile_X2Y17_FrameData_O),
    .FrameStrobe(Tile_X2Y18_FrameStrobe_O),
    .FrameStrobe_O(Tile_X2Y17_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
nonlinear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X3Y17_Emulate_Bitstream)
    )
`endif
    Tile_X3Y17_nonlinear_LMDPL
    (
    .from_NA(Tile_X3Y18_to_NA),
    .from_NB(Tile_X3Y18_to_NB),
    .from_NC(Tile_X3Y18_to_NC),
    .from_ND(Tile_X3Y18_to_ND),
    .from_NF(Tile_X3Y18_to_NF),
    .from_NG(Tile_X3Y18_to_NG),
    .from_NH(Tile_X3Y18_to_NH),
    .from_NI(Tile_X3Y18_to_NI),
    .from_EA(Tile_X2Y17_to_EA),
    .from_EB(Tile_X2Y17_to_EB),
    .from_EC(Tile_X2Y17_to_EC),
    .from_ED(Tile_X2Y17_to_ED),
    .from_EF(Tile_X2Y17_to_EF),
    .from_EG(Tile_X2Y17_to_EG),
    .from_EH(Tile_X2Y17_to_EH),
    .from_EI(Tile_X2Y17_to_EI),
    .from_SA(Tile_X3Y16_to_SA),
    .from_SB(Tile_X3Y16_to_SB),
    .from_SC(Tile_X3Y16_to_SC),
    .from_SD(Tile_X3Y16_to_SD),
    .from_SF(Tile_X3Y16_to_SF),
    .from_SG(Tile_X3Y16_to_SG),
    .from_SH(Tile_X3Y16_to_SH),
    .from_SI(Tile_X3Y16_to_SI),
    .from_WA(Tile_X4Y17_to_WA),
    .from_WB(Tile_X4Y17_to_WB),
    .from_WC(Tile_X4Y17_to_WC),
    .from_WD(Tile_X4Y17_to_WD),
    .from_WF(Tile_X4Y17_to_WF),
    .from_WG(Tile_X4Y17_to_WG),
    .from_WH(Tile_X4Y17_to_WH),
    .from_WI(Tile_X4Y17_to_WI),
    .to_EA(Tile_X3Y17_to_EA),
    .to_EB(Tile_X3Y17_to_EB),
    .to_EC(Tile_X3Y17_to_EC),
    .to_ED(Tile_X3Y17_to_ED),
    .to_EF(Tile_X3Y17_to_EF),
    .to_EG(Tile_X3Y17_to_EG),
    .to_EH(Tile_X3Y17_to_EH),
    .to_EI(Tile_X3Y17_to_EI),
    .to_WA(Tile_X3Y17_to_WA),
    .to_WB(Tile_X3Y17_to_WB),
    .to_WC(Tile_X3Y17_to_WC),
    .to_WD(Tile_X3Y17_to_WD),
    .to_WF(Tile_X3Y17_to_WF),
    .to_WG(Tile_X3Y17_to_WG),
    .to_WH(Tile_X3Y17_to_WH),
    .to_WI(Tile_X3Y17_to_WI),
    .to_NA(Tile_X3Y17_to_NA),
    .to_NB(Tile_X3Y17_to_NB),
    .to_NC(Tile_X3Y17_to_NC),
    .to_ND(Tile_X3Y17_to_ND),
    .to_NF(Tile_X3Y17_to_NF),
    .to_NG(Tile_X3Y17_to_NG),
    .to_NH(Tile_X3Y17_to_NH),
    .to_NI(Tile_X3Y17_to_NI),
    .to_SA(Tile_X3Y17_to_SA),
    .to_SB(Tile_X3Y17_to_SB),
    .to_SC(Tile_X3Y17_to_SC),
    .to_SD(Tile_X3Y17_to_SD),
    .to_SF(Tile_X3Y17_to_SF),
    .to_SG(Tile_X3Y17_to_SG),
    .to_SH(Tile_X3Y17_to_SH),
    .to_SI(Tile_X3Y17_to_SI),
    .R_t(Tile_X3Y17_R_t),
    .R_f(Tile_X3Y17_R_f),
    .F_masked1(Tile_X3Y17_F_masked1),
    .F_masked2(Tile_X3Y17_F_masked2),
    .UserCLK(Tile_X3Y18_UserCLKo),
    .UserCLKo(Tile_X3Y17_UserCLKo),
    .rst(Tile_X3Y18_rsto),
    .rsto(Tile_X3Y17_rsto),
    .FrameData(Tile_X2Y17_FrameData_O),
    .FrameData_O(Tile_X3Y17_FrameData_O),
    .FrameStrobe(Tile_X3Y18_FrameStrobe_O),
    .FrameStrobe_O(Tile_X3Y17_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X4Y17_Emulate_Bitstream)
    )
`endif
    Tile_X4Y17_linear_LMDPL
    (
    .from_NA(Tile_X4Y18_to_NA),
    .from_NB(Tile_X4Y18_to_NB),
    .from_NC(Tile_X4Y18_to_NC),
    .from_ND(Tile_X4Y18_to_ND),
    .from_NF(Tile_X4Y18_to_NF),
    .from_NG(Tile_X4Y18_to_NG),
    .from_NH(Tile_X4Y18_to_NH),
    .from_NI(Tile_X4Y18_to_NI),
    .from_EA(Tile_X3Y17_to_EA),
    .from_EB(Tile_X3Y17_to_EB),
    .from_EC(Tile_X3Y17_to_EC),
    .from_ED(Tile_X3Y17_to_ED),
    .from_EF(Tile_X3Y17_to_EF),
    .from_EG(Tile_X3Y17_to_EG),
    .from_EH(Tile_X3Y17_to_EH),
    .from_EI(Tile_X3Y17_to_EI),
    .from_SA(Tile_X4Y16_to_SA),
    .from_SB(Tile_X4Y16_to_SB),
    .from_SC(Tile_X4Y16_to_SC),
    .from_SD(Tile_X4Y16_to_SD),
    .from_SF(Tile_X4Y16_to_SF),
    .from_SG(Tile_X4Y16_to_SG),
    .from_SH(Tile_X4Y16_to_SH),
    .from_SI(Tile_X4Y16_to_SI),
    .from_WA(Tile_X5Y17_to_WA),
    .from_WB(Tile_X5Y17_to_WB),
    .from_WC(Tile_X5Y17_to_WC),
    .from_WD(Tile_X5Y17_to_WD),
    .from_WF(Tile_X5Y17_to_WF),
    .from_WG(Tile_X5Y17_to_WG),
    .from_WH(Tile_X5Y17_to_WH),
    .from_WI(Tile_X5Y17_to_WI),
    .to_EA(Tile_X4Y17_to_EA),
    .to_EB(Tile_X4Y17_to_EB),
    .to_EC(Tile_X4Y17_to_EC),
    .to_ED(Tile_X4Y17_to_ED),
    .to_EF(Tile_X4Y17_to_EF),
    .to_EG(Tile_X4Y17_to_EG),
    .to_EH(Tile_X4Y17_to_EH),
    .to_EI(Tile_X4Y17_to_EI),
    .to_WA(Tile_X4Y17_to_WA),
    .to_WB(Tile_X4Y17_to_WB),
    .to_WC(Tile_X4Y17_to_WC),
    .to_WD(Tile_X4Y17_to_WD),
    .to_WF(Tile_X4Y17_to_WF),
    .to_WG(Tile_X4Y17_to_WG),
    .to_WH(Tile_X4Y17_to_WH),
    .to_WI(Tile_X4Y17_to_WI),
    .to_NA(Tile_X4Y17_to_NA),
    .to_NB(Tile_X4Y17_to_NB),
    .to_NC(Tile_X4Y17_to_NC),
    .to_ND(Tile_X4Y17_to_ND),
    .to_NF(Tile_X4Y17_to_NF),
    .to_NG(Tile_X4Y17_to_NG),
    .to_NH(Tile_X4Y17_to_NH),
    .to_NI(Tile_X4Y17_to_NI),
    .to_SA(Tile_X4Y17_to_SA),
    .to_SB(Tile_X4Y17_to_SB),
    .to_SC(Tile_X4Y17_to_SC),
    .to_SD(Tile_X4Y17_to_SD),
    .to_SF(Tile_X4Y17_to_SF),
    .to_SG(Tile_X4Y17_to_SG),
    .to_SH(Tile_X4Y17_to_SH),
    .to_SI(Tile_X4Y17_to_SI),
    .F_masked1(Tile_X4Y17_F_masked1),
    .F_masked2(Tile_X4Y17_F_masked2),
    .UserCLK(Tile_X4Y18_UserCLKo),
    .UserCLKo(Tile_X4Y17_UserCLKo),
    .rst(Tile_X4Y18_rsto),
    .rsto(Tile_X4Y17_rsto),
    .FrameData(Tile_X3Y17_FrameData_O),
    .FrameData_O(Tile_X4Y17_FrameData_O),
    .FrameStrobe(Tile_X4Y18_FrameStrobe_O),
    .FrameStrobe_O(Tile_X4Y17_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X5Y17_Emulate_Bitstream)
    )
`endif
    Tile_X5Y17_linear_LMDPL
    (
    .from_NA(Tile_X5Y18_to_NA),
    .from_NB(Tile_X5Y18_to_NB),
    .from_NC(Tile_X5Y18_to_NC),
    .from_ND(Tile_X5Y18_to_ND),
    .from_NF(Tile_X5Y18_to_NF),
    .from_NG(Tile_X5Y18_to_NG),
    .from_NH(Tile_X5Y18_to_NH),
    .from_NI(Tile_X5Y18_to_NI),
    .from_EA(Tile_X4Y17_to_EA),
    .from_EB(Tile_X4Y17_to_EB),
    .from_EC(Tile_X4Y17_to_EC),
    .from_ED(Tile_X4Y17_to_ED),
    .from_EF(Tile_X4Y17_to_EF),
    .from_EG(Tile_X4Y17_to_EG),
    .from_EH(Tile_X4Y17_to_EH),
    .from_EI(Tile_X4Y17_to_EI),
    .from_SA(Tile_X5Y16_to_SA),
    .from_SB(Tile_X5Y16_to_SB),
    .from_SC(Tile_X5Y16_to_SC),
    .from_SD(Tile_X5Y16_to_SD),
    .from_SF(Tile_X5Y16_to_SF),
    .from_SG(Tile_X5Y16_to_SG),
    .from_SH(Tile_X5Y16_to_SH),
    .from_SI(Tile_X5Y16_to_SI),
    .from_WA(Tile_X6Y17_to_WA),
    .from_WB(Tile_X6Y17_to_WB),
    .from_WC(Tile_X6Y17_to_WC),
    .from_WD(Tile_X6Y17_to_WD),
    .from_WF(Tile_X6Y17_to_WF),
    .from_WG(Tile_X6Y17_to_WG),
    .from_WH(Tile_X6Y17_to_WH),
    .from_WI(Tile_X6Y17_to_WI),
    .to_EA(Tile_X5Y17_to_EA),
    .to_EB(Tile_X5Y17_to_EB),
    .to_EC(Tile_X5Y17_to_EC),
    .to_ED(Tile_X5Y17_to_ED),
    .to_EF(Tile_X5Y17_to_EF),
    .to_EG(Tile_X5Y17_to_EG),
    .to_EH(Tile_X5Y17_to_EH),
    .to_EI(Tile_X5Y17_to_EI),
    .to_WA(Tile_X5Y17_to_WA),
    .to_WB(Tile_X5Y17_to_WB),
    .to_WC(Tile_X5Y17_to_WC),
    .to_WD(Tile_X5Y17_to_WD),
    .to_WF(Tile_X5Y17_to_WF),
    .to_WG(Tile_X5Y17_to_WG),
    .to_WH(Tile_X5Y17_to_WH),
    .to_WI(Tile_X5Y17_to_WI),
    .to_NA(Tile_X5Y17_to_NA),
    .to_NB(Tile_X5Y17_to_NB),
    .to_NC(Tile_X5Y17_to_NC),
    .to_ND(Tile_X5Y17_to_ND),
    .to_NF(Tile_X5Y17_to_NF),
    .to_NG(Tile_X5Y17_to_NG),
    .to_NH(Tile_X5Y17_to_NH),
    .to_NI(Tile_X5Y17_to_NI),
    .to_SA(Tile_X5Y17_to_SA),
    .to_SB(Tile_X5Y17_to_SB),
    .to_SC(Tile_X5Y17_to_SC),
    .to_SD(Tile_X5Y17_to_SD),
    .to_SF(Tile_X5Y17_to_SF),
    .to_SG(Tile_X5Y17_to_SG),
    .to_SH(Tile_X5Y17_to_SH),
    .to_SI(Tile_X5Y17_to_SI),
    .F_masked1(Tile_X5Y17_F_masked1),
    .F_masked2(Tile_X5Y17_F_masked2),
    .UserCLK(Tile_X5Y18_UserCLKo),
    .UserCLKo(Tile_X5Y17_UserCLKo),
    .rst(Tile_X5Y18_rsto),
    .rsto(Tile_X5Y17_rsto),
    .FrameData(Tile_X4Y17_FrameData_O),
    .FrameData_O(Tile_X5Y17_FrameData_O),
    .FrameStrobe(Tile_X5Y18_FrameStrobe_O),
    .FrameStrobe_O(Tile_X5Y17_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
nonlinear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X6Y17_Emulate_Bitstream)
    )
`endif
    Tile_X6Y17_nonlinear_LMDPL
    (
    .from_NA(Tile_X6Y18_to_NA),
    .from_NB(Tile_X6Y18_to_NB),
    .from_NC(Tile_X6Y18_to_NC),
    .from_ND(Tile_X6Y18_to_ND),
    .from_NF(Tile_X6Y18_to_NF),
    .from_NG(Tile_X6Y18_to_NG),
    .from_NH(Tile_X6Y18_to_NH),
    .from_NI(Tile_X6Y18_to_NI),
    .from_EA(Tile_X5Y17_to_EA),
    .from_EB(Tile_X5Y17_to_EB),
    .from_EC(Tile_X5Y17_to_EC),
    .from_ED(Tile_X5Y17_to_ED),
    .from_EF(Tile_X5Y17_to_EF),
    .from_EG(Tile_X5Y17_to_EG),
    .from_EH(Tile_X5Y17_to_EH),
    .from_EI(Tile_X5Y17_to_EI),
    .from_SA(Tile_X6Y16_to_SA),
    .from_SB(Tile_X6Y16_to_SB),
    .from_SC(Tile_X6Y16_to_SC),
    .from_SD(Tile_X6Y16_to_SD),
    .from_SF(Tile_X6Y16_to_SF),
    .from_SG(Tile_X6Y16_to_SG),
    .from_SH(Tile_X6Y16_to_SH),
    .from_SI(Tile_X6Y16_to_SI),
    .from_WA(Tile_X7Y17_to_WA),
    .from_WB(Tile_X7Y17_to_WB),
    .from_WC(Tile_X7Y17_to_WC),
    .from_WD(Tile_X7Y17_to_WD),
    .from_WF(Tile_X7Y17_to_WF),
    .from_WG(Tile_X7Y17_to_WG),
    .from_WH(Tile_X7Y17_to_WH),
    .from_WI(Tile_X7Y17_to_WI),
    .to_EA(Tile_X6Y17_to_EA),
    .to_EB(Tile_X6Y17_to_EB),
    .to_EC(Tile_X6Y17_to_EC),
    .to_ED(Tile_X6Y17_to_ED),
    .to_EF(Tile_X6Y17_to_EF),
    .to_EG(Tile_X6Y17_to_EG),
    .to_EH(Tile_X6Y17_to_EH),
    .to_EI(Tile_X6Y17_to_EI),
    .to_WA(Tile_X6Y17_to_WA),
    .to_WB(Tile_X6Y17_to_WB),
    .to_WC(Tile_X6Y17_to_WC),
    .to_WD(Tile_X6Y17_to_WD),
    .to_WF(Tile_X6Y17_to_WF),
    .to_WG(Tile_X6Y17_to_WG),
    .to_WH(Tile_X6Y17_to_WH),
    .to_WI(Tile_X6Y17_to_WI),
    .to_NA(Tile_X6Y17_to_NA),
    .to_NB(Tile_X6Y17_to_NB),
    .to_NC(Tile_X6Y17_to_NC),
    .to_ND(Tile_X6Y17_to_ND),
    .to_NF(Tile_X6Y17_to_NF),
    .to_NG(Tile_X6Y17_to_NG),
    .to_NH(Tile_X6Y17_to_NH),
    .to_NI(Tile_X6Y17_to_NI),
    .to_SA(Tile_X6Y17_to_SA),
    .to_SB(Tile_X6Y17_to_SB),
    .to_SC(Tile_X6Y17_to_SC),
    .to_SD(Tile_X6Y17_to_SD),
    .to_SF(Tile_X6Y17_to_SF),
    .to_SG(Tile_X6Y17_to_SG),
    .to_SH(Tile_X6Y17_to_SH),
    .to_SI(Tile_X6Y17_to_SI),
    .R_t(Tile_X6Y17_R_t),
    .R_f(Tile_X6Y17_R_f),
    .F_masked1(Tile_X6Y17_F_masked1),
    .F_masked2(Tile_X6Y17_F_masked2),
    .UserCLK(Tile_X6Y18_UserCLKo),
    .UserCLKo(Tile_X6Y17_UserCLKo),
    .rst(Tile_X6Y18_rsto),
    .rsto(Tile_X6Y17_rsto),
    .FrameData(Tile_X5Y17_FrameData_O),
    .FrameData_O(Tile_X6Y17_FrameData_O),
    .FrameStrobe(Tile_X6Y18_FrameStrobe_O),
    .FrameStrobe_O(Tile_X6Y17_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X7Y17_Emulate_Bitstream)
    )
`endif
    Tile_X7Y17_linear_LMDPL
    (
    .from_NA(Tile_X7Y18_to_NA),
    .from_NB(Tile_X7Y18_to_NB),
    .from_NC(Tile_X7Y18_to_NC),
    .from_ND(Tile_X7Y18_to_ND),
    .from_NF(Tile_X7Y18_to_NF),
    .from_NG(Tile_X7Y18_to_NG),
    .from_NH(Tile_X7Y18_to_NH),
    .from_NI(Tile_X7Y18_to_NI),
    .from_EA(Tile_X6Y17_to_EA),
    .from_EB(Tile_X6Y17_to_EB),
    .from_EC(Tile_X6Y17_to_EC),
    .from_ED(Tile_X6Y17_to_ED),
    .from_EF(Tile_X6Y17_to_EF),
    .from_EG(Tile_X6Y17_to_EG),
    .from_EH(Tile_X6Y17_to_EH),
    .from_EI(Tile_X6Y17_to_EI),
    .from_SA(Tile_X7Y16_to_SA),
    .from_SB(Tile_X7Y16_to_SB),
    .from_SC(Tile_X7Y16_to_SC),
    .from_SD(Tile_X7Y16_to_SD),
    .from_SF(Tile_X7Y16_to_SF),
    .from_SG(Tile_X7Y16_to_SG),
    .from_SH(Tile_X7Y16_to_SH),
    .from_SI(Tile_X7Y16_to_SI),
    .from_WA(Tile_X8Y17_to_WA),
    .from_WB(Tile_X8Y17_to_WB),
    .from_WC(Tile_X8Y17_to_WC),
    .from_WD(Tile_X8Y17_to_WD),
    .from_WF(Tile_X8Y17_to_WF),
    .from_WG(Tile_X8Y17_to_WG),
    .from_WH(Tile_X8Y17_to_WH),
    .from_WI(Tile_X8Y17_to_WI),
    .to_EA(Tile_X7Y17_to_EA),
    .to_EB(Tile_X7Y17_to_EB),
    .to_EC(Tile_X7Y17_to_EC),
    .to_ED(Tile_X7Y17_to_ED),
    .to_EF(Tile_X7Y17_to_EF),
    .to_EG(Tile_X7Y17_to_EG),
    .to_EH(Tile_X7Y17_to_EH),
    .to_EI(Tile_X7Y17_to_EI),
    .to_WA(Tile_X7Y17_to_WA),
    .to_WB(Tile_X7Y17_to_WB),
    .to_WC(Tile_X7Y17_to_WC),
    .to_WD(Tile_X7Y17_to_WD),
    .to_WF(Tile_X7Y17_to_WF),
    .to_WG(Tile_X7Y17_to_WG),
    .to_WH(Tile_X7Y17_to_WH),
    .to_WI(Tile_X7Y17_to_WI),
    .to_NA(Tile_X7Y17_to_NA),
    .to_NB(Tile_X7Y17_to_NB),
    .to_NC(Tile_X7Y17_to_NC),
    .to_ND(Tile_X7Y17_to_ND),
    .to_NF(Tile_X7Y17_to_NF),
    .to_NG(Tile_X7Y17_to_NG),
    .to_NH(Tile_X7Y17_to_NH),
    .to_NI(Tile_X7Y17_to_NI),
    .to_SA(Tile_X7Y17_to_SA),
    .to_SB(Tile_X7Y17_to_SB),
    .to_SC(Tile_X7Y17_to_SC),
    .to_SD(Tile_X7Y17_to_SD),
    .to_SF(Tile_X7Y17_to_SF),
    .to_SG(Tile_X7Y17_to_SG),
    .to_SH(Tile_X7Y17_to_SH),
    .to_SI(Tile_X7Y17_to_SI),
    .F_masked1(Tile_X7Y17_F_masked1),
    .F_masked2(Tile_X7Y17_F_masked2),
    .UserCLK(Tile_X7Y18_UserCLKo),
    .UserCLKo(Tile_X7Y17_UserCLKo),
    .rst(Tile_X7Y18_rsto),
    .rsto(Tile_X7Y17_rsto),
    .FrameData(Tile_X6Y17_FrameData_O),
    .FrameData_O(Tile_X7Y17_FrameData_O),
    .FrameStrobe(Tile_X7Y18_FrameStrobe_O),
    .FrameStrobe_O(Tile_X7Y17_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
ctrl_to_sec
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X8Y17_Emulate_Bitstream)
    )
`endif
    Tile_X8Y17_ctrl_to_sec
    (
    .from_NA(Tile_X8Y18_to_NA),
    .from_NB(Tile_X8Y18_to_NB),
    .from_NC(Tile_X8Y18_to_NC),
    .from_ND(Tile_X8Y18_to_ND),
    .from_NF(Tile_X8Y18_to_NF),
    .from_NG(Tile_X8Y18_to_NG),
    .from_NH(Tile_X8Y18_to_NH),
    .from_NI(Tile_X8Y18_to_NI),
    .from_EA(Tile_X7Y17_to_EA),
    .from_EB(Tile_X7Y17_to_EB),
    .from_EC(Tile_X7Y17_to_EC),
    .from_ED(Tile_X7Y17_to_ED),
    .from_EF(Tile_X7Y17_to_EF),
    .from_EG(Tile_X7Y17_to_EG),
    .from_EH(Tile_X7Y17_to_EH),
    .from_EI(Tile_X7Y17_to_EI),
    .from_SA(Tile_X8Y16_to_SA),
    .from_SB(Tile_X8Y16_to_SB),
    .from_SC(Tile_X8Y16_to_SC),
    .from_SD(Tile_X8Y16_to_SD),
    .from_SF(Tile_X8Y16_to_SF),
    .from_SG(Tile_X8Y16_to_SG),
    .from_SH(Tile_X8Y16_to_SH),
    .from_SI(Tile_X8Y16_to_SI),
    .from_WA_1s(Tile_X9Y17_to_WA_1s),
    .from_WB_1s(Tile_X9Y17_to_WB_1s),
    .from_WC_1s(Tile_X9Y17_to_WC_1s),
    .from_WD_1s(Tile_X9Y17_to_WD_1s),
    .from_WF_1s(Tile_X9Y17_to_WF_1s),
    .from_WG_1s(Tile_X9Y17_to_WG_1s),
    .from_WH_1s(Tile_X9Y17_to_WH_1s),
    .from_WI_1s(Tile_X9Y17_to_WI_1s),
    .to_WA(Tile_X8Y17_to_WA),
    .to_WB(Tile_X8Y17_to_WB),
    .to_WC(Tile_X8Y17_to_WC),
    .to_WD(Tile_X8Y17_to_WD),
    .to_WF(Tile_X8Y17_to_WF),
    .to_WG(Tile_X8Y17_to_WG),
    .to_WH(Tile_X8Y17_to_WH),
    .to_WI(Tile_X8Y17_to_WI),
    .to_NA(Tile_X8Y17_to_NA),
    .to_NB(Tile_X8Y17_to_NB),
    .to_NC(Tile_X8Y17_to_NC),
    .to_ND(Tile_X8Y17_to_ND),
    .to_NF(Tile_X8Y17_to_NF),
    .to_NG(Tile_X8Y17_to_NG),
    .to_NH(Tile_X8Y17_to_NH),
    .to_NI(Tile_X8Y17_to_NI),
    .to_SA(Tile_X8Y17_to_SA),
    .to_SB(Tile_X8Y17_to_SB),
    .to_SC(Tile_X8Y17_to_SC),
    .to_SD(Tile_X8Y17_to_SD),
    .to_SF(Tile_X8Y17_to_SF),
    .to_SG(Tile_X8Y17_to_SG),
    .to_SH(Tile_X8Y17_to_SH),
    .to_SI(Tile_X8Y17_to_SI),
    .UserCLK(Tile_X8Y18_UserCLKo),
    .UserCLKo(Tile_X8Y17_UserCLKo),
    .rst(Tile_X8Y18_rsto),
    .rsto(Tile_X8Y17_rsto),
    .FrameData(Tile_X7Y17_FrameData_O),
    .FrameData_O(Tile_X8Y17_FrameData_O),
    .FrameStrobe(Tile_X8Y18_FrameStrobe_O),
    .FrameStrobe_O(Tile_X8Y17_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
combined_WDDL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X9Y17_Emulate_Bitstream)
    )
`endif
    Tile_X9Y17_combined_WDDL
    (
    .from_NA_1s(Tile_X9Y18_to_NA_1s),
    .from_NB_1s(Tile_X9Y18_to_NB_1s),
    .from_NC_1s(Tile_X9Y18_to_NC_1s),
    .from_ND_1s(Tile_X9Y18_to_ND_1s),
    .from_NF_1s(Tile_X9Y18_to_NF_1s),
    .from_NG_1s(Tile_X9Y18_to_NG_1s),
    .from_NH_1s(Tile_X9Y18_to_NH_1s),
    .from_NI_1s(Tile_X9Y18_to_NI_1s),
    .from_SA_1s(Tile_X9Y16_to_SA_1s),
    .from_SB_1s(Tile_X9Y16_to_SB_1s),
    .from_SC_1s(Tile_X9Y16_to_SC_1s),
    .from_SD_1s(Tile_X9Y16_to_SD_1s),
    .from_SF_1s(Tile_X9Y16_to_SF_1s),
    .from_SG_1s(Tile_X9Y16_to_SG_1s),
    .from_SH_1s(Tile_X9Y16_to_SH_1s),
    .from_SI_1s(Tile_X9Y16_to_SI_1s),
    .from_WA_1s(Tile_X10Y17_to_WA_1s),
    .from_WB_1s(Tile_X10Y17_to_WB_1s),
    .from_WC_1s(Tile_X10Y17_to_WC_1s),
    .from_WD_1s(Tile_X10Y17_to_WD_1s),
    .from_WF_1s(Tile_X10Y17_to_WF_1s),
    .from_WG_1s(Tile_X10Y17_to_WG_1s),
    .from_WH_1s(Tile_X10Y17_to_WH_1s),
    .from_WI_1s(Tile_X10Y17_to_WI_1s),
    .to_EA_1s(Tile_X9Y17_to_EA_1s),
    .to_EB_1s(Tile_X9Y17_to_EB_1s),
    .to_EC_1s(Tile_X9Y17_to_EC_1s),
    .to_ED_1s(Tile_X9Y17_to_ED_1s),
    .to_EF_1s(Tile_X9Y17_to_EF_1s),
    .to_EG_1s(Tile_X9Y17_to_EG_1s),
    .to_EH_1s(Tile_X9Y17_to_EH_1s),
    .to_EI_1s(Tile_X9Y17_to_EI_1s),
    .to_WA_1s(Tile_X9Y17_to_WA_1s),
    .to_WB_1s(Tile_X9Y17_to_WB_1s),
    .to_WC_1s(Tile_X9Y17_to_WC_1s),
    .to_WD_1s(Tile_X9Y17_to_WD_1s),
    .to_WF_1s(Tile_X9Y17_to_WF_1s),
    .to_WG_1s(Tile_X9Y17_to_WG_1s),
    .to_WH_1s(Tile_X9Y17_to_WH_1s),
    .to_WI_1s(Tile_X9Y17_to_WI_1s),
    .to_NA_1s(Tile_X9Y17_to_NA_1s),
    .to_NB_1s(Tile_X9Y17_to_NB_1s),
    .to_NC_1s(Tile_X9Y17_to_NC_1s),
    .to_ND_1s(Tile_X9Y17_to_ND_1s),
    .to_NF_1s(Tile_X9Y17_to_NF_1s),
    .to_NG_1s(Tile_X9Y17_to_NG_1s),
    .to_NH_1s(Tile_X9Y17_to_NH_1s),
    .to_NI_1s(Tile_X9Y17_to_NI_1s),
    .to_SA_1s(Tile_X9Y17_to_SA_1s),
    .to_SB_1s(Tile_X9Y17_to_SB_1s),
    .to_SC_1s(Tile_X9Y17_to_SC_1s),
    .to_SD_1s(Tile_X9Y17_to_SD_1s),
    .to_SF_1s(Tile_X9Y17_to_SF_1s),
    .to_SG_1s(Tile_X9Y17_to_SG_1s),
    .to_SH_1s(Tile_X9Y17_to_SH_1s),
    .to_SI_1s(Tile_X9Y17_to_SI_1s),
    .F_ctrl(Tile_X9Y17_F_ctrl),
    .UserCLK(Tile_X9Y18_UserCLKo),
    .UserCLKo(Tile_X9Y17_UserCLKo),
    .rst(Tile_X9Y18_rsto),
    .rsto(Tile_X9Y17_rsto),
    .FrameData(Tile_X8Y17_FrameData_O),
    .FrameData_O(Tile_X9Y17_FrameData_O),
    .FrameStrobe(Tile_X9Y18_FrameStrobe_O),
    .FrameStrobe_O(Tile_X9Y17_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
ctrl_IO
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X10Y17_Emulate_Bitstream)
    )
`endif
    Tile_X10Y17_ctrl_IO
    (
    .from_EA_1s(Tile_X9Y17_to_EA_1s),
    .from_EB_1s(Tile_X9Y17_to_EB_1s),
    .from_EC_1s(Tile_X9Y17_to_EC_1s),
    .from_ED_1s(Tile_X9Y17_to_ED_1s),
    .from_EF_1s(Tile_X9Y17_to_EF_1s),
    .from_EG_1s(Tile_X9Y17_to_EG_1s),
    .from_EH_1s(Tile_X9Y17_to_EH_1s),
    .from_EI_1s(Tile_X9Y17_to_EI_1s),
    .to_WA_1s(Tile_X10Y17_to_WA_1s),
    .to_WB_1s(Tile_X10Y17_to_WB_1s),
    .to_WC_1s(Tile_X10Y17_to_WC_1s),
    .to_WD_1s(Tile_X10Y17_to_WD_1s),
    .to_WF_1s(Tile_X10Y17_to_WF_1s),
    .to_WG_1s(Tile_X10Y17_to_WG_1s),
    .to_WH_1s(Tile_X10Y17_to_WH_1s),
    .to_WI_1s(Tile_X10Y17_to_WI_1s),
    .A_O_top_0_t(Tile_X10Y17_A_O_top_0_t),
    .A_O_top_0_f(Tile_X10Y17_A_O_top_0_f),
    .A_prech2(Tile_X10Y17_A_prech2),
    .A_DR_fault(Tile_X10Y17_A_DR_fault),
    .A_I_top_0_t(Tile_X10Y17_A_I_top_0_t),
    .A_I_top_0_f(Tile_X10Y17_A_I_top_0_f),
    .A_T_top(Tile_X10Y17_A_T_top),
    .A_F_ctrl(Tile_X10Y17_A_F_ctrl),
    .UserCLK(Tile_X10Y18_UserCLKo),
    .UserCLKo(Tile_X10Y17_UserCLKo),
    .rst(Tile_X10Y18_rsto),
    .rsto(Tile_X10Y17_rsto),
    .FrameData(Tile_X9Y17_FrameData_O),
    .FrameData_O(Tile_X10Y17_FrameData_O),
    .FrameStrobe(Tile_X10Y18_FrameStrobe_O),
    .FrameStrobe_O(Tile_X10Y17_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
W_IO_custom
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X0Y18_Emulate_Bitstream)
    )
`endif
    Tile_X0Y18_W_IO_custom
    (
    .from_NA(Tile_X0Y19_to_NA),
    .from_NB(Tile_X0Y19_to_NB),
    .from_NC(Tile_X0Y19_to_NC),
    .from_ND(Tile_X0Y19_to_ND),
    .from_NF(Tile_X0Y19_to_NF),
    .from_NG(Tile_X0Y19_to_NG),
    .from_NH(Tile_X0Y19_to_NH),
    .from_NI(Tile_X0Y19_to_NI),
    .from_SA(Tile_X0Y17_to_SA),
    .from_SB(Tile_X0Y17_to_SB),
    .from_SC(Tile_X0Y17_to_SC),
    .from_SD(Tile_X0Y17_to_SD),
    .from_SF(Tile_X0Y17_to_SF),
    .from_SG(Tile_X0Y17_to_SG),
    .from_SH(Tile_X0Y17_to_SH),
    .from_SI(Tile_X0Y17_to_SI),
    .from_WA(Tile_X1Y18_to_WA),
    .from_WB(Tile_X1Y18_to_WB),
    .from_WC(Tile_X1Y18_to_WC),
    .from_WD(Tile_X1Y18_to_WD),
    .from_WF(Tile_X1Y18_to_WF),
    .from_WG(Tile_X1Y18_to_WG),
    .from_WH(Tile_X1Y18_to_WH),
    .from_WI(Tile_X1Y18_to_WI),
    .to_EA(Tile_X0Y18_to_EA),
    .to_EB(Tile_X0Y18_to_EB),
    .to_EC(Tile_X0Y18_to_EC),
    .to_ED(Tile_X0Y18_to_ED),
    .to_EF(Tile_X0Y18_to_EF),
    .to_EG(Tile_X0Y18_to_EG),
    .to_EH(Tile_X0Y18_to_EH),
    .to_EI(Tile_X0Y18_to_EI),
    .to_NA(Tile_X0Y18_to_NA),
    .to_NB(Tile_X0Y18_to_NB),
    .to_NC(Tile_X0Y18_to_NC),
    .to_ND(Tile_X0Y18_to_ND),
    .to_NF(Tile_X0Y18_to_NF),
    .to_NG(Tile_X0Y18_to_NG),
    .to_NH(Tile_X0Y18_to_NH),
    .to_NI(Tile_X0Y18_to_NI),
    .to_SA(Tile_X0Y18_to_SA),
    .to_SB(Tile_X0Y18_to_SB),
    .to_SC(Tile_X0Y18_to_SC),
    .to_SD(Tile_X0Y18_to_SD),
    .to_SF(Tile_X0Y18_to_SF),
    .to_SG(Tile_X0Y18_to_SG),
    .to_SH(Tile_X0Y18_to_SH),
    .to_SI(Tile_X0Y18_to_SI),
    .A_O_top_0_t(Tile_X0Y18_A_O_top_0_t),
    .A_O_top_0_f(Tile_X0Y18_A_O_top_0_f),
    .A_O_top_1_t(Tile_X0Y18_A_O_top_1_t),
    .A_O_top_1_f(Tile_X0Y18_A_O_top_1_f),
    .A_prech1(Tile_X0Y18_A_prech1),
    .A_prech2(Tile_X0Y18_A_prech2),
    .A_DR_fault(Tile_X0Y18_A_DR_fault),
    .A_I_top_0_t(Tile_X0Y18_A_I_top_0_t),
    .A_I_top_0_f(Tile_X0Y18_A_I_top_0_f),
    .A_I_top_1_t(Tile_X0Y18_A_I_top_1_t),
    .A_I_top_1_f(Tile_X0Y18_A_I_top_1_f),
    .A_T_top(Tile_X0Y18_A_T_top),
    .A_F_masked1(Tile_X0Y18_A_F_masked1),
    .A_F_masked2(Tile_X0Y18_A_F_masked2),
    .A_config_C_bit0(Tile_X0Y18_A_config_C_bit0),
    .A_config_C_bit1(Tile_X0Y18_A_config_C_bit1),
    .A_config_C_bit2(Tile_X0Y18_A_config_C_bit2),
    .A_config_C_bit3(Tile_X0Y18_A_config_C_bit3),
    .B_config_C_bit0(Tile_X0Y18_B_config_C_bit0),
    .B_config_C_bit1(Tile_X0Y18_B_config_C_bit1),
    .B_config_C_bit2(Tile_X0Y18_B_config_C_bit2),
    .B_config_C_bit3(Tile_X0Y18_B_config_C_bit3),
    .UserCLK(Tile_X0Y19_UserCLKo),
    .UserCLKo(Tile_X0Y18_UserCLKo),
    .rst(Tile_X0Y19_rsto),
    .rsto(Tile_X0Y18_rsto),
    .FrameData(Tile_Y18_FrameData),
    .FrameData_O(Tile_X0Y18_FrameData_O),
    .FrameStrobe(Tile_X0Y19_FrameStrobe_O),
    .FrameStrobe_O(Tile_X0Y18_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X1Y18_Emulate_Bitstream)
    )
`endif
    Tile_X1Y18_linear_LMDPL
    (
    .from_NA(Tile_X1Y19_to_NA),
    .from_NB(Tile_X1Y19_to_NB),
    .from_NC(Tile_X1Y19_to_NC),
    .from_ND(Tile_X1Y19_to_ND),
    .from_NF(Tile_X1Y19_to_NF),
    .from_NG(Tile_X1Y19_to_NG),
    .from_NH(Tile_X1Y19_to_NH),
    .from_NI(Tile_X1Y19_to_NI),
    .from_EA(Tile_X0Y18_to_EA),
    .from_EB(Tile_X0Y18_to_EB),
    .from_EC(Tile_X0Y18_to_EC),
    .from_ED(Tile_X0Y18_to_ED),
    .from_EF(Tile_X0Y18_to_EF),
    .from_EG(Tile_X0Y18_to_EG),
    .from_EH(Tile_X0Y18_to_EH),
    .from_EI(Tile_X0Y18_to_EI),
    .from_SA(Tile_X1Y17_to_SA),
    .from_SB(Tile_X1Y17_to_SB),
    .from_SC(Tile_X1Y17_to_SC),
    .from_SD(Tile_X1Y17_to_SD),
    .from_SF(Tile_X1Y17_to_SF),
    .from_SG(Tile_X1Y17_to_SG),
    .from_SH(Tile_X1Y17_to_SH),
    .from_SI(Tile_X1Y17_to_SI),
    .from_WA(Tile_X2Y18_to_WA),
    .from_WB(Tile_X2Y18_to_WB),
    .from_WC(Tile_X2Y18_to_WC),
    .from_WD(Tile_X2Y18_to_WD),
    .from_WF(Tile_X2Y18_to_WF),
    .from_WG(Tile_X2Y18_to_WG),
    .from_WH(Tile_X2Y18_to_WH),
    .from_WI(Tile_X2Y18_to_WI),
    .to_EA(Tile_X1Y18_to_EA),
    .to_EB(Tile_X1Y18_to_EB),
    .to_EC(Tile_X1Y18_to_EC),
    .to_ED(Tile_X1Y18_to_ED),
    .to_EF(Tile_X1Y18_to_EF),
    .to_EG(Tile_X1Y18_to_EG),
    .to_EH(Tile_X1Y18_to_EH),
    .to_EI(Tile_X1Y18_to_EI),
    .to_WA(Tile_X1Y18_to_WA),
    .to_WB(Tile_X1Y18_to_WB),
    .to_WC(Tile_X1Y18_to_WC),
    .to_WD(Tile_X1Y18_to_WD),
    .to_WF(Tile_X1Y18_to_WF),
    .to_WG(Tile_X1Y18_to_WG),
    .to_WH(Tile_X1Y18_to_WH),
    .to_WI(Tile_X1Y18_to_WI),
    .to_NA(Tile_X1Y18_to_NA),
    .to_NB(Tile_X1Y18_to_NB),
    .to_NC(Tile_X1Y18_to_NC),
    .to_ND(Tile_X1Y18_to_ND),
    .to_NF(Tile_X1Y18_to_NF),
    .to_NG(Tile_X1Y18_to_NG),
    .to_NH(Tile_X1Y18_to_NH),
    .to_NI(Tile_X1Y18_to_NI),
    .to_SA(Tile_X1Y18_to_SA),
    .to_SB(Tile_X1Y18_to_SB),
    .to_SC(Tile_X1Y18_to_SC),
    .to_SD(Tile_X1Y18_to_SD),
    .to_SF(Tile_X1Y18_to_SF),
    .to_SG(Tile_X1Y18_to_SG),
    .to_SH(Tile_X1Y18_to_SH),
    .to_SI(Tile_X1Y18_to_SI),
    .F_masked1(Tile_X1Y18_F_masked1),
    .F_masked2(Tile_X1Y18_F_masked2),
    .UserCLK(Tile_X1Y19_UserCLKo),
    .UserCLKo(Tile_X1Y18_UserCLKo),
    .rst(Tile_X1Y19_rsto),
    .rsto(Tile_X1Y18_rsto),
    .FrameData(Tile_X0Y18_FrameData_O),
    .FrameData_O(Tile_X1Y18_FrameData_O),
    .FrameStrobe(Tile_X1Y19_FrameStrobe_O),
    .FrameStrobe_O(Tile_X1Y18_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X2Y18_Emulate_Bitstream)
    )
`endif
    Tile_X2Y18_linear_LMDPL
    (
    .from_NA(Tile_X2Y19_to_NA),
    .from_NB(Tile_X2Y19_to_NB),
    .from_NC(Tile_X2Y19_to_NC),
    .from_ND(Tile_X2Y19_to_ND),
    .from_NF(Tile_X2Y19_to_NF),
    .from_NG(Tile_X2Y19_to_NG),
    .from_NH(Tile_X2Y19_to_NH),
    .from_NI(Tile_X2Y19_to_NI),
    .from_EA(Tile_X1Y18_to_EA),
    .from_EB(Tile_X1Y18_to_EB),
    .from_EC(Tile_X1Y18_to_EC),
    .from_ED(Tile_X1Y18_to_ED),
    .from_EF(Tile_X1Y18_to_EF),
    .from_EG(Tile_X1Y18_to_EG),
    .from_EH(Tile_X1Y18_to_EH),
    .from_EI(Tile_X1Y18_to_EI),
    .from_SA(Tile_X2Y17_to_SA),
    .from_SB(Tile_X2Y17_to_SB),
    .from_SC(Tile_X2Y17_to_SC),
    .from_SD(Tile_X2Y17_to_SD),
    .from_SF(Tile_X2Y17_to_SF),
    .from_SG(Tile_X2Y17_to_SG),
    .from_SH(Tile_X2Y17_to_SH),
    .from_SI(Tile_X2Y17_to_SI),
    .from_WA(Tile_X3Y18_to_WA),
    .from_WB(Tile_X3Y18_to_WB),
    .from_WC(Tile_X3Y18_to_WC),
    .from_WD(Tile_X3Y18_to_WD),
    .from_WF(Tile_X3Y18_to_WF),
    .from_WG(Tile_X3Y18_to_WG),
    .from_WH(Tile_X3Y18_to_WH),
    .from_WI(Tile_X3Y18_to_WI),
    .to_EA(Tile_X2Y18_to_EA),
    .to_EB(Tile_X2Y18_to_EB),
    .to_EC(Tile_X2Y18_to_EC),
    .to_ED(Tile_X2Y18_to_ED),
    .to_EF(Tile_X2Y18_to_EF),
    .to_EG(Tile_X2Y18_to_EG),
    .to_EH(Tile_X2Y18_to_EH),
    .to_EI(Tile_X2Y18_to_EI),
    .to_WA(Tile_X2Y18_to_WA),
    .to_WB(Tile_X2Y18_to_WB),
    .to_WC(Tile_X2Y18_to_WC),
    .to_WD(Tile_X2Y18_to_WD),
    .to_WF(Tile_X2Y18_to_WF),
    .to_WG(Tile_X2Y18_to_WG),
    .to_WH(Tile_X2Y18_to_WH),
    .to_WI(Tile_X2Y18_to_WI),
    .to_NA(Tile_X2Y18_to_NA),
    .to_NB(Tile_X2Y18_to_NB),
    .to_NC(Tile_X2Y18_to_NC),
    .to_ND(Tile_X2Y18_to_ND),
    .to_NF(Tile_X2Y18_to_NF),
    .to_NG(Tile_X2Y18_to_NG),
    .to_NH(Tile_X2Y18_to_NH),
    .to_NI(Tile_X2Y18_to_NI),
    .to_SA(Tile_X2Y18_to_SA),
    .to_SB(Tile_X2Y18_to_SB),
    .to_SC(Tile_X2Y18_to_SC),
    .to_SD(Tile_X2Y18_to_SD),
    .to_SF(Tile_X2Y18_to_SF),
    .to_SG(Tile_X2Y18_to_SG),
    .to_SH(Tile_X2Y18_to_SH),
    .to_SI(Tile_X2Y18_to_SI),
    .F_masked1(Tile_X2Y18_F_masked1),
    .F_masked2(Tile_X2Y18_F_masked2),
    .UserCLK(Tile_X2Y19_UserCLKo),
    .UserCLKo(Tile_X2Y18_UserCLKo),
    .rst(Tile_X2Y19_rsto),
    .rsto(Tile_X2Y18_rsto),
    .FrameData(Tile_X1Y18_FrameData_O),
    .FrameData_O(Tile_X2Y18_FrameData_O),
    .FrameStrobe(Tile_X2Y19_FrameStrobe_O),
    .FrameStrobe_O(Tile_X2Y18_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
nonlinear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X3Y18_Emulate_Bitstream)
    )
`endif
    Tile_X3Y18_nonlinear_LMDPL
    (
    .from_NA(Tile_X3Y19_to_NA),
    .from_NB(Tile_X3Y19_to_NB),
    .from_NC(Tile_X3Y19_to_NC),
    .from_ND(Tile_X3Y19_to_ND),
    .from_NF(Tile_X3Y19_to_NF),
    .from_NG(Tile_X3Y19_to_NG),
    .from_NH(Tile_X3Y19_to_NH),
    .from_NI(Tile_X3Y19_to_NI),
    .from_EA(Tile_X2Y18_to_EA),
    .from_EB(Tile_X2Y18_to_EB),
    .from_EC(Tile_X2Y18_to_EC),
    .from_ED(Tile_X2Y18_to_ED),
    .from_EF(Tile_X2Y18_to_EF),
    .from_EG(Tile_X2Y18_to_EG),
    .from_EH(Tile_X2Y18_to_EH),
    .from_EI(Tile_X2Y18_to_EI),
    .from_SA(Tile_X3Y17_to_SA),
    .from_SB(Tile_X3Y17_to_SB),
    .from_SC(Tile_X3Y17_to_SC),
    .from_SD(Tile_X3Y17_to_SD),
    .from_SF(Tile_X3Y17_to_SF),
    .from_SG(Tile_X3Y17_to_SG),
    .from_SH(Tile_X3Y17_to_SH),
    .from_SI(Tile_X3Y17_to_SI),
    .from_WA(Tile_X4Y18_to_WA),
    .from_WB(Tile_X4Y18_to_WB),
    .from_WC(Tile_X4Y18_to_WC),
    .from_WD(Tile_X4Y18_to_WD),
    .from_WF(Tile_X4Y18_to_WF),
    .from_WG(Tile_X4Y18_to_WG),
    .from_WH(Tile_X4Y18_to_WH),
    .from_WI(Tile_X4Y18_to_WI),
    .to_EA(Tile_X3Y18_to_EA),
    .to_EB(Tile_X3Y18_to_EB),
    .to_EC(Tile_X3Y18_to_EC),
    .to_ED(Tile_X3Y18_to_ED),
    .to_EF(Tile_X3Y18_to_EF),
    .to_EG(Tile_X3Y18_to_EG),
    .to_EH(Tile_X3Y18_to_EH),
    .to_EI(Tile_X3Y18_to_EI),
    .to_WA(Tile_X3Y18_to_WA),
    .to_WB(Tile_X3Y18_to_WB),
    .to_WC(Tile_X3Y18_to_WC),
    .to_WD(Tile_X3Y18_to_WD),
    .to_WF(Tile_X3Y18_to_WF),
    .to_WG(Tile_X3Y18_to_WG),
    .to_WH(Tile_X3Y18_to_WH),
    .to_WI(Tile_X3Y18_to_WI),
    .to_NA(Tile_X3Y18_to_NA),
    .to_NB(Tile_X3Y18_to_NB),
    .to_NC(Tile_X3Y18_to_NC),
    .to_ND(Tile_X3Y18_to_ND),
    .to_NF(Tile_X3Y18_to_NF),
    .to_NG(Tile_X3Y18_to_NG),
    .to_NH(Tile_X3Y18_to_NH),
    .to_NI(Tile_X3Y18_to_NI),
    .to_SA(Tile_X3Y18_to_SA),
    .to_SB(Tile_X3Y18_to_SB),
    .to_SC(Tile_X3Y18_to_SC),
    .to_SD(Tile_X3Y18_to_SD),
    .to_SF(Tile_X3Y18_to_SF),
    .to_SG(Tile_X3Y18_to_SG),
    .to_SH(Tile_X3Y18_to_SH),
    .to_SI(Tile_X3Y18_to_SI),
    .R_t(Tile_X3Y18_R_t),
    .R_f(Tile_X3Y18_R_f),
    .F_masked1(Tile_X3Y18_F_masked1),
    .F_masked2(Tile_X3Y18_F_masked2),
    .UserCLK(Tile_X3Y19_UserCLKo),
    .UserCLKo(Tile_X3Y18_UserCLKo),
    .rst(Tile_X3Y19_rsto),
    .rsto(Tile_X3Y18_rsto),
    .FrameData(Tile_X2Y18_FrameData_O),
    .FrameData_O(Tile_X3Y18_FrameData_O),
    .FrameStrobe(Tile_X3Y19_FrameStrobe_O),
    .FrameStrobe_O(Tile_X3Y18_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X4Y18_Emulate_Bitstream)
    )
`endif
    Tile_X4Y18_linear_LMDPL
    (
    .from_NA(Tile_X4Y19_to_NA),
    .from_NB(Tile_X4Y19_to_NB),
    .from_NC(Tile_X4Y19_to_NC),
    .from_ND(Tile_X4Y19_to_ND),
    .from_NF(Tile_X4Y19_to_NF),
    .from_NG(Tile_X4Y19_to_NG),
    .from_NH(Tile_X4Y19_to_NH),
    .from_NI(Tile_X4Y19_to_NI),
    .from_EA(Tile_X3Y18_to_EA),
    .from_EB(Tile_X3Y18_to_EB),
    .from_EC(Tile_X3Y18_to_EC),
    .from_ED(Tile_X3Y18_to_ED),
    .from_EF(Tile_X3Y18_to_EF),
    .from_EG(Tile_X3Y18_to_EG),
    .from_EH(Tile_X3Y18_to_EH),
    .from_EI(Tile_X3Y18_to_EI),
    .from_SA(Tile_X4Y17_to_SA),
    .from_SB(Tile_X4Y17_to_SB),
    .from_SC(Tile_X4Y17_to_SC),
    .from_SD(Tile_X4Y17_to_SD),
    .from_SF(Tile_X4Y17_to_SF),
    .from_SG(Tile_X4Y17_to_SG),
    .from_SH(Tile_X4Y17_to_SH),
    .from_SI(Tile_X4Y17_to_SI),
    .from_WA(Tile_X5Y18_to_WA),
    .from_WB(Tile_X5Y18_to_WB),
    .from_WC(Tile_X5Y18_to_WC),
    .from_WD(Tile_X5Y18_to_WD),
    .from_WF(Tile_X5Y18_to_WF),
    .from_WG(Tile_X5Y18_to_WG),
    .from_WH(Tile_X5Y18_to_WH),
    .from_WI(Tile_X5Y18_to_WI),
    .to_EA(Tile_X4Y18_to_EA),
    .to_EB(Tile_X4Y18_to_EB),
    .to_EC(Tile_X4Y18_to_EC),
    .to_ED(Tile_X4Y18_to_ED),
    .to_EF(Tile_X4Y18_to_EF),
    .to_EG(Tile_X4Y18_to_EG),
    .to_EH(Tile_X4Y18_to_EH),
    .to_EI(Tile_X4Y18_to_EI),
    .to_WA(Tile_X4Y18_to_WA),
    .to_WB(Tile_X4Y18_to_WB),
    .to_WC(Tile_X4Y18_to_WC),
    .to_WD(Tile_X4Y18_to_WD),
    .to_WF(Tile_X4Y18_to_WF),
    .to_WG(Tile_X4Y18_to_WG),
    .to_WH(Tile_X4Y18_to_WH),
    .to_WI(Tile_X4Y18_to_WI),
    .to_NA(Tile_X4Y18_to_NA),
    .to_NB(Tile_X4Y18_to_NB),
    .to_NC(Tile_X4Y18_to_NC),
    .to_ND(Tile_X4Y18_to_ND),
    .to_NF(Tile_X4Y18_to_NF),
    .to_NG(Tile_X4Y18_to_NG),
    .to_NH(Tile_X4Y18_to_NH),
    .to_NI(Tile_X4Y18_to_NI),
    .to_SA(Tile_X4Y18_to_SA),
    .to_SB(Tile_X4Y18_to_SB),
    .to_SC(Tile_X4Y18_to_SC),
    .to_SD(Tile_X4Y18_to_SD),
    .to_SF(Tile_X4Y18_to_SF),
    .to_SG(Tile_X4Y18_to_SG),
    .to_SH(Tile_X4Y18_to_SH),
    .to_SI(Tile_X4Y18_to_SI),
    .F_masked1(Tile_X4Y18_F_masked1),
    .F_masked2(Tile_X4Y18_F_masked2),
    .UserCLK(Tile_X4Y19_UserCLKo),
    .UserCLKo(Tile_X4Y18_UserCLKo),
    .rst(Tile_X4Y19_rsto),
    .rsto(Tile_X4Y18_rsto),
    .FrameData(Tile_X3Y18_FrameData_O),
    .FrameData_O(Tile_X4Y18_FrameData_O),
    .FrameStrobe(Tile_X4Y19_FrameStrobe_O),
    .FrameStrobe_O(Tile_X4Y18_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X5Y18_Emulate_Bitstream)
    )
`endif
    Tile_X5Y18_linear_LMDPL
    (
    .from_NA(Tile_X5Y19_to_NA),
    .from_NB(Tile_X5Y19_to_NB),
    .from_NC(Tile_X5Y19_to_NC),
    .from_ND(Tile_X5Y19_to_ND),
    .from_NF(Tile_X5Y19_to_NF),
    .from_NG(Tile_X5Y19_to_NG),
    .from_NH(Tile_X5Y19_to_NH),
    .from_NI(Tile_X5Y19_to_NI),
    .from_EA(Tile_X4Y18_to_EA),
    .from_EB(Tile_X4Y18_to_EB),
    .from_EC(Tile_X4Y18_to_EC),
    .from_ED(Tile_X4Y18_to_ED),
    .from_EF(Tile_X4Y18_to_EF),
    .from_EG(Tile_X4Y18_to_EG),
    .from_EH(Tile_X4Y18_to_EH),
    .from_EI(Tile_X4Y18_to_EI),
    .from_SA(Tile_X5Y17_to_SA),
    .from_SB(Tile_X5Y17_to_SB),
    .from_SC(Tile_X5Y17_to_SC),
    .from_SD(Tile_X5Y17_to_SD),
    .from_SF(Tile_X5Y17_to_SF),
    .from_SG(Tile_X5Y17_to_SG),
    .from_SH(Tile_X5Y17_to_SH),
    .from_SI(Tile_X5Y17_to_SI),
    .from_WA(Tile_X6Y18_to_WA),
    .from_WB(Tile_X6Y18_to_WB),
    .from_WC(Tile_X6Y18_to_WC),
    .from_WD(Tile_X6Y18_to_WD),
    .from_WF(Tile_X6Y18_to_WF),
    .from_WG(Tile_X6Y18_to_WG),
    .from_WH(Tile_X6Y18_to_WH),
    .from_WI(Tile_X6Y18_to_WI),
    .to_EA(Tile_X5Y18_to_EA),
    .to_EB(Tile_X5Y18_to_EB),
    .to_EC(Tile_X5Y18_to_EC),
    .to_ED(Tile_X5Y18_to_ED),
    .to_EF(Tile_X5Y18_to_EF),
    .to_EG(Tile_X5Y18_to_EG),
    .to_EH(Tile_X5Y18_to_EH),
    .to_EI(Tile_X5Y18_to_EI),
    .to_WA(Tile_X5Y18_to_WA),
    .to_WB(Tile_X5Y18_to_WB),
    .to_WC(Tile_X5Y18_to_WC),
    .to_WD(Tile_X5Y18_to_WD),
    .to_WF(Tile_X5Y18_to_WF),
    .to_WG(Tile_X5Y18_to_WG),
    .to_WH(Tile_X5Y18_to_WH),
    .to_WI(Tile_X5Y18_to_WI),
    .to_NA(Tile_X5Y18_to_NA),
    .to_NB(Tile_X5Y18_to_NB),
    .to_NC(Tile_X5Y18_to_NC),
    .to_ND(Tile_X5Y18_to_ND),
    .to_NF(Tile_X5Y18_to_NF),
    .to_NG(Tile_X5Y18_to_NG),
    .to_NH(Tile_X5Y18_to_NH),
    .to_NI(Tile_X5Y18_to_NI),
    .to_SA(Tile_X5Y18_to_SA),
    .to_SB(Tile_X5Y18_to_SB),
    .to_SC(Tile_X5Y18_to_SC),
    .to_SD(Tile_X5Y18_to_SD),
    .to_SF(Tile_X5Y18_to_SF),
    .to_SG(Tile_X5Y18_to_SG),
    .to_SH(Tile_X5Y18_to_SH),
    .to_SI(Tile_X5Y18_to_SI),
    .F_masked1(Tile_X5Y18_F_masked1),
    .F_masked2(Tile_X5Y18_F_masked2),
    .UserCLK(Tile_X5Y19_UserCLKo),
    .UserCLKo(Tile_X5Y18_UserCLKo),
    .rst(Tile_X5Y19_rsto),
    .rsto(Tile_X5Y18_rsto),
    .FrameData(Tile_X4Y18_FrameData_O),
    .FrameData_O(Tile_X5Y18_FrameData_O),
    .FrameStrobe(Tile_X5Y19_FrameStrobe_O),
    .FrameStrobe_O(Tile_X5Y18_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
nonlinear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X6Y18_Emulate_Bitstream)
    )
`endif
    Tile_X6Y18_nonlinear_LMDPL
    (
    .from_NA(Tile_X6Y19_to_NA),
    .from_NB(Tile_X6Y19_to_NB),
    .from_NC(Tile_X6Y19_to_NC),
    .from_ND(Tile_X6Y19_to_ND),
    .from_NF(Tile_X6Y19_to_NF),
    .from_NG(Tile_X6Y19_to_NG),
    .from_NH(Tile_X6Y19_to_NH),
    .from_NI(Tile_X6Y19_to_NI),
    .from_EA(Tile_X5Y18_to_EA),
    .from_EB(Tile_X5Y18_to_EB),
    .from_EC(Tile_X5Y18_to_EC),
    .from_ED(Tile_X5Y18_to_ED),
    .from_EF(Tile_X5Y18_to_EF),
    .from_EG(Tile_X5Y18_to_EG),
    .from_EH(Tile_X5Y18_to_EH),
    .from_EI(Tile_X5Y18_to_EI),
    .from_SA(Tile_X6Y17_to_SA),
    .from_SB(Tile_X6Y17_to_SB),
    .from_SC(Tile_X6Y17_to_SC),
    .from_SD(Tile_X6Y17_to_SD),
    .from_SF(Tile_X6Y17_to_SF),
    .from_SG(Tile_X6Y17_to_SG),
    .from_SH(Tile_X6Y17_to_SH),
    .from_SI(Tile_X6Y17_to_SI),
    .from_WA(Tile_X7Y18_to_WA),
    .from_WB(Tile_X7Y18_to_WB),
    .from_WC(Tile_X7Y18_to_WC),
    .from_WD(Tile_X7Y18_to_WD),
    .from_WF(Tile_X7Y18_to_WF),
    .from_WG(Tile_X7Y18_to_WG),
    .from_WH(Tile_X7Y18_to_WH),
    .from_WI(Tile_X7Y18_to_WI),
    .to_EA(Tile_X6Y18_to_EA),
    .to_EB(Tile_X6Y18_to_EB),
    .to_EC(Tile_X6Y18_to_EC),
    .to_ED(Tile_X6Y18_to_ED),
    .to_EF(Tile_X6Y18_to_EF),
    .to_EG(Tile_X6Y18_to_EG),
    .to_EH(Tile_X6Y18_to_EH),
    .to_EI(Tile_X6Y18_to_EI),
    .to_WA(Tile_X6Y18_to_WA),
    .to_WB(Tile_X6Y18_to_WB),
    .to_WC(Tile_X6Y18_to_WC),
    .to_WD(Tile_X6Y18_to_WD),
    .to_WF(Tile_X6Y18_to_WF),
    .to_WG(Tile_X6Y18_to_WG),
    .to_WH(Tile_X6Y18_to_WH),
    .to_WI(Tile_X6Y18_to_WI),
    .to_NA(Tile_X6Y18_to_NA),
    .to_NB(Tile_X6Y18_to_NB),
    .to_NC(Tile_X6Y18_to_NC),
    .to_ND(Tile_X6Y18_to_ND),
    .to_NF(Tile_X6Y18_to_NF),
    .to_NG(Tile_X6Y18_to_NG),
    .to_NH(Tile_X6Y18_to_NH),
    .to_NI(Tile_X6Y18_to_NI),
    .to_SA(Tile_X6Y18_to_SA),
    .to_SB(Tile_X6Y18_to_SB),
    .to_SC(Tile_X6Y18_to_SC),
    .to_SD(Tile_X6Y18_to_SD),
    .to_SF(Tile_X6Y18_to_SF),
    .to_SG(Tile_X6Y18_to_SG),
    .to_SH(Tile_X6Y18_to_SH),
    .to_SI(Tile_X6Y18_to_SI),
    .R_t(Tile_X6Y18_R_t),
    .R_f(Tile_X6Y18_R_f),
    .F_masked1(Tile_X6Y18_F_masked1),
    .F_masked2(Tile_X6Y18_F_masked2),
    .UserCLK(Tile_X6Y19_UserCLKo),
    .UserCLKo(Tile_X6Y18_UserCLKo),
    .rst(Tile_X6Y19_rsto),
    .rsto(Tile_X6Y18_rsto),
    .FrameData(Tile_X5Y18_FrameData_O),
    .FrameData_O(Tile_X6Y18_FrameData_O),
    .FrameStrobe(Tile_X6Y19_FrameStrobe_O),
    .FrameStrobe_O(Tile_X6Y18_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X7Y18_Emulate_Bitstream)
    )
`endif
    Tile_X7Y18_linear_LMDPL
    (
    .from_NA(Tile_X7Y19_to_NA),
    .from_NB(Tile_X7Y19_to_NB),
    .from_NC(Tile_X7Y19_to_NC),
    .from_ND(Tile_X7Y19_to_ND),
    .from_NF(Tile_X7Y19_to_NF),
    .from_NG(Tile_X7Y19_to_NG),
    .from_NH(Tile_X7Y19_to_NH),
    .from_NI(Tile_X7Y19_to_NI),
    .from_EA(Tile_X6Y18_to_EA),
    .from_EB(Tile_X6Y18_to_EB),
    .from_EC(Tile_X6Y18_to_EC),
    .from_ED(Tile_X6Y18_to_ED),
    .from_EF(Tile_X6Y18_to_EF),
    .from_EG(Tile_X6Y18_to_EG),
    .from_EH(Tile_X6Y18_to_EH),
    .from_EI(Tile_X6Y18_to_EI),
    .from_SA(Tile_X7Y17_to_SA),
    .from_SB(Tile_X7Y17_to_SB),
    .from_SC(Tile_X7Y17_to_SC),
    .from_SD(Tile_X7Y17_to_SD),
    .from_SF(Tile_X7Y17_to_SF),
    .from_SG(Tile_X7Y17_to_SG),
    .from_SH(Tile_X7Y17_to_SH),
    .from_SI(Tile_X7Y17_to_SI),
    .from_WA(Tile_X8Y18_to_WA),
    .from_WB(Tile_X8Y18_to_WB),
    .from_WC(Tile_X8Y18_to_WC),
    .from_WD(Tile_X8Y18_to_WD),
    .from_WF(Tile_X8Y18_to_WF),
    .from_WG(Tile_X8Y18_to_WG),
    .from_WH(Tile_X8Y18_to_WH),
    .from_WI(Tile_X8Y18_to_WI),
    .to_EA(Tile_X7Y18_to_EA),
    .to_EB(Tile_X7Y18_to_EB),
    .to_EC(Tile_X7Y18_to_EC),
    .to_ED(Tile_X7Y18_to_ED),
    .to_EF(Tile_X7Y18_to_EF),
    .to_EG(Tile_X7Y18_to_EG),
    .to_EH(Tile_X7Y18_to_EH),
    .to_EI(Tile_X7Y18_to_EI),
    .to_WA(Tile_X7Y18_to_WA),
    .to_WB(Tile_X7Y18_to_WB),
    .to_WC(Tile_X7Y18_to_WC),
    .to_WD(Tile_X7Y18_to_WD),
    .to_WF(Tile_X7Y18_to_WF),
    .to_WG(Tile_X7Y18_to_WG),
    .to_WH(Tile_X7Y18_to_WH),
    .to_WI(Tile_X7Y18_to_WI),
    .to_NA(Tile_X7Y18_to_NA),
    .to_NB(Tile_X7Y18_to_NB),
    .to_NC(Tile_X7Y18_to_NC),
    .to_ND(Tile_X7Y18_to_ND),
    .to_NF(Tile_X7Y18_to_NF),
    .to_NG(Tile_X7Y18_to_NG),
    .to_NH(Tile_X7Y18_to_NH),
    .to_NI(Tile_X7Y18_to_NI),
    .to_SA(Tile_X7Y18_to_SA),
    .to_SB(Tile_X7Y18_to_SB),
    .to_SC(Tile_X7Y18_to_SC),
    .to_SD(Tile_X7Y18_to_SD),
    .to_SF(Tile_X7Y18_to_SF),
    .to_SG(Tile_X7Y18_to_SG),
    .to_SH(Tile_X7Y18_to_SH),
    .to_SI(Tile_X7Y18_to_SI),
    .F_masked1(Tile_X7Y18_F_masked1),
    .F_masked2(Tile_X7Y18_F_masked2),
    .UserCLK(Tile_X7Y19_UserCLKo),
    .UserCLKo(Tile_X7Y18_UserCLKo),
    .rst(Tile_X7Y19_rsto),
    .rsto(Tile_X7Y18_rsto),
    .FrameData(Tile_X6Y18_FrameData_O),
    .FrameData_O(Tile_X7Y18_FrameData_O),
    .FrameStrobe(Tile_X7Y19_FrameStrobe_O),
    .FrameStrobe_O(Tile_X7Y18_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
ctrl_to_sec
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X8Y18_Emulate_Bitstream)
    )
`endif
    Tile_X8Y18_ctrl_to_sec
    (
    .from_NA(Tile_X8Y19_to_NA),
    .from_NB(Tile_X8Y19_to_NB),
    .from_NC(Tile_X8Y19_to_NC),
    .from_ND(Tile_X8Y19_to_ND),
    .from_NF(Tile_X8Y19_to_NF),
    .from_NG(Tile_X8Y19_to_NG),
    .from_NH(Tile_X8Y19_to_NH),
    .from_NI(Tile_X8Y19_to_NI),
    .from_EA(Tile_X7Y18_to_EA),
    .from_EB(Tile_X7Y18_to_EB),
    .from_EC(Tile_X7Y18_to_EC),
    .from_ED(Tile_X7Y18_to_ED),
    .from_EF(Tile_X7Y18_to_EF),
    .from_EG(Tile_X7Y18_to_EG),
    .from_EH(Tile_X7Y18_to_EH),
    .from_EI(Tile_X7Y18_to_EI),
    .from_SA(Tile_X8Y17_to_SA),
    .from_SB(Tile_X8Y17_to_SB),
    .from_SC(Tile_X8Y17_to_SC),
    .from_SD(Tile_X8Y17_to_SD),
    .from_SF(Tile_X8Y17_to_SF),
    .from_SG(Tile_X8Y17_to_SG),
    .from_SH(Tile_X8Y17_to_SH),
    .from_SI(Tile_X8Y17_to_SI),
    .from_WA_1s(Tile_X9Y18_to_WA_1s),
    .from_WB_1s(Tile_X9Y18_to_WB_1s),
    .from_WC_1s(Tile_X9Y18_to_WC_1s),
    .from_WD_1s(Tile_X9Y18_to_WD_1s),
    .from_WF_1s(Tile_X9Y18_to_WF_1s),
    .from_WG_1s(Tile_X9Y18_to_WG_1s),
    .from_WH_1s(Tile_X9Y18_to_WH_1s),
    .from_WI_1s(Tile_X9Y18_to_WI_1s),
    .to_WA(Tile_X8Y18_to_WA),
    .to_WB(Tile_X8Y18_to_WB),
    .to_WC(Tile_X8Y18_to_WC),
    .to_WD(Tile_X8Y18_to_WD),
    .to_WF(Tile_X8Y18_to_WF),
    .to_WG(Tile_X8Y18_to_WG),
    .to_WH(Tile_X8Y18_to_WH),
    .to_WI(Tile_X8Y18_to_WI),
    .to_NA(Tile_X8Y18_to_NA),
    .to_NB(Tile_X8Y18_to_NB),
    .to_NC(Tile_X8Y18_to_NC),
    .to_ND(Tile_X8Y18_to_ND),
    .to_NF(Tile_X8Y18_to_NF),
    .to_NG(Tile_X8Y18_to_NG),
    .to_NH(Tile_X8Y18_to_NH),
    .to_NI(Tile_X8Y18_to_NI),
    .to_SA(Tile_X8Y18_to_SA),
    .to_SB(Tile_X8Y18_to_SB),
    .to_SC(Tile_X8Y18_to_SC),
    .to_SD(Tile_X8Y18_to_SD),
    .to_SF(Tile_X8Y18_to_SF),
    .to_SG(Tile_X8Y18_to_SG),
    .to_SH(Tile_X8Y18_to_SH),
    .to_SI(Tile_X8Y18_to_SI),
    .UserCLK(Tile_X8Y19_UserCLKo),
    .UserCLKo(Tile_X8Y18_UserCLKo),
    .rst(Tile_X8Y19_rsto),
    .rsto(Tile_X8Y18_rsto),
    .FrameData(Tile_X7Y18_FrameData_O),
    .FrameData_O(Tile_X8Y18_FrameData_O),
    .FrameStrobe(Tile_X8Y19_FrameStrobe_O),
    .FrameStrobe_O(Tile_X8Y18_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
combined_WDDL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X9Y18_Emulate_Bitstream)
    )
`endif
    Tile_X9Y18_combined_WDDL
    (
    .from_NA_1s(Tile_X9Y19_to_NA_1s),
    .from_NB_1s(Tile_X9Y19_to_NB_1s),
    .from_NC_1s(Tile_X9Y19_to_NC_1s),
    .from_ND_1s(Tile_X9Y19_to_ND_1s),
    .from_NF_1s(Tile_X9Y19_to_NF_1s),
    .from_NG_1s(Tile_X9Y19_to_NG_1s),
    .from_NH_1s(Tile_X9Y19_to_NH_1s),
    .from_NI_1s(Tile_X9Y19_to_NI_1s),
    .from_SA_1s(Tile_X9Y17_to_SA_1s),
    .from_SB_1s(Tile_X9Y17_to_SB_1s),
    .from_SC_1s(Tile_X9Y17_to_SC_1s),
    .from_SD_1s(Tile_X9Y17_to_SD_1s),
    .from_SF_1s(Tile_X9Y17_to_SF_1s),
    .from_SG_1s(Tile_X9Y17_to_SG_1s),
    .from_SH_1s(Tile_X9Y17_to_SH_1s),
    .from_SI_1s(Tile_X9Y17_to_SI_1s),
    .from_WA_1s(Tile_X10Y18_to_WA_1s),
    .from_WB_1s(Tile_X10Y18_to_WB_1s),
    .from_WC_1s(Tile_X10Y18_to_WC_1s),
    .from_WD_1s(Tile_X10Y18_to_WD_1s),
    .from_WF_1s(Tile_X10Y18_to_WF_1s),
    .from_WG_1s(Tile_X10Y18_to_WG_1s),
    .from_WH_1s(Tile_X10Y18_to_WH_1s),
    .from_WI_1s(Tile_X10Y18_to_WI_1s),
    .to_EA_1s(Tile_X9Y18_to_EA_1s),
    .to_EB_1s(Tile_X9Y18_to_EB_1s),
    .to_EC_1s(Tile_X9Y18_to_EC_1s),
    .to_ED_1s(Tile_X9Y18_to_ED_1s),
    .to_EF_1s(Tile_X9Y18_to_EF_1s),
    .to_EG_1s(Tile_X9Y18_to_EG_1s),
    .to_EH_1s(Tile_X9Y18_to_EH_1s),
    .to_EI_1s(Tile_X9Y18_to_EI_1s),
    .to_WA_1s(Tile_X9Y18_to_WA_1s),
    .to_WB_1s(Tile_X9Y18_to_WB_1s),
    .to_WC_1s(Tile_X9Y18_to_WC_1s),
    .to_WD_1s(Tile_X9Y18_to_WD_1s),
    .to_WF_1s(Tile_X9Y18_to_WF_1s),
    .to_WG_1s(Tile_X9Y18_to_WG_1s),
    .to_WH_1s(Tile_X9Y18_to_WH_1s),
    .to_WI_1s(Tile_X9Y18_to_WI_1s),
    .to_NA_1s(Tile_X9Y18_to_NA_1s),
    .to_NB_1s(Tile_X9Y18_to_NB_1s),
    .to_NC_1s(Tile_X9Y18_to_NC_1s),
    .to_ND_1s(Tile_X9Y18_to_ND_1s),
    .to_NF_1s(Tile_X9Y18_to_NF_1s),
    .to_NG_1s(Tile_X9Y18_to_NG_1s),
    .to_NH_1s(Tile_X9Y18_to_NH_1s),
    .to_NI_1s(Tile_X9Y18_to_NI_1s),
    .to_SA_1s(Tile_X9Y18_to_SA_1s),
    .to_SB_1s(Tile_X9Y18_to_SB_1s),
    .to_SC_1s(Tile_X9Y18_to_SC_1s),
    .to_SD_1s(Tile_X9Y18_to_SD_1s),
    .to_SF_1s(Tile_X9Y18_to_SF_1s),
    .to_SG_1s(Tile_X9Y18_to_SG_1s),
    .to_SH_1s(Tile_X9Y18_to_SH_1s),
    .to_SI_1s(Tile_X9Y18_to_SI_1s),
    .F_ctrl(Tile_X9Y18_F_ctrl),
    .UserCLK(Tile_X9Y19_UserCLKo),
    .UserCLKo(Tile_X9Y18_UserCLKo),
    .rst(Tile_X9Y19_rsto),
    .rsto(Tile_X9Y18_rsto),
    .FrameData(Tile_X8Y18_FrameData_O),
    .FrameData_O(Tile_X9Y18_FrameData_O),
    .FrameStrobe(Tile_X9Y19_FrameStrobe_O),
    .FrameStrobe_O(Tile_X9Y18_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
ctrl_IO
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X10Y18_Emulate_Bitstream)
    )
`endif
    Tile_X10Y18_ctrl_IO
    (
    .from_EA_1s(Tile_X9Y18_to_EA_1s),
    .from_EB_1s(Tile_X9Y18_to_EB_1s),
    .from_EC_1s(Tile_X9Y18_to_EC_1s),
    .from_ED_1s(Tile_X9Y18_to_ED_1s),
    .from_EF_1s(Tile_X9Y18_to_EF_1s),
    .from_EG_1s(Tile_X9Y18_to_EG_1s),
    .from_EH_1s(Tile_X9Y18_to_EH_1s),
    .from_EI_1s(Tile_X9Y18_to_EI_1s),
    .to_WA_1s(Tile_X10Y18_to_WA_1s),
    .to_WB_1s(Tile_X10Y18_to_WB_1s),
    .to_WC_1s(Tile_X10Y18_to_WC_1s),
    .to_WD_1s(Tile_X10Y18_to_WD_1s),
    .to_WF_1s(Tile_X10Y18_to_WF_1s),
    .to_WG_1s(Tile_X10Y18_to_WG_1s),
    .to_WH_1s(Tile_X10Y18_to_WH_1s),
    .to_WI_1s(Tile_X10Y18_to_WI_1s),
    .A_O_top_0_t(Tile_X10Y18_A_O_top_0_t),
    .A_O_top_0_f(Tile_X10Y18_A_O_top_0_f),
    .A_prech2(Tile_X10Y18_A_prech2),
    .A_DR_fault(Tile_X10Y18_A_DR_fault),
    .A_I_top_0_t(Tile_X10Y18_A_I_top_0_t),
    .A_I_top_0_f(Tile_X10Y18_A_I_top_0_f),
    .A_T_top(Tile_X10Y18_A_T_top),
    .A_F_ctrl(Tile_X10Y18_A_F_ctrl),
    .UserCLK(Tile_X10Y19_UserCLKo),
    .UserCLKo(Tile_X10Y18_UserCLKo),
    .rst(Tile_X10Y19_rsto),
    .rsto(Tile_X10Y18_rsto),
    .FrameData(Tile_X9Y18_FrameData_O),
    .FrameData_O(Tile_X10Y18_FrameData_O),
    .FrameStrobe(Tile_X10Y19_FrameStrobe_O),
    .FrameStrobe_O(Tile_X10Y18_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
W_IO_custom
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X0Y19_Emulate_Bitstream)
    )
`endif
    Tile_X0Y19_W_IO_custom
    (
    .from_NA(Tile_X0Y20_to_NA),
    .from_NB(Tile_X0Y20_to_NB),
    .from_NC(Tile_X0Y20_to_NC),
    .from_ND(Tile_X0Y20_to_ND),
    .from_NF(Tile_X0Y20_to_NF),
    .from_NG(Tile_X0Y20_to_NG),
    .from_NH(Tile_X0Y20_to_NH),
    .from_NI(Tile_X0Y20_to_NI),
    .from_SA(Tile_X0Y18_to_SA),
    .from_SB(Tile_X0Y18_to_SB),
    .from_SC(Tile_X0Y18_to_SC),
    .from_SD(Tile_X0Y18_to_SD),
    .from_SF(Tile_X0Y18_to_SF),
    .from_SG(Tile_X0Y18_to_SG),
    .from_SH(Tile_X0Y18_to_SH),
    .from_SI(Tile_X0Y18_to_SI),
    .from_WA(Tile_X1Y19_to_WA),
    .from_WB(Tile_X1Y19_to_WB),
    .from_WC(Tile_X1Y19_to_WC),
    .from_WD(Tile_X1Y19_to_WD),
    .from_WF(Tile_X1Y19_to_WF),
    .from_WG(Tile_X1Y19_to_WG),
    .from_WH(Tile_X1Y19_to_WH),
    .from_WI(Tile_X1Y19_to_WI),
    .to_EA(Tile_X0Y19_to_EA),
    .to_EB(Tile_X0Y19_to_EB),
    .to_EC(Tile_X0Y19_to_EC),
    .to_ED(Tile_X0Y19_to_ED),
    .to_EF(Tile_X0Y19_to_EF),
    .to_EG(Tile_X0Y19_to_EG),
    .to_EH(Tile_X0Y19_to_EH),
    .to_EI(Tile_X0Y19_to_EI),
    .to_NA(Tile_X0Y19_to_NA),
    .to_NB(Tile_X0Y19_to_NB),
    .to_NC(Tile_X0Y19_to_NC),
    .to_ND(Tile_X0Y19_to_ND),
    .to_NF(Tile_X0Y19_to_NF),
    .to_NG(Tile_X0Y19_to_NG),
    .to_NH(Tile_X0Y19_to_NH),
    .to_NI(Tile_X0Y19_to_NI),
    .to_SA(Tile_X0Y19_to_SA),
    .to_SB(Tile_X0Y19_to_SB),
    .to_SC(Tile_X0Y19_to_SC),
    .to_SD(Tile_X0Y19_to_SD),
    .to_SF(Tile_X0Y19_to_SF),
    .to_SG(Tile_X0Y19_to_SG),
    .to_SH(Tile_X0Y19_to_SH),
    .to_SI(Tile_X0Y19_to_SI),
    .A_O_top_0_t(Tile_X0Y19_A_O_top_0_t),
    .A_O_top_0_f(Tile_X0Y19_A_O_top_0_f),
    .A_O_top_1_t(Tile_X0Y19_A_O_top_1_t),
    .A_O_top_1_f(Tile_X0Y19_A_O_top_1_f),
    .A_prech1(Tile_X0Y19_A_prech1),
    .A_prech2(Tile_X0Y19_A_prech2),
    .A_DR_fault(Tile_X0Y19_A_DR_fault),
    .A_I_top_0_t(Tile_X0Y19_A_I_top_0_t),
    .A_I_top_0_f(Tile_X0Y19_A_I_top_0_f),
    .A_I_top_1_t(Tile_X0Y19_A_I_top_1_t),
    .A_I_top_1_f(Tile_X0Y19_A_I_top_1_f),
    .A_T_top(Tile_X0Y19_A_T_top),
    .A_F_masked1(Tile_X0Y19_A_F_masked1),
    .A_F_masked2(Tile_X0Y19_A_F_masked2),
    .A_config_C_bit0(Tile_X0Y19_A_config_C_bit0),
    .A_config_C_bit1(Tile_X0Y19_A_config_C_bit1),
    .A_config_C_bit2(Tile_X0Y19_A_config_C_bit2),
    .A_config_C_bit3(Tile_X0Y19_A_config_C_bit3),
    .B_config_C_bit0(Tile_X0Y19_B_config_C_bit0),
    .B_config_C_bit1(Tile_X0Y19_B_config_C_bit1),
    .B_config_C_bit2(Tile_X0Y19_B_config_C_bit2),
    .B_config_C_bit3(Tile_X0Y19_B_config_C_bit3),
    .UserCLK(Tile_X0Y20_UserCLKo),
    .UserCLKo(Tile_X0Y19_UserCLKo),
    .rst(Tile_X0Y20_rsto),
    .rsto(Tile_X0Y19_rsto),
    .FrameData(Tile_Y19_FrameData),
    .FrameData_O(Tile_X0Y19_FrameData_O),
    .FrameStrobe(Tile_X0Y20_FrameStrobe_O),
    .FrameStrobe_O(Tile_X0Y19_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X1Y19_Emulate_Bitstream)
    )
`endif
    Tile_X1Y19_linear_LMDPL
    (
    .from_NA(Tile_X1Y20_to_NA),
    .from_NB(Tile_X1Y20_to_NB),
    .from_NC(Tile_X1Y20_to_NC),
    .from_ND(Tile_X1Y20_to_ND),
    .from_NF(Tile_X1Y20_to_NF),
    .from_NG(Tile_X1Y20_to_NG),
    .from_NH(Tile_X1Y20_to_NH),
    .from_NI(Tile_X1Y20_to_NI),
    .from_EA(Tile_X0Y19_to_EA),
    .from_EB(Tile_X0Y19_to_EB),
    .from_EC(Tile_X0Y19_to_EC),
    .from_ED(Tile_X0Y19_to_ED),
    .from_EF(Tile_X0Y19_to_EF),
    .from_EG(Tile_X0Y19_to_EG),
    .from_EH(Tile_X0Y19_to_EH),
    .from_EI(Tile_X0Y19_to_EI),
    .from_SA(Tile_X1Y18_to_SA),
    .from_SB(Tile_X1Y18_to_SB),
    .from_SC(Tile_X1Y18_to_SC),
    .from_SD(Tile_X1Y18_to_SD),
    .from_SF(Tile_X1Y18_to_SF),
    .from_SG(Tile_X1Y18_to_SG),
    .from_SH(Tile_X1Y18_to_SH),
    .from_SI(Tile_X1Y18_to_SI),
    .from_WA(Tile_X2Y19_to_WA),
    .from_WB(Tile_X2Y19_to_WB),
    .from_WC(Tile_X2Y19_to_WC),
    .from_WD(Tile_X2Y19_to_WD),
    .from_WF(Tile_X2Y19_to_WF),
    .from_WG(Tile_X2Y19_to_WG),
    .from_WH(Tile_X2Y19_to_WH),
    .from_WI(Tile_X2Y19_to_WI),
    .to_EA(Tile_X1Y19_to_EA),
    .to_EB(Tile_X1Y19_to_EB),
    .to_EC(Tile_X1Y19_to_EC),
    .to_ED(Tile_X1Y19_to_ED),
    .to_EF(Tile_X1Y19_to_EF),
    .to_EG(Tile_X1Y19_to_EG),
    .to_EH(Tile_X1Y19_to_EH),
    .to_EI(Tile_X1Y19_to_EI),
    .to_WA(Tile_X1Y19_to_WA),
    .to_WB(Tile_X1Y19_to_WB),
    .to_WC(Tile_X1Y19_to_WC),
    .to_WD(Tile_X1Y19_to_WD),
    .to_WF(Tile_X1Y19_to_WF),
    .to_WG(Tile_X1Y19_to_WG),
    .to_WH(Tile_X1Y19_to_WH),
    .to_WI(Tile_X1Y19_to_WI),
    .to_NA(Tile_X1Y19_to_NA),
    .to_NB(Tile_X1Y19_to_NB),
    .to_NC(Tile_X1Y19_to_NC),
    .to_ND(Tile_X1Y19_to_ND),
    .to_NF(Tile_X1Y19_to_NF),
    .to_NG(Tile_X1Y19_to_NG),
    .to_NH(Tile_X1Y19_to_NH),
    .to_NI(Tile_X1Y19_to_NI),
    .to_SA(Tile_X1Y19_to_SA),
    .to_SB(Tile_X1Y19_to_SB),
    .to_SC(Tile_X1Y19_to_SC),
    .to_SD(Tile_X1Y19_to_SD),
    .to_SF(Tile_X1Y19_to_SF),
    .to_SG(Tile_X1Y19_to_SG),
    .to_SH(Tile_X1Y19_to_SH),
    .to_SI(Tile_X1Y19_to_SI),
    .F_masked1(Tile_X1Y19_F_masked1),
    .F_masked2(Tile_X1Y19_F_masked2),
    .UserCLK(Tile_X1Y20_UserCLKo),
    .UserCLKo(Tile_X1Y19_UserCLKo),
    .rst(Tile_X1Y20_rsto),
    .rsto(Tile_X1Y19_rsto),
    .FrameData(Tile_X0Y19_FrameData_O),
    .FrameData_O(Tile_X1Y19_FrameData_O),
    .FrameStrobe(Tile_X1Y20_FrameStrobe_O),
    .FrameStrobe_O(Tile_X1Y19_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X2Y19_Emulate_Bitstream)
    )
`endif
    Tile_X2Y19_linear_LMDPL
    (
    .from_NA(Tile_X2Y20_to_NA),
    .from_NB(Tile_X2Y20_to_NB),
    .from_NC(Tile_X2Y20_to_NC),
    .from_ND(Tile_X2Y20_to_ND),
    .from_NF(Tile_X2Y20_to_NF),
    .from_NG(Tile_X2Y20_to_NG),
    .from_NH(Tile_X2Y20_to_NH),
    .from_NI(Tile_X2Y20_to_NI),
    .from_EA(Tile_X1Y19_to_EA),
    .from_EB(Tile_X1Y19_to_EB),
    .from_EC(Tile_X1Y19_to_EC),
    .from_ED(Tile_X1Y19_to_ED),
    .from_EF(Tile_X1Y19_to_EF),
    .from_EG(Tile_X1Y19_to_EG),
    .from_EH(Tile_X1Y19_to_EH),
    .from_EI(Tile_X1Y19_to_EI),
    .from_SA(Tile_X2Y18_to_SA),
    .from_SB(Tile_X2Y18_to_SB),
    .from_SC(Tile_X2Y18_to_SC),
    .from_SD(Tile_X2Y18_to_SD),
    .from_SF(Tile_X2Y18_to_SF),
    .from_SG(Tile_X2Y18_to_SG),
    .from_SH(Tile_X2Y18_to_SH),
    .from_SI(Tile_X2Y18_to_SI),
    .from_WA(Tile_X3Y19_to_WA),
    .from_WB(Tile_X3Y19_to_WB),
    .from_WC(Tile_X3Y19_to_WC),
    .from_WD(Tile_X3Y19_to_WD),
    .from_WF(Tile_X3Y19_to_WF),
    .from_WG(Tile_X3Y19_to_WG),
    .from_WH(Tile_X3Y19_to_WH),
    .from_WI(Tile_X3Y19_to_WI),
    .to_EA(Tile_X2Y19_to_EA),
    .to_EB(Tile_X2Y19_to_EB),
    .to_EC(Tile_X2Y19_to_EC),
    .to_ED(Tile_X2Y19_to_ED),
    .to_EF(Tile_X2Y19_to_EF),
    .to_EG(Tile_X2Y19_to_EG),
    .to_EH(Tile_X2Y19_to_EH),
    .to_EI(Tile_X2Y19_to_EI),
    .to_WA(Tile_X2Y19_to_WA),
    .to_WB(Tile_X2Y19_to_WB),
    .to_WC(Tile_X2Y19_to_WC),
    .to_WD(Tile_X2Y19_to_WD),
    .to_WF(Tile_X2Y19_to_WF),
    .to_WG(Tile_X2Y19_to_WG),
    .to_WH(Tile_X2Y19_to_WH),
    .to_WI(Tile_X2Y19_to_WI),
    .to_NA(Tile_X2Y19_to_NA),
    .to_NB(Tile_X2Y19_to_NB),
    .to_NC(Tile_X2Y19_to_NC),
    .to_ND(Tile_X2Y19_to_ND),
    .to_NF(Tile_X2Y19_to_NF),
    .to_NG(Tile_X2Y19_to_NG),
    .to_NH(Tile_X2Y19_to_NH),
    .to_NI(Tile_X2Y19_to_NI),
    .to_SA(Tile_X2Y19_to_SA),
    .to_SB(Tile_X2Y19_to_SB),
    .to_SC(Tile_X2Y19_to_SC),
    .to_SD(Tile_X2Y19_to_SD),
    .to_SF(Tile_X2Y19_to_SF),
    .to_SG(Tile_X2Y19_to_SG),
    .to_SH(Tile_X2Y19_to_SH),
    .to_SI(Tile_X2Y19_to_SI),
    .F_masked1(Tile_X2Y19_F_masked1),
    .F_masked2(Tile_X2Y19_F_masked2),
    .UserCLK(Tile_X2Y20_UserCLKo),
    .UserCLKo(Tile_X2Y19_UserCLKo),
    .rst(Tile_X2Y20_rsto),
    .rsto(Tile_X2Y19_rsto),
    .FrameData(Tile_X1Y19_FrameData_O),
    .FrameData_O(Tile_X2Y19_FrameData_O),
    .FrameStrobe(Tile_X2Y20_FrameStrobe_O),
    .FrameStrobe_O(Tile_X2Y19_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
nonlinear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X3Y19_Emulate_Bitstream)
    )
`endif
    Tile_X3Y19_nonlinear_LMDPL
    (
    .from_NA(Tile_X3Y20_to_NA),
    .from_NB(Tile_X3Y20_to_NB),
    .from_NC(Tile_X3Y20_to_NC),
    .from_ND(Tile_X3Y20_to_ND),
    .from_NF(Tile_X3Y20_to_NF),
    .from_NG(Tile_X3Y20_to_NG),
    .from_NH(Tile_X3Y20_to_NH),
    .from_NI(Tile_X3Y20_to_NI),
    .from_EA(Tile_X2Y19_to_EA),
    .from_EB(Tile_X2Y19_to_EB),
    .from_EC(Tile_X2Y19_to_EC),
    .from_ED(Tile_X2Y19_to_ED),
    .from_EF(Tile_X2Y19_to_EF),
    .from_EG(Tile_X2Y19_to_EG),
    .from_EH(Tile_X2Y19_to_EH),
    .from_EI(Tile_X2Y19_to_EI),
    .from_SA(Tile_X3Y18_to_SA),
    .from_SB(Tile_X3Y18_to_SB),
    .from_SC(Tile_X3Y18_to_SC),
    .from_SD(Tile_X3Y18_to_SD),
    .from_SF(Tile_X3Y18_to_SF),
    .from_SG(Tile_X3Y18_to_SG),
    .from_SH(Tile_X3Y18_to_SH),
    .from_SI(Tile_X3Y18_to_SI),
    .from_WA(Tile_X4Y19_to_WA),
    .from_WB(Tile_X4Y19_to_WB),
    .from_WC(Tile_X4Y19_to_WC),
    .from_WD(Tile_X4Y19_to_WD),
    .from_WF(Tile_X4Y19_to_WF),
    .from_WG(Tile_X4Y19_to_WG),
    .from_WH(Tile_X4Y19_to_WH),
    .from_WI(Tile_X4Y19_to_WI),
    .to_EA(Tile_X3Y19_to_EA),
    .to_EB(Tile_X3Y19_to_EB),
    .to_EC(Tile_X3Y19_to_EC),
    .to_ED(Tile_X3Y19_to_ED),
    .to_EF(Tile_X3Y19_to_EF),
    .to_EG(Tile_X3Y19_to_EG),
    .to_EH(Tile_X3Y19_to_EH),
    .to_EI(Tile_X3Y19_to_EI),
    .to_WA(Tile_X3Y19_to_WA),
    .to_WB(Tile_X3Y19_to_WB),
    .to_WC(Tile_X3Y19_to_WC),
    .to_WD(Tile_X3Y19_to_WD),
    .to_WF(Tile_X3Y19_to_WF),
    .to_WG(Tile_X3Y19_to_WG),
    .to_WH(Tile_X3Y19_to_WH),
    .to_WI(Tile_X3Y19_to_WI),
    .to_NA(Tile_X3Y19_to_NA),
    .to_NB(Tile_X3Y19_to_NB),
    .to_NC(Tile_X3Y19_to_NC),
    .to_ND(Tile_X3Y19_to_ND),
    .to_NF(Tile_X3Y19_to_NF),
    .to_NG(Tile_X3Y19_to_NG),
    .to_NH(Tile_X3Y19_to_NH),
    .to_NI(Tile_X3Y19_to_NI),
    .to_SA(Tile_X3Y19_to_SA),
    .to_SB(Tile_X3Y19_to_SB),
    .to_SC(Tile_X3Y19_to_SC),
    .to_SD(Tile_X3Y19_to_SD),
    .to_SF(Tile_X3Y19_to_SF),
    .to_SG(Tile_X3Y19_to_SG),
    .to_SH(Tile_X3Y19_to_SH),
    .to_SI(Tile_X3Y19_to_SI),
    .R_t(Tile_X3Y19_R_t),
    .R_f(Tile_X3Y19_R_f),
    .F_masked1(Tile_X3Y19_F_masked1),
    .F_masked2(Tile_X3Y19_F_masked2),
    .UserCLK(Tile_X3Y20_UserCLKo),
    .UserCLKo(Tile_X3Y19_UserCLKo),
    .rst(Tile_X3Y20_rsto),
    .rsto(Tile_X3Y19_rsto),
    .FrameData(Tile_X2Y19_FrameData_O),
    .FrameData_O(Tile_X3Y19_FrameData_O),
    .FrameStrobe(Tile_X3Y20_FrameStrobe_O),
    .FrameStrobe_O(Tile_X3Y19_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X4Y19_Emulate_Bitstream)
    )
`endif
    Tile_X4Y19_linear_LMDPL
    (
    .from_NA(Tile_X4Y20_to_NA),
    .from_NB(Tile_X4Y20_to_NB),
    .from_NC(Tile_X4Y20_to_NC),
    .from_ND(Tile_X4Y20_to_ND),
    .from_NF(Tile_X4Y20_to_NF),
    .from_NG(Tile_X4Y20_to_NG),
    .from_NH(Tile_X4Y20_to_NH),
    .from_NI(Tile_X4Y20_to_NI),
    .from_EA(Tile_X3Y19_to_EA),
    .from_EB(Tile_X3Y19_to_EB),
    .from_EC(Tile_X3Y19_to_EC),
    .from_ED(Tile_X3Y19_to_ED),
    .from_EF(Tile_X3Y19_to_EF),
    .from_EG(Tile_X3Y19_to_EG),
    .from_EH(Tile_X3Y19_to_EH),
    .from_EI(Tile_X3Y19_to_EI),
    .from_SA(Tile_X4Y18_to_SA),
    .from_SB(Tile_X4Y18_to_SB),
    .from_SC(Tile_X4Y18_to_SC),
    .from_SD(Tile_X4Y18_to_SD),
    .from_SF(Tile_X4Y18_to_SF),
    .from_SG(Tile_X4Y18_to_SG),
    .from_SH(Tile_X4Y18_to_SH),
    .from_SI(Tile_X4Y18_to_SI),
    .from_WA(Tile_X5Y19_to_WA),
    .from_WB(Tile_X5Y19_to_WB),
    .from_WC(Tile_X5Y19_to_WC),
    .from_WD(Tile_X5Y19_to_WD),
    .from_WF(Tile_X5Y19_to_WF),
    .from_WG(Tile_X5Y19_to_WG),
    .from_WH(Tile_X5Y19_to_WH),
    .from_WI(Tile_X5Y19_to_WI),
    .to_EA(Tile_X4Y19_to_EA),
    .to_EB(Tile_X4Y19_to_EB),
    .to_EC(Tile_X4Y19_to_EC),
    .to_ED(Tile_X4Y19_to_ED),
    .to_EF(Tile_X4Y19_to_EF),
    .to_EG(Tile_X4Y19_to_EG),
    .to_EH(Tile_X4Y19_to_EH),
    .to_EI(Tile_X4Y19_to_EI),
    .to_WA(Tile_X4Y19_to_WA),
    .to_WB(Tile_X4Y19_to_WB),
    .to_WC(Tile_X4Y19_to_WC),
    .to_WD(Tile_X4Y19_to_WD),
    .to_WF(Tile_X4Y19_to_WF),
    .to_WG(Tile_X4Y19_to_WG),
    .to_WH(Tile_X4Y19_to_WH),
    .to_WI(Tile_X4Y19_to_WI),
    .to_NA(Tile_X4Y19_to_NA),
    .to_NB(Tile_X4Y19_to_NB),
    .to_NC(Tile_X4Y19_to_NC),
    .to_ND(Tile_X4Y19_to_ND),
    .to_NF(Tile_X4Y19_to_NF),
    .to_NG(Tile_X4Y19_to_NG),
    .to_NH(Tile_X4Y19_to_NH),
    .to_NI(Tile_X4Y19_to_NI),
    .to_SA(Tile_X4Y19_to_SA),
    .to_SB(Tile_X4Y19_to_SB),
    .to_SC(Tile_X4Y19_to_SC),
    .to_SD(Tile_X4Y19_to_SD),
    .to_SF(Tile_X4Y19_to_SF),
    .to_SG(Tile_X4Y19_to_SG),
    .to_SH(Tile_X4Y19_to_SH),
    .to_SI(Tile_X4Y19_to_SI),
    .F_masked1(Tile_X4Y19_F_masked1),
    .F_masked2(Tile_X4Y19_F_masked2),
    .UserCLK(Tile_X4Y20_UserCLKo),
    .UserCLKo(Tile_X4Y19_UserCLKo),
    .rst(Tile_X4Y20_rsto),
    .rsto(Tile_X4Y19_rsto),
    .FrameData(Tile_X3Y19_FrameData_O),
    .FrameData_O(Tile_X4Y19_FrameData_O),
    .FrameStrobe(Tile_X4Y20_FrameStrobe_O),
    .FrameStrobe_O(Tile_X4Y19_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X5Y19_Emulate_Bitstream)
    )
`endif
    Tile_X5Y19_linear_LMDPL
    (
    .from_NA(Tile_X5Y20_to_NA),
    .from_NB(Tile_X5Y20_to_NB),
    .from_NC(Tile_X5Y20_to_NC),
    .from_ND(Tile_X5Y20_to_ND),
    .from_NF(Tile_X5Y20_to_NF),
    .from_NG(Tile_X5Y20_to_NG),
    .from_NH(Tile_X5Y20_to_NH),
    .from_NI(Tile_X5Y20_to_NI),
    .from_EA(Tile_X4Y19_to_EA),
    .from_EB(Tile_X4Y19_to_EB),
    .from_EC(Tile_X4Y19_to_EC),
    .from_ED(Tile_X4Y19_to_ED),
    .from_EF(Tile_X4Y19_to_EF),
    .from_EG(Tile_X4Y19_to_EG),
    .from_EH(Tile_X4Y19_to_EH),
    .from_EI(Tile_X4Y19_to_EI),
    .from_SA(Tile_X5Y18_to_SA),
    .from_SB(Tile_X5Y18_to_SB),
    .from_SC(Tile_X5Y18_to_SC),
    .from_SD(Tile_X5Y18_to_SD),
    .from_SF(Tile_X5Y18_to_SF),
    .from_SG(Tile_X5Y18_to_SG),
    .from_SH(Tile_X5Y18_to_SH),
    .from_SI(Tile_X5Y18_to_SI),
    .from_WA(Tile_X6Y19_to_WA),
    .from_WB(Tile_X6Y19_to_WB),
    .from_WC(Tile_X6Y19_to_WC),
    .from_WD(Tile_X6Y19_to_WD),
    .from_WF(Tile_X6Y19_to_WF),
    .from_WG(Tile_X6Y19_to_WG),
    .from_WH(Tile_X6Y19_to_WH),
    .from_WI(Tile_X6Y19_to_WI),
    .to_EA(Tile_X5Y19_to_EA),
    .to_EB(Tile_X5Y19_to_EB),
    .to_EC(Tile_X5Y19_to_EC),
    .to_ED(Tile_X5Y19_to_ED),
    .to_EF(Tile_X5Y19_to_EF),
    .to_EG(Tile_X5Y19_to_EG),
    .to_EH(Tile_X5Y19_to_EH),
    .to_EI(Tile_X5Y19_to_EI),
    .to_WA(Tile_X5Y19_to_WA),
    .to_WB(Tile_X5Y19_to_WB),
    .to_WC(Tile_X5Y19_to_WC),
    .to_WD(Tile_X5Y19_to_WD),
    .to_WF(Tile_X5Y19_to_WF),
    .to_WG(Tile_X5Y19_to_WG),
    .to_WH(Tile_X5Y19_to_WH),
    .to_WI(Tile_X5Y19_to_WI),
    .to_NA(Tile_X5Y19_to_NA),
    .to_NB(Tile_X5Y19_to_NB),
    .to_NC(Tile_X5Y19_to_NC),
    .to_ND(Tile_X5Y19_to_ND),
    .to_NF(Tile_X5Y19_to_NF),
    .to_NG(Tile_X5Y19_to_NG),
    .to_NH(Tile_X5Y19_to_NH),
    .to_NI(Tile_X5Y19_to_NI),
    .to_SA(Tile_X5Y19_to_SA),
    .to_SB(Tile_X5Y19_to_SB),
    .to_SC(Tile_X5Y19_to_SC),
    .to_SD(Tile_X5Y19_to_SD),
    .to_SF(Tile_X5Y19_to_SF),
    .to_SG(Tile_X5Y19_to_SG),
    .to_SH(Tile_X5Y19_to_SH),
    .to_SI(Tile_X5Y19_to_SI),
    .F_masked1(Tile_X5Y19_F_masked1),
    .F_masked2(Tile_X5Y19_F_masked2),
    .UserCLK(Tile_X5Y20_UserCLKo),
    .UserCLKo(Tile_X5Y19_UserCLKo),
    .rst(Tile_X5Y20_rsto),
    .rsto(Tile_X5Y19_rsto),
    .FrameData(Tile_X4Y19_FrameData_O),
    .FrameData_O(Tile_X5Y19_FrameData_O),
    .FrameStrobe(Tile_X5Y20_FrameStrobe_O),
    .FrameStrobe_O(Tile_X5Y19_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
nonlinear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X6Y19_Emulate_Bitstream)
    )
`endif
    Tile_X6Y19_nonlinear_LMDPL
    (
    .from_NA(Tile_X6Y20_to_NA),
    .from_NB(Tile_X6Y20_to_NB),
    .from_NC(Tile_X6Y20_to_NC),
    .from_ND(Tile_X6Y20_to_ND),
    .from_NF(Tile_X6Y20_to_NF),
    .from_NG(Tile_X6Y20_to_NG),
    .from_NH(Tile_X6Y20_to_NH),
    .from_NI(Tile_X6Y20_to_NI),
    .from_EA(Tile_X5Y19_to_EA),
    .from_EB(Tile_X5Y19_to_EB),
    .from_EC(Tile_X5Y19_to_EC),
    .from_ED(Tile_X5Y19_to_ED),
    .from_EF(Tile_X5Y19_to_EF),
    .from_EG(Tile_X5Y19_to_EG),
    .from_EH(Tile_X5Y19_to_EH),
    .from_EI(Tile_X5Y19_to_EI),
    .from_SA(Tile_X6Y18_to_SA),
    .from_SB(Tile_X6Y18_to_SB),
    .from_SC(Tile_X6Y18_to_SC),
    .from_SD(Tile_X6Y18_to_SD),
    .from_SF(Tile_X6Y18_to_SF),
    .from_SG(Tile_X6Y18_to_SG),
    .from_SH(Tile_X6Y18_to_SH),
    .from_SI(Tile_X6Y18_to_SI),
    .from_WA(Tile_X7Y19_to_WA),
    .from_WB(Tile_X7Y19_to_WB),
    .from_WC(Tile_X7Y19_to_WC),
    .from_WD(Tile_X7Y19_to_WD),
    .from_WF(Tile_X7Y19_to_WF),
    .from_WG(Tile_X7Y19_to_WG),
    .from_WH(Tile_X7Y19_to_WH),
    .from_WI(Tile_X7Y19_to_WI),
    .to_EA(Tile_X6Y19_to_EA),
    .to_EB(Tile_X6Y19_to_EB),
    .to_EC(Tile_X6Y19_to_EC),
    .to_ED(Tile_X6Y19_to_ED),
    .to_EF(Tile_X6Y19_to_EF),
    .to_EG(Tile_X6Y19_to_EG),
    .to_EH(Tile_X6Y19_to_EH),
    .to_EI(Tile_X6Y19_to_EI),
    .to_WA(Tile_X6Y19_to_WA),
    .to_WB(Tile_X6Y19_to_WB),
    .to_WC(Tile_X6Y19_to_WC),
    .to_WD(Tile_X6Y19_to_WD),
    .to_WF(Tile_X6Y19_to_WF),
    .to_WG(Tile_X6Y19_to_WG),
    .to_WH(Tile_X6Y19_to_WH),
    .to_WI(Tile_X6Y19_to_WI),
    .to_NA(Tile_X6Y19_to_NA),
    .to_NB(Tile_X6Y19_to_NB),
    .to_NC(Tile_X6Y19_to_NC),
    .to_ND(Tile_X6Y19_to_ND),
    .to_NF(Tile_X6Y19_to_NF),
    .to_NG(Tile_X6Y19_to_NG),
    .to_NH(Tile_X6Y19_to_NH),
    .to_NI(Tile_X6Y19_to_NI),
    .to_SA(Tile_X6Y19_to_SA),
    .to_SB(Tile_X6Y19_to_SB),
    .to_SC(Tile_X6Y19_to_SC),
    .to_SD(Tile_X6Y19_to_SD),
    .to_SF(Tile_X6Y19_to_SF),
    .to_SG(Tile_X6Y19_to_SG),
    .to_SH(Tile_X6Y19_to_SH),
    .to_SI(Tile_X6Y19_to_SI),
    .R_t(Tile_X6Y19_R_t),
    .R_f(Tile_X6Y19_R_f),
    .F_masked1(Tile_X6Y19_F_masked1),
    .F_masked2(Tile_X6Y19_F_masked2),
    .UserCLK(Tile_X6Y20_UserCLKo),
    .UserCLKo(Tile_X6Y19_UserCLKo),
    .rst(Tile_X6Y20_rsto),
    .rsto(Tile_X6Y19_rsto),
    .FrameData(Tile_X5Y19_FrameData_O),
    .FrameData_O(Tile_X6Y19_FrameData_O),
    .FrameStrobe(Tile_X6Y20_FrameStrobe_O),
    .FrameStrobe_O(Tile_X6Y19_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X7Y19_Emulate_Bitstream)
    )
`endif
    Tile_X7Y19_linear_LMDPL
    (
    .from_NA(Tile_X7Y20_to_NA),
    .from_NB(Tile_X7Y20_to_NB),
    .from_NC(Tile_X7Y20_to_NC),
    .from_ND(Tile_X7Y20_to_ND),
    .from_NF(Tile_X7Y20_to_NF),
    .from_NG(Tile_X7Y20_to_NG),
    .from_NH(Tile_X7Y20_to_NH),
    .from_NI(Tile_X7Y20_to_NI),
    .from_EA(Tile_X6Y19_to_EA),
    .from_EB(Tile_X6Y19_to_EB),
    .from_EC(Tile_X6Y19_to_EC),
    .from_ED(Tile_X6Y19_to_ED),
    .from_EF(Tile_X6Y19_to_EF),
    .from_EG(Tile_X6Y19_to_EG),
    .from_EH(Tile_X6Y19_to_EH),
    .from_EI(Tile_X6Y19_to_EI),
    .from_SA(Tile_X7Y18_to_SA),
    .from_SB(Tile_X7Y18_to_SB),
    .from_SC(Tile_X7Y18_to_SC),
    .from_SD(Tile_X7Y18_to_SD),
    .from_SF(Tile_X7Y18_to_SF),
    .from_SG(Tile_X7Y18_to_SG),
    .from_SH(Tile_X7Y18_to_SH),
    .from_SI(Tile_X7Y18_to_SI),
    .from_WA(Tile_X8Y19_to_WA),
    .from_WB(Tile_X8Y19_to_WB),
    .from_WC(Tile_X8Y19_to_WC),
    .from_WD(Tile_X8Y19_to_WD),
    .from_WF(Tile_X8Y19_to_WF),
    .from_WG(Tile_X8Y19_to_WG),
    .from_WH(Tile_X8Y19_to_WH),
    .from_WI(Tile_X8Y19_to_WI),
    .to_EA(Tile_X7Y19_to_EA),
    .to_EB(Tile_X7Y19_to_EB),
    .to_EC(Tile_X7Y19_to_EC),
    .to_ED(Tile_X7Y19_to_ED),
    .to_EF(Tile_X7Y19_to_EF),
    .to_EG(Tile_X7Y19_to_EG),
    .to_EH(Tile_X7Y19_to_EH),
    .to_EI(Tile_X7Y19_to_EI),
    .to_WA(Tile_X7Y19_to_WA),
    .to_WB(Tile_X7Y19_to_WB),
    .to_WC(Tile_X7Y19_to_WC),
    .to_WD(Tile_X7Y19_to_WD),
    .to_WF(Tile_X7Y19_to_WF),
    .to_WG(Tile_X7Y19_to_WG),
    .to_WH(Tile_X7Y19_to_WH),
    .to_WI(Tile_X7Y19_to_WI),
    .to_NA(Tile_X7Y19_to_NA),
    .to_NB(Tile_X7Y19_to_NB),
    .to_NC(Tile_X7Y19_to_NC),
    .to_ND(Tile_X7Y19_to_ND),
    .to_NF(Tile_X7Y19_to_NF),
    .to_NG(Tile_X7Y19_to_NG),
    .to_NH(Tile_X7Y19_to_NH),
    .to_NI(Tile_X7Y19_to_NI),
    .to_SA(Tile_X7Y19_to_SA),
    .to_SB(Tile_X7Y19_to_SB),
    .to_SC(Tile_X7Y19_to_SC),
    .to_SD(Tile_X7Y19_to_SD),
    .to_SF(Tile_X7Y19_to_SF),
    .to_SG(Tile_X7Y19_to_SG),
    .to_SH(Tile_X7Y19_to_SH),
    .to_SI(Tile_X7Y19_to_SI),
    .F_masked1(Tile_X7Y19_F_masked1),
    .F_masked2(Tile_X7Y19_F_masked2),
    .UserCLK(Tile_X7Y20_UserCLKo),
    .UserCLKo(Tile_X7Y19_UserCLKo),
    .rst(Tile_X7Y20_rsto),
    .rsto(Tile_X7Y19_rsto),
    .FrameData(Tile_X6Y19_FrameData_O),
    .FrameData_O(Tile_X7Y19_FrameData_O),
    .FrameStrobe(Tile_X7Y20_FrameStrobe_O),
    .FrameStrobe_O(Tile_X7Y19_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
ctrl_to_sec
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X8Y19_Emulate_Bitstream)
    )
`endif
    Tile_X8Y19_ctrl_to_sec
    (
    .from_NA(Tile_X8Y20_to_NA),
    .from_NB(Tile_X8Y20_to_NB),
    .from_NC(Tile_X8Y20_to_NC),
    .from_ND(Tile_X8Y20_to_ND),
    .from_NF(Tile_X8Y20_to_NF),
    .from_NG(Tile_X8Y20_to_NG),
    .from_NH(Tile_X8Y20_to_NH),
    .from_NI(Tile_X8Y20_to_NI),
    .from_EA(Tile_X7Y19_to_EA),
    .from_EB(Tile_X7Y19_to_EB),
    .from_EC(Tile_X7Y19_to_EC),
    .from_ED(Tile_X7Y19_to_ED),
    .from_EF(Tile_X7Y19_to_EF),
    .from_EG(Tile_X7Y19_to_EG),
    .from_EH(Tile_X7Y19_to_EH),
    .from_EI(Tile_X7Y19_to_EI),
    .from_SA(Tile_X8Y18_to_SA),
    .from_SB(Tile_X8Y18_to_SB),
    .from_SC(Tile_X8Y18_to_SC),
    .from_SD(Tile_X8Y18_to_SD),
    .from_SF(Tile_X8Y18_to_SF),
    .from_SG(Tile_X8Y18_to_SG),
    .from_SH(Tile_X8Y18_to_SH),
    .from_SI(Tile_X8Y18_to_SI),
    .from_WA_1s(Tile_X9Y19_to_WA_1s),
    .from_WB_1s(Tile_X9Y19_to_WB_1s),
    .from_WC_1s(Tile_X9Y19_to_WC_1s),
    .from_WD_1s(Tile_X9Y19_to_WD_1s),
    .from_WF_1s(Tile_X9Y19_to_WF_1s),
    .from_WG_1s(Tile_X9Y19_to_WG_1s),
    .from_WH_1s(Tile_X9Y19_to_WH_1s),
    .from_WI_1s(Tile_X9Y19_to_WI_1s),
    .to_WA(Tile_X8Y19_to_WA),
    .to_WB(Tile_X8Y19_to_WB),
    .to_WC(Tile_X8Y19_to_WC),
    .to_WD(Tile_X8Y19_to_WD),
    .to_WF(Tile_X8Y19_to_WF),
    .to_WG(Tile_X8Y19_to_WG),
    .to_WH(Tile_X8Y19_to_WH),
    .to_WI(Tile_X8Y19_to_WI),
    .to_NA(Tile_X8Y19_to_NA),
    .to_NB(Tile_X8Y19_to_NB),
    .to_NC(Tile_X8Y19_to_NC),
    .to_ND(Tile_X8Y19_to_ND),
    .to_NF(Tile_X8Y19_to_NF),
    .to_NG(Tile_X8Y19_to_NG),
    .to_NH(Tile_X8Y19_to_NH),
    .to_NI(Tile_X8Y19_to_NI),
    .to_SA(Tile_X8Y19_to_SA),
    .to_SB(Tile_X8Y19_to_SB),
    .to_SC(Tile_X8Y19_to_SC),
    .to_SD(Tile_X8Y19_to_SD),
    .to_SF(Tile_X8Y19_to_SF),
    .to_SG(Tile_X8Y19_to_SG),
    .to_SH(Tile_X8Y19_to_SH),
    .to_SI(Tile_X8Y19_to_SI),
    .UserCLK(Tile_X8Y20_UserCLKo),
    .UserCLKo(Tile_X8Y19_UserCLKo),
    .rst(Tile_X8Y20_rsto),
    .rsto(Tile_X8Y19_rsto),
    .FrameData(Tile_X7Y19_FrameData_O),
    .FrameData_O(Tile_X8Y19_FrameData_O),
    .FrameStrobe(Tile_X8Y20_FrameStrobe_O),
    .FrameStrobe_O(Tile_X8Y19_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
combined_WDDL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X9Y19_Emulate_Bitstream)
    )
`endif
    Tile_X9Y19_combined_WDDL
    (
    .from_NA_1s(Tile_X9Y20_to_NA_1s),
    .from_NB_1s(Tile_X9Y20_to_NB_1s),
    .from_NC_1s(Tile_X9Y20_to_NC_1s),
    .from_ND_1s(Tile_X9Y20_to_ND_1s),
    .from_NF_1s(Tile_X9Y20_to_NF_1s),
    .from_NG_1s(Tile_X9Y20_to_NG_1s),
    .from_NH_1s(Tile_X9Y20_to_NH_1s),
    .from_NI_1s(Tile_X9Y20_to_NI_1s),
    .from_SA_1s(Tile_X9Y18_to_SA_1s),
    .from_SB_1s(Tile_X9Y18_to_SB_1s),
    .from_SC_1s(Tile_X9Y18_to_SC_1s),
    .from_SD_1s(Tile_X9Y18_to_SD_1s),
    .from_SF_1s(Tile_X9Y18_to_SF_1s),
    .from_SG_1s(Tile_X9Y18_to_SG_1s),
    .from_SH_1s(Tile_X9Y18_to_SH_1s),
    .from_SI_1s(Tile_X9Y18_to_SI_1s),
    .from_WA_1s(Tile_X10Y19_to_WA_1s),
    .from_WB_1s(Tile_X10Y19_to_WB_1s),
    .from_WC_1s(Tile_X10Y19_to_WC_1s),
    .from_WD_1s(Tile_X10Y19_to_WD_1s),
    .from_WF_1s(Tile_X10Y19_to_WF_1s),
    .from_WG_1s(Tile_X10Y19_to_WG_1s),
    .from_WH_1s(Tile_X10Y19_to_WH_1s),
    .from_WI_1s(Tile_X10Y19_to_WI_1s),
    .to_EA_1s(Tile_X9Y19_to_EA_1s),
    .to_EB_1s(Tile_X9Y19_to_EB_1s),
    .to_EC_1s(Tile_X9Y19_to_EC_1s),
    .to_ED_1s(Tile_X9Y19_to_ED_1s),
    .to_EF_1s(Tile_X9Y19_to_EF_1s),
    .to_EG_1s(Tile_X9Y19_to_EG_1s),
    .to_EH_1s(Tile_X9Y19_to_EH_1s),
    .to_EI_1s(Tile_X9Y19_to_EI_1s),
    .to_WA_1s(Tile_X9Y19_to_WA_1s),
    .to_WB_1s(Tile_X9Y19_to_WB_1s),
    .to_WC_1s(Tile_X9Y19_to_WC_1s),
    .to_WD_1s(Tile_X9Y19_to_WD_1s),
    .to_WF_1s(Tile_X9Y19_to_WF_1s),
    .to_WG_1s(Tile_X9Y19_to_WG_1s),
    .to_WH_1s(Tile_X9Y19_to_WH_1s),
    .to_WI_1s(Tile_X9Y19_to_WI_1s),
    .to_NA_1s(Tile_X9Y19_to_NA_1s),
    .to_NB_1s(Tile_X9Y19_to_NB_1s),
    .to_NC_1s(Tile_X9Y19_to_NC_1s),
    .to_ND_1s(Tile_X9Y19_to_ND_1s),
    .to_NF_1s(Tile_X9Y19_to_NF_1s),
    .to_NG_1s(Tile_X9Y19_to_NG_1s),
    .to_NH_1s(Tile_X9Y19_to_NH_1s),
    .to_NI_1s(Tile_X9Y19_to_NI_1s),
    .to_SA_1s(Tile_X9Y19_to_SA_1s),
    .to_SB_1s(Tile_X9Y19_to_SB_1s),
    .to_SC_1s(Tile_X9Y19_to_SC_1s),
    .to_SD_1s(Tile_X9Y19_to_SD_1s),
    .to_SF_1s(Tile_X9Y19_to_SF_1s),
    .to_SG_1s(Tile_X9Y19_to_SG_1s),
    .to_SH_1s(Tile_X9Y19_to_SH_1s),
    .to_SI_1s(Tile_X9Y19_to_SI_1s),
    .F_ctrl(Tile_X9Y19_F_ctrl),
    .UserCLK(Tile_X9Y20_UserCLKo),
    .UserCLKo(Tile_X9Y19_UserCLKo),
    .rst(Tile_X9Y20_rsto),
    .rsto(Tile_X9Y19_rsto),
    .FrameData(Tile_X8Y19_FrameData_O),
    .FrameData_O(Tile_X9Y19_FrameData_O),
    .FrameStrobe(Tile_X9Y20_FrameStrobe_O),
    .FrameStrobe_O(Tile_X9Y19_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
ctrl_IO
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X10Y19_Emulate_Bitstream)
    )
`endif
    Tile_X10Y19_ctrl_IO
    (
    .from_EA_1s(Tile_X9Y19_to_EA_1s),
    .from_EB_1s(Tile_X9Y19_to_EB_1s),
    .from_EC_1s(Tile_X9Y19_to_EC_1s),
    .from_ED_1s(Tile_X9Y19_to_ED_1s),
    .from_EF_1s(Tile_X9Y19_to_EF_1s),
    .from_EG_1s(Tile_X9Y19_to_EG_1s),
    .from_EH_1s(Tile_X9Y19_to_EH_1s),
    .from_EI_1s(Tile_X9Y19_to_EI_1s),
    .to_WA_1s(Tile_X10Y19_to_WA_1s),
    .to_WB_1s(Tile_X10Y19_to_WB_1s),
    .to_WC_1s(Tile_X10Y19_to_WC_1s),
    .to_WD_1s(Tile_X10Y19_to_WD_1s),
    .to_WF_1s(Tile_X10Y19_to_WF_1s),
    .to_WG_1s(Tile_X10Y19_to_WG_1s),
    .to_WH_1s(Tile_X10Y19_to_WH_1s),
    .to_WI_1s(Tile_X10Y19_to_WI_1s),
    .A_O_top_0_t(Tile_X10Y19_A_O_top_0_t),
    .A_O_top_0_f(Tile_X10Y19_A_O_top_0_f),
    .A_prech2(Tile_X10Y19_A_prech2),
    .A_DR_fault(Tile_X10Y19_A_DR_fault),
    .A_I_top_0_t(Tile_X10Y19_A_I_top_0_t),
    .A_I_top_0_f(Tile_X10Y19_A_I_top_0_f),
    .A_T_top(Tile_X10Y19_A_T_top),
    .A_F_ctrl(Tile_X10Y19_A_F_ctrl),
    .UserCLK(Tile_X10Y20_UserCLKo),
    .UserCLKo(Tile_X10Y19_UserCLKo),
    .rst(Tile_X10Y20_rsto),
    .rsto(Tile_X10Y19_rsto),
    .FrameData(Tile_X9Y19_FrameData_O),
    .FrameData_O(Tile_X10Y19_FrameData_O),
    .FrameStrobe(Tile_X10Y20_FrameStrobe_O),
    .FrameStrobe_O(Tile_X10Y19_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
W_IO_custom
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X0Y20_Emulate_Bitstream)
    )
`endif
    Tile_X0Y20_W_IO_custom
    (
    .from_NA(Tile_X0Y21_to_NA),
    .from_NB(Tile_X0Y21_to_NB),
    .from_NC(Tile_X0Y21_to_NC),
    .from_ND(Tile_X0Y21_to_ND),
    .from_NF(Tile_X0Y21_to_NF),
    .from_NG(Tile_X0Y21_to_NG),
    .from_NH(Tile_X0Y21_to_NH),
    .from_NI(Tile_X0Y21_to_NI),
    .from_SA(Tile_X0Y19_to_SA),
    .from_SB(Tile_X0Y19_to_SB),
    .from_SC(Tile_X0Y19_to_SC),
    .from_SD(Tile_X0Y19_to_SD),
    .from_SF(Tile_X0Y19_to_SF),
    .from_SG(Tile_X0Y19_to_SG),
    .from_SH(Tile_X0Y19_to_SH),
    .from_SI(Tile_X0Y19_to_SI),
    .from_WA(Tile_X1Y20_to_WA),
    .from_WB(Tile_X1Y20_to_WB),
    .from_WC(Tile_X1Y20_to_WC),
    .from_WD(Tile_X1Y20_to_WD),
    .from_WF(Tile_X1Y20_to_WF),
    .from_WG(Tile_X1Y20_to_WG),
    .from_WH(Tile_X1Y20_to_WH),
    .from_WI(Tile_X1Y20_to_WI),
    .to_EA(Tile_X0Y20_to_EA),
    .to_EB(Tile_X0Y20_to_EB),
    .to_EC(Tile_X0Y20_to_EC),
    .to_ED(Tile_X0Y20_to_ED),
    .to_EF(Tile_X0Y20_to_EF),
    .to_EG(Tile_X0Y20_to_EG),
    .to_EH(Tile_X0Y20_to_EH),
    .to_EI(Tile_X0Y20_to_EI),
    .to_NA(Tile_X0Y20_to_NA),
    .to_NB(Tile_X0Y20_to_NB),
    .to_NC(Tile_X0Y20_to_NC),
    .to_ND(Tile_X0Y20_to_ND),
    .to_NF(Tile_X0Y20_to_NF),
    .to_NG(Tile_X0Y20_to_NG),
    .to_NH(Tile_X0Y20_to_NH),
    .to_NI(Tile_X0Y20_to_NI),
    .to_SA(Tile_X0Y20_to_SA),
    .to_SB(Tile_X0Y20_to_SB),
    .to_SC(Tile_X0Y20_to_SC),
    .to_SD(Tile_X0Y20_to_SD),
    .to_SF(Tile_X0Y20_to_SF),
    .to_SG(Tile_X0Y20_to_SG),
    .to_SH(Tile_X0Y20_to_SH),
    .to_SI(Tile_X0Y20_to_SI),
    .A_O_top_0_t(Tile_X0Y20_A_O_top_0_t),
    .A_O_top_0_f(Tile_X0Y20_A_O_top_0_f),
    .A_O_top_1_t(Tile_X0Y20_A_O_top_1_t),
    .A_O_top_1_f(Tile_X0Y20_A_O_top_1_f),
    .A_prech1(Tile_X0Y20_A_prech1),
    .A_prech2(Tile_X0Y20_A_prech2),
    .A_DR_fault(Tile_X0Y20_A_DR_fault),
    .A_I_top_0_t(Tile_X0Y20_A_I_top_0_t),
    .A_I_top_0_f(Tile_X0Y20_A_I_top_0_f),
    .A_I_top_1_t(Tile_X0Y20_A_I_top_1_t),
    .A_I_top_1_f(Tile_X0Y20_A_I_top_1_f),
    .A_T_top(Tile_X0Y20_A_T_top),
    .A_F_masked1(Tile_X0Y20_A_F_masked1),
    .A_F_masked2(Tile_X0Y20_A_F_masked2),
    .A_config_C_bit0(Tile_X0Y20_A_config_C_bit0),
    .A_config_C_bit1(Tile_X0Y20_A_config_C_bit1),
    .A_config_C_bit2(Tile_X0Y20_A_config_C_bit2),
    .A_config_C_bit3(Tile_X0Y20_A_config_C_bit3),
    .B_config_C_bit0(Tile_X0Y20_B_config_C_bit0),
    .B_config_C_bit1(Tile_X0Y20_B_config_C_bit1),
    .B_config_C_bit2(Tile_X0Y20_B_config_C_bit2),
    .B_config_C_bit3(Tile_X0Y20_B_config_C_bit3),
    .UserCLK(Tile_X0Y21_UserCLKo),
    .UserCLKo(Tile_X0Y20_UserCLKo),
    .rst(Tile_X0Y21_rsto),
    .rsto(Tile_X0Y20_rsto),
    .FrameData(Tile_Y20_FrameData),
    .FrameData_O(Tile_X0Y20_FrameData_O),
    .FrameStrobe(Tile_X0Y21_FrameStrobe_O),
    .FrameStrobe_O(Tile_X0Y20_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X1Y20_Emulate_Bitstream)
    )
`endif
    Tile_X1Y20_linear_LMDPL
    (
    .from_NA(Tile_X1Y21_to_NA),
    .from_NB(Tile_X1Y21_to_NB),
    .from_NC(Tile_X1Y21_to_NC),
    .from_ND(Tile_X1Y21_to_ND),
    .from_NF(Tile_X1Y21_to_NF),
    .from_NG(Tile_X1Y21_to_NG),
    .from_NH(Tile_X1Y21_to_NH),
    .from_NI(Tile_X1Y21_to_NI),
    .from_EA(Tile_X0Y20_to_EA),
    .from_EB(Tile_X0Y20_to_EB),
    .from_EC(Tile_X0Y20_to_EC),
    .from_ED(Tile_X0Y20_to_ED),
    .from_EF(Tile_X0Y20_to_EF),
    .from_EG(Tile_X0Y20_to_EG),
    .from_EH(Tile_X0Y20_to_EH),
    .from_EI(Tile_X0Y20_to_EI),
    .from_SA(Tile_X1Y19_to_SA),
    .from_SB(Tile_X1Y19_to_SB),
    .from_SC(Tile_X1Y19_to_SC),
    .from_SD(Tile_X1Y19_to_SD),
    .from_SF(Tile_X1Y19_to_SF),
    .from_SG(Tile_X1Y19_to_SG),
    .from_SH(Tile_X1Y19_to_SH),
    .from_SI(Tile_X1Y19_to_SI),
    .from_WA(Tile_X2Y20_to_WA),
    .from_WB(Tile_X2Y20_to_WB),
    .from_WC(Tile_X2Y20_to_WC),
    .from_WD(Tile_X2Y20_to_WD),
    .from_WF(Tile_X2Y20_to_WF),
    .from_WG(Tile_X2Y20_to_WG),
    .from_WH(Tile_X2Y20_to_WH),
    .from_WI(Tile_X2Y20_to_WI),
    .to_EA(Tile_X1Y20_to_EA),
    .to_EB(Tile_X1Y20_to_EB),
    .to_EC(Tile_X1Y20_to_EC),
    .to_ED(Tile_X1Y20_to_ED),
    .to_EF(Tile_X1Y20_to_EF),
    .to_EG(Tile_X1Y20_to_EG),
    .to_EH(Tile_X1Y20_to_EH),
    .to_EI(Tile_X1Y20_to_EI),
    .to_WA(Tile_X1Y20_to_WA),
    .to_WB(Tile_X1Y20_to_WB),
    .to_WC(Tile_X1Y20_to_WC),
    .to_WD(Tile_X1Y20_to_WD),
    .to_WF(Tile_X1Y20_to_WF),
    .to_WG(Tile_X1Y20_to_WG),
    .to_WH(Tile_X1Y20_to_WH),
    .to_WI(Tile_X1Y20_to_WI),
    .to_NA(Tile_X1Y20_to_NA),
    .to_NB(Tile_X1Y20_to_NB),
    .to_NC(Tile_X1Y20_to_NC),
    .to_ND(Tile_X1Y20_to_ND),
    .to_NF(Tile_X1Y20_to_NF),
    .to_NG(Tile_X1Y20_to_NG),
    .to_NH(Tile_X1Y20_to_NH),
    .to_NI(Tile_X1Y20_to_NI),
    .to_SA(Tile_X1Y20_to_SA),
    .to_SB(Tile_X1Y20_to_SB),
    .to_SC(Tile_X1Y20_to_SC),
    .to_SD(Tile_X1Y20_to_SD),
    .to_SF(Tile_X1Y20_to_SF),
    .to_SG(Tile_X1Y20_to_SG),
    .to_SH(Tile_X1Y20_to_SH),
    .to_SI(Tile_X1Y20_to_SI),
    .F_masked1(Tile_X1Y20_F_masked1),
    .F_masked2(Tile_X1Y20_F_masked2),
    .UserCLK(Tile_X1Y21_UserCLKo),
    .UserCLKo(Tile_X1Y20_UserCLKo),
    .rst(Tile_X1Y21_rsto),
    .rsto(Tile_X1Y20_rsto),
    .FrameData(Tile_X0Y20_FrameData_O),
    .FrameData_O(Tile_X1Y20_FrameData_O),
    .FrameStrobe(Tile_X1Y21_FrameStrobe_O),
    .FrameStrobe_O(Tile_X1Y20_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X2Y20_Emulate_Bitstream)
    )
`endif
    Tile_X2Y20_linear_LMDPL
    (
    .from_NA(Tile_X2Y21_to_NA),
    .from_NB(Tile_X2Y21_to_NB),
    .from_NC(Tile_X2Y21_to_NC),
    .from_ND(Tile_X2Y21_to_ND),
    .from_NF(Tile_X2Y21_to_NF),
    .from_NG(Tile_X2Y21_to_NG),
    .from_NH(Tile_X2Y21_to_NH),
    .from_NI(Tile_X2Y21_to_NI),
    .from_EA(Tile_X1Y20_to_EA),
    .from_EB(Tile_X1Y20_to_EB),
    .from_EC(Tile_X1Y20_to_EC),
    .from_ED(Tile_X1Y20_to_ED),
    .from_EF(Tile_X1Y20_to_EF),
    .from_EG(Tile_X1Y20_to_EG),
    .from_EH(Tile_X1Y20_to_EH),
    .from_EI(Tile_X1Y20_to_EI),
    .from_SA(Tile_X2Y19_to_SA),
    .from_SB(Tile_X2Y19_to_SB),
    .from_SC(Tile_X2Y19_to_SC),
    .from_SD(Tile_X2Y19_to_SD),
    .from_SF(Tile_X2Y19_to_SF),
    .from_SG(Tile_X2Y19_to_SG),
    .from_SH(Tile_X2Y19_to_SH),
    .from_SI(Tile_X2Y19_to_SI),
    .from_WA(Tile_X3Y20_to_WA),
    .from_WB(Tile_X3Y20_to_WB),
    .from_WC(Tile_X3Y20_to_WC),
    .from_WD(Tile_X3Y20_to_WD),
    .from_WF(Tile_X3Y20_to_WF),
    .from_WG(Tile_X3Y20_to_WG),
    .from_WH(Tile_X3Y20_to_WH),
    .from_WI(Tile_X3Y20_to_WI),
    .to_EA(Tile_X2Y20_to_EA),
    .to_EB(Tile_X2Y20_to_EB),
    .to_EC(Tile_X2Y20_to_EC),
    .to_ED(Tile_X2Y20_to_ED),
    .to_EF(Tile_X2Y20_to_EF),
    .to_EG(Tile_X2Y20_to_EG),
    .to_EH(Tile_X2Y20_to_EH),
    .to_EI(Tile_X2Y20_to_EI),
    .to_WA(Tile_X2Y20_to_WA),
    .to_WB(Tile_X2Y20_to_WB),
    .to_WC(Tile_X2Y20_to_WC),
    .to_WD(Tile_X2Y20_to_WD),
    .to_WF(Tile_X2Y20_to_WF),
    .to_WG(Tile_X2Y20_to_WG),
    .to_WH(Tile_X2Y20_to_WH),
    .to_WI(Tile_X2Y20_to_WI),
    .to_NA(Tile_X2Y20_to_NA),
    .to_NB(Tile_X2Y20_to_NB),
    .to_NC(Tile_X2Y20_to_NC),
    .to_ND(Tile_X2Y20_to_ND),
    .to_NF(Tile_X2Y20_to_NF),
    .to_NG(Tile_X2Y20_to_NG),
    .to_NH(Tile_X2Y20_to_NH),
    .to_NI(Tile_X2Y20_to_NI),
    .to_SA(Tile_X2Y20_to_SA),
    .to_SB(Tile_X2Y20_to_SB),
    .to_SC(Tile_X2Y20_to_SC),
    .to_SD(Tile_X2Y20_to_SD),
    .to_SF(Tile_X2Y20_to_SF),
    .to_SG(Tile_X2Y20_to_SG),
    .to_SH(Tile_X2Y20_to_SH),
    .to_SI(Tile_X2Y20_to_SI),
    .F_masked1(Tile_X2Y20_F_masked1),
    .F_masked2(Tile_X2Y20_F_masked2),
    .UserCLK(Tile_X2Y21_UserCLKo),
    .UserCLKo(Tile_X2Y20_UserCLKo),
    .rst(Tile_X2Y21_rsto),
    .rsto(Tile_X2Y20_rsto),
    .FrameData(Tile_X1Y20_FrameData_O),
    .FrameData_O(Tile_X2Y20_FrameData_O),
    .FrameStrobe(Tile_X2Y21_FrameStrobe_O),
    .FrameStrobe_O(Tile_X2Y20_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
nonlinear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X3Y20_Emulate_Bitstream)
    )
`endif
    Tile_X3Y20_nonlinear_LMDPL
    (
    .from_NA(Tile_X3Y21_to_NA),
    .from_NB(Tile_X3Y21_to_NB),
    .from_NC(Tile_X3Y21_to_NC),
    .from_ND(Tile_X3Y21_to_ND),
    .from_NF(Tile_X3Y21_to_NF),
    .from_NG(Tile_X3Y21_to_NG),
    .from_NH(Tile_X3Y21_to_NH),
    .from_NI(Tile_X3Y21_to_NI),
    .from_EA(Tile_X2Y20_to_EA),
    .from_EB(Tile_X2Y20_to_EB),
    .from_EC(Tile_X2Y20_to_EC),
    .from_ED(Tile_X2Y20_to_ED),
    .from_EF(Tile_X2Y20_to_EF),
    .from_EG(Tile_X2Y20_to_EG),
    .from_EH(Tile_X2Y20_to_EH),
    .from_EI(Tile_X2Y20_to_EI),
    .from_SA(Tile_X3Y19_to_SA),
    .from_SB(Tile_X3Y19_to_SB),
    .from_SC(Tile_X3Y19_to_SC),
    .from_SD(Tile_X3Y19_to_SD),
    .from_SF(Tile_X3Y19_to_SF),
    .from_SG(Tile_X3Y19_to_SG),
    .from_SH(Tile_X3Y19_to_SH),
    .from_SI(Tile_X3Y19_to_SI),
    .from_WA(Tile_X4Y20_to_WA),
    .from_WB(Tile_X4Y20_to_WB),
    .from_WC(Tile_X4Y20_to_WC),
    .from_WD(Tile_X4Y20_to_WD),
    .from_WF(Tile_X4Y20_to_WF),
    .from_WG(Tile_X4Y20_to_WG),
    .from_WH(Tile_X4Y20_to_WH),
    .from_WI(Tile_X4Y20_to_WI),
    .to_EA(Tile_X3Y20_to_EA),
    .to_EB(Tile_X3Y20_to_EB),
    .to_EC(Tile_X3Y20_to_EC),
    .to_ED(Tile_X3Y20_to_ED),
    .to_EF(Tile_X3Y20_to_EF),
    .to_EG(Tile_X3Y20_to_EG),
    .to_EH(Tile_X3Y20_to_EH),
    .to_EI(Tile_X3Y20_to_EI),
    .to_WA(Tile_X3Y20_to_WA),
    .to_WB(Tile_X3Y20_to_WB),
    .to_WC(Tile_X3Y20_to_WC),
    .to_WD(Tile_X3Y20_to_WD),
    .to_WF(Tile_X3Y20_to_WF),
    .to_WG(Tile_X3Y20_to_WG),
    .to_WH(Tile_X3Y20_to_WH),
    .to_WI(Tile_X3Y20_to_WI),
    .to_NA(Tile_X3Y20_to_NA),
    .to_NB(Tile_X3Y20_to_NB),
    .to_NC(Tile_X3Y20_to_NC),
    .to_ND(Tile_X3Y20_to_ND),
    .to_NF(Tile_X3Y20_to_NF),
    .to_NG(Tile_X3Y20_to_NG),
    .to_NH(Tile_X3Y20_to_NH),
    .to_NI(Tile_X3Y20_to_NI),
    .to_SA(Tile_X3Y20_to_SA),
    .to_SB(Tile_X3Y20_to_SB),
    .to_SC(Tile_X3Y20_to_SC),
    .to_SD(Tile_X3Y20_to_SD),
    .to_SF(Tile_X3Y20_to_SF),
    .to_SG(Tile_X3Y20_to_SG),
    .to_SH(Tile_X3Y20_to_SH),
    .to_SI(Tile_X3Y20_to_SI),
    .R_t(Tile_X3Y20_R_t),
    .R_f(Tile_X3Y20_R_f),
    .F_masked1(Tile_X3Y20_F_masked1),
    .F_masked2(Tile_X3Y20_F_masked2),
    .UserCLK(Tile_X3Y21_UserCLKo),
    .UserCLKo(Tile_X3Y20_UserCLKo),
    .rst(Tile_X3Y21_rsto),
    .rsto(Tile_X3Y20_rsto),
    .FrameData(Tile_X2Y20_FrameData_O),
    .FrameData_O(Tile_X3Y20_FrameData_O),
    .FrameStrobe(Tile_X3Y21_FrameStrobe_O),
    .FrameStrobe_O(Tile_X3Y20_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X4Y20_Emulate_Bitstream)
    )
`endif
    Tile_X4Y20_linear_LMDPL
    (
    .from_NA(Tile_X4Y21_to_NA),
    .from_NB(Tile_X4Y21_to_NB),
    .from_NC(Tile_X4Y21_to_NC),
    .from_ND(Tile_X4Y21_to_ND),
    .from_NF(Tile_X4Y21_to_NF),
    .from_NG(Tile_X4Y21_to_NG),
    .from_NH(Tile_X4Y21_to_NH),
    .from_NI(Tile_X4Y21_to_NI),
    .from_EA(Tile_X3Y20_to_EA),
    .from_EB(Tile_X3Y20_to_EB),
    .from_EC(Tile_X3Y20_to_EC),
    .from_ED(Tile_X3Y20_to_ED),
    .from_EF(Tile_X3Y20_to_EF),
    .from_EG(Tile_X3Y20_to_EG),
    .from_EH(Tile_X3Y20_to_EH),
    .from_EI(Tile_X3Y20_to_EI),
    .from_SA(Tile_X4Y19_to_SA),
    .from_SB(Tile_X4Y19_to_SB),
    .from_SC(Tile_X4Y19_to_SC),
    .from_SD(Tile_X4Y19_to_SD),
    .from_SF(Tile_X4Y19_to_SF),
    .from_SG(Tile_X4Y19_to_SG),
    .from_SH(Tile_X4Y19_to_SH),
    .from_SI(Tile_X4Y19_to_SI),
    .from_WA(Tile_X5Y20_to_WA),
    .from_WB(Tile_X5Y20_to_WB),
    .from_WC(Tile_X5Y20_to_WC),
    .from_WD(Tile_X5Y20_to_WD),
    .from_WF(Tile_X5Y20_to_WF),
    .from_WG(Tile_X5Y20_to_WG),
    .from_WH(Tile_X5Y20_to_WH),
    .from_WI(Tile_X5Y20_to_WI),
    .to_EA(Tile_X4Y20_to_EA),
    .to_EB(Tile_X4Y20_to_EB),
    .to_EC(Tile_X4Y20_to_EC),
    .to_ED(Tile_X4Y20_to_ED),
    .to_EF(Tile_X4Y20_to_EF),
    .to_EG(Tile_X4Y20_to_EG),
    .to_EH(Tile_X4Y20_to_EH),
    .to_EI(Tile_X4Y20_to_EI),
    .to_WA(Tile_X4Y20_to_WA),
    .to_WB(Tile_X4Y20_to_WB),
    .to_WC(Tile_X4Y20_to_WC),
    .to_WD(Tile_X4Y20_to_WD),
    .to_WF(Tile_X4Y20_to_WF),
    .to_WG(Tile_X4Y20_to_WG),
    .to_WH(Tile_X4Y20_to_WH),
    .to_WI(Tile_X4Y20_to_WI),
    .to_NA(Tile_X4Y20_to_NA),
    .to_NB(Tile_X4Y20_to_NB),
    .to_NC(Tile_X4Y20_to_NC),
    .to_ND(Tile_X4Y20_to_ND),
    .to_NF(Tile_X4Y20_to_NF),
    .to_NG(Tile_X4Y20_to_NG),
    .to_NH(Tile_X4Y20_to_NH),
    .to_NI(Tile_X4Y20_to_NI),
    .to_SA(Tile_X4Y20_to_SA),
    .to_SB(Tile_X4Y20_to_SB),
    .to_SC(Tile_X4Y20_to_SC),
    .to_SD(Tile_X4Y20_to_SD),
    .to_SF(Tile_X4Y20_to_SF),
    .to_SG(Tile_X4Y20_to_SG),
    .to_SH(Tile_X4Y20_to_SH),
    .to_SI(Tile_X4Y20_to_SI),
    .F_masked1(Tile_X4Y20_F_masked1),
    .F_masked2(Tile_X4Y20_F_masked2),
    .UserCLK(Tile_X4Y21_UserCLKo),
    .UserCLKo(Tile_X4Y20_UserCLKo),
    .rst(Tile_X4Y21_rsto),
    .rsto(Tile_X4Y20_rsto),
    .FrameData(Tile_X3Y20_FrameData_O),
    .FrameData_O(Tile_X4Y20_FrameData_O),
    .FrameStrobe(Tile_X4Y21_FrameStrobe_O),
    .FrameStrobe_O(Tile_X4Y20_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X5Y20_Emulate_Bitstream)
    )
`endif
    Tile_X5Y20_linear_LMDPL
    (
    .from_NA(Tile_X5Y21_to_NA),
    .from_NB(Tile_X5Y21_to_NB),
    .from_NC(Tile_X5Y21_to_NC),
    .from_ND(Tile_X5Y21_to_ND),
    .from_NF(Tile_X5Y21_to_NF),
    .from_NG(Tile_X5Y21_to_NG),
    .from_NH(Tile_X5Y21_to_NH),
    .from_NI(Tile_X5Y21_to_NI),
    .from_EA(Tile_X4Y20_to_EA),
    .from_EB(Tile_X4Y20_to_EB),
    .from_EC(Tile_X4Y20_to_EC),
    .from_ED(Tile_X4Y20_to_ED),
    .from_EF(Tile_X4Y20_to_EF),
    .from_EG(Tile_X4Y20_to_EG),
    .from_EH(Tile_X4Y20_to_EH),
    .from_EI(Tile_X4Y20_to_EI),
    .from_SA(Tile_X5Y19_to_SA),
    .from_SB(Tile_X5Y19_to_SB),
    .from_SC(Tile_X5Y19_to_SC),
    .from_SD(Tile_X5Y19_to_SD),
    .from_SF(Tile_X5Y19_to_SF),
    .from_SG(Tile_X5Y19_to_SG),
    .from_SH(Tile_X5Y19_to_SH),
    .from_SI(Tile_X5Y19_to_SI),
    .from_WA(Tile_X6Y20_to_WA),
    .from_WB(Tile_X6Y20_to_WB),
    .from_WC(Tile_X6Y20_to_WC),
    .from_WD(Tile_X6Y20_to_WD),
    .from_WF(Tile_X6Y20_to_WF),
    .from_WG(Tile_X6Y20_to_WG),
    .from_WH(Tile_X6Y20_to_WH),
    .from_WI(Tile_X6Y20_to_WI),
    .to_EA(Tile_X5Y20_to_EA),
    .to_EB(Tile_X5Y20_to_EB),
    .to_EC(Tile_X5Y20_to_EC),
    .to_ED(Tile_X5Y20_to_ED),
    .to_EF(Tile_X5Y20_to_EF),
    .to_EG(Tile_X5Y20_to_EG),
    .to_EH(Tile_X5Y20_to_EH),
    .to_EI(Tile_X5Y20_to_EI),
    .to_WA(Tile_X5Y20_to_WA),
    .to_WB(Tile_X5Y20_to_WB),
    .to_WC(Tile_X5Y20_to_WC),
    .to_WD(Tile_X5Y20_to_WD),
    .to_WF(Tile_X5Y20_to_WF),
    .to_WG(Tile_X5Y20_to_WG),
    .to_WH(Tile_X5Y20_to_WH),
    .to_WI(Tile_X5Y20_to_WI),
    .to_NA(Tile_X5Y20_to_NA),
    .to_NB(Tile_X5Y20_to_NB),
    .to_NC(Tile_X5Y20_to_NC),
    .to_ND(Tile_X5Y20_to_ND),
    .to_NF(Tile_X5Y20_to_NF),
    .to_NG(Tile_X5Y20_to_NG),
    .to_NH(Tile_X5Y20_to_NH),
    .to_NI(Tile_X5Y20_to_NI),
    .to_SA(Tile_X5Y20_to_SA),
    .to_SB(Tile_X5Y20_to_SB),
    .to_SC(Tile_X5Y20_to_SC),
    .to_SD(Tile_X5Y20_to_SD),
    .to_SF(Tile_X5Y20_to_SF),
    .to_SG(Tile_X5Y20_to_SG),
    .to_SH(Tile_X5Y20_to_SH),
    .to_SI(Tile_X5Y20_to_SI),
    .F_masked1(Tile_X5Y20_F_masked1),
    .F_masked2(Tile_X5Y20_F_masked2),
    .UserCLK(Tile_X5Y21_UserCLKo),
    .UserCLKo(Tile_X5Y20_UserCLKo),
    .rst(Tile_X5Y21_rsto),
    .rsto(Tile_X5Y20_rsto),
    .FrameData(Tile_X4Y20_FrameData_O),
    .FrameData_O(Tile_X5Y20_FrameData_O),
    .FrameStrobe(Tile_X5Y21_FrameStrobe_O),
    .FrameStrobe_O(Tile_X5Y20_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
nonlinear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X6Y20_Emulate_Bitstream)
    )
`endif
    Tile_X6Y20_nonlinear_LMDPL
    (
    .from_NA(Tile_X6Y21_to_NA),
    .from_NB(Tile_X6Y21_to_NB),
    .from_NC(Tile_X6Y21_to_NC),
    .from_ND(Tile_X6Y21_to_ND),
    .from_NF(Tile_X6Y21_to_NF),
    .from_NG(Tile_X6Y21_to_NG),
    .from_NH(Tile_X6Y21_to_NH),
    .from_NI(Tile_X6Y21_to_NI),
    .from_EA(Tile_X5Y20_to_EA),
    .from_EB(Tile_X5Y20_to_EB),
    .from_EC(Tile_X5Y20_to_EC),
    .from_ED(Tile_X5Y20_to_ED),
    .from_EF(Tile_X5Y20_to_EF),
    .from_EG(Tile_X5Y20_to_EG),
    .from_EH(Tile_X5Y20_to_EH),
    .from_EI(Tile_X5Y20_to_EI),
    .from_SA(Tile_X6Y19_to_SA),
    .from_SB(Tile_X6Y19_to_SB),
    .from_SC(Tile_X6Y19_to_SC),
    .from_SD(Tile_X6Y19_to_SD),
    .from_SF(Tile_X6Y19_to_SF),
    .from_SG(Tile_X6Y19_to_SG),
    .from_SH(Tile_X6Y19_to_SH),
    .from_SI(Tile_X6Y19_to_SI),
    .from_WA(Tile_X7Y20_to_WA),
    .from_WB(Tile_X7Y20_to_WB),
    .from_WC(Tile_X7Y20_to_WC),
    .from_WD(Tile_X7Y20_to_WD),
    .from_WF(Tile_X7Y20_to_WF),
    .from_WG(Tile_X7Y20_to_WG),
    .from_WH(Tile_X7Y20_to_WH),
    .from_WI(Tile_X7Y20_to_WI),
    .to_EA(Tile_X6Y20_to_EA),
    .to_EB(Tile_X6Y20_to_EB),
    .to_EC(Tile_X6Y20_to_EC),
    .to_ED(Tile_X6Y20_to_ED),
    .to_EF(Tile_X6Y20_to_EF),
    .to_EG(Tile_X6Y20_to_EG),
    .to_EH(Tile_X6Y20_to_EH),
    .to_EI(Tile_X6Y20_to_EI),
    .to_WA(Tile_X6Y20_to_WA),
    .to_WB(Tile_X6Y20_to_WB),
    .to_WC(Tile_X6Y20_to_WC),
    .to_WD(Tile_X6Y20_to_WD),
    .to_WF(Tile_X6Y20_to_WF),
    .to_WG(Tile_X6Y20_to_WG),
    .to_WH(Tile_X6Y20_to_WH),
    .to_WI(Tile_X6Y20_to_WI),
    .to_NA(Tile_X6Y20_to_NA),
    .to_NB(Tile_X6Y20_to_NB),
    .to_NC(Tile_X6Y20_to_NC),
    .to_ND(Tile_X6Y20_to_ND),
    .to_NF(Tile_X6Y20_to_NF),
    .to_NG(Tile_X6Y20_to_NG),
    .to_NH(Tile_X6Y20_to_NH),
    .to_NI(Tile_X6Y20_to_NI),
    .to_SA(Tile_X6Y20_to_SA),
    .to_SB(Tile_X6Y20_to_SB),
    .to_SC(Tile_X6Y20_to_SC),
    .to_SD(Tile_X6Y20_to_SD),
    .to_SF(Tile_X6Y20_to_SF),
    .to_SG(Tile_X6Y20_to_SG),
    .to_SH(Tile_X6Y20_to_SH),
    .to_SI(Tile_X6Y20_to_SI),
    .R_t(Tile_X6Y20_R_t),
    .R_f(Tile_X6Y20_R_f),
    .F_masked1(Tile_X6Y20_F_masked1),
    .F_masked2(Tile_X6Y20_F_masked2),
    .UserCLK(Tile_X6Y21_UserCLKo),
    .UserCLKo(Tile_X6Y20_UserCLKo),
    .rst(Tile_X6Y21_rsto),
    .rsto(Tile_X6Y20_rsto),
    .FrameData(Tile_X5Y20_FrameData_O),
    .FrameData_O(Tile_X6Y20_FrameData_O),
    .FrameStrobe(Tile_X6Y21_FrameStrobe_O),
    .FrameStrobe_O(Tile_X6Y20_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X7Y20_Emulate_Bitstream)
    )
`endif
    Tile_X7Y20_linear_LMDPL
    (
    .from_NA(Tile_X7Y21_to_NA),
    .from_NB(Tile_X7Y21_to_NB),
    .from_NC(Tile_X7Y21_to_NC),
    .from_ND(Tile_X7Y21_to_ND),
    .from_NF(Tile_X7Y21_to_NF),
    .from_NG(Tile_X7Y21_to_NG),
    .from_NH(Tile_X7Y21_to_NH),
    .from_NI(Tile_X7Y21_to_NI),
    .from_EA(Tile_X6Y20_to_EA),
    .from_EB(Tile_X6Y20_to_EB),
    .from_EC(Tile_X6Y20_to_EC),
    .from_ED(Tile_X6Y20_to_ED),
    .from_EF(Tile_X6Y20_to_EF),
    .from_EG(Tile_X6Y20_to_EG),
    .from_EH(Tile_X6Y20_to_EH),
    .from_EI(Tile_X6Y20_to_EI),
    .from_SA(Tile_X7Y19_to_SA),
    .from_SB(Tile_X7Y19_to_SB),
    .from_SC(Tile_X7Y19_to_SC),
    .from_SD(Tile_X7Y19_to_SD),
    .from_SF(Tile_X7Y19_to_SF),
    .from_SG(Tile_X7Y19_to_SG),
    .from_SH(Tile_X7Y19_to_SH),
    .from_SI(Tile_X7Y19_to_SI),
    .from_WA(Tile_X8Y20_to_WA),
    .from_WB(Tile_X8Y20_to_WB),
    .from_WC(Tile_X8Y20_to_WC),
    .from_WD(Tile_X8Y20_to_WD),
    .from_WF(Tile_X8Y20_to_WF),
    .from_WG(Tile_X8Y20_to_WG),
    .from_WH(Tile_X8Y20_to_WH),
    .from_WI(Tile_X8Y20_to_WI),
    .to_EA(Tile_X7Y20_to_EA),
    .to_EB(Tile_X7Y20_to_EB),
    .to_EC(Tile_X7Y20_to_EC),
    .to_ED(Tile_X7Y20_to_ED),
    .to_EF(Tile_X7Y20_to_EF),
    .to_EG(Tile_X7Y20_to_EG),
    .to_EH(Tile_X7Y20_to_EH),
    .to_EI(Tile_X7Y20_to_EI),
    .to_WA(Tile_X7Y20_to_WA),
    .to_WB(Tile_X7Y20_to_WB),
    .to_WC(Tile_X7Y20_to_WC),
    .to_WD(Tile_X7Y20_to_WD),
    .to_WF(Tile_X7Y20_to_WF),
    .to_WG(Tile_X7Y20_to_WG),
    .to_WH(Tile_X7Y20_to_WH),
    .to_WI(Tile_X7Y20_to_WI),
    .to_NA(Tile_X7Y20_to_NA),
    .to_NB(Tile_X7Y20_to_NB),
    .to_NC(Tile_X7Y20_to_NC),
    .to_ND(Tile_X7Y20_to_ND),
    .to_NF(Tile_X7Y20_to_NF),
    .to_NG(Tile_X7Y20_to_NG),
    .to_NH(Tile_X7Y20_to_NH),
    .to_NI(Tile_X7Y20_to_NI),
    .to_SA(Tile_X7Y20_to_SA),
    .to_SB(Tile_X7Y20_to_SB),
    .to_SC(Tile_X7Y20_to_SC),
    .to_SD(Tile_X7Y20_to_SD),
    .to_SF(Tile_X7Y20_to_SF),
    .to_SG(Tile_X7Y20_to_SG),
    .to_SH(Tile_X7Y20_to_SH),
    .to_SI(Tile_X7Y20_to_SI),
    .F_masked1(Tile_X7Y20_F_masked1),
    .F_masked2(Tile_X7Y20_F_masked2),
    .UserCLK(Tile_X7Y21_UserCLKo),
    .UserCLKo(Tile_X7Y20_UserCLKo),
    .rst(Tile_X7Y21_rsto),
    .rsto(Tile_X7Y20_rsto),
    .FrameData(Tile_X6Y20_FrameData_O),
    .FrameData_O(Tile_X7Y20_FrameData_O),
    .FrameStrobe(Tile_X7Y21_FrameStrobe_O),
    .FrameStrobe_O(Tile_X7Y20_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
ctrl_to_sec
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X8Y20_Emulate_Bitstream)
    )
`endif
    Tile_X8Y20_ctrl_to_sec
    (
    .from_NA(Tile_X8Y21_to_NA),
    .from_NB(Tile_X8Y21_to_NB),
    .from_NC(Tile_X8Y21_to_NC),
    .from_ND(Tile_X8Y21_to_ND),
    .from_NF(Tile_X8Y21_to_NF),
    .from_NG(Tile_X8Y21_to_NG),
    .from_NH(Tile_X8Y21_to_NH),
    .from_NI(Tile_X8Y21_to_NI),
    .from_EA(Tile_X7Y20_to_EA),
    .from_EB(Tile_X7Y20_to_EB),
    .from_EC(Tile_X7Y20_to_EC),
    .from_ED(Tile_X7Y20_to_ED),
    .from_EF(Tile_X7Y20_to_EF),
    .from_EG(Tile_X7Y20_to_EG),
    .from_EH(Tile_X7Y20_to_EH),
    .from_EI(Tile_X7Y20_to_EI),
    .from_SA(Tile_X8Y19_to_SA),
    .from_SB(Tile_X8Y19_to_SB),
    .from_SC(Tile_X8Y19_to_SC),
    .from_SD(Tile_X8Y19_to_SD),
    .from_SF(Tile_X8Y19_to_SF),
    .from_SG(Tile_X8Y19_to_SG),
    .from_SH(Tile_X8Y19_to_SH),
    .from_SI(Tile_X8Y19_to_SI),
    .from_WA_1s(Tile_X9Y20_to_WA_1s),
    .from_WB_1s(Tile_X9Y20_to_WB_1s),
    .from_WC_1s(Tile_X9Y20_to_WC_1s),
    .from_WD_1s(Tile_X9Y20_to_WD_1s),
    .from_WF_1s(Tile_X9Y20_to_WF_1s),
    .from_WG_1s(Tile_X9Y20_to_WG_1s),
    .from_WH_1s(Tile_X9Y20_to_WH_1s),
    .from_WI_1s(Tile_X9Y20_to_WI_1s),
    .to_WA(Tile_X8Y20_to_WA),
    .to_WB(Tile_X8Y20_to_WB),
    .to_WC(Tile_X8Y20_to_WC),
    .to_WD(Tile_X8Y20_to_WD),
    .to_WF(Tile_X8Y20_to_WF),
    .to_WG(Tile_X8Y20_to_WG),
    .to_WH(Tile_X8Y20_to_WH),
    .to_WI(Tile_X8Y20_to_WI),
    .to_NA(Tile_X8Y20_to_NA),
    .to_NB(Tile_X8Y20_to_NB),
    .to_NC(Tile_X8Y20_to_NC),
    .to_ND(Tile_X8Y20_to_ND),
    .to_NF(Tile_X8Y20_to_NF),
    .to_NG(Tile_X8Y20_to_NG),
    .to_NH(Tile_X8Y20_to_NH),
    .to_NI(Tile_X8Y20_to_NI),
    .to_SA(Tile_X8Y20_to_SA),
    .to_SB(Tile_X8Y20_to_SB),
    .to_SC(Tile_X8Y20_to_SC),
    .to_SD(Tile_X8Y20_to_SD),
    .to_SF(Tile_X8Y20_to_SF),
    .to_SG(Tile_X8Y20_to_SG),
    .to_SH(Tile_X8Y20_to_SH),
    .to_SI(Tile_X8Y20_to_SI),
    .UserCLK(Tile_X8Y21_UserCLKo),
    .UserCLKo(Tile_X8Y20_UserCLKo),
    .rst(Tile_X8Y21_rsto),
    .rsto(Tile_X8Y20_rsto),
    .FrameData(Tile_X7Y20_FrameData_O),
    .FrameData_O(Tile_X8Y20_FrameData_O),
    .FrameStrobe(Tile_X8Y21_FrameStrobe_O),
    .FrameStrobe_O(Tile_X8Y20_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
combined_WDDL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X9Y20_Emulate_Bitstream)
    )
`endif
    Tile_X9Y20_combined_WDDL
    (
    .from_NA_1s(Tile_X9Y21_to_NA_1s),
    .from_NB_1s(Tile_X9Y21_to_NB_1s),
    .from_NC_1s(Tile_X9Y21_to_NC_1s),
    .from_ND_1s(Tile_X9Y21_to_ND_1s),
    .from_NF_1s(Tile_X9Y21_to_NF_1s),
    .from_NG_1s(Tile_X9Y21_to_NG_1s),
    .from_NH_1s(Tile_X9Y21_to_NH_1s),
    .from_NI_1s(Tile_X9Y21_to_NI_1s),
    .from_SA_1s(Tile_X9Y19_to_SA_1s),
    .from_SB_1s(Tile_X9Y19_to_SB_1s),
    .from_SC_1s(Tile_X9Y19_to_SC_1s),
    .from_SD_1s(Tile_X9Y19_to_SD_1s),
    .from_SF_1s(Tile_X9Y19_to_SF_1s),
    .from_SG_1s(Tile_X9Y19_to_SG_1s),
    .from_SH_1s(Tile_X9Y19_to_SH_1s),
    .from_SI_1s(Tile_X9Y19_to_SI_1s),
    .from_WA_1s(Tile_X10Y20_to_WA_1s),
    .from_WB_1s(Tile_X10Y20_to_WB_1s),
    .from_WC_1s(Tile_X10Y20_to_WC_1s),
    .from_WD_1s(Tile_X10Y20_to_WD_1s),
    .from_WF_1s(Tile_X10Y20_to_WF_1s),
    .from_WG_1s(Tile_X10Y20_to_WG_1s),
    .from_WH_1s(Tile_X10Y20_to_WH_1s),
    .from_WI_1s(Tile_X10Y20_to_WI_1s),
    .to_EA_1s(Tile_X9Y20_to_EA_1s),
    .to_EB_1s(Tile_X9Y20_to_EB_1s),
    .to_EC_1s(Tile_X9Y20_to_EC_1s),
    .to_ED_1s(Tile_X9Y20_to_ED_1s),
    .to_EF_1s(Tile_X9Y20_to_EF_1s),
    .to_EG_1s(Tile_X9Y20_to_EG_1s),
    .to_EH_1s(Tile_X9Y20_to_EH_1s),
    .to_EI_1s(Tile_X9Y20_to_EI_1s),
    .to_WA_1s(Tile_X9Y20_to_WA_1s),
    .to_WB_1s(Tile_X9Y20_to_WB_1s),
    .to_WC_1s(Tile_X9Y20_to_WC_1s),
    .to_WD_1s(Tile_X9Y20_to_WD_1s),
    .to_WF_1s(Tile_X9Y20_to_WF_1s),
    .to_WG_1s(Tile_X9Y20_to_WG_1s),
    .to_WH_1s(Tile_X9Y20_to_WH_1s),
    .to_WI_1s(Tile_X9Y20_to_WI_1s),
    .to_NA_1s(Tile_X9Y20_to_NA_1s),
    .to_NB_1s(Tile_X9Y20_to_NB_1s),
    .to_NC_1s(Tile_X9Y20_to_NC_1s),
    .to_ND_1s(Tile_X9Y20_to_ND_1s),
    .to_NF_1s(Tile_X9Y20_to_NF_1s),
    .to_NG_1s(Tile_X9Y20_to_NG_1s),
    .to_NH_1s(Tile_X9Y20_to_NH_1s),
    .to_NI_1s(Tile_X9Y20_to_NI_1s),
    .to_SA_1s(Tile_X9Y20_to_SA_1s),
    .to_SB_1s(Tile_X9Y20_to_SB_1s),
    .to_SC_1s(Tile_X9Y20_to_SC_1s),
    .to_SD_1s(Tile_X9Y20_to_SD_1s),
    .to_SF_1s(Tile_X9Y20_to_SF_1s),
    .to_SG_1s(Tile_X9Y20_to_SG_1s),
    .to_SH_1s(Tile_X9Y20_to_SH_1s),
    .to_SI_1s(Tile_X9Y20_to_SI_1s),
    .F_ctrl(Tile_X9Y20_F_ctrl),
    .UserCLK(Tile_X9Y21_UserCLKo),
    .UserCLKo(Tile_X9Y20_UserCLKo),
    .rst(Tile_X9Y21_rsto),
    .rsto(Tile_X9Y20_rsto),
    .FrameData(Tile_X8Y20_FrameData_O),
    .FrameData_O(Tile_X9Y20_FrameData_O),
    .FrameStrobe(Tile_X9Y21_FrameStrobe_O),
    .FrameStrobe_O(Tile_X9Y20_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
ctrl_IO
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X10Y20_Emulate_Bitstream)
    )
`endif
    Tile_X10Y20_ctrl_IO
    (
    .from_EA_1s(Tile_X9Y20_to_EA_1s),
    .from_EB_1s(Tile_X9Y20_to_EB_1s),
    .from_EC_1s(Tile_X9Y20_to_EC_1s),
    .from_ED_1s(Tile_X9Y20_to_ED_1s),
    .from_EF_1s(Tile_X9Y20_to_EF_1s),
    .from_EG_1s(Tile_X9Y20_to_EG_1s),
    .from_EH_1s(Tile_X9Y20_to_EH_1s),
    .from_EI_1s(Tile_X9Y20_to_EI_1s),
    .to_WA_1s(Tile_X10Y20_to_WA_1s),
    .to_WB_1s(Tile_X10Y20_to_WB_1s),
    .to_WC_1s(Tile_X10Y20_to_WC_1s),
    .to_WD_1s(Tile_X10Y20_to_WD_1s),
    .to_WF_1s(Tile_X10Y20_to_WF_1s),
    .to_WG_1s(Tile_X10Y20_to_WG_1s),
    .to_WH_1s(Tile_X10Y20_to_WH_1s),
    .to_WI_1s(Tile_X10Y20_to_WI_1s),
    .A_O_top_0_t(Tile_X10Y20_A_O_top_0_t),
    .A_O_top_0_f(Tile_X10Y20_A_O_top_0_f),
    .A_prech2(Tile_X10Y20_A_prech2),
    .A_DR_fault(Tile_X10Y20_A_DR_fault),
    .A_I_top_0_t(Tile_X10Y20_A_I_top_0_t),
    .A_I_top_0_f(Tile_X10Y20_A_I_top_0_f),
    .A_T_top(Tile_X10Y20_A_T_top),
    .A_F_ctrl(Tile_X10Y20_A_F_ctrl),
    .UserCLK(Tile_X10Y21_UserCLKo),
    .UserCLKo(Tile_X10Y20_UserCLKo),
    .rst(Tile_X10Y21_rsto),
    .rsto(Tile_X10Y20_rsto),
    .FrameData(Tile_X9Y20_FrameData_O),
    .FrameData_O(Tile_X10Y20_FrameData_O),
    .FrameStrobe(Tile_X10Y21_FrameStrobe_O),
    .FrameStrobe_O(Tile_X10Y20_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
W_IO_custom
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X0Y21_Emulate_Bitstream)
    )
`endif
    Tile_X0Y21_W_IO_custom
    (
    .from_NA(Tile_X0Y22_to_NA),
    .from_NB(Tile_X0Y22_to_NB),
    .from_NC(Tile_X0Y22_to_NC),
    .from_ND(Tile_X0Y22_to_ND),
    .from_NF(Tile_X0Y22_to_NF),
    .from_NG(Tile_X0Y22_to_NG),
    .from_NH(Tile_X0Y22_to_NH),
    .from_NI(Tile_X0Y22_to_NI),
    .from_SA(Tile_X0Y20_to_SA),
    .from_SB(Tile_X0Y20_to_SB),
    .from_SC(Tile_X0Y20_to_SC),
    .from_SD(Tile_X0Y20_to_SD),
    .from_SF(Tile_X0Y20_to_SF),
    .from_SG(Tile_X0Y20_to_SG),
    .from_SH(Tile_X0Y20_to_SH),
    .from_SI(Tile_X0Y20_to_SI),
    .from_WA(Tile_X1Y21_to_WA),
    .from_WB(Tile_X1Y21_to_WB),
    .from_WC(Tile_X1Y21_to_WC),
    .from_WD(Tile_X1Y21_to_WD),
    .from_WF(Tile_X1Y21_to_WF),
    .from_WG(Tile_X1Y21_to_WG),
    .from_WH(Tile_X1Y21_to_WH),
    .from_WI(Tile_X1Y21_to_WI),
    .to_EA(Tile_X0Y21_to_EA),
    .to_EB(Tile_X0Y21_to_EB),
    .to_EC(Tile_X0Y21_to_EC),
    .to_ED(Tile_X0Y21_to_ED),
    .to_EF(Tile_X0Y21_to_EF),
    .to_EG(Tile_X0Y21_to_EG),
    .to_EH(Tile_X0Y21_to_EH),
    .to_EI(Tile_X0Y21_to_EI),
    .to_NA(Tile_X0Y21_to_NA),
    .to_NB(Tile_X0Y21_to_NB),
    .to_NC(Tile_X0Y21_to_NC),
    .to_ND(Tile_X0Y21_to_ND),
    .to_NF(Tile_X0Y21_to_NF),
    .to_NG(Tile_X0Y21_to_NG),
    .to_NH(Tile_X0Y21_to_NH),
    .to_NI(Tile_X0Y21_to_NI),
    .to_SA(Tile_X0Y21_to_SA),
    .to_SB(Tile_X0Y21_to_SB),
    .to_SC(Tile_X0Y21_to_SC),
    .to_SD(Tile_X0Y21_to_SD),
    .to_SF(Tile_X0Y21_to_SF),
    .to_SG(Tile_X0Y21_to_SG),
    .to_SH(Tile_X0Y21_to_SH),
    .to_SI(Tile_X0Y21_to_SI),
    .A_O_top_0_t(Tile_X0Y21_A_O_top_0_t),
    .A_O_top_0_f(Tile_X0Y21_A_O_top_0_f),
    .A_O_top_1_t(Tile_X0Y21_A_O_top_1_t),
    .A_O_top_1_f(Tile_X0Y21_A_O_top_1_f),
    .A_prech1(Tile_X0Y21_A_prech1),
    .A_prech2(Tile_X0Y21_A_prech2),
    .A_DR_fault(Tile_X0Y21_A_DR_fault),
    .A_I_top_0_t(Tile_X0Y21_A_I_top_0_t),
    .A_I_top_0_f(Tile_X0Y21_A_I_top_0_f),
    .A_I_top_1_t(Tile_X0Y21_A_I_top_1_t),
    .A_I_top_1_f(Tile_X0Y21_A_I_top_1_f),
    .A_T_top(Tile_X0Y21_A_T_top),
    .A_F_masked1(Tile_X0Y21_A_F_masked1),
    .A_F_masked2(Tile_X0Y21_A_F_masked2),
    .A_config_C_bit0(Tile_X0Y21_A_config_C_bit0),
    .A_config_C_bit1(Tile_X0Y21_A_config_C_bit1),
    .A_config_C_bit2(Tile_X0Y21_A_config_C_bit2),
    .A_config_C_bit3(Tile_X0Y21_A_config_C_bit3),
    .B_config_C_bit0(Tile_X0Y21_B_config_C_bit0),
    .B_config_C_bit1(Tile_X0Y21_B_config_C_bit1),
    .B_config_C_bit2(Tile_X0Y21_B_config_C_bit2),
    .B_config_C_bit3(Tile_X0Y21_B_config_C_bit3),
    .UserCLK(Tile_X0Y22_UserCLKo),
    .UserCLKo(Tile_X0Y21_UserCLKo),
    .rst(Tile_X0Y22_rsto),
    .rsto(Tile_X0Y21_rsto),
    .FrameData(Tile_Y21_FrameData),
    .FrameData_O(Tile_X0Y21_FrameData_O),
    .FrameStrobe(Tile_X0Y22_FrameStrobe_O),
    .FrameStrobe_O(Tile_X0Y21_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X1Y21_Emulate_Bitstream)
    )
`endif
    Tile_X1Y21_linear_LMDPL
    (
    .from_NA(Tile_X1Y22_to_NA),
    .from_NB(Tile_X1Y22_to_NB),
    .from_NC(Tile_X1Y22_to_NC),
    .from_ND(Tile_X1Y22_to_ND),
    .from_NF(Tile_X1Y22_to_NF),
    .from_NG(Tile_X1Y22_to_NG),
    .from_NH(Tile_X1Y22_to_NH),
    .from_NI(Tile_X1Y22_to_NI),
    .from_EA(Tile_X0Y21_to_EA),
    .from_EB(Tile_X0Y21_to_EB),
    .from_EC(Tile_X0Y21_to_EC),
    .from_ED(Tile_X0Y21_to_ED),
    .from_EF(Tile_X0Y21_to_EF),
    .from_EG(Tile_X0Y21_to_EG),
    .from_EH(Tile_X0Y21_to_EH),
    .from_EI(Tile_X0Y21_to_EI),
    .from_SA(Tile_X1Y20_to_SA),
    .from_SB(Tile_X1Y20_to_SB),
    .from_SC(Tile_X1Y20_to_SC),
    .from_SD(Tile_X1Y20_to_SD),
    .from_SF(Tile_X1Y20_to_SF),
    .from_SG(Tile_X1Y20_to_SG),
    .from_SH(Tile_X1Y20_to_SH),
    .from_SI(Tile_X1Y20_to_SI),
    .from_WA(Tile_X2Y21_to_WA),
    .from_WB(Tile_X2Y21_to_WB),
    .from_WC(Tile_X2Y21_to_WC),
    .from_WD(Tile_X2Y21_to_WD),
    .from_WF(Tile_X2Y21_to_WF),
    .from_WG(Tile_X2Y21_to_WG),
    .from_WH(Tile_X2Y21_to_WH),
    .from_WI(Tile_X2Y21_to_WI),
    .to_EA(Tile_X1Y21_to_EA),
    .to_EB(Tile_X1Y21_to_EB),
    .to_EC(Tile_X1Y21_to_EC),
    .to_ED(Tile_X1Y21_to_ED),
    .to_EF(Tile_X1Y21_to_EF),
    .to_EG(Tile_X1Y21_to_EG),
    .to_EH(Tile_X1Y21_to_EH),
    .to_EI(Tile_X1Y21_to_EI),
    .to_WA(Tile_X1Y21_to_WA),
    .to_WB(Tile_X1Y21_to_WB),
    .to_WC(Tile_X1Y21_to_WC),
    .to_WD(Tile_X1Y21_to_WD),
    .to_WF(Tile_X1Y21_to_WF),
    .to_WG(Tile_X1Y21_to_WG),
    .to_WH(Tile_X1Y21_to_WH),
    .to_WI(Tile_X1Y21_to_WI),
    .to_NA(Tile_X1Y21_to_NA),
    .to_NB(Tile_X1Y21_to_NB),
    .to_NC(Tile_X1Y21_to_NC),
    .to_ND(Tile_X1Y21_to_ND),
    .to_NF(Tile_X1Y21_to_NF),
    .to_NG(Tile_X1Y21_to_NG),
    .to_NH(Tile_X1Y21_to_NH),
    .to_NI(Tile_X1Y21_to_NI),
    .to_SA(Tile_X1Y21_to_SA),
    .to_SB(Tile_X1Y21_to_SB),
    .to_SC(Tile_X1Y21_to_SC),
    .to_SD(Tile_X1Y21_to_SD),
    .to_SF(Tile_X1Y21_to_SF),
    .to_SG(Tile_X1Y21_to_SG),
    .to_SH(Tile_X1Y21_to_SH),
    .to_SI(Tile_X1Y21_to_SI),
    .F_masked1(Tile_X1Y21_F_masked1),
    .F_masked2(Tile_X1Y21_F_masked2),
    .UserCLK(Tile_X1Y22_UserCLKo),
    .UserCLKo(Tile_X1Y21_UserCLKo),
    .rst(Tile_X1Y22_rsto),
    .rsto(Tile_X1Y21_rsto),
    .FrameData(Tile_X0Y21_FrameData_O),
    .FrameData_O(Tile_X1Y21_FrameData_O),
    .FrameStrobe(Tile_X1Y22_FrameStrobe_O),
    .FrameStrobe_O(Tile_X1Y21_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X2Y21_Emulate_Bitstream)
    )
`endif
    Tile_X2Y21_linear_LMDPL
    (
    .from_NA(Tile_X2Y22_to_NA),
    .from_NB(Tile_X2Y22_to_NB),
    .from_NC(Tile_X2Y22_to_NC),
    .from_ND(Tile_X2Y22_to_ND),
    .from_NF(Tile_X2Y22_to_NF),
    .from_NG(Tile_X2Y22_to_NG),
    .from_NH(Tile_X2Y22_to_NH),
    .from_NI(Tile_X2Y22_to_NI),
    .from_EA(Tile_X1Y21_to_EA),
    .from_EB(Tile_X1Y21_to_EB),
    .from_EC(Tile_X1Y21_to_EC),
    .from_ED(Tile_X1Y21_to_ED),
    .from_EF(Tile_X1Y21_to_EF),
    .from_EG(Tile_X1Y21_to_EG),
    .from_EH(Tile_X1Y21_to_EH),
    .from_EI(Tile_X1Y21_to_EI),
    .from_SA(Tile_X2Y20_to_SA),
    .from_SB(Tile_X2Y20_to_SB),
    .from_SC(Tile_X2Y20_to_SC),
    .from_SD(Tile_X2Y20_to_SD),
    .from_SF(Tile_X2Y20_to_SF),
    .from_SG(Tile_X2Y20_to_SG),
    .from_SH(Tile_X2Y20_to_SH),
    .from_SI(Tile_X2Y20_to_SI),
    .from_WA(Tile_X3Y21_to_WA),
    .from_WB(Tile_X3Y21_to_WB),
    .from_WC(Tile_X3Y21_to_WC),
    .from_WD(Tile_X3Y21_to_WD),
    .from_WF(Tile_X3Y21_to_WF),
    .from_WG(Tile_X3Y21_to_WG),
    .from_WH(Tile_X3Y21_to_WH),
    .from_WI(Tile_X3Y21_to_WI),
    .to_EA(Tile_X2Y21_to_EA),
    .to_EB(Tile_X2Y21_to_EB),
    .to_EC(Tile_X2Y21_to_EC),
    .to_ED(Tile_X2Y21_to_ED),
    .to_EF(Tile_X2Y21_to_EF),
    .to_EG(Tile_X2Y21_to_EG),
    .to_EH(Tile_X2Y21_to_EH),
    .to_EI(Tile_X2Y21_to_EI),
    .to_WA(Tile_X2Y21_to_WA),
    .to_WB(Tile_X2Y21_to_WB),
    .to_WC(Tile_X2Y21_to_WC),
    .to_WD(Tile_X2Y21_to_WD),
    .to_WF(Tile_X2Y21_to_WF),
    .to_WG(Tile_X2Y21_to_WG),
    .to_WH(Tile_X2Y21_to_WH),
    .to_WI(Tile_X2Y21_to_WI),
    .to_NA(Tile_X2Y21_to_NA),
    .to_NB(Tile_X2Y21_to_NB),
    .to_NC(Tile_X2Y21_to_NC),
    .to_ND(Tile_X2Y21_to_ND),
    .to_NF(Tile_X2Y21_to_NF),
    .to_NG(Tile_X2Y21_to_NG),
    .to_NH(Tile_X2Y21_to_NH),
    .to_NI(Tile_X2Y21_to_NI),
    .to_SA(Tile_X2Y21_to_SA),
    .to_SB(Tile_X2Y21_to_SB),
    .to_SC(Tile_X2Y21_to_SC),
    .to_SD(Tile_X2Y21_to_SD),
    .to_SF(Tile_X2Y21_to_SF),
    .to_SG(Tile_X2Y21_to_SG),
    .to_SH(Tile_X2Y21_to_SH),
    .to_SI(Tile_X2Y21_to_SI),
    .F_masked1(Tile_X2Y21_F_masked1),
    .F_masked2(Tile_X2Y21_F_masked2),
    .UserCLK(Tile_X2Y22_UserCLKo),
    .UserCLKo(Tile_X2Y21_UserCLKo),
    .rst(Tile_X2Y22_rsto),
    .rsto(Tile_X2Y21_rsto),
    .FrameData(Tile_X1Y21_FrameData_O),
    .FrameData_O(Tile_X2Y21_FrameData_O),
    .FrameStrobe(Tile_X2Y22_FrameStrobe_O),
    .FrameStrobe_O(Tile_X2Y21_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
nonlinear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X3Y21_Emulate_Bitstream)
    )
`endif
    Tile_X3Y21_nonlinear_LMDPL
    (
    .from_NA(Tile_X3Y22_to_NA),
    .from_NB(Tile_X3Y22_to_NB),
    .from_NC(Tile_X3Y22_to_NC),
    .from_ND(Tile_X3Y22_to_ND),
    .from_NF(Tile_X3Y22_to_NF),
    .from_NG(Tile_X3Y22_to_NG),
    .from_NH(Tile_X3Y22_to_NH),
    .from_NI(Tile_X3Y22_to_NI),
    .from_EA(Tile_X2Y21_to_EA),
    .from_EB(Tile_X2Y21_to_EB),
    .from_EC(Tile_X2Y21_to_EC),
    .from_ED(Tile_X2Y21_to_ED),
    .from_EF(Tile_X2Y21_to_EF),
    .from_EG(Tile_X2Y21_to_EG),
    .from_EH(Tile_X2Y21_to_EH),
    .from_EI(Tile_X2Y21_to_EI),
    .from_SA(Tile_X3Y20_to_SA),
    .from_SB(Tile_X3Y20_to_SB),
    .from_SC(Tile_X3Y20_to_SC),
    .from_SD(Tile_X3Y20_to_SD),
    .from_SF(Tile_X3Y20_to_SF),
    .from_SG(Tile_X3Y20_to_SG),
    .from_SH(Tile_X3Y20_to_SH),
    .from_SI(Tile_X3Y20_to_SI),
    .from_WA(Tile_X4Y21_to_WA),
    .from_WB(Tile_X4Y21_to_WB),
    .from_WC(Tile_X4Y21_to_WC),
    .from_WD(Tile_X4Y21_to_WD),
    .from_WF(Tile_X4Y21_to_WF),
    .from_WG(Tile_X4Y21_to_WG),
    .from_WH(Tile_X4Y21_to_WH),
    .from_WI(Tile_X4Y21_to_WI),
    .to_EA(Tile_X3Y21_to_EA),
    .to_EB(Tile_X3Y21_to_EB),
    .to_EC(Tile_X3Y21_to_EC),
    .to_ED(Tile_X3Y21_to_ED),
    .to_EF(Tile_X3Y21_to_EF),
    .to_EG(Tile_X3Y21_to_EG),
    .to_EH(Tile_X3Y21_to_EH),
    .to_EI(Tile_X3Y21_to_EI),
    .to_WA(Tile_X3Y21_to_WA),
    .to_WB(Tile_X3Y21_to_WB),
    .to_WC(Tile_X3Y21_to_WC),
    .to_WD(Tile_X3Y21_to_WD),
    .to_WF(Tile_X3Y21_to_WF),
    .to_WG(Tile_X3Y21_to_WG),
    .to_WH(Tile_X3Y21_to_WH),
    .to_WI(Tile_X3Y21_to_WI),
    .to_NA(Tile_X3Y21_to_NA),
    .to_NB(Tile_X3Y21_to_NB),
    .to_NC(Tile_X3Y21_to_NC),
    .to_ND(Tile_X3Y21_to_ND),
    .to_NF(Tile_X3Y21_to_NF),
    .to_NG(Tile_X3Y21_to_NG),
    .to_NH(Tile_X3Y21_to_NH),
    .to_NI(Tile_X3Y21_to_NI),
    .to_SA(Tile_X3Y21_to_SA),
    .to_SB(Tile_X3Y21_to_SB),
    .to_SC(Tile_X3Y21_to_SC),
    .to_SD(Tile_X3Y21_to_SD),
    .to_SF(Tile_X3Y21_to_SF),
    .to_SG(Tile_X3Y21_to_SG),
    .to_SH(Tile_X3Y21_to_SH),
    .to_SI(Tile_X3Y21_to_SI),
    .R_t(Tile_X3Y21_R_t),
    .R_f(Tile_X3Y21_R_f),
    .F_masked1(Tile_X3Y21_F_masked1),
    .F_masked2(Tile_X3Y21_F_masked2),
    .UserCLK(Tile_X3Y22_UserCLKo),
    .UserCLKo(Tile_X3Y21_UserCLKo),
    .rst(Tile_X3Y22_rsto),
    .rsto(Tile_X3Y21_rsto),
    .FrameData(Tile_X2Y21_FrameData_O),
    .FrameData_O(Tile_X3Y21_FrameData_O),
    .FrameStrobe(Tile_X3Y22_FrameStrobe_O),
    .FrameStrobe_O(Tile_X3Y21_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X4Y21_Emulate_Bitstream)
    )
`endif
    Tile_X4Y21_linear_LMDPL
    (
    .from_NA(Tile_X4Y22_to_NA),
    .from_NB(Tile_X4Y22_to_NB),
    .from_NC(Tile_X4Y22_to_NC),
    .from_ND(Tile_X4Y22_to_ND),
    .from_NF(Tile_X4Y22_to_NF),
    .from_NG(Tile_X4Y22_to_NG),
    .from_NH(Tile_X4Y22_to_NH),
    .from_NI(Tile_X4Y22_to_NI),
    .from_EA(Tile_X3Y21_to_EA),
    .from_EB(Tile_X3Y21_to_EB),
    .from_EC(Tile_X3Y21_to_EC),
    .from_ED(Tile_X3Y21_to_ED),
    .from_EF(Tile_X3Y21_to_EF),
    .from_EG(Tile_X3Y21_to_EG),
    .from_EH(Tile_X3Y21_to_EH),
    .from_EI(Tile_X3Y21_to_EI),
    .from_SA(Tile_X4Y20_to_SA),
    .from_SB(Tile_X4Y20_to_SB),
    .from_SC(Tile_X4Y20_to_SC),
    .from_SD(Tile_X4Y20_to_SD),
    .from_SF(Tile_X4Y20_to_SF),
    .from_SG(Tile_X4Y20_to_SG),
    .from_SH(Tile_X4Y20_to_SH),
    .from_SI(Tile_X4Y20_to_SI),
    .from_WA(Tile_X5Y21_to_WA),
    .from_WB(Tile_X5Y21_to_WB),
    .from_WC(Tile_X5Y21_to_WC),
    .from_WD(Tile_X5Y21_to_WD),
    .from_WF(Tile_X5Y21_to_WF),
    .from_WG(Tile_X5Y21_to_WG),
    .from_WH(Tile_X5Y21_to_WH),
    .from_WI(Tile_X5Y21_to_WI),
    .to_EA(Tile_X4Y21_to_EA),
    .to_EB(Tile_X4Y21_to_EB),
    .to_EC(Tile_X4Y21_to_EC),
    .to_ED(Tile_X4Y21_to_ED),
    .to_EF(Tile_X4Y21_to_EF),
    .to_EG(Tile_X4Y21_to_EG),
    .to_EH(Tile_X4Y21_to_EH),
    .to_EI(Tile_X4Y21_to_EI),
    .to_WA(Tile_X4Y21_to_WA),
    .to_WB(Tile_X4Y21_to_WB),
    .to_WC(Tile_X4Y21_to_WC),
    .to_WD(Tile_X4Y21_to_WD),
    .to_WF(Tile_X4Y21_to_WF),
    .to_WG(Tile_X4Y21_to_WG),
    .to_WH(Tile_X4Y21_to_WH),
    .to_WI(Tile_X4Y21_to_WI),
    .to_NA(Tile_X4Y21_to_NA),
    .to_NB(Tile_X4Y21_to_NB),
    .to_NC(Tile_X4Y21_to_NC),
    .to_ND(Tile_X4Y21_to_ND),
    .to_NF(Tile_X4Y21_to_NF),
    .to_NG(Tile_X4Y21_to_NG),
    .to_NH(Tile_X4Y21_to_NH),
    .to_NI(Tile_X4Y21_to_NI),
    .to_SA(Tile_X4Y21_to_SA),
    .to_SB(Tile_X4Y21_to_SB),
    .to_SC(Tile_X4Y21_to_SC),
    .to_SD(Tile_X4Y21_to_SD),
    .to_SF(Tile_X4Y21_to_SF),
    .to_SG(Tile_X4Y21_to_SG),
    .to_SH(Tile_X4Y21_to_SH),
    .to_SI(Tile_X4Y21_to_SI),
    .F_masked1(Tile_X4Y21_F_masked1),
    .F_masked2(Tile_X4Y21_F_masked2),
    .UserCLK(Tile_X4Y22_UserCLKo),
    .UserCLKo(Tile_X4Y21_UserCLKo),
    .rst(Tile_X4Y22_rsto),
    .rsto(Tile_X4Y21_rsto),
    .FrameData(Tile_X3Y21_FrameData_O),
    .FrameData_O(Tile_X4Y21_FrameData_O),
    .FrameStrobe(Tile_X4Y22_FrameStrobe_O),
    .FrameStrobe_O(Tile_X4Y21_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X5Y21_Emulate_Bitstream)
    )
`endif
    Tile_X5Y21_linear_LMDPL
    (
    .from_NA(Tile_X5Y22_to_NA),
    .from_NB(Tile_X5Y22_to_NB),
    .from_NC(Tile_X5Y22_to_NC),
    .from_ND(Tile_X5Y22_to_ND),
    .from_NF(Tile_X5Y22_to_NF),
    .from_NG(Tile_X5Y22_to_NG),
    .from_NH(Tile_X5Y22_to_NH),
    .from_NI(Tile_X5Y22_to_NI),
    .from_EA(Tile_X4Y21_to_EA),
    .from_EB(Tile_X4Y21_to_EB),
    .from_EC(Tile_X4Y21_to_EC),
    .from_ED(Tile_X4Y21_to_ED),
    .from_EF(Tile_X4Y21_to_EF),
    .from_EG(Tile_X4Y21_to_EG),
    .from_EH(Tile_X4Y21_to_EH),
    .from_EI(Tile_X4Y21_to_EI),
    .from_SA(Tile_X5Y20_to_SA),
    .from_SB(Tile_X5Y20_to_SB),
    .from_SC(Tile_X5Y20_to_SC),
    .from_SD(Tile_X5Y20_to_SD),
    .from_SF(Tile_X5Y20_to_SF),
    .from_SG(Tile_X5Y20_to_SG),
    .from_SH(Tile_X5Y20_to_SH),
    .from_SI(Tile_X5Y20_to_SI),
    .from_WA(Tile_X6Y21_to_WA),
    .from_WB(Tile_X6Y21_to_WB),
    .from_WC(Tile_X6Y21_to_WC),
    .from_WD(Tile_X6Y21_to_WD),
    .from_WF(Tile_X6Y21_to_WF),
    .from_WG(Tile_X6Y21_to_WG),
    .from_WH(Tile_X6Y21_to_WH),
    .from_WI(Tile_X6Y21_to_WI),
    .to_EA(Tile_X5Y21_to_EA),
    .to_EB(Tile_X5Y21_to_EB),
    .to_EC(Tile_X5Y21_to_EC),
    .to_ED(Tile_X5Y21_to_ED),
    .to_EF(Tile_X5Y21_to_EF),
    .to_EG(Tile_X5Y21_to_EG),
    .to_EH(Tile_X5Y21_to_EH),
    .to_EI(Tile_X5Y21_to_EI),
    .to_WA(Tile_X5Y21_to_WA),
    .to_WB(Tile_X5Y21_to_WB),
    .to_WC(Tile_X5Y21_to_WC),
    .to_WD(Tile_X5Y21_to_WD),
    .to_WF(Tile_X5Y21_to_WF),
    .to_WG(Tile_X5Y21_to_WG),
    .to_WH(Tile_X5Y21_to_WH),
    .to_WI(Tile_X5Y21_to_WI),
    .to_NA(Tile_X5Y21_to_NA),
    .to_NB(Tile_X5Y21_to_NB),
    .to_NC(Tile_X5Y21_to_NC),
    .to_ND(Tile_X5Y21_to_ND),
    .to_NF(Tile_X5Y21_to_NF),
    .to_NG(Tile_X5Y21_to_NG),
    .to_NH(Tile_X5Y21_to_NH),
    .to_NI(Tile_X5Y21_to_NI),
    .to_SA(Tile_X5Y21_to_SA),
    .to_SB(Tile_X5Y21_to_SB),
    .to_SC(Tile_X5Y21_to_SC),
    .to_SD(Tile_X5Y21_to_SD),
    .to_SF(Tile_X5Y21_to_SF),
    .to_SG(Tile_X5Y21_to_SG),
    .to_SH(Tile_X5Y21_to_SH),
    .to_SI(Tile_X5Y21_to_SI),
    .F_masked1(Tile_X5Y21_F_masked1),
    .F_masked2(Tile_X5Y21_F_masked2),
    .UserCLK(Tile_X5Y22_UserCLKo),
    .UserCLKo(Tile_X5Y21_UserCLKo),
    .rst(Tile_X5Y22_rsto),
    .rsto(Tile_X5Y21_rsto),
    .FrameData(Tile_X4Y21_FrameData_O),
    .FrameData_O(Tile_X5Y21_FrameData_O),
    .FrameStrobe(Tile_X5Y22_FrameStrobe_O),
    .FrameStrobe_O(Tile_X5Y21_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
nonlinear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X6Y21_Emulate_Bitstream)
    )
`endif
    Tile_X6Y21_nonlinear_LMDPL
    (
    .from_NA(Tile_X6Y22_to_NA),
    .from_NB(Tile_X6Y22_to_NB),
    .from_NC(Tile_X6Y22_to_NC),
    .from_ND(Tile_X6Y22_to_ND),
    .from_NF(Tile_X6Y22_to_NF),
    .from_NG(Tile_X6Y22_to_NG),
    .from_NH(Tile_X6Y22_to_NH),
    .from_NI(Tile_X6Y22_to_NI),
    .from_EA(Tile_X5Y21_to_EA),
    .from_EB(Tile_X5Y21_to_EB),
    .from_EC(Tile_X5Y21_to_EC),
    .from_ED(Tile_X5Y21_to_ED),
    .from_EF(Tile_X5Y21_to_EF),
    .from_EG(Tile_X5Y21_to_EG),
    .from_EH(Tile_X5Y21_to_EH),
    .from_EI(Tile_X5Y21_to_EI),
    .from_SA(Tile_X6Y20_to_SA),
    .from_SB(Tile_X6Y20_to_SB),
    .from_SC(Tile_X6Y20_to_SC),
    .from_SD(Tile_X6Y20_to_SD),
    .from_SF(Tile_X6Y20_to_SF),
    .from_SG(Tile_X6Y20_to_SG),
    .from_SH(Tile_X6Y20_to_SH),
    .from_SI(Tile_X6Y20_to_SI),
    .from_WA(Tile_X7Y21_to_WA),
    .from_WB(Tile_X7Y21_to_WB),
    .from_WC(Tile_X7Y21_to_WC),
    .from_WD(Tile_X7Y21_to_WD),
    .from_WF(Tile_X7Y21_to_WF),
    .from_WG(Tile_X7Y21_to_WG),
    .from_WH(Tile_X7Y21_to_WH),
    .from_WI(Tile_X7Y21_to_WI),
    .to_EA(Tile_X6Y21_to_EA),
    .to_EB(Tile_X6Y21_to_EB),
    .to_EC(Tile_X6Y21_to_EC),
    .to_ED(Tile_X6Y21_to_ED),
    .to_EF(Tile_X6Y21_to_EF),
    .to_EG(Tile_X6Y21_to_EG),
    .to_EH(Tile_X6Y21_to_EH),
    .to_EI(Tile_X6Y21_to_EI),
    .to_WA(Tile_X6Y21_to_WA),
    .to_WB(Tile_X6Y21_to_WB),
    .to_WC(Tile_X6Y21_to_WC),
    .to_WD(Tile_X6Y21_to_WD),
    .to_WF(Tile_X6Y21_to_WF),
    .to_WG(Tile_X6Y21_to_WG),
    .to_WH(Tile_X6Y21_to_WH),
    .to_WI(Tile_X6Y21_to_WI),
    .to_NA(Tile_X6Y21_to_NA),
    .to_NB(Tile_X6Y21_to_NB),
    .to_NC(Tile_X6Y21_to_NC),
    .to_ND(Tile_X6Y21_to_ND),
    .to_NF(Tile_X6Y21_to_NF),
    .to_NG(Tile_X6Y21_to_NG),
    .to_NH(Tile_X6Y21_to_NH),
    .to_NI(Tile_X6Y21_to_NI),
    .to_SA(Tile_X6Y21_to_SA),
    .to_SB(Tile_X6Y21_to_SB),
    .to_SC(Tile_X6Y21_to_SC),
    .to_SD(Tile_X6Y21_to_SD),
    .to_SF(Tile_X6Y21_to_SF),
    .to_SG(Tile_X6Y21_to_SG),
    .to_SH(Tile_X6Y21_to_SH),
    .to_SI(Tile_X6Y21_to_SI),
    .R_t(Tile_X6Y21_R_t),
    .R_f(Tile_X6Y21_R_f),
    .F_masked1(Tile_X6Y21_F_masked1),
    .F_masked2(Tile_X6Y21_F_masked2),
    .UserCLK(Tile_X6Y22_UserCLKo),
    .UserCLKo(Tile_X6Y21_UserCLKo),
    .rst(Tile_X6Y22_rsto),
    .rsto(Tile_X6Y21_rsto),
    .FrameData(Tile_X5Y21_FrameData_O),
    .FrameData_O(Tile_X6Y21_FrameData_O),
    .FrameStrobe(Tile_X6Y22_FrameStrobe_O),
    .FrameStrobe_O(Tile_X6Y21_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X7Y21_Emulate_Bitstream)
    )
`endif
    Tile_X7Y21_linear_LMDPL
    (
    .from_NA(Tile_X7Y22_to_NA),
    .from_NB(Tile_X7Y22_to_NB),
    .from_NC(Tile_X7Y22_to_NC),
    .from_ND(Tile_X7Y22_to_ND),
    .from_NF(Tile_X7Y22_to_NF),
    .from_NG(Tile_X7Y22_to_NG),
    .from_NH(Tile_X7Y22_to_NH),
    .from_NI(Tile_X7Y22_to_NI),
    .from_EA(Tile_X6Y21_to_EA),
    .from_EB(Tile_X6Y21_to_EB),
    .from_EC(Tile_X6Y21_to_EC),
    .from_ED(Tile_X6Y21_to_ED),
    .from_EF(Tile_X6Y21_to_EF),
    .from_EG(Tile_X6Y21_to_EG),
    .from_EH(Tile_X6Y21_to_EH),
    .from_EI(Tile_X6Y21_to_EI),
    .from_SA(Tile_X7Y20_to_SA),
    .from_SB(Tile_X7Y20_to_SB),
    .from_SC(Tile_X7Y20_to_SC),
    .from_SD(Tile_X7Y20_to_SD),
    .from_SF(Tile_X7Y20_to_SF),
    .from_SG(Tile_X7Y20_to_SG),
    .from_SH(Tile_X7Y20_to_SH),
    .from_SI(Tile_X7Y20_to_SI),
    .from_WA(Tile_X8Y21_to_WA),
    .from_WB(Tile_X8Y21_to_WB),
    .from_WC(Tile_X8Y21_to_WC),
    .from_WD(Tile_X8Y21_to_WD),
    .from_WF(Tile_X8Y21_to_WF),
    .from_WG(Tile_X8Y21_to_WG),
    .from_WH(Tile_X8Y21_to_WH),
    .from_WI(Tile_X8Y21_to_WI),
    .to_EA(Tile_X7Y21_to_EA),
    .to_EB(Tile_X7Y21_to_EB),
    .to_EC(Tile_X7Y21_to_EC),
    .to_ED(Tile_X7Y21_to_ED),
    .to_EF(Tile_X7Y21_to_EF),
    .to_EG(Tile_X7Y21_to_EG),
    .to_EH(Tile_X7Y21_to_EH),
    .to_EI(Tile_X7Y21_to_EI),
    .to_WA(Tile_X7Y21_to_WA),
    .to_WB(Tile_X7Y21_to_WB),
    .to_WC(Tile_X7Y21_to_WC),
    .to_WD(Tile_X7Y21_to_WD),
    .to_WF(Tile_X7Y21_to_WF),
    .to_WG(Tile_X7Y21_to_WG),
    .to_WH(Tile_X7Y21_to_WH),
    .to_WI(Tile_X7Y21_to_WI),
    .to_NA(Tile_X7Y21_to_NA),
    .to_NB(Tile_X7Y21_to_NB),
    .to_NC(Tile_X7Y21_to_NC),
    .to_ND(Tile_X7Y21_to_ND),
    .to_NF(Tile_X7Y21_to_NF),
    .to_NG(Tile_X7Y21_to_NG),
    .to_NH(Tile_X7Y21_to_NH),
    .to_NI(Tile_X7Y21_to_NI),
    .to_SA(Tile_X7Y21_to_SA),
    .to_SB(Tile_X7Y21_to_SB),
    .to_SC(Tile_X7Y21_to_SC),
    .to_SD(Tile_X7Y21_to_SD),
    .to_SF(Tile_X7Y21_to_SF),
    .to_SG(Tile_X7Y21_to_SG),
    .to_SH(Tile_X7Y21_to_SH),
    .to_SI(Tile_X7Y21_to_SI),
    .F_masked1(Tile_X7Y21_F_masked1),
    .F_masked2(Tile_X7Y21_F_masked2),
    .UserCLK(Tile_X7Y22_UserCLKo),
    .UserCLKo(Tile_X7Y21_UserCLKo),
    .rst(Tile_X7Y22_rsto),
    .rsto(Tile_X7Y21_rsto),
    .FrameData(Tile_X6Y21_FrameData_O),
    .FrameData_O(Tile_X7Y21_FrameData_O),
    .FrameStrobe(Tile_X7Y22_FrameStrobe_O),
    .FrameStrobe_O(Tile_X7Y21_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
ctrl_to_sec
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X8Y21_Emulate_Bitstream)
    )
`endif
    Tile_X8Y21_ctrl_to_sec
    (
    .from_NA(Tile_X8Y22_to_NA),
    .from_NB(Tile_X8Y22_to_NB),
    .from_NC(Tile_X8Y22_to_NC),
    .from_ND(Tile_X8Y22_to_ND),
    .from_NF(Tile_X8Y22_to_NF),
    .from_NG(Tile_X8Y22_to_NG),
    .from_NH(Tile_X8Y22_to_NH),
    .from_NI(Tile_X8Y22_to_NI),
    .from_EA(Tile_X7Y21_to_EA),
    .from_EB(Tile_X7Y21_to_EB),
    .from_EC(Tile_X7Y21_to_EC),
    .from_ED(Tile_X7Y21_to_ED),
    .from_EF(Tile_X7Y21_to_EF),
    .from_EG(Tile_X7Y21_to_EG),
    .from_EH(Tile_X7Y21_to_EH),
    .from_EI(Tile_X7Y21_to_EI),
    .from_SA(Tile_X8Y20_to_SA),
    .from_SB(Tile_X8Y20_to_SB),
    .from_SC(Tile_X8Y20_to_SC),
    .from_SD(Tile_X8Y20_to_SD),
    .from_SF(Tile_X8Y20_to_SF),
    .from_SG(Tile_X8Y20_to_SG),
    .from_SH(Tile_X8Y20_to_SH),
    .from_SI(Tile_X8Y20_to_SI),
    .from_WA_1s(Tile_X9Y21_to_WA_1s),
    .from_WB_1s(Tile_X9Y21_to_WB_1s),
    .from_WC_1s(Tile_X9Y21_to_WC_1s),
    .from_WD_1s(Tile_X9Y21_to_WD_1s),
    .from_WF_1s(Tile_X9Y21_to_WF_1s),
    .from_WG_1s(Tile_X9Y21_to_WG_1s),
    .from_WH_1s(Tile_X9Y21_to_WH_1s),
    .from_WI_1s(Tile_X9Y21_to_WI_1s),
    .to_WA(Tile_X8Y21_to_WA),
    .to_WB(Tile_X8Y21_to_WB),
    .to_WC(Tile_X8Y21_to_WC),
    .to_WD(Tile_X8Y21_to_WD),
    .to_WF(Tile_X8Y21_to_WF),
    .to_WG(Tile_X8Y21_to_WG),
    .to_WH(Tile_X8Y21_to_WH),
    .to_WI(Tile_X8Y21_to_WI),
    .to_NA(Tile_X8Y21_to_NA),
    .to_NB(Tile_X8Y21_to_NB),
    .to_NC(Tile_X8Y21_to_NC),
    .to_ND(Tile_X8Y21_to_ND),
    .to_NF(Tile_X8Y21_to_NF),
    .to_NG(Tile_X8Y21_to_NG),
    .to_NH(Tile_X8Y21_to_NH),
    .to_NI(Tile_X8Y21_to_NI),
    .to_SA(Tile_X8Y21_to_SA),
    .to_SB(Tile_X8Y21_to_SB),
    .to_SC(Tile_X8Y21_to_SC),
    .to_SD(Tile_X8Y21_to_SD),
    .to_SF(Tile_X8Y21_to_SF),
    .to_SG(Tile_X8Y21_to_SG),
    .to_SH(Tile_X8Y21_to_SH),
    .to_SI(Tile_X8Y21_to_SI),
    .UserCLK(Tile_X8Y22_UserCLKo),
    .UserCLKo(Tile_X8Y21_UserCLKo),
    .rst(Tile_X8Y22_rsto),
    .rsto(Tile_X8Y21_rsto),
    .FrameData(Tile_X7Y21_FrameData_O),
    .FrameData_O(Tile_X8Y21_FrameData_O),
    .FrameStrobe(Tile_X8Y22_FrameStrobe_O),
    .FrameStrobe_O(Tile_X8Y21_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
combined_WDDL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X9Y21_Emulate_Bitstream)
    )
`endif
    Tile_X9Y21_combined_WDDL
    (
    .from_NA_1s(Tile_X9Y22_to_NA_1s),
    .from_NB_1s(Tile_X9Y22_to_NB_1s),
    .from_NC_1s(Tile_X9Y22_to_NC_1s),
    .from_ND_1s(Tile_X9Y22_to_ND_1s),
    .from_NF_1s(Tile_X9Y22_to_NF_1s),
    .from_NG_1s(Tile_X9Y22_to_NG_1s),
    .from_NH_1s(Tile_X9Y22_to_NH_1s),
    .from_NI_1s(Tile_X9Y22_to_NI_1s),
    .from_SA_1s(Tile_X9Y20_to_SA_1s),
    .from_SB_1s(Tile_X9Y20_to_SB_1s),
    .from_SC_1s(Tile_X9Y20_to_SC_1s),
    .from_SD_1s(Tile_X9Y20_to_SD_1s),
    .from_SF_1s(Tile_X9Y20_to_SF_1s),
    .from_SG_1s(Tile_X9Y20_to_SG_1s),
    .from_SH_1s(Tile_X9Y20_to_SH_1s),
    .from_SI_1s(Tile_X9Y20_to_SI_1s),
    .from_WA_1s(Tile_X10Y21_to_WA_1s),
    .from_WB_1s(Tile_X10Y21_to_WB_1s),
    .from_WC_1s(Tile_X10Y21_to_WC_1s),
    .from_WD_1s(Tile_X10Y21_to_WD_1s),
    .from_WF_1s(Tile_X10Y21_to_WF_1s),
    .from_WG_1s(Tile_X10Y21_to_WG_1s),
    .from_WH_1s(Tile_X10Y21_to_WH_1s),
    .from_WI_1s(Tile_X10Y21_to_WI_1s),
    .to_EA_1s(Tile_X9Y21_to_EA_1s),
    .to_EB_1s(Tile_X9Y21_to_EB_1s),
    .to_EC_1s(Tile_X9Y21_to_EC_1s),
    .to_ED_1s(Tile_X9Y21_to_ED_1s),
    .to_EF_1s(Tile_X9Y21_to_EF_1s),
    .to_EG_1s(Tile_X9Y21_to_EG_1s),
    .to_EH_1s(Tile_X9Y21_to_EH_1s),
    .to_EI_1s(Tile_X9Y21_to_EI_1s),
    .to_WA_1s(Tile_X9Y21_to_WA_1s),
    .to_WB_1s(Tile_X9Y21_to_WB_1s),
    .to_WC_1s(Tile_X9Y21_to_WC_1s),
    .to_WD_1s(Tile_X9Y21_to_WD_1s),
    .to_WF_1s(Tile_X9Y21_to_WF_1s),
    .to_WG_1s(Tile_X9Y21_to_WG_1s),
    .to_WH_1s(Tile_X9Y21_to_WH_1s),
    .to_WI_1s(Tile_X9Y21_to_WI_1s),
    .to_NA_1s(Tile_X9Y21_to_NA_1s),
    .to_NB_1s(Tile_X9Y21_to_NB_1s),
    .to_NC_1s(Tile_X9Y21_to_NC_1s),
    .to_ND_1s(Tile_X9Y21_to_ND_1s),
    .to_NF_1s(Tile_X9Y21_to_NF_1s),
    .to_NG_1s(Tile_X9Y21_to_NG_1s),
    .to_NH_1s(Tile_X9Y21_to_NH_1s),
    .to_NI_1s(Tile_X9Y21_to_NI_1s),
    .to_SA_1s(Tile_X9Y21_to_SA_1s),
    .to_SB_1s(Tile_X9Y21_to_SB_1s),
    .to_SC_1s(Tile_X9Y21_to_SC_1s),
    .to_SD_1s(Tile_X9Y21_to_SD_1s),
    .to_SF_1s(Tile_X9Y21_to_SF_1s),
    .to_SG_1s(Tile_X9Y21_to_SG_1s),
    .to_SH_1s(Tile_X9Y21_to_SH_1s),
    .to_SI_1s(Tile_X9Y21_to_SI_1s),
    .F_ctrl(Tile_X9Y21_F_ctrl),
    .UserCLK(Tile_X9Y22_UserCLKo),
    .UserCLKo(Tile_X9Y21_UserCLKo),
    .rst(Tile_X9Y22_rsto),
    .rsto(Tile_X9Y21_rsto),
    .FrameData(Tile_X8Y21_FrameData_O),
    .FrameData_O(Tile_X9Y21_FrameData_O),
    .FrameStrobe(Tile_X9Y22_FrameStrobe_O),
    .FrameStrobe_O(Tile_X9Y21_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
ctrl_IO
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X10Y21_Emulate_Bitstream)
    )
`endif
    Tile_X10Y21_ctrl_IO
    (
    .from_EA_1s(Tile_X9Y21_to_EA_1s),
    .from_EB_1s(Tile_X9Y21_to_EB_1s),
    .from_EC_1s(Tile_X9Y21_to_EC_1s),
    .from_ED_1s(Tile_X9Y21_to_ED_1s),
    .from_EF_1s(Tile_X9Y21_to_EF_1s),
    .from_EG_1s(Tile_X9Y21_to_EG_1s),
    .from_EH_1s(Tile_X9Y21_to_EH_1s),
    .from_EI_1s(Tile_X9Y21_to_EI_1s),
    .to_WA_1s(Tile_X10Y21_to_WA_1s),
    .to_WB_1s(Tile_X10Y21_to_WB_1s),
    .to_WC_1s(Tile_X10Y21_to_WC_1s),
    .to_WD_1s(Tile_X10Y21_to_WD_1s),
    .to_WF_1s(Tile_X10Y21_to_WF_1s),
    .to_WG_1s(Tile_X10Y21_to_WG_1s),
    .to_WH_1s(Tile_X10Y21_to_WH_1s),
    .to_WI_1s(Tile_X10Y21_to_WI_1s),
    .A_O_top_0_t(Tile_X10Y21_A_O_top_0_t),
    .A_O_top_0_f(Tile_X10Y21_A_O_top_0_f),
    .A_prech2(Tile_X10Y21_A_prech2),
    .A_DR_fault(Tile_X10Y21_A_DR_fault),
    .A_I_top_0_t(Tile_X10Y21_A_I_top_0_t),
    .A_I_top_0_f(Tile_X10Y21_A_I_top_0_f),
    .A_T_top(Tile_X10Y21_A_T_top),
    .A_F_ctrl(Tile_X10Y21_A_F_ctrl),
    .UserCLK(Tile_X10Y22_UserCLKo),
    .UserCLKo(Tile_X10Y21_UserCLKo),
    .rst(Tile_X10Y22_rsto),
    .rsto(Tile_X10Y21_rsto),
    .FrameData(Tile_X9Y21_FrameData_O),
    .FrameData_O(Tile_X10Y21_FrameData_O),
    .FrameStrobe(Tile_X10Y22_FrameStrobe_O),
    .FrameStrobe_O(Tile_X10Y21_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
W_IO_custom
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X0Y22_Emulate_Bitstream)
    )
`endif
    Tile_X0Y22_W_IO_custom
    (
    .from_NA(Tile_X0Y23_to_NA),
    .from_NB(Tile_X0Y23_to_NB),
    .from_NC(Tile_X0Y23_to_NC),
    .from_ND(Tile_X0Y23_to_ND),
    .from_NF(Tile_X0Y23_to_NF),
    .from_NG(Tile_X0Y23_to_NG),
    .from_NH(Tile_X0Y23_to_NH),
    .from_NI(Tile_X0Y23_to_NI),
    .from_SA(Tile_X0Y21_to_SA),
    .from_SB(Tile_X0Y21_to_SB),
    .from_SC(Tile_X0Y21_to_SC),
    .from_SD(Tile_X0Y21_to_SD),
    .from_SF(Tile_X0Y21_to_SF),
    .from_SG(Tile_X0Y21_to_SG),
    .from_SH(Tile_X0Y21_to_SH),
    .from_SI(Tile_X0Y21_to_SI),
    .from_WA(Tile_X1Y22_to_WA),
    .from_WB(Tile_X1Y22_to_WB),
    .from_WC(Tile_X1Y22_to_WC),
    .from_WD(Tile_X1Y22_to_WD),
    .from_WF(Tile_X1Y22_to_WF),
    .from_WG(Tile_X1Y22_to_WG),
    .from_WH(Tile_X1Y22_to_WH),
    .from_WI(Tile_X1Y22_to_WI),
    .to_EA(Tile_X0Y22_to_EA),
    .to_EB(Tile_X0Y22_to_EB),
    .to_EC(Tile_X0Y22_to_EC),
    .to_ED(Tile_X0Y22_to_ED),
    .to_EF(Tile_X0Y22_to_EF),
    .to_EG(Tile_X0Y22_to_EG),
    .to_EH(Tile_X0Y22_to_EH),
    .to_EI(Tile_X0Y22_to_EI),
    .to_NA(Tile_X0Y22_to_NA),
    .to_NB(Tile_X0Y22_to_NB),
    .to_NC(Tile_X0Y22_to_NC),
    .to_ND(Tile_X0Y22_to_ND),
    .to_NF(Tile_X0Y22_to_NF),
    .to_NG(Tile_X0Y22_to_NG),
    .to_NH(Tile_X0Y22_to_NH),
    .to_NI(Tile_X0Y22_to_NI),
    .to_SA(Tile_X0Y22_to_SA),
    .to_SB(Tile_X0Y22_to_SB),
    .to_SC(Tile_X0Y22_to_SC),
    .to_SD(Tile_X0Y22_to_SD),
    .to_SF(Tile_X0Y22_to_SF),
    .to_SG(Tile_X0Y22_to_SG),
    .to_SH(Tile_X0Y22_to_SH),
    .to_SI(Tile_X0Y22_to_SI),
    .A_O_top_0_t(Tile_X0Y22_A_O_top_0_t),
    .A_O_top_0_f(Tile_X0Y22_A_O_top_0_f),
    .A_O_top_1_t(Tile_X0Y22_A_O_top_1_t),
    .A_O_top_1_f(Tile_X0Y22_A_O_top_1_f),
    .A_prech1(Tile_X0Y22_A_prech1),
    .A_prech2(Tile_X0Y22_A_prech2),
    .A_DR_fault(Tile_X0Y22_A_DR_fault),
    .A_I_top_0_t(Tile_X0Y22_A_I_top_0_t),
    .A_I_top_0_f(Tile_X0Y22_A_I_top_0_f),
    .A_I_top_1_t(Tile_X0Y22_A_I_top_1_t),
    .A_I_top_1_f(Tile_X0Y22_A_I_top_1_f),
    .A_T_top(Tile_X0Y22_A_T_top),
    .A_F_masked1(Tile_X0Y22_A_F_masked1),
    .A_F_masked2(Tile_X0Y22_A_F_masked2),
    .A_config_C_bit0(Tile_X0Y22_A_config_C_bit0),
    .A_config_C_bit1(Tile_X0Y22_A_config_C_bit1),
    .A_config_C_bit2(Tile_X0Y22_A_config_C_bit2),
    .A_config_C_bit3(Tile_X0Y22_A_config_C_bit3),
    .B_config_C_bit0(Tile_X0Y22_B_config_C_bit0),
    .B_config_C_bit1(Tile_X0Y22_B_config_C_bit1),
    .B_config_C_bit2(Tile_X0Y22_B_config_C_bit2),
    .B_config_C_bit3(Tile_X0Y22_B_config_C_bit3),
    .UserCLK(Tile_X0Y23_UserCLKo),
    .UserCLKo(Tile_X0Y22_UserCLKo),
    .rst(Tile_X0Y23_rsto),
    .rsto(Tile_X0Y22_rsto),
    .FrameData(Tile_Y22_FrameData),
    .FrameData_O(Tile_X0Y22_FrameData_O),
    .FrameStrobe(Tile_X0Y23_FrameStrobe_O),
    .FrameStrobe_O(Tile_X0Y22_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X1Y22_Emulate_Bitstream)
    )
`endif
    Tile_X1Y22_linear_LMDPL
    (
    .from_NA(Tile_X1Y23_to_NA),
    .from_NB(Tile_X1Y23_to_NB),
    .from_NC(Tile_X1Y23_to_NC),
    .from_ND(Tile_X1Y23_to_ND),
    .from_NF(Tile_X1Y23_to_NF),
    .from_NG(Tile_X1Y23_to_NG),
    .from_NH(Tile_X1Y23_to_NH),
    .from_NI(Tile_X1Y23_to_NI),
    .from_EA(Tile_X0Y22_to_EA),
    .from_EB(Tile_X0Y22_to_EB),
    .from_EC(Tile_X0Y22_to_EC),
    .from_ED(Tile_X0Y22_to_ED),
    .from_EF(Tile_X0Y22_to_EF),
    .from_EG(Tile_X0Y22_to_EG),
    .from_EH(Tile_X0Y22_to_EH),
    .from_EI(Tile_X0Y22_to_EI),
    .from_SA(Tile_X1Y21_to_SA),
    .from_SB(Tile_X1Y21_to_SB),
    .from_SC(Tile_X1Y21_to_SC),
    .from_SD(Tile_X1Y21_to_SD),
    .from_SF(Tile_X1Y21_to_SF),
    .from_SG(Tile_X1Y21_to_SG),
    .from_SH(Tile_X1Y21_to_SH),
    .from_SI(Tile_X1Y21_to_SI),
    .from_WA(Tile_X2Y22_to_WA),
    .from_WB(Tile_X2Y22_to_WB),
    .from_WC(Tile_X2Y22_to_WC),
    .from_WD(Tile_X2Y22_to_WD),
    .from_WF(Tile_X2Y22_to_WF),
    .from_WG(Tile_X2Y22_to_WG),
    .from_WH(Tile_X2Y22_to_WH),
    .from_WI(Tile_X2Y22_to_WI),
    .to_EA(Tile_X1Y22_to_EA),
    .to_EB(Tile_X1Y22_to_EB),
    .to_EC(Tile_X1Y22_to_EC),
    .to_ED(Tile_X1Y22_to_ED),
    .to_EF(Tile_X1Y22_to_EF),
    .to_EG(Tile_X1Y22_to_EG),
    .to_EH(Tile_X1Y22_to_EH),
    .to_EI(Tile_X1Y22_to_EI),
    .to_WA(Tile_X1Y22_to_WA),
    .to_WB(Tile_X1Y22_to_WB),
    .to_WC(Tile_X1Y22_to_WC),
    .to_WD(Tile_X1Y22_to_WD),
    .to_WF(Tile_X1Y22_to_WF),
    .to_WG(Tile_X1Y22_to_WG),
    .to_WH(Tile_X1Y22_to_WH),
    .to_WI(Tile_X1Y22_to_WI),
    .to_NA(Tile_X1Y22_to_NA),
    .to_NB(Tile_X1Y22_to_NB),
    .to_NC(Tile_X1Y22_to_NC),
    .to_ND(Tile_X1Y22_to_ND),
    .to_NF(Tile_X1Y22_to_NF),
    .to_NG(Tile_X1Y22_to_NG),
    .to_NH(Tile_X1Y22_to_NH),
    .to_NI(Tile_X1Y22_to_NI),
    .to_SA(Tile_X1Y22_to_SA),
    .to_SB(Tile_X1Y22_to_SB),
    .to_SC(Tile_X1Y22_to_SC),
    .to_SD(Tile_X1Y22_to_SD),
    .to_SF(Tile_X1Y22_to_SF),
    .to_SG(Tile_X1Y22_to_SG),
    .to_SH(Tile_X1Y22_to_SH),
    .to_SI(Tile_X1Y22_to_SI),
    .F_masked1(Tile_X1Y22_F_masked1),
    .F_masked2(Tile_X1Y22_F_masked2),
    .UserCLK(Tile_X1Y23_UserCLKo),
    .UserCLKo(Tile_X1Y22_UserCLKo),
    .rst(Tile_X1Y23_rsto),
    .rsto(Tile_X1Y22_rsto),
    .FrameData(Tile_X0Y22_FrameData_O),
    .FrameData_O(Tile_X1Y22_FrameData_O),
    .FrameStrobe(Tile_X1Y23_FrameStrobe_O),
    .FrameStrobe_O(Tile_X1Y22_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X2Y22_Emulate_Bitstream)
    )
`endif
    Tile_X2Y22_linear_LMDPL
    (
    .from_NA(Tile_X2Y23_to_NA),
    .from_NB(Tile_X2Y23_to_NB),
    .from_NC(Tile_X2Y23_to_NC),
    .from_ND(Tile_X2Y23_to_ND),
    .from_NF(Tile_X2Y23_to_NF),
    .from_NG(Tile_X2Y23_to_NG),
    .from_NH(Tile_X2Y23_to_NH),
    .from_NI(Tile_X2Y23_to_NI),
    .from_EA(Tile_X1Y22_to_EA),
    .from_EB(Tile_X1Y22_to_EB),
    .from_EC(Tile_X1Y22_to_EC),
    .from_ED(Tile_X1Y22_to_ED),
    .from_EF(Tile_X1Y22_to_EF),
    .from_EG(Tile_X1Y22_to_EG),
    .from_EH(Tile_X1Y22_to_EH),
    .from_EI(Tile_X1Y22_to_EI),
    .from_SA(Tile_X2Y21_to_SA),
    .from_SB(Tile_X2Y21_to_SB),
    .from_SC(Tile_X2Y21_to_SC),
    .from_SD(Tile_X2Y21_to_SD),
    .from_SF(Tile_X2Y21_to_SF),
    .from_SG(Tile_X2Y21_to_SG),
    .from_SH(Tile_X2Y21_to_SH),
    .from_SI(Tile_X2Y21_to_SI),
    .from_WA(Tile_X3Y22_to_WA),
    .from_WB(Tile_X3Y22_to_WB),
    .from_WC(Tile_X3Y22_to_WC),
    .from_WD(Tile_X3Y22_to_WD),
    .from_WF(Tile_X3Y22_to_WF),
    .from_WG(Tile_X3Y22_to_WG),
    .from_WH(Tile_X3Y22_to_WH),
    .from_WI(Tile_X3Y22_to_WI),
    .to_EA(Tile_X2Y22_to_EA),
    .to_EB(Tile_X2Y22_to_EB),
    .to_EC(Tile_X2Y22_to_EC),
    .to_ED(Tile_X2Y22_to_ED),
    .to_EF(Tile_X2Y22_to_EF),
    .to_EG(Tile_X2Y22_to_EG),
    .to_EH(Tile_X2Y22_to_EH),
    .to_EI(Tile_X2Y22_to_EI),
    .to_WA(Tile_X2Y22_to_WA),
    .to_WB(Tile_X2Y22_to_WB),
    .to_WC(Tile_X2Y22_to_WC),
    .to_WD(Tile_X2Y22_to_WD),
    .to_WF(Tile_X2Y22_to_WF),
    .to_WG(Tile_X2Y22_to_WG),
    .to_WH(Tile_X2Y22_to_WH),
    .to_WI(Tile_X2Y22_to_WI),
    .to_NA(Tile_X2Y22_to_NA),
    .to_NB(Tile_X2Y22_to_NB),
    .to_NC(Tile_X2Y22_to_NC),
    .to_ND(Tile_X2Y22_to_ND),
    .to_NF(Tile_X2Y22_to_NF),
    .to_NG(Tile_X2Y22_to_NG),
    .to_NH(Tile_X2Y22_to_NH),
    .to_NI(Tile_X2Y22_to_NI),
    .to_SA(Tile_X2Y22_to_SA),
    .to_SB(Tile_X2Y22_to_SB),
    .to_SC(Tile_X2Y22_to_SC),
    .to_SD(Tile_X2Y22_to_SD),
    .to_SF(Tile_X2Y22_to_SF),
    .to_SG(Tile_X2Y22_to_SG),
    .to_SH(Tile_X2Y22_to_SH),
    .to_SI(Tile_X2Y22_to_SI),
    .F_masked1(Tile_X2Y22_F_masked1),
    .F_masked2(Tile_X2Y22_F_masked2),
    .UserCLK(Tile_X2Y23_UserCLKo),
    .UserCLKo(Tile_X2Y22_UserCLKo),
    .rst(Tile_X2Y23_rsto),
    .rsto(Tile_X2Y22_rsto),
    .FrameData(Tile_X1Y22_FrameData_O),
    .FrameData_O(Tile_X2Y22_FrameData_O),
    .FrameStrobe(Tile_X2Y23_FrameStrobe_O),
    .FrameStrobe_O(Tile_X2Y22_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
nonlinear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X3Y22_Emulate_Bitstream)
    )
`endif
    Tile_X3Y22_nonlinear_LMDPL
    (
    .from_NA(Tile_X3Y23_to_NA),
    .from_NB(Tile_X3Y23_to_NB),
    .from_NC(Tile_X3Y23_to_NC),
    .from_ND(Tile_X3Y23_to_ND),
    .from_NF(Tile_X3Y23_to_NF),
    .from_NG(Tile_X3Y23_to_NG),
    .from_NH(Tile_X3Y23_to_NH),
    .from_NI(Tile_X3Y23_to_NI),
    .from_EA(Tile_X2Y22_to_EA),
    .from_EB(Tile_X2Y22_to_EB),
    .from_EC(Tile_X2Y22_to_EC),
    .from_ED(Tile_X2Y22_to_ED),
    .from_EF(Tile_X2Y22_to_EF),
    .from_EG(Tile_X2Y22_to_EG),
    .from_EH(Tile_X2Y22_to_EH),
    .from_EI(Tile_X2Y22_to_EI),
    .from_SA(Tile_X3Y21_to_SA),
    .from_SB(Tile_X3Y21_to_SB),
    .from_SC(Tile_X3Y21_to_SC),
    .from_SD(Tile_X3Y21_to_SD),
    .from_SF(Tile_X3Y21_to_SF),
    .from_SG(Tile_X3Y21_to_SG),
    .from_SH(Tile_X3Y21_to_SH),
    .from_SI(Tile_X3Y21_to_SI),
    .from_WA(Tile_X4Y22_to_WA),
    .from_WB(Tile_X4Y22_to_WB),
    .from_WC(Tile_X4Y22_to_WC),
    .from_WD(Tile_X4Y22_to_WD),
    .from_WF(Tile_X4Y22_to_WF),
    .from_WG(Tile_X4Y22_to_WG),
    .from_WH(Tile_X4Y22_to_WH),
    .from_WI(Tile_X4Y22_to_WI),
    .to_EA(Tile_X3Y22_to_EA),
    .to_EB(Tile_X3Y22_to_EB),
    .to_EC(Tile_X3Y22_to_EC),
    .to_ED(Tile_X3Y22_to_ED),
    .to_EF(Tile_X3Y22_to_EF),
    .to_EG(Tile_X3Y22_to_EG),
    .to_EH(Tile_X3Y22_to_EH),
    .to_EI(Tile_X3Y22_to_EI),
    .to_WA(Tile_X3Y22_to_WA),
    .to_WB(Tile_X3Y22_to_WB),
    .to_WC(Tile_X3Y22_to_WC),
    .to_WD(Tile_X3Y22_to_WD),
    .to_WF(Tile_X3Y22_to_WF),
    .to_WG(Tile_X3Y22_to_WG),
    .to_WH(Tile_X3Y22_to_WH),
    .to_WI(Tile_X3Y22_to_WI),
    .to_NA(Tile_X3Y22_to_NA),
    .to_NB(Tile_X3Y22_to_NB),
    .to_NC(Tile_X3Y22_to_NC),
    .to_ND(Tile_X3Y22_to_ND),
    .to_NF(Tile_X3Y22_to_NF),
    .to_NG(Tile_X3Y22_to_NG),
    .to_NH(Tile_X3Y22_to_NH),
    .to_NI(Tile_X3Y22_to_NI),
    .to_SA(Tile_X3Y22_to_SA),
    .to_SB(Tile_X3Y22_to_SB),
    .to_SC(Tile_X3Y22_to_SC),
    .to_SD(Tile_X3Y22_to_SD),
    .to_SF(Tile_X3Y22_to_SF),
    .to_SG(Tile_X3Y22_to_SG),
    .to_SH(Tile_X3Y22_to_SH),
    .to_SI(Tile_X3Y22_to_SI),
    .R_t(Tile_X3Y22_R_t),
    .R_f(Tile_X3Y22_R_f),
    .F_masked1(Tile_X3Y22_F_masked1),
    .F_masked2(Tile_X3Y22_F_masked2),
    .UserCLK(Tile_X3Y23_UserCLKo),
    .UserCLKo(Tile_X3Y22_UserCLKo),
    .rst(Tile_X3Y23_rsto),
    .rsto(Tile_X3Y22_rsto),
    .FrameData(Tile_X2Y22_FrameData_O),
    .FrameData_O(Tile_X3Y22_FrameData_O),
    .FrameStrobe(Tile_X3Y23_FrameStrobe_O),
    .FrameStrobe_O(Tile_X3Y22_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X4Y22_Emulate_Bitstream)
    )
`endif
    Tile_X4Y22_linear_LMDPL
    (
    .from_NA(Tile_X4Y23_to_NA),
    .from_NB(Tile_X4Y23_to_NB),
    .from_NC(Tile_X4Y23_to_NC),
    .from_ND(Tile_X4Y23_to_ND),
    .from_NF(Tile_X4Y23_to_NF),
    .from_NG(Tile_X4Y23_to_NG),
    .from_NH(Tile_X4Y23_to_NH),
    .from_NI(Tile_X4Y23_to_NI),
    .from_EA(Tile_X3Y22_to_EA),
    .from_EB(Tile_X3Y22_to_EB),
    .from_EC(Tile_X3Y22_to_EC),
    .from_ED(Tile_X3Y22_to_ED),
    .from_EF(Tile_X3Y22_to_EF),
    .from_EG(Tile_X3Y22_to_EG),
    .from_EH(Tile_X3Y22_to_EH),
    .from_EI(Tile_X3Y22_to_EI),
    .from_SA(Tile_X4Y21_to_SA),
    .from_SB(Tile_X4Y21_to_SB),
    .from_SC(Tile_X4Y21_to_SC),
    .from_SD(Tile_X4Y21_to_SD),
    .from_SF(Tile_X4Y21_to_SF),
    .from_SG(Tile_X4Y21_to_SG),
    .from_SH(Tile_X4Y21_to_SH),
    .from_SI(Tile_X4Y21_to_SI),
    .from_WA(Tile_X5Y22_to_WA),
    .from_WB(Tile_X5Y22_to_WB),
    .from_WC(Tile_X5Y22_to_WC),
    .from_WD(Tile_X5Y22_to_WD),
    .from_WF(Tile_X5Y22_to_WF),
    .from_WG(Tile_X5Y22_to_WG),
    .from_WH(Tile_X5Y22_to_WH),
    .from_WI(Tile_X5Y22_to_WI),
    .to_EA(Tile_X4Y22_to_EA),
    .to_EB(Tile_X4Y22_to_EB),
    .to_EC(Tile_X4Y22_to_EC),
    .to_ED(Tile_X4Y22_to_ED),
    .to_EF(Tile_X4Y22_to_EF),
    .to_EG(Tile_X4Y22_to_EG),
    .to_EH(Tile_X4Y22_to_EH),
    .to_EI(Tile_X4Y22_to_EI),
    .to_WA(Tile_X4Y22_to_WA),
    .to_WB(Tile_X4Y22_to_WB),
    .to_WC(Tile_X4Y22_to_WC),
    .to_WD(Tile_X4Y22_to_WD),
    .to_WF(Tile_X4Y22_to_WF),
    .to_WG(Tile_X4Y22_to_WG),
    .to_WH(Tile_X4Y22_to_WH),
    .to_WI(Tile_X4Y22_to_WI),
    .to_NA(Tile_X4Y22_to_NA),
    .to_NB(Tile_X4Y22_to_NB),
    .to_NC(Tile_X4Y22_to_NC),
    .to_ND(Tile_X4Y22_to_ND),
    .to_NF(Tile_X4Y22_to_NF),
    .to_NG(Tile_X4Y22_to_NG),
    .to_NH(Tile_X4Y22_to_NH),
    .to_NI(Tile_X4Y22_to_NI),
    .to_SA(Tile_X4Y22_to_SA),
    .to_SB(Tile_X4Y22_to_SB),
    .to_SC(Tile_X4Y22_to_SC),
    .to_SD(Tile_X4Y22_to_SD),
    .to_SF(Tile_X4Y22_to_SF),
    .to_SG(Tile_X4Y22_to_SG),
    .to_SH(Tile_X4Y22_to_SH),
    .to_SI(Tile_X4Y22_to_SI),
    .F_masked1(Tile_X4Y22_F_masked1),
    .F_masked2(Tile_X4Y22_F_masked2),
    .UserCLK(Tile_X4Y23_UserCLKo),
    .UserCLKo(Tile_X4Y22_UserCLKo),
    .rst(Tile_X4Y23_rsto),
    .rsto(Tile_X4Y22_rsto),
    .FrameData(Tile_X3Y22_FrameData_O),
    .FrameData_O(Tile_X4Y22_FrameData_O),
    .FrameStrobe(Tile_X4Y23_FrameStrobe_O),
    .FrameStrobe_O(Tile_X4Y22_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X5Y22_Emulate_Bitstream)
    )
`endif
    Tile_X5Y22_linear_LMDPL
    (
    .from_NA(Tile_X5Y23_to_NA),
    .from_NB(Tile_X5Y23_to_NB),
    .from_NC(Tile_X5Y23_to_NC),
    .from_ND(Tile_X5Y23_to_ND),
    .from_NF(Tile_X5Y23_to_NF),
    .from_NG(Tile_X5Y23_to_NG),
    .from_NH(Tile_X5Y23_to_NH),
    .from_NI(Tile_X5Y23_to_NI),
    .from_EA(Tile_X4Y22_to_EA),
    .from_EB(Tile_X4Y22_to_EB),
    .from_EC(Tile_X4Y22_to_EC),
    .from_ED(Tile_X4Y22_to_ED),
    .from_EF(Tile_X4Y22_to_EF),
    .from_EG(Tile_X4Y22_to_EG),
    .from_EH(Tile_X4Y22_to_EH),
    .from_EI(Tile_X4Y22_to_EI),
    .from_SA(Tile_X5Y21_to_SA),
    .from_SB(Tile_X5Y21_to_SB),
    .from_SC(Tile_X5Y21_to_SC),
    .from_SD(Tile_X5Y21_to_SD),
    .from_SF(Tile_X5Y21_to_SF),
    .from_SG(Tile_X5Y21_to_SG),
    .from_SH(Tile_X5Y21_to_SH),
    .from_SI(Tile_X5Y21_to_SI),
    .from_WA(Tile_X6Y22_to_WA),
    .from_WB(Tile_X6Y22_to_WB),
    .from_WC(Tile_X6Y22_to_WC),
    .from_WD(Tile_X6Y22_to_WD),
    .from_WF(Tile_X6Y22_to_WF),
    .from_WG(Tile_X6Y22_to_WG),
    .from_WH(Tile_X6Y22_to_WH),
    .from_WI(Tile_X6Y22_to_WI),
    .to_EA(Tile_X5Y22_to_EA),
    .to_EB(Tile_X5Y22_to_EB),
    .to_EC(Tile_X5Y22_to_EC),
    .to_ED(Tile_X5Y22_to_ED),
    .to_EF(Tile_X5Y22_to_EF),
    .to_EG(Tile_X5Y22_to_EG),
    .to_EH(Tile_X5Y22_to_EH),
    .to_EI(Tile_X5Y22_to_EI),
    .to_WA(Tile_X5Y22_to_WA),
    .to_WB(Tile_X5Y22_to_WB),
    .to_WC(Tile_X5Y22_to_WC),
    .to_WD(Tile_X5Y22_to_WD),
    .to_WF(Tile_X5Y22_to_WF),
    .to_WG(Tile_X5Y22_to_WG),
    .to_WH(Tile_X5Y22_to_WH),
    .to_WI(Tile_X5Y22_to_WI),
    .to_NA(Tile_X5Y22_to_NA),
    .to_NB(Tile_X5Y22_to_NB),
    .to_NC(Tile_X5Y22_to_NC),
    .to_ND(Tile_X5Y22_to_ND),
    .to_NF(Tile_X5Y22_to_NF),
    .to_NG(Tile_X5Y22_to_NG),
    .to_NH(Tile_X5Y22_to_NH),
    .to_NI(Tile_X5Y22_to_NI),
    .to_SA(Tile_X5Y22_to_SA),
    .to_SB(Tile_X5Y22_to_SB),
    .to_SC(Tile_X5Y22_to_SC),
    .to_SD(Tile_X5Y22_to_SD),
    .to_SF(Tile_X5Y22_to_SF),
    .to_SG(Tile_X5Y22_to_SG),
    .to_SH(Tile_X5Y22_to_SH),
    .to_SI(Tile_X5Y22_to_SI),
    .F_masked1(Tile_X5Y22_F_masked1),
    .F_masked2(Tile_X5Y22_F_masked2),
    .UserCLK(Tile_X5Y23_UserCLKo),
    .UserCLKo(Tile_X5Y22_UserCLKo),
    .rst(Tile_X5Y23_rsto),
    .rsto(Tile_X5Y22_rsto),
    .FrameData(Tile_X4Y22_FrameData_O),
    .FrameData_O(Tile_X5Y22_FrameData_O),
    .FrameStrobe(Tile_X5Y23_FrameStrobe_O),
    .FrameStrobe_O(Tile_X5Y22_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
nonlinear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X6Y22_Emulate_Bitstream)
    )
`endif
    Tile_X6Y22_nonlinear_LMDPL
    (
    .from_NA(Tile_X6Y23_to_NA),
    .from_NB(Tile_X6Y23_to_NB),
    .from_NC(Tile_X6Y23_to_NC),
    .from_ND(Tile_X6Y23_to_ND),
    .from_NF(Tile_X6Y23_to_NF),
    .from_NG(Tile_X6Y23_to_NG),
    .from_NH(Tile_X6Y23_to_NH),
    .from_NI(Tile_X6Y23_to_NI),
    .from_EA(Tile_X5Y22_to_EA),
    .from_EB(Tile_X5Y22_to_EB),
    .from_EC(Tile_X5Y22_to_EC),
    .from_ED(Tile_X5Y22_to_ED),
    .from_EF(Tile_X5Y22_to_EF),
    .from_EG(Tile_X5Y22_to_EG),
    .from_EH(Tile_X5Y22_to_EH),
    .from_EI(Tile_X5Y22_to_EI),
    .from_SA(Tile_X6Y21_to_SA),
    .from_SB(Tile_X6Y21_to_SB),
    .from_SC(Tile_X6Y21_to_SC),
    .from_SD(Tile_X6Y21_to_SD),
    .from_SF(Tile_X6Y21_to_SF),
    .from_SG(Tile_X6Y21_to_SG),
    .from_SH(Tile_X6Y21_to_SH),
    .from_SI(Tile_X6Y21_to_SI),
    .from_WA(Tile_X7Y22_to_WA),
    .from_WB(Tile_X7Y22_to_WB),
    .from_WC(Tile_X7Y22_to_WC),
    .from_WD(Tile_X7Y22_to_WD),
    .from_WF(Tile_X7Y22_to_WF),
    .from_WG(Tile_X7Y22_to_WG),
    .from_WH(Tile_X7Y22_to_WH),
    .from_WI(Tile_X7Y22_to_WI),
    .to_EA(Tile_X6Y22_to_EA),
    .to_EB(Tile_X6Y22_to_EB),
    .to_EC(Tile_X6Y22_to_EC),
    .to_ED(Tile_X6Y22_to_ED),
    .to_EF(Tile_X6Y22_to_EF),
    .to_EG(Tile_X6Y22_to_EG),
    .to_EH(Tile_X6Y22_to_EH),
    .to_EI(Tile_X6Y22_to_EI),
    .to_WA(Tile_X6Y22_to_WA),
    .to_WB(Tile_X6Y22_to_WB),
    .to_WC(Tile_X6Y22_to_WC),
    .to_WD(Tile_X6Y22_to_WD),
    .to_WF(Tile_X6Y22_to_WF),
    .to_WG(Tile_X6Y22_to_WG),
    .to_WH(Tile_X6Y22_to_WH),
    .to_WI(Tile_X6Y22_to_WI),
    .to_NA(Tile_X6Y22_to_NA),
    .to_NB(Tile_X6Y22_to_NB),
    .to_NC(Tile_X6Y22_to_NC),
    .to_ND(Tile_X6Y22_to_ND),
    .to_NF(Tile_X6Y22_to_NF),
    .to_NG(Tile_X6Y22_to_NG),
    .to_NH(Tile_X6Y22_to_NH),
    .to_NI(Tile_X6Y22_to_NI),
    .to_SA(Tile_X6Y22_to_SA),
    .to_SB(Tile_X6Y22_to_SB),
    .to_SC(Tile_X6Y22_to_SC),
    .to_SD(Tile_X6Y22_to_SD),
    .to_SF(Tile_X6Y22_to_SF),
    .to_SG(Tile_X6Y22_to_SG),
    .to_SH(Tile_X6Y22_to_SH),
    .to_SI(Tile_X6Y22_to_SI),
    .R_t(Tile_X6Y22_R_t),
    .R_f(Tile_X6Y22_R_f),
    .F_masked1(Tile_X6Y22_F_masked1),
    .F_masked2(Tile_X6Y22_F_masked2),
    .UserCLK(Tile_X6Y23_UserCLKo),
    .UserCLKo(Tile_X6Y22_UserCLKo),
    .rst(Tile_X6Y23_rsto),
    .rsto(Tile_X6Y22_rsto),
    .FrameData(Tile_X5Y22_FrameData_O),
    .FrameData_O(Tile_X6Y22_FrameData_O),
    .FrameStrobe(Tile_X6Y23_FrameStrobe_O),
    .FrameStrobe_O(Tile_X6Y22_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X7Y22_Emulate_Bitstream)
    )
`endif
    Tile_X7Y22_linear_LMDPL
    (
    .from_NA(Tile_X7Y23_to_NA),
    .from_NB(Tile_X7Y23_to_NB),
    .from_NC(Tile_X7Y23_to_NC),
    .from_ND(Tile_X7Y23_to_ND),
    .from_NF(Tile_X7Y23_to_NF),
    .from_NG(Tile_X7Y23_to_NG),
    .from_NH(Tile_X7Y23_to_NH),
    .from_NI(Tile_X7Y23_to_NI),
    .from_EA(Tile_X6Y22_to_EA),
    .from_EB(Tile_X6Y22_to_EB),
    .from_EC(Tile_X6Y22_to_EC),
    .from_ED(Tile_X6Y22_to_ED),
    .from_EF(Tile_X6Y22_to_EF),
    .from_EG(Tile_X6Y22_to_EG),
    .from_EH(Tile_X6Y22_to_EH),
    .from_EI(Tile_X6Y22_to_EI),
    .from_SA(Tile_X7Y21_to_SA),
    .from_SB(Tile_X7Y21_to_SB),
    .from_SC(Tile_X7Y21_to_SC),
    .from_SD(Tile_X7Y21_to_SD),
    .from_SF(Tile_X7Y21_to_SF),
    .from_SG(Tile_X7Y21_to_SG),
    .from_SH(Tile_X7Y21_to_SH),
    .from_SI(Tile_X7Y21_to_SI),
    .from_WA(Tile_X8Y22_to_WA),
    .from_WB(Tile_X8Y22_to_WB),
    .from_WC(Tile_X8Y22_to_WC),
    .from_WD(Tile_X8Y22_to_WD),
    .from_WF(Tile_X8Y22_to_WF),
    .from_WG(Tile_X8Y22_to_WG),
    .from_WH(Tile_X8Y22_to_WH),
    .from_WI(Tile_X8Y22_to_WI),
    .to_EA(Tile_X7Y22_to_EA),
    .to_EB(Tile_X7Y22_to_EB),
    .to_EC(Tile_X7Y22_to_EC),
    .to_ED(Tile_X7Y22_to_ED),
    .to_EF(Tile_X7Y22_to_EF),
    .to_EG(Tile_X7Y22_to_EG),
    .to_EH(Tile_X7Y22_to_EH),
    .to_EI(Tile_X7Y22_to_EI),
    .to_WA(Tile_X7Y22_to_WA),
    .to_WB(Tile_X7Y22_to_WB),
    .to_WC(Tile_X7Y22_to_WC),
    .to_WD(Tile_X7Y22_to_WD),
    .to_WF(Tile_X7Y22_to_WF),
    .to_WG(Tile_X7Y22_to_WG),
    .to_WH(Tile_X7Y22_to_WH),
    .to_WI(Tile_X7Y22_to_WI),
    .to_NA(Tile_X7Y22_to_NA),
    .to_NB(Tile_X7Y22_to_NB),
    .to_NC(Tile_X7Y22_to_NC),
    .to_ND(Tile_X7Y22_to_ND),
    .to_NF(Tile_X7Y22_to_NF),
    .to_NG(Tile_X7Y22_to_NG),
    .to_NH(Tile_X7Y22_to_NH),
    .to_NI(Tile_X7Y22_to_NI),
    .to_SA(Tile_X7Y22_to_SA),
    .to_SB(Tile_X7Y22_to_SB),
    .to_SC(Tile_X7Y22_to_SC),
    .to_SD(Tile_X7Y22_to_SD),
    .to_SF(Tile_X7Y22_to_SF),
    .to_SG(Tile_X7Y22_to_SG),
    .to_SH(Tile_X7Y22_to_SH),
    .to_SI(Tile_X7Y22_to_SI),
    .F_masked1(Tile_X7Y22_F_masked1),
    .F_masked2(Tile_X7Y22_F_masked2),
    .UserCLK(Tile_X7Y23_UserCLKo),
    .UserCLKo(Tile_X7Y22_UserCLKo),
    .rst(Tile_X7Y23_rsto),
    .rsto(Tile_X7Y22_rsto),
    .FrameData(Tile_X6Y22_FrameData_O),
    .FrameData_O(Tile_X7Y22_FrameData_O),
    .FrameStrobe(Tile_X7Y23_FrameStrobe_O),
    .FrameStrobe_O(Tile_X7Y22_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
ctrl_to_sec
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X8Y22_Emulate_Bitstream)
    )
`endif
    Tile_X8Y22_ctrl_to_sec
    (
    .from_NA(Tile_X8Y23_to_NA),
    .from_NB(Tile_X8Y23_to_NB),
    .from_NC(Tile_X8Y23_to_NC),
    .from_ND(Tile_X8Y23_to_ND),
    .from_NF(Tile_X8Y23_to_NF),
    .from_NG(Tile_X8Y23_to_NG),
    .from_NH(Tile_X8Y23_to_NH),
    .from_NI(Tile_X8Y23_to_NI),
    .from_EA(Tile_X7Y22_to_EA),
    .from_EB(Tile_X7Y22_to_EB),
    .from_EC(Tile_X7Y22_to_EC),
    .from_ED(Tile_X7Y22_to_ED),
    .from_EF(Tile_X7Y22_to_EF),
    .from_EG(Tile_X7Y22_to_EG),
    .from_EH(Tile_X7Y22_to_EH),
    .from_EI(Tile_X7Y22_to_EI),
    .from_SA(Tile_X8Y21_to_SA),
    .from_SB(Tile_X8Y21_to_SB),
    .from_SC(Tile_X8Y21_to_SC),
    .from_SD(Tile_X8Y21_to_SD),
    .from_SF(Tile_X8Y21_to_SF),
    .from_SG(Tile_X8Y21_to_SG),
    .from_SH(Tile_X8Y21_to_SH),
    .from_SI(Tile_X8Y21_to_SI),
    .from_WA_1s(Tile_X9Y22_to_WA_1s),
    .from_WB_1s(Tile_X9Y22_to_WB_1s),
    .from_WC_1s(Tile_X9Y22_to_WC_1s),
    .from_WD_1s(Tile_X9Y22_to_WD_1s),
    .from_WF_1s(Tile_X9Y22_to_WF_1s),
    .from_WG_1s(Tile_X9Y22_to_WG_1s),
    .from_WH_1s(Tile_X9Y22_to_WH_1s),
    .from_WI_1s(Tile_X9Y22_to_WI_1s),
    .to_WA(Tile_X8Y22_to_WA),
    .to_WB(Tile_X8Y22_to_WB),
    .to_WC(Tile_X8Y22_to_WC),
    .to_WD(Tile_X8Y22_to_WD),
    .to_WF(Tile_X8Y22_to_WF),
    .to_WG(Tile_X8Y22_to_WG),
    .to_WH(Tile_X8Y22_to_WH),
    .to_WI(Tile_X8Y22_to_WI),
    .to_NA(Tile_X8Y22_to_NA),
    .to_NB(Tile_X8Y22_to_NB),
    .to_NC(Tile_X8Y22_to_NC),
    .to_ND(Tile_X8Y22_to_ND),
    .to_NF(Tile_X8Y22_to_NF),
    .to_NG(Tile_X8Y22_to_NG),
    .to_NH(Tile_X8Y22_to_NH),
    .to_NI(Tile_X8Y22_to_NI),
    .to_SA(Tile_X8Y22_to_SA),
    .to_SB(Tile_X8Y22_to_SB),
    .to_SC(Tile_X8Y22_to_SC),
    .to_SD(Tile_X8Y22_to_SD),
    .to_SF(Tile_X8Y22_to_SF),
    .to_SG(Tile_X8Y22_to_SG),
    .to_SH(Tile_X8Y22_to_SH),
    .to_SI(Tile_X8Y22_to_SI),
    .UserCLK(Tile_X8Y23_UserCLKo),
    .UserCLKo(Tile_X8Y22_UserCLKo),
    .rst(Tile_X8Y23_rsto),
    .rsto(Tile_X8Y22_rsto),
    .FrameData(Tile_X7Y22_FrameData_O),
    .FrameData_O(Tile_X8Y22_FrameData_O),
    .FrameStrobe(Tile_X8Y23_FrameStrobe_O),
    .FrameStrobe_O(Tile_X8Y22_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
combined_WDDL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X9Y22_Emulate_Bitstream)
    )
`endif
    Tile_X9Y22_combined_WDDL
    (
    .from_NA_1s(Tile_X9Y23_to_NA_1s),
    .from_NB_1s(Tile_X9Y23_to_NB_1s),
    .from_NC_1s(Tile_X9Y23_to_NC_1s),
    .from_ND_1s(Tile_X9Y23_to_ND_1s),
    .from_NF_1s(Tile_X9Y23_to_NF_1s),
    .from_NG_1s(Tile_X9Y23_to_NG_1s),
    .from_NH_1s(Tile_X9Y23_to_NH_1s),
    .from_NI_1s(Tile_X9Y23_to_NI_1s),
    .from_SA_1s(Tile_X9Y21_to_SA_1s),
    .from_SB_1s(Tile_X9Y21_to_SB_1s),
    .from_SC_1s(Tile_X9Y21_to_SC_1s),
    .from_SD_1s(Tile_X9Y21_to_SD_1s),
    .from_SF_1s(Tile_X9Y21_to_SF_1s),
    .from_SG_1s(Tile_X9Y21_to_SG_1s),
    .from_SH_1s(Tile_X9Y21_to_SH_1s),
    .from_SI_1s(Tile_X9Y21_to_SI_1s),
    .from_WA_1s(Tile_X10Y22_to_WA_1s),
    .from_WB_1s(Tile_X10Y22_to_WB_1s),
    .from_WC_1s(Tile_X10Y22_to_WC_1s),
    .from_WD_1s(Tile_X10Y22_to_WD_1s),
    .from_WF_1s(Tile_X10Y22_to_WF_1s),
    .from_WG_1s(Tile_X10Y22_to_WG_1s),
    .from_WH_1s(Tile_X10Y22_to_WH_1s),
    .from_WI_1s(Tile_X10Y22_to_WI_1s),
    .to_EA_1s(Tile_X9Y22_to_EA_1s),
    .to_EB_1s(Tile_X9Y22_to_EB_1s),
    .to_EC_1s(Tile_X9Y22_to_EC_1s),
    .to_ED_1s(Tile_X9Y22_to_ED_1s),
    .to_EF_1s(Tile_X9Y22_to_EF_1s),
    .to_EG_1s(Tile_X9Y22_to_EG_1s),
    .to_EH_1s(Tile_X9Y22_to_EH_1s),
    .to_EI_1s(Tile_X9Y22_to_EI_1s),
    .to_WA_1s(Tile_X9Y22_to_WA_1s),
    .to_WB_1s(Tile_X9Y22_to_WB_1s),
    .to_WC_1s(Tile_X9Y22_to_WC_1s),
    .to_WD_1s(Tile_X9Y22_to_WD_1s),
    .to_WF_1s(Tile_X9Y22_to_WF_1s),
    .to_WG_1s(Tile_X9Y22_to_WG_1s),
    .to_WH_1s(Tile_X9Y22_to_WH_1s),
    .to_WI_1s(Tile_X9Y22_to_WI_1s),
    .to_NA_1s(Tile_X9Y22_to_NA_1s),
    .to_NB_1s(Tile_X9Y22_to_NB_1s),
    .to_NC_1s(Tile_X9Y22_to_NC_1s),
    .to_ND_1s(Tile_X9Y22_to_ND_1s),
    .to_NF_1s(Tile_X9Y22_to_NF_1s),
    .to_NG_1s(Tile_X9Y22_to_NG_1s),
    .to_NH_1s(Tile_X9Y22_to_NH_1s),
    .to_NI_1s(Tile_X9Y22_to_NI_1s),
    .to_SA_1s(Tile_X9Y22_to_SA_1s),
    .to_SB_1s(Tile_X9Y22_to_SB_1s),
    .to_SC_1s(Tile_X9Y22_to_SC_1s),
    .to_SD_1s(Tile_X9Y22_to_SD_1s),
    .to_SF_1s(Tile_X9Y22_to_SF_1s),
    .to_SG_1s(Tile_X9Y22_to_SG_1s),
    .to_SH_1s(Tile_X9Y22_to_SH_1s),
    .to_SI_1s(Tile_X9Y22_to_SI_1s),
    .F_ctrl(Tile_X9Y22_F_ctrl),
    .UserCLK(Tile_X9Y23_UserCLKo),
    .UserCLKo(Tile_X9Y22_UserCLKo),
    .rst(Tile_X9Y23_rsto),
    .rsto(Tile_X9Y22_rsto),
    .FrameData(Tile_X8Y22_FrameData_O),
    .FrameData_O(Tile_X9Y22_FrameData_O),
    .FrameStrobe(Tile_X9Y23_FrameStrobe_O),
    .FrameStrobe_O(Tile_X9Y22_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
ctrl_IO
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X10Y22_Emulate_Bitstream)
    )
`endif
    Tile_X10Y22_ctrl_IO
    (
    .from_EA_1s(Tile_X9Y22_to_EA_1s),
    .from_EB_1s(Tile_X9Y22_to_EB_1s),
    .from_EC_1s(Tile_X9Y22_to_EC_1s),
    .from_ED_1s(Tile_X9Y22_to_ED_1s),
    .from_EF_1s(Tile_X9Y22_to_EF_1s),
    .from_EG_1s(Tile_X9Y22_to_EG_1s),
    .from_EH_1s(Tile_X9Y22_to_EH_1s),
    .from_EI_1s(Tile_X9Y22_to_EI_1s),
    .to_WA_1s(Tile_X10Y22_to_WA_1s),
    .to_WB_1s(Tile_X10Y22_to_WB_1s),
    .to_WC_1s(Tile_X10Y22_to_WC_1s),
    .to_WD_1s(Tile_X10Y22_to_WD_1s),
    .to_WF_1s(Tile_X10Y22_to_WF_1s),
    .to_WG_1s(Tile_X10Y22_to_WG_1s),
    .to_WH_1s(Tile_X10Y22_to_WH_1s),
    .to_WI_1s(Tile_X10Y22_to_WI_1s),
    .A_O_top_0_t(Tile_X10Y22_A_O_top_0_t),
    .A_O_top_0_f(Tile_X10Y22_A_O_top_0_f),
    .A_prech2(Tile_X10Y22_A_prech2),
    .A_DR_fault(Tile_X10Y22_A_DR_fault),
    .A_I_top_0_t(Tile_X10Y22_A_I_top_0_t),
    .A_I_top_0_f(Tile_X10Y22_A_I_top_0_f),
    .A_T_top(Tile_X10Y22_A_T_top),
    .A_F_ctrl(Tile_X10Y22_A_F_ctrl),
    .UserCLK(Tile_X10Y23_UserCLKo),
    .UserCLKo(Tile_X10Y22_UserCLKo),
    .rst(Tile_X10Y23_rsto),
    .rsto(Tile_X10Y22_rsto),
    .FrameData(Tile_X9Y22_FrameData_O),
    .FrameData_O(Tile_X10Y22_FrameData_O),
    .FrameStrobe(Tile_X10Y23_FrameStrobe_O),
    .FrameStrobe_O(Tile_X10Y22_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
W_IO_custom
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X0Y23_Emulate_Bitstream)
    )
`endif
    Tile_X0Y23_W_IO_custom
    (
    .from_NA(Tile_X0Y24_to_NA),
    .from_NB(Tile_X0Y24_to_NB),
    .from_NC(Tile_X0Y24_to_NC),
    .from_ND(Tile_X0Y24_to_ND),
    .from_NF(Tile_X0Y24_to_NF),
    .from_NG(Tile_X0Y24_to_NG),
    .from_NH(Tile_X0Y24_to_NH),
    .from_NI(Tile_X0Y24_to_NI),
    .from_SA(Tile_X0Y22_to_SA),
    .from_SB(Tile_X0Y22_to_SB),
    .from_SC(Tile_X0Y22_to_SC),
    .from_SD(Tile_X0Y22_to_SD),
    .from_SF(Tile_X0Y22_to_SF),
    .from_SG(Tile_X0Y22_to_SG),
    .from_SH(Tile_X0Y22_to_SH),
    .from_SI(Tile_X0Y22_to_SI),
    .from_WA(Tile_X1Y23_to_WA),
    .from_WB(Tile_X1Y23_to_WB),
    .from_WC(Tile_X1Y23_to_WC),
    .from_WD(Tile_X1Y23_to_WD),
    .from_WF(Tile_X1Y23_to_WF),
    .from_WG(Tile_X1Y23_to_WG),
    .from_WH(Tile_X1Y23_to_WH),
    .from_WI(Tile_X1Y23_to_WI),
    .to_EA(Tile_X0Y23_to_EA),
    .to_EB(Tile_X0Y23_to_EB),
    .to_EC(Tile_X0Y23_to_EC),
    .to_ED(Tile_X0Y23_to_ED),
    .to_EF(Tile_X0Y23_to_EF),
    .to_EG(Tile_X0Y23_to_EG),
    .to_EH(Tile_X0Y23_to_EH),
    .to_EI(Tile_X0Y23_to_EI),
    .to_NA(Tile_X0Y23_to_NA),
    .to_NB(Tile_X0Y23_to_NB),
    .to_NC(Tile_X0Y23_to_NC),
    .to_ND(Tile_X0Y23_to_ND),
    .to_NF(Tile_X0Y23_to_NF),
    .to_NG(Tile_X0Y23_to_NG),
    .to_NH(Tile_X0Y23_to_NH),
    .to_NI(Tile_X0Y23_to_NI),
    .to_SA(Tile_X0Y23_to_SA),
    .to_SB(Tile_X0Y23_to_SB),
    .to_SC(Tile_X0Y23_to_SC),
    .to_SD(Tile_X0Y23_to_SD),
    .to_SF(Tile_X0Y23_to_SF),
    .to_SG(Tile_X0Y23_to_SG),
    .to_SH(Tile_X0Y23_to_SH),
    .to_SI(Tile_X0Y23_to_SI),
    .A_O_top_0_t(Tile_X0Y23_A_O_top_0_t),
    .A_O_top_0_f(Tile_X0Y23_A_O_top_0_f),
    .A_O_top_1_t(Tile_X0Y23_A_O_top_1_t),
    .A_O_top_1_f(Tile_X0Y23_A_O_top_1_f),
    .A_prech1(Tile_X0Y23_A_prech1),
    .A_prech2(Tile_X0Y23_A_prech2),
    .A_DR_fault(Tile_X0Y23_A_DR_fault),
    .A_I_top_0_t(Tile_X0Y23_A_I_top_0_t),
    .A_I_top_0_f(Tile_X0Y23_A_I_top_0_f),
    .A_I_top_1_t(Tile_X0Y23_A_I_top_1_t),
    .A_I_top_1_f(Tile_X0Y23_A_I_top_1_f),
    .A_T_top(Tile_X0Y23_A_T_top),
    .A_F_masked1(Tile_X0Y23_A_F_masked1),
    .A_F_masked2(Tile_X0Y23_A_F_masked2),
    .A_config_C_bit0(Tile_X0Y23_A_config_C_bit0),
    .A_config_C_bit1(Tile_X0Y23_A_config_C_bit1),
    .A_config_C_bit2(Tile_X0Y23_A_config_C_bit2),
    .A_config_C_bit3(Tile_X0Y23_A_config_C_bit3),
    .B_config_C_bit0(Tile_X0Y23_B_config_C_bit0),
    .B_config_C_bit1(Tile_X0Y23_B_config_C_bit1),
    .B_config_C_bit2(Tile_X0Y23_B_config_C_bit2),
    .B_config_C_bit3(Tile_X0Y23_B_config_C_bit3),
    .UserCLK(Tile_X0Y24_UserCLKo),
    .UserCLKo(Tile_X0Y23_UserCLKo),
    .rst(Tile_X0Y24_rsto),
    .rsto(Tile_X0Y23_rsto),
    .FrameData(Tile_Y23_FrameData),
    .FrameData_O(Tile_X0Y23_FrameData_O),
    .FrameStrobe(Tile_X0Y24_FrameStrobe_O),
    .FrameStrobe_O(Tile_X0Y23_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X1Y23_Emulate_Bitstream)
    )
`endif
    Tile_X1Y23_linear_LMDPL
    (
    .from_NA(Tile_X1Y24_to_NA),
    .from_NB(Tile_X1Y24_to_NB),
    .from_NC(Tile_X1Y24_to_NC),
    .from_ND(Tile_X1Y24_to_ND),
    .from_NF(Tile_X1Y24_to_NF),
    .from_NG(Tile_X1Y24_to_NG),
    .from_NH(Tile_X1Y24_to_NH),
    .from_NI(Tile_X1Y24_to_NI),
    .from_EA(Tile_X0Y23_to_EA),
    .from_EB(Tile_X0Y23_to_EB),
    .from_EC(Tile_X0Y23_to_EC),
    .from_ED(Tile_X0Y23_to_ED),
    .from_EF(Tile_X0Y23_to_EF),
    .from_EG(Tile_X0Y23_to_EG),
    .from_EH(Tile_X0Y23_to_EH),
    .from_EI(Tile_X0Y23_to_EI),
    .from_SA(Tile_X1Y22_to_SA),
    .from_SB(Tile_X1Y22_to_SB),
    .from_SC(Tile_X1Y22_to_SC),
    .from_SD(Tile_X1Y22_to_SD),
    .from_SF(Tile_X1Y22_to_SF),
    .from_SG(Tile_X1Y22_to_SG),
    .from_SH(Tile_X1Y22_to_SH),
    .from_SI(Tile_X1Y22_to_SI),
    .from_WA(Tile_X2Y23_to_WA),
    .from_WB(Tile_X2Y23_to_WB),
    .from_WC(Tile_X2Y23_to_WC),
    .from_WD(Tile_X2Y23_to_WD),
    .from_WF(Tile_X2Y23_to_WF),
    .from_WG(Tile_X2Y23_to_WG),
    .from_WH(Tile_X2Y23_to_WH),
    .from_WI(Tile_X2Y23_to_WI),
    .to_EA(Tile_X1Y23_to_EA),
    .to_EB(Tile_X1Y23_to_EB),
    .to_EC(Tile_X1Y23_to_EC),
    .to_ED(Tile_X1Y23_to_ED),
    .to_EF(Tile_X1Y23_to_EF),
    .to_EG(Tile_X1Y23_to_EG),
    .to_EH(Tile_X1Y23_to_EH),
    .to_EI(Tile_X1Y23_to_EI),
    .to_WA(Tile_X1Y23_to_WA),
    .to_WB(Tile_X1Y23_to_WB),
    .to_WC(Tile_X1Y23_to_WC),
    .to_WD(Tile_X1Y23_to_WD),
    .to_WF(Tile_X1Y23_to_WF),
    .to_WG(Tile_X1Y23_to_WG),
    .to_WH(Tile_X1Y23_to_WH),
    .to_WI(Tile_X1Y23_to_WI),
    .to_NA(Tile_X1Y23_to_NA),
    .to_NB(Tile_X1Y23_to_NB),
    .to_NC(Tile_X1Y23_to_NC),
    .to_ND(Tile_X1Y23_to_ND),
    .to_NF(Tile_X1Y23_to_NF),
    .to_NG(Tile_X1Y23_to_NG),
    .to_NH(Tile_X1Y23_to_NH),
    .to_NI(Tile_X1Y23_to_NI),
    .to_SA(Tile_X1Y23_to_SA),
    .to_SB(Tile_X1Y23_to_SB),
    .to_SC(Tile_X1Y23_to_SC),
    .to_SD(Tile_X1Y23_to_SD),
    .to_SF(Tile_X1Y23_to_SF),
    .to_SG(Tile_X1Y23_to_SG),
    .to_SH(Tile_X1Y23_to_SH),
    .to_SI(Tile_X1Y23_to_SI),
    .F_masked1(Tile_X1Y23_F_masked1),
    .F_masked2(Tile_X1Y23_F_masked2),
    .UserCLK(Tile_X1Y24_UserCLKo),
    .UserCLKo(Tile_X1Y23_UserCLKo),
    .rst(Tile_X1Y24_rsto),
    .rsto(Tile_X1Y23_rsto),
    .FrameData(Tile_X0Y23_FrameData_O),
    .FrameData_O(Tile_X1Y23_FrameData_O),
    .FrameStrobe(Tile_X1Y24_FrameStrobe_O),
    .FrameStrobe_O(Tile_X1Y23_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X2Y23_Emulate_Bitstream)
    )
`endif
    Tile_X2Y23_linear_LMDPL
    (
    .from_NA(Tile_X2Y24_to_NA),
    .from_NB(Tile_X2Y24_to_NB),
    .from_NC(Tile_X2Y24_to_NC),
    .from_ND(Tile_X2Y24_to_ND),
    .from_NF(Tile_X2Y24_to_NF),
    .from_NG(Tile_X2Y24_to_NG),
    .from_NH(Tile_X2Y24_to_NH),
    .from_NI(Tile_X2Y24_to_NI),
    .from_EA(Tile_X1Y23_to_EA),
    .from_EB(Tile_X1Y23_to_EB),
    .from_EC(Tile_X1Y23_to_EC),
    .from_ED(Tile_X1Y23_to_ED),
    .from_EF(Tile_X1Y23_to_EF),
    .from_EG(Tile_X1Y23_to_EG),
    .from_EH(Tile_X1Y23_to_EH),
    .from_EI(Tile_X1Y23_to_EI),
    .from_SA(Tile_X2Y22_to_SA),
    .from_SB(Tile_X2Y22_to_SB),
    .from_SC(Tile_X2Y22_to_SC),
    .from_SD(Tile_X2Y22_to_SD),
    .from_SF(Tile_X2Y22_to_SF),
    .from_SG(Tile_X2Y22_to_SG),
    .from_SH(Tile_X2Y22_to_SH),
    .from_SI(Tile_X2Y22_to_SI),
    .from_WA(Tile_X3Y23_to_WA),
    .from_WB(Tile_X3Y23_to_WB),
    .from_WC(Tile_X3Y23_to_WC),
    .from_WD(Tile_X3Y23_to_WD),
    .from_WF(Tile_X3Y23_to_WF),
    .from_WG(Tile_X3Y23_to_WG),
    .from_WH(Tile_X3Y23_to_WH),
    .from_WI(Tile_X3Y23_to_WI),
    .to_EA(Tile_X2Y23_to_EA),
    .to_EB(Tile_X2Y23_to_EB),
    .to_EC(Tile_X2Y23_to_EC),
    .to_ED(Tile_X2Y23_to_ED),
    .to_EF(Tile_X2Y23_to_EF),
    .to_EG(Tile_X2Y23_to_EG),
    .to_EH(Tile_X2Y23_to_EH),
    .to_EI(Tile_X2Y23_to_EI),
    .to_WA(Tile_X2Y23_to_WA),
    .to_WB(Tile_X2Y23_to_WB),
    .to_WC(Tile_X2Y23_to_WC),
    .to_WD(Tile_X2Y23_to_WD),
    .to_WF(Tile_X2Y23_to_WF),
    .to_WG(Tile_X2Y23_to_WG),
    .to_WH(Tile_X2Y23_to_WH),
    .to_WI(Tile_X2Y23_to_WI),
    .to_NA(Tile_X2Y23_to_NA),
    .to_NB(Tile_X2Y23_to_NB),
    .to_NC(Tile_X2Y23_to_NC),
    .to_ND(Tile_X2Y23_to_ND),
    .to_NF(Tile_X2Y23_to_NF),
    .to_NG(Tile_X2Y23_to_NG),
    .to_NH(Tile_X2Y23_to_NH),
    .to_NI(Tile_X2Y23_to_NI),
    .to_SA(Tile_X2Y23_to_SA),
    .to_SB(Tile_X2Y23_to_SB),
    .to_SC(Tile_X2Y23_to_SC),
    .to_SD(Tile_X2Y23_to_SD),
    .to_SF(Tile_X2Y23_to_SF),
    .to_SG(Tile_X2Y23_to_SG),
    .to_SH(Tile_X2Y23_to_SH),
    .to_SI(Tile_X2Y23_to_SI),
    .F_masked1(Tile_X2Y23_F_masked1),
    .F_masked2(Tile_X2Y23_F_masked2),
    .UserCLK(Tile_X2Y24_UserCLKo),
    .UserCLKo(Tile_X2Y23_UserCLKo),
    .rst(Tile_X2Y24_rsto),
    .rsto(Tile_X2Y23_rsto),
    .FrameData(Tile_X1Y23_FrameData_O),
    .FrameData_O(Tile_X2Y23_FrameData_O),
    .FrameStrobe(Tile_X2Y24_FrameStrobe_O),
    .FrameStrobe_O(Tile_X2Y23_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
nonlinear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X3Y23_Emulate_Bitstream)
    )
`endif
    Tile_X3Y23_nonlinear_LMDPL
    (
    .from_NA(Tile_X3Y24_to_NA),
    .from_NB(Tile_X3Y24_to_NB),
    .from_NC(Tile_X3Y24_to_NC),
    .from_ND(Tile_X3Y24_to_ND),
    .from_NF(Tile_X3Y24_to_NF),
    .from_NG(Tile_X3Y24_to_NG),
    .from_NH(Tile_X3Y24_to_NH),
    .from_NI(Tile_X3Y24_to_NI),
    .from_EA(Tile_X2Y23_to_EA),
    .from_EB(Tile_X2Y23_to_EB),
    .from_EC(Tile_X2Y23_to_EC),
    .from_ED(Tile_X2Y23_to_ED),
    .from_EF(Tile_X2Y23_to_EF),
    .from_EG(Tile_X2Y23_to_EG),
    .from_EH(Tile_X2Y23_to_EH),
    .from_EI(Tile_X2Y23_to_EI),
    .from_SA(Tile_X3Y22_to_SA),
    .from_SB(Tile_X3Y22_to_SB),
    .from_SC(Tile_X3Y22_to_SC),
    .from_SD(Tile_X3Y22_to_SD),
    .from_SF(Tile_X3Y22_to_SF),
    .from_SG(Tile_X3Y22_to_SG),
    .from_SH(Tile_X3Y22_to_SH),
    .from_SI(Tile_X3Y22_to_SI),
    .from_WA(Tile_X4Y23_to_WA),
    .from_WB(Tile_X4Y23_to_WB),
    .from_WC(Tile_X4Y23_to_WC),
    .from_WD(Tile_X4Y23_to_WD),
    .from_WF(Tile_X4Y23_to_WF),
    .from_WG(Tile_X4Y23_to_WG),
    .from_WH(Tile_X4Y23_to_WH),
    .from_WI(Tile_X4Y23_to_WI),
    .to_EA(Tile_X3Y23_to_EA),
    .to_EB(Tile_X3Y23_to_EB),
    .to_EC(Tile_X3Y23_to_EC),
    .to_ED(Tile_X3Y23_to_ED),
    .to_EF(Tile_X3Y23_to_EF),
    .to_EG(Tile_X3Y23_to_EG),
    .to_EH(Tile_X3Y23_to_EH),
    .to_EI(Tile_X3Y23_to_EI),
    .to_WA(Tile_X3Y23_to_WA),
    .to_WB(Tile_X3Y23_to_WB),
    .to_WC(Tile_X3Y23_to_WC),
    .to_WD(Tile_X3Y23_to_WD),
    .to_WF(Tile_X3Y23_to_WF),
    .to_WG(Tile_X3Y23_to_WG),
    .to_WH(Tile_X3Y23_to_WH),
    .to_WI(Tile_X3Y23_to_WI),
    .to_NA(Tile_X3Y23_to_NA),
    .to_NB(Tile_X3Y23_to_NB),
    .to_NC(Tile_X3Y23_to_NC),
    .to_ND(Tile_X3Y23_to_ND),
    .to_NF(Tile_X3Y23_to_NF),
    .to_NG(Tile_X3Y23_to_NG),
    .to_NH(Tile_X3Y23_to_NH),
    .to_NI(Tile_X3Y23_to_NI),
    .to_SA(Tile_X3Y23_to_SA),
    .to_SB(Tile_X3Y23_to_SB),
    .to_SC(Tile_X3Y23_to_SC),
    .to_SD(Tile_X3Y23_to_SD),
    .to_SF(Tile_X3Y23_to_SF),
    .to_SG(Tile_X3Y23_to_SG),
    .to_SH(Tile_X3Y23_to_SH),
    .to_SI(Tile_X3Y23_to_SI),
    .R_t(Tile_X3Y23_R_t),
    .R_f(Tile_X3Y23_R_f),
    .F_masked1(Tile_X3Y23_F_masked1),
    .F_masked2(Tile_X3Y23_F_masked2),
    .UserCLK(Tile_X3Y24_UserCLKo),
    .UserCLKo(Tile_X3Y23_UserCLKo),
    .rst(Tile_X3Y24_rsto),
    .rsto(Tile_X3Y23_rsto),
    .FrameData(Tile_X2Y23_FrameData_O),
    .FrameData_O(Tile_X3Y23_FrameData_O),
    .FrameStrobe(Tile_X3Y24_FrameStrobe_O),
    .FrameStrobe_O(Tile_X3Y23_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X4Y23_Emulate_Bitstream)
    )
`endif
    Tile_X4Y23_linear_LMDPL
    (
    .from_NA(Tile_X4Y24_to_NA),
    .from_NB(Tile_X4Y24_to_NB),
    .from_NC(Tile_X4Y24_to_NC),
    .from_ND(Tile_X4Y24_to_ND),
    .from_NF(Tile_X4Y24_to_NF),
    .from_NG(Tile_X4Y24_to_NG),
    .from_NH(Tile_X4Y24_to_NH),
    .from_NI(Tile_X4Y24_to_NI),
    .from_EA(Tile_X3Y23_to_EA),
    .from_EB(Tile_X3Y23_to_EB),
    .from_EC(Tile_X3Y23_to_EC),
    .from_ED(Tile_X3Y23_to_ED),
    .from_EF(Tile_X3Y23_to_EF),
    .from_EG(Tile_X3Y23_to_EG),
    .from_EH(Tile_X3Y23_to_EH),
    .from_EI(Tile_X3Y23_to_EI),
    .from_SA(Tile_X4Y22_to_SA),
    .from_SB(Tile_X4Y22_to_SB),
    .from_SC(Tile_X4Y22_to_SC),
    .from_SD(Tile_X4Y22_to_SD),
    .from_SF(Tile_X4Y22_to_SF),
    .from_SG(Tile_X4Y22_to_SG),
    .from_SH(Tile_X4Y22_to_SH),
    .from_SI(Tile_X4Y22_to_SI),
    .from_WA(Tile_X5Y23_to_WA),
    .from_WB(Tile_X5Y23_to_WB),
    .from_WC(Tile_X5Y23_to_WC),
    .from_WD(Tile_X5Y23_to_WD),
    .from_WF(Tile_X5Y23_to_WF),
    .from_WG(Tile_X5Y23_to_WG),
    .from_WH(Tile_X5Y23_to_WH),
    .from_WI(Tile_X5Y23_to_WI),
    .to_EA(Tile_X4Y23_to_EA),
    .to_EB(Tile_X4Y23_to_EB),
    .to_EC(Tile_X4Y23_to_EC),
    .to_ED(Tile_X4Y23_to_ED),
    .to_EF(Tile_X4Y23_to_EF),
    .to_EG(Tile_X4Y23_to_EG),
    .to_EH(Tile_X4Y23_to_EH),
    .to_EI(Tile_X4Y23_to_EI),
    .to_WA(Tile_X4Y23_to_WA),
    .to_WB(Tile_X4Y23_to_WB),
    .to_WC(Tile_X4Y23_to_WC),
    .to_WD(Tile_X4Y23_to_WD),
    .to_WF(Tile_X4Y23_to_WF),
    .to_WG(Tile_X4Y23_to_WG),
    .to_WH(Tile_X4Y23_to_WH),
    .to_WI(Tile_X4Y23_to_WI),
    .to_NA(Tile_X4Y23_to_NA),
    .to_NB(Tile_X4Y23_to_NB),
    .to_NC(Tile_X4Y23_to_NC),
    .to_ND(Tile_X4Y23_to_ND),
    .to_NF(Tile_X4Y23_to_NF),
    .to_NG(Tile_X4Y23_to_NG),
    .to_NH(Tile_X4Y23_to_NH),
    .to_NI(Tile_X4Y23_to_NI),
    .to_SA(Tile_X4Y23_to_SA),
    .to_SB(Tile_X4Y23_to_SB),
    .to_SC(Tile_X4Y23_to_SC),
    .to_SD(Tile_X4Y23_to_SD),
    .to_SF(Tile_X4Y23_to_SF),
    .to_SG(Tile_X4Y23_to_SG),
    .to_SH(Tile_X4Y23_to_SH),
    .to_SI(Tile_X4Y23_to_SI),
    .F_masked1(Tile_X4Y23_F_masked1),
    .F_masked2(Tile_X4Y23_F_masked2),
    .UserCLK(Tile_X4Y24_UserCLKo),
    .UserCLKo(Tile_X4Y23_UserCLKo),
    .rst(Tile_X4Y24_rsto),
    .rsto(Tile_X4Y23_rsto),
    .FrameData(Tile_X3Y23_FrameData_O),
    .FrameData_O(Tile_X4Y23_FrameData_O),
    .FrameStrobe(Tile_X4Y24_FrameStrobe_O),
    .FrameStrobe_O(Tile_X4Y23_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X5Y23_Emulate_Bitstream)
    )
`endif
    Tile_X5Y23_linear_LMDPL
    (
    .from_NA(Tile_X5Y24_to_NA),
    .from_NB(Tile_X5Y24_to_NB),
    .from_NC(Tile_X5Y24_to_NC),
    .from_ND(Tile_X5Y24_to_ND),
    .from_NF(Tile_X5Y24_to_NF),
    .from_NG(Tile_X5Y24_to_NG),
    .from_NH(Tile_X5Y24_to_NH),
    .from_NI(Tile_X5Y24_to_NI),
    .from_EA(Tile_X4Y23_to_EA),
    .from_EB(Tile_X4Y23_to_EB),
    .from_EC(Tile_X4Y23_to_EC),
    .from_ED(Tile_X4Y23_to_ED),
    .from_EF(Tile_X4Y23_to_EF),
    .from_EG(Tile_X4Y23_to_EG),
    .from_EH(Tile_X4Y23_to_EH),
    .from_EI(Tile_X4Y23_to_EI),
    .from_SA(Tile_X5Y22_to_SA),
    .from_SB(Tile_X5Y22_to_SB),
    .from_SC(Tile_X5Y22_to_SC),
    .from_SD(Tile_X5Y22_to_SD),
    .from_SF(Tile_X5Y22_to_SF),
    .from_SG(Tile_X5Y22_to_SG),
    .from_SH(Tile_X5Y22_to_SH),
    .from_SI(Tile_X5Y22_to_SI),
    .from_WA(Tile_X6Y23_to_WA),
    .from_WB(Tile_X6Y23_to_WB),
    .from_WC(Tile_X6Y23_to_WC),
    .from_WD(Tile_X6Y23_to_WD),
    .from_WF(Tile_X6Y23_to_WF),
    .from_WG(Tile_X6Y23_to_WG),
    .from_WH(Tile_X6Y23_to_WH),
    .from_WI(Tile_X6Y23_to_WI),
    .to_EA(Tile_X5Y23_to_EA),
    .to_EB(Tile_X5Y23_to_EB),
    .to_EC(Tile_X5Y23_to_EC),
    .to_ED(Tile_X5Y23_to_ED),
    .to_EF(Tile_X5Y23_to_EF),
    .to_EG(Tile_X5Y23_to_EG),
    .to_EH(Tile_X5Y23_to_EH),
    .to_EI(Tile_X5Y23_to_EI),
    .to_WA(Tile_X5Y23_to_WA),
    .to_WB(Tile_X5Y23_to_WB),
    .to_WC(Tile_X5Y23_to_WC),
    .to_WD(Tile_X5Y23_to_WD),
    .to_WF(Tile_X5Y23_to_WF),
    .to_WG(Tile_X5Y23_to_WG),
    .to_WH(Tile_X5Y23_to_WH),
    .to_WI(Tile_X5Y23_to_WI),
    .to_NA(Tile_X5Y23_to_NA),
    .to_NB(Tile_X5Y23_to_NB),
    .to_NC(Tile_X5Y23_to_NC),
    .to_ND(Tile_X5Y23_to_ND),
    .to_NF(Tile_X5Y23_to_NF),
    .to_NG(Tile_X5Y23_to_NG),
    .to_NH(Tile_X5Y23_to_NH),
    .to_NI(Tile_X5Y23_to_NI),
    .to_SA(Tile_X5Y23_to_SA),
    .to_SB(Tile_X5Y23_to_SB),
    .to_SC(Tile_X5Y23_to_SC),
    .to_SD(Tile_X5Y23_to_SD),
    .to_SF(Tile_X5Y23_to_SF),
    .to_SG(Tile_X5Y23_to_SG),
    .to_SH(Tile_X5Y23_to_SH),
    .to_SI(Tile_X5Y23_to_SI),
    .F_masked1(Tile_X5Y23_F_masked1),
    .F_masked2(Tile_X5Y23_F_masked2),
    .UserCLK(Tile_X5Y24_UserCLKo),
    .UserCLKo(Tile_X5Y23_UserCLKo),
    .rst(Tile_X5Y24_rsto),
    .rsto(Tile_X5Y23_rsto),
    .FrameData(Tile_X4Y23_FrameData_O),
    .FrameData_O(Tile_X5Y23_FrameData_O),
    .FrameStrobe(Tile_X5Y24_FrameStrobe_O),
    .FrameStrobe_O(Tile_X5Y23_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
nonlinear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X6Y23_Emulate_Bitstream)
    )
`endif
    Tile_X6Y23_nonlinear_LMDPL
    (
    .from_NA(Tile_X6Y24_to_NA),
    .from_NB(Tile_X6Y24_to_NB),
    .from_NC(Tile_X6Y24_to_NC),
    .from_ND(Tile_X6Y24_to_ND),
    .from_NF(Tile_X6Y24_to_NF),
    .from_NG(Tile_X6Y24_to_NG),
    .from_NH(Tile_X6Y24_to_NH),
    .from_NI(Tile_X6Y24_to_NI),
    .from_EA(Tile_X5Y23_to_EA),
    .from_EB(Tile_X5Y23_to_EB),
    .from_EC(Tile_X5Y23_to_EC),
    .from_ED(Tile_X5Y23_to_ED),
    .from_EF(Tile_X5Y23_to_EF),
    .from_EG(Tile_X5Y23_to_EG),
    .from_EH(Tile_X5Y23_to_EH),
    .from_EI(Tile_X5Y23_to_EI),
    .from_SA(Tile_X6Y22_to_SA),
    .from_SB(Tile_X6Y22_to_SB),
    .from_SC(Tile_X6Y22_to_SC),
    .from_SD(Tile_X6Y22_to_SD),
    .from_SF(Tile_X6Y22_to_SF),
    .from_SG(Tile_X6Y22_to_SG),
    .from_SH(Tile_X6Y22_to_SH),
    .from_SI(Tile_X6Y22_to_SI),
    .from_WA(Tile_X7Y23_to_WA),
    .from_WB(Tile_X7Y23_to_WB),
    .from_WC(Tile_X7Y23_to_WC),
    .from_WD(Tile_X7Y23_to_WD),
    .from_WF(Tile_X7Y23_to_WF),
    .from_WG(Tile_X7Y23_to_WG),
    .from_WH(Tile_X7Y23_to_WH),
    .from_WI(Tile_X7Y23_to_WI),
    .to_EA(Tile_X6Y23_to_EA),
    .to_EB(Tile_X6Y23_to_EB),
    .to_EC(Tile_X6Y23_to_EC),
    .to_ED(Tile_X6Y23_to_ED),
    .to_EF(Tile_X6Y23_to_EF),
    .to_EG(Tile_X6Y23_to_EG),
    .to_EH(Tile_X6Y23_to_EH),
    .to_EI(Tile_X6Y23_to_EI),
    .to_WA(Tile_X6Y23_to_WA),
    .to_WB(Tile_X6Y23_to_WB),
    .to_WC(Tile_X6Y23_to_WC),
    .to_WD(Tile_X6Y23_to_WD),
    .to_WF(Tile_X6Y23_to_WF),
    .to_WG(Tile_X6Y23_to_WG),
    .to_WH(Tile_X6Y23_to_WH),
    .to_WI(Tile_X6Y23_to_WI),
    .to_NA(Tile_X6Y23_to_NA),
    .to_NB(Tile_X6Y23_to_NB),
    .to_NC(Tile_X6Y23_to_NC),
    .to_ND(Tile_X6Y23_to_ND),
    .to_NF(Tile_X6Y23_to_NF),
    .to_NG(Tile_X6Y23_to_NG),
    .to_NH(Tile_X6Y23_to_NH),
    .to_NI(Tile_X6Y23_to_NI),
    .to_SA(Tile_X6Y23_to_SA),
    .to_SB(Tile_X6Y23_to_SB),
    .to_SC(Tile_X6Y23_to_SC),
    .to_SD(Tile_X6Y23_to_SD),
    .to_SF(Tile_X6Y23_to_SF),
    .to_SG(Tile_X6Y23_to_SG),
    .to_SH(Tile_X6Y23_to_SH),
    .to_SI(Tile_X6Y23_to_SI),
    .R_t(Tile_X6Y23_R_t),
    .R_f(Tile_X6Y23_R_f),
    .F_masked1(Tile_X6Y23_F_masked1),
    .F_masked2(Tile_X6Y23_F_masked2),
    .UserCLK(Tile_X6Y24_UserCLKo),
    .UserCLKo(Tile_X6Y23_UserCLKo),
    .rst(Tile_X6Y24_rsto),
    .rsto(Tile_X6Y23_rsto),
    .FrameData(Tile_X5Y23_FrameData_O),
    .FrameData_O(Tile_X6Y23_FrameData_O),
    .FrameStrobe(Tile_X6Y24_FrameStrobe_O),
    .FrameStrobe_O(Tile_X6Y23_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
linear_LMDPL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X7Y23_Emulate_Bitstream)
    )
`endif
    Tile_X7Y23_linear_LMDPL
    (
    .from_NA(Tile_X7Y24_to_NA),
    .from_NB(Tile_X7Y24_to_NB),
    .from_NC(Tile_X7Y24_to_NC),
    .from_ND(Tile_X7Y24_to_ND),
    .from_NF(Tile_X7Y24_to_NF),
    .from_NG(Tile_X7Y24_to_NG),
    .from_NH(Tile_X7Y24_to_NH),
    .from_NI(Tile_X7Y24_to_NI),
    .from_EA(Tile_X6Y23_to_EA),
    .from_EB(Tile_X6Y23_to_EB),
    .from_EC(Tile_X6Y23_to_EC),
    .from_ED(Tile_X6Y23_to_ED),
    .from_EF(Tile_X6Y23_to_EF),
    .from_EG(Tile_X6Y23_to_EG),
    .from_EH(Tile_X6Y23_to_EH),
    .from_EI(Tile_X6Y23_to_EI),
    .from_SA(Tile_X7Y22_to_SA),
    .from_SB(Tile_X7Y22_to_SB),
    .from_SC(Tile_X7Y22_to_SC),
    .from_SD(Tile_X7Y22_to_SD),
    .from_SF(Tile_X7Y22_to_SF),
    .from_SG(Tile_X7Y22_to_SG),
    .from_SH(Tile_X7Y22_to_SH),
    .from_SI(Tile_X7Y22_to_SI),
    .from_WA(Tile_X8Y23_to_WA),
    .from_WB(Tile_X8Y23_to_WB),
    .from_WC(Tile_X8Y23_to_WC),
    .from_WD(Tile_X8Y23_to_WD),
    .from_WF(Tile_X8Y23_to_WF),
    .from_WG(Tile_X8Y23_to_WG),
    .from_WH(Tile_X8Y23_to_WH),
    .from_WI(Tile_X8Y23_to_WI),
    .to_EA(Tile_X7Y23_to_EA),
    .to_EB(Tile_X7Y23_to_EB),
    .to_EC(Tile_X7Y23_to_EC),
    .to_ED(Tile_X7Y23_to_ED),
    .to_EF(Tile_X7Y23_to_EF),
    .to_EG(Tile_X7Y23_to_EG),
    .to_EH(Tile_X7Y23_to_EH),
    .to_EI(Tile_X7Y23_to_EI),
    .to_WA(Tile_X7Y23_to_WA),
    .to_WB(Tile_X7Y23_to_WB),
    .to_WC(Tile_X7Y23_to_WC),
    .to_WD(Tile_X7Y23_to_WD),
    .to_WF(Tile_X7Y23_to_WF),
    .to_WG(Tile_X7Y23_to_WG),
    .to_WH(Tile_X7Y23_to_WH),
    .to_WI(Tile_X7Y23_to_WI),
    .to_NA(Tile_X7Y23_to_NA),
    .to_NB(Tile_X7Y23_to_NB),
    .to_NC(Tile_X7Y23_to_NC),
    .to_ND(Tile_X7Y23_to_ND),
    .to_NF(Tile_X7Y23_to_NF),
    .to_NG(Tile_X7Y23_to_NG),
    .to_NH(Tile_X7Y23_to_NH),
    .to_NI(Tile_X7Y23_to_NI),
    .to_SA(Tile_X7Y23_to_SA),
    .to_SB(Tile_X7Y23_to_SB),
    .to_SC(Tile_X7Y23_to_SC),
    .to_SD(Tile_X7Y23_to_SD),
    .to_SF(Tile_X7Y23_to_SF),
    .to_SG(Tile_X7Y23_to_SG),
    .to_SH(Tile_X7Y23_to_SH),
    .to_SI(Tile_X7Y23_to_SI),
    .F_masked1(Tile_X7Y23_F_masked1),
    .F_masked2(Tile_X7Y23_F_masked2),
    .UserCLK(Tile_X7Y24_UserCLKo),
    .UserCLKo(Tile_X7Y23_UserCLKo),
    .rst(Tile_X7Y24_rsto),
    .rsto(Tile_X7Y23_rsto),
    .FrameData(Tile_X6Y23_FrameData_O),
    .FrameData_O(Tile_X7Y23_FrameData_O),
    .FrameStrobe(Tile_X7Y24_FrameStrobe_O),
    .FrameStrobe_O(Tile_X7Y23_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
ctrl_to_sec
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X8Y23_Emulate_Bitstream)
    )
`endif
    Tile_X8Y23_ctrl_to_sec
    (
    .from_NA(Tile_X8Y24_to_NA),
    .from_NB(Tile_X8Y24_to_NB),
    .from_NC(Tile_X8Y24_to_NC),
    .from_ND(Tile_X8Y24_to_ND),
    .from_NF(Tile_X8Y24_to_NF),
    .from_NG(Tile_X8Y24_to_NG),
    .from_NH(Tile_X8Y24_to_NH),
    .from_NI(Tile_X8Y24_to_NI),
    .from_EA(Tile_X7Y23_to_EA),
    .from_EB(Tile_X7Y23_to_EB),
    .from_EC(Tile_X7Y23_to_EC),
    .from_ED(Tile_X7Y23_to_ED),
    .from_EF(Tile_X7Y23_to_EF),
    .from_EG(Tile_X7Y23_to_EG),
    .from_EH(Tile_X7Y23_to_EH),
    .from_EI(Tile_X7Y23_to_EI),
    .from_SA(Tile_X8Y22_to_SA),
    .from_SB(Tile_X8Y22_to_SB),
    .from_SC(Tile_X8Y22_to_SC),
    .from_SD(Tile_X8Y22_to_SD),
    .from_SF(Tile_X8Y22_to_SF),
    .from_SG(Tile_X8Y22_to_SG),
    .from_SH(Tile_X8Y22_to_SH),
    .from_SI(Tile_X8Y22_to_SI),
    .from_WA_1s(Tile_X9Y23_to_WA_1s),
    .from_WB_1s(Tile_X9Y23_to_WB_1s),
    .from_WC_1s(Tile_X9Y23_to_WC_1s),
    .from_WD_1s(Tile_X9Y23_to_WD_1s),
    .from_WF_1s(Tile_X9Y23_to_WF_1s),
    .from_WG_1s(Tile_X9Y23_to_WG_1s),
    .from_WH_1s(Tile_X9Y23_to_WH_1s),
    .from_WI_1s(Tile_X9Y23_to_WI_1s),
    .to_WA(Tile_X8Y23_to_WA),
    .to_WB(Tile_X8Y23_to_WB),
    .to_WC(Tile_X8Y23_to_WC),
    .to_WD(Tile_X8Y23_to_WD),
    .to_WF(Tile_X8Y23_to_WF),
    .to_WG(Tile_X8Y23_to_WG),
    .to_WH(Tile_X8Y23_to_WH),
    .to_WI(Tile_X8Y23_to_WI),
    .to_NA(Tile_X8Y23_to_NA),
    .to_NB(Tile_X8Y23_to_NB),
    .to_NC(Tile_X8Y23_to_NC),
    .to_ND(Tile_X8Y23_to_ND),
    .to_NF(Tile_X8Y23_to_NF),
    .to_NG(Tile_X8Y23_to_NG),
    .to_NH(Tile_X8Y23_to_NH),
    .to_NI(Tile_X8Y23_to_NI),
    .to_SA(Tile_X8Y23_to_SA),
    .to_SB(Tile_X8Y23_to_SB),
    .to_SC(Tile_X8Y23_to_SC),
    .to_SD(Tile_X8Y23_to_SD),
    .to_SF(Tile_X8Y23_to_SF),
    .to_SG(Tile_X8Y23_to_SG),
    .to_SH(Tile_X8Y23_to_SH),
    .to_SI(Tile_X8Y23_to_SI),
    .UserCLK(Tile_X8Y24_UserCLKo),
    .UserCLKo(Tile_X8Y23_UserCLKo),
    .rst(Tile_X8Y24_rsto),
    .rsto(Tile_X8Y23_rsto),
    .FrameData(Tile_X7Y23_FrameData_O),
    .FrameData_O(Tile_X8Y23_FrameData_O),
    .FrameStrobe(Tile_X8Y24_FrameStrobe_O),
    .FrameStrobe_O(Tile_X8Y23_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
combined_WDDL
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X9Y23_Emulate_Bitstream)
    )
`endif
    Tile_X9Y23_combined_WDDL
    (
    .from_NA_1s(Tile_X9Y24_to_NA_1s),
    .from_NB_1s(Tile_X9Y24_to_NB_1s),
    .from_NC_1s(Tile_X9Y24_to_NC_1s),
    .from_ND_1s(Tile_X9Y24_to_ND_1s),
    .from_NF_1s(Tile_X9Y24_to_NF_1s),
    .from_NG_1s(Tile_X9Y24_to_NG_1s),
    .from_NH_1s(Tile_X9Y24_to_NH_1s),
    .from_NI_1s(Tile_X9Y24_to_NI_1s),
    .from_SA_1s(Tile_X9Y22_to_SA_1s),
    .from_SB_1s(Tile_X9Y22_to_SB_1s),
    .from_SC_1s(Tile_X9Y22_to_SC_1s),
    .from_SD_1s(Tile_X9Y22_to_SD_1s),
    .from_SF_1s(Tile_X9Y22_to_SF_1s),
    .from_SG_1s(Tile_X9Y22_to_SG_1s),
    .from_SH_1s(Tile_X9Y22_to_SH_1s),
    .from_SI_1s(Tile_X9Y22_to_SI_1s),
    .from_WA_1s(Tile_X10Y23_to_WA_1s),
    .from_WB_1s(Tile_X10Y23_to_WB_1s),
    .from_WC_1s(Tile_X10Y23_to_WC_1s),
    .from_WD_1s(Tile_X10Y23_to_WD_1s),
    .from_WF_1s(Tile_X10Y23_to_WF_1s),
    .from_WG_1s(Tile_X10Y23_to_WG_1s),
    .from_WH_1s(Tile_X10Y23_to_WH_1s),
    .from_WI_1s(Tile_X10Y23_to_WI_1s),
    .to_EA_1s(Tile_X9Y23_to_EA_1s),
    .to_EB_1s(Tile_X9Y23_to_EB_1s),
    .to_EC_1s(Tile_X9Y23_to_EC_1s),
    .to_ED_1s(Tile_X9Y23_to_ED_1s),
    .to_EF_1s(Tile_X9Y23_to_EF_1s),
    .to_EG_1s(Tile_X9Y23_to_EG_1s),
    .to_EH_1s(Tile_X9Y23_to_EH_1s),
    .to_EI_1s(Tile_X9Y23_to_EI_1s),
    .to_WA_1s(Tile_X9Y23_to_WA_1s),
    .to_WB_1s(Tile_X9Y23_to_WB_1s),
    .to_WC_1s(Tile_X9Y23_to_WC_1s),
    .to_WD_1s(Tile_X9Y23_to_WD_1s),
    .to_WF_1s(Tile_X9Y23_to_WF_1s),
    .to_WG_1s(Tile_X9Y23_to_WG_1s),
    .to_WH_1s(Tile_X9Y23_to_WH_1s),
    .to_WI_1s(Tile_X9Y23_to_WI_1s),
    .to_NA_1s(Tile_X9Y23_to_NA_1s),
    .to_NB_1s(Tile_X9Y23_to_NB_1s),
    .to_NC_1s(Tile_X9Y23_to_NC_1s),
    .to_ND_1s(Tile_X9Y23_to_ND_1s),
    .to_NF_1s(Tile_X9Y23_to_NF_1s),
    .to_NG_1s(Tile_X9Y23_to_NG_1s),
    .to_NH_1s(Tile_X9Y23_to_NH_1s),
    .to_NI_1s(Tile_X9Y23_to_NI_1s),
    .to_SA_1s(Tile_X9Y23_to_SA_1s),
    .to_SB_1s(Tile_X9Y23_to_SB_1s),
    .to_SC_1s(Tile_X9Y23_to_SC_1s),
    .to_SD_1s(Tile_X9Y23_to_SD_1s),
    .to_SF_1s(Tile_X9Y23_to_SF_1s),
    .to_SG_1s(Tile_X9Y23_to_SG_1s),
    .to_SH_1s(Tile_X9Y23_to_SH_1s),
    .to_SI_1s(Tile_X9Y23_to_SI_1s),
    .F_ctrl(Tile_X9Y23_F_ctrl),
    .UserCLK(Tile_X9Y24_UserCLKo),
    .UserCLKo(Tile_X9Y23_UserCLKo),
    .rst(Tile_X9Y24_rsto),
    .rsto(Tile_X9Y23_rsto),
    .FrameData(Tile_X8Y23_FrameData_O),
    .FrameData_O(Tile_X9Y23_FrameData_O),
    .FrameStrobe(Tile_X9Y24_FrameStrobe_O),
    .FrameStrobe_O(Tile_X9Y23_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
ctrl_IO
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X10Y23_Emulate_Bitstream)
    )
`endif
    Tile_X10Y23_ctrl_IO
    (
    .from_EA_1s(Tile_X9Y23_to_EA_1s),
    .from_EB_1s(Tile_X9Y23_to_EB_1s),
    .from_EC_1s(Tile_X9Y23_to_EC_1s),
    .from_ED_1s(Tile_X9Y23_to_ED_1s),
    .from_EF_1s(Tile_X9Y23_to_EF_1s),
    .from_EG_1s(Tile_X9Y23_to_EG_1s),
    .from_EH_1s(Tile_X9Y23_to_EH_1s),
    .from_EI_1s(Tile_X9Y23_to_EI_1s),
    .to_WA_1s(Tile_X10Y23_to_WA_1s),
    .to_WB_1s(Tile_X10Y23_to_WB_1s),
    .to_WC_1s(Tile_X10Y23_to_WC_1s),
    .to_WD_1s(Tile_X10Y23_to_WD_1s),
    .to_WF_1s(Tile_X10Y23_to_WF_1s),
    .to_WG_1s(Tile_X10Y23_to_WG_1s),
    .to_WH_1s(Tile_X10Y23_to_WH_1s),
    .to_WI_1s(Tile_X10Y23_to_WI_1s),
    .A_O_top_0_t(Tile_X10Y23_A_O_top_0_t),
    .A_O_top_0_f(Tile_X10Y23_A_O_top_0_f),
    .A_prech2(Tile_X10Y23_A_prech2),
    .A_DR_fault(Tile_X10Y23_A_DR_fault),
    .A_I_top_0_t(Tile_X10Y23_A_I_top_0_t),
    .A_I_top_0_f(Tile_X10Y23_A_I_top_0_f),
    .A_T_top(Tile_X10Y23_A_T_top),
    .A_F_ctrl(Tile_X10Y23_A_F_ctrl),
    .UserCLK(Tile_X10Y24_UserCLKo),
    .UserCLKo(Tile_X10Y23_UserCLKo),
    .rst(Tile_X10Y24_rsto),
    .rsto(Tile_X10Y23_rsto),
    .FrameData(Tile_X9Y23_FrameData_O),
    .FrameData_O(Tile_X10Y23_FrameData_O),
    .FrameStrobe(Tile_X10Y24_FrameStrobe_O),
    .FrameStrobe_O(Tile_X10Y23_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
S_term_custom Tile_X0Y24_S_term_custom (
    .from_SA(Tile_X0Y23_to_SA),
    .from_SB(Tile_X0Y23_to_SB),
    .from_SC(Tile_X0Y23_to_SC),
    .from_SD(Tile_X0Y23_to_SD),
    .from_SF(Tile_X0Y23_to_SF),
    .from_SG(Tile_X0Y23_to_SG),
    .from_SH(Tile_X0Y23_to_SH),
    .from_SI(Tile_X0Y23_to_SI),
    .to_NA(Tile_X0Y24_to_NA),
    .to_NB(Tile_X0Y24_to_NB),
    .to_NC(Tile_X0Y24_to_NC),
    .to_ND(Tile_X0Y24_to_ND),
    .to_NF(Tile_X0Y24_to_NF),
    .to_NG(Tile_X0Y24_to_NG),
    .to_NH(Tile_X0Y24_to_NH),
    .to_NI(Tile_X0Y24_to_NI),
    .UserCLK(UserCLK),
    .UserCLKo(Tile_X0Y24_UserCLKo),
    .rst(rst),
    .rsto(Tile_X0Y24_rsto),
    .FrameStrobe(Tile_X0_FrameStrobe),
    .FrameStrobe_O(Tile_X0Y24_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
S_term_custom Tile_X1Y24_S_term_custom (
    .from_SA(Tile_X1Y23_to_SA),
    .from_SB(Tile_X1Y23_to_SB),
    .from_SC(Tile_X1Y23_to_SC),
    .from_SD(Tile_X1Y23_to_SD),
    .from_SF(Tile_X1Y23_to_SF),
    .from_SG(Tile_X1Y23_to_SG),
    .from_SH(Tile_X1Y23_to_SH),
    .from_SI(Tile_X1Y23_to_SI),
    .to_NA(Tile_X1Y24_to_NA),
    .to_NB(Tile_X1Y24_to_NB),
    .to_NC(Tile_X1Y24_to_NC),
    .to_ND(Tile_X1Y24_to_ND),
    .to_NF(Tile_X1Y24_to_NF),
    .to_NG(Tile_X1Y24_to_NG),
    .to_NH(Tile_X1Y24_to_NH),
    .to_NI(Tile_X1Y24_to_NI),
    .UserCLK(UserCLK),
    .UserCLKo(Tile_X1Y24_UserCLKo),
    .rst(rst),
    .rsto(Tile_X1Y24_rsto),
    .FrameStrobe(Tile_X1_FrameStrobe),
    .FrameStrobe_O(Tile_X1Y24_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
S_term_custom Tile_X2Y24_S_term_custom (
    .from_SA(Tile_X2Y23_to_SA),
    .from_SB(Tile_X2Y23_to_SB),
    .from_SC(Tile_X2Y23_to_SC),
    .from_SD(Tile_X2Y23_to_SD),
    .from_SF(Tile_X2Y23_to_SF),
    .from_SG(Tile_X2Y23_to_SG),
    .from_SH(Tile_X2Y23_to_SH),
    .from_SI(Tile_X2Y23_to_SI),
    .to_NA(Tile_X2Y24_to_NA),
    .to_NB(Tile_X2Y24_to_NB),
    .to_NC(Tile_X2Y24_to_NC),
    .to_ND(Tile_X2Y24_to_ND),
    .to_NF(Tile_X2Y24_to_NF),
    .to_NG(Tile_X2Y24_to_NG),
    .to_NH(Tile_X2Y24_to_NH),
    .to_NI(Tile_X2Y24_to_NI),
    .UserCLK(UserCLK),
    .UserCLKo(Tile_X2Y24_UserCLKo),
    .rst(rst),
    .rsto(Tile_X2Y24_rsto),
    .FrameStrobe(Tile_X2_FrameStrobe),
    .FrameStrobe_O(Tile_X2Y24_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
S_term_custom Tile_X3Y24_S_term_custom (
    .from_SA(Tile_X3Y23_to_SA),
    .from_SB(Tile_X3Y23_to_SB),
    .from_SC(Tile_X3Y23_to_SC),
    .from_SD(Tile_X3Y23_to_SD),
    .from_SF(Tile_X3Y23_to_SF),
    .from_SG(Tile_X3Y23_to_SG),
    .from_SH(Tile_X3Y23_to_SH),
    .from_SI(Tile_X3Y23_to_SI),
    .to_NA(Tile_X3Y24_to_NA),
    .to_NB(Tile_X3Y24_to_NB),
    .to_NC(Tile_X3Y24_to_NC),
    .to_ND(Tile_X3Y24_to_ND),
    .to_NF(Tile_X3Y24_to_NF),
    .to_NG(Tile_X3Y24_to_NG),
    .to_NH(Tile_X3Y24_to_NH),
    .to_NI(Tile_X3Y24_to_NI),
    .UserCLK(UserCLK),
    .UserCLKo(Tile_X3Y24_UserCLKo),
    .rst(rst),
    .rsto(Tile_X3Y24_rsto),
    .FrameStrobe(Tile_X3_FrameStrobe),
    .FrameStrobe_O(Tile_X3Y24_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
S_term_custom Tile_X4Y24_S_term_custom (
    .from_SA(Tile_X4Y23_to_SA),
    .from_SB(Tile_X4Y23_to_SB),
    .from_SC(Tile_X4Y23_to_SC),
    .from_SD(Tile_X4Y23_to_SD),
    .from_SF(Tile_X4Y23_to_SF),
    .from_SG(Tile_X4Y23_to_SG),
    .from_SH(Tile_X4Y23_to_SH),
    .from_SI(Tile_X4Y23_to_SI),
    .to_NA(Tile_X4Y24_to_NA),
    .to_NB(Tile_X4Y24_to_NB),
    .to_NC(Tile_X4Y24_to_NC),
    .to_ND(Tile_X4Y24_to_ND),
    .to_NF(Tile_X4Y24_to_NF),
    .to_NG(Tile_X4Y24_to_NG),
    .to_NH(Tile_X4Y24_to_NH),
    .to_NI(Tile_X4Y24_to_NI),
    .UserCLK(UserCLK),
    .UserCLKo(Tile_X4Y24_UserCLKo),
    .rst(rst),
    .rsto(Tile_X4Y24_rsto),
    .FrameStrobe(Tile_X4_FrameStrobe),
    .FrameStrobe_O(Tile_X4Y24_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
S_term_custom Tile_X5Y24_S_term_custom (
    .from_SA(Tile_X5Y23_to_SA),
    .from_SB(Tile_X5Y23_to_SB),
    .from_SC(Tile_X5Y23_to_SC),
    .from_SD(Tile_X5Y23_to_SD),
    .from_SF(Tile_X5Y23_to_SF),
    .from_SG(Tile_X5Y23_to_SG),
    .from_SH(Tile_X5Y23_to_SH),
    .from_SI(Tile_X5Y23_to_SI),
    .to_NA(Tile_X5Y24_to_NA),
    .to_NB(Tile_X5Y24_to_NB),
    .to_NC(Tile_X5Y24_to_NC),
    .to_ND(Tile_X5Y24_to_ND),
    .to_NF(Tile_X5Y24_to_NF),
    .to_NG(Tile_X5Y24_to_NG),
    .to_NH(Tile_X5Y24_to_NH),
    .to_NI(Tile_X5Y24_to_NI),
    .UserCLK(UserCLK),
    .UserCLKo(Tile_X5Y24_UserCLKo),
    .rst(rst),
    .rsto(Tile_X5Y24_rsto),
    .FrameStrobe(Tile_X5_FrameStrobe),
    .FrameStrobe_O(Tile_X5Y24_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
S_term_custom Tile_X6Y24_S_term_custom (
    .from_SA(Tile_X6Y23_to_SA),
    .from_SB(Tile_X6Y23_to_SB),
    .from_SC(Tile_X6Y23_to_SC),
    .from_SD(Tile_X6Y23_to_SD),
    .from_SF(Tile_X6Y23_to_SF),
    .from_SG(Tile_X6Y23_to_SG),
    .from_SH(Tile_X6Y23_to_SH),
    .from_SI(Tile_X6Y23_to_SI),
    .to_NA(Tile_X6Y24_to_NA),
    .to_NB(Tile_X6Y24_to_NB),
    .to_NC(Tile_X6Y24_to_NC),
    .to_ND(Tile_X6Y24_to_ND),
    .to_NF(Tile_X6Y24_to_NF),
    .to_NG(Tile_X6Y24_to_NG),
    .to_NH(Tile_X6Y24_to_NH),
    .to_NI(Tile_X6Y24_to_NI),
    .UserCLK(UserCLK),
    .UserCLKo(Tile_X6Y24_UserCLKo),
    .rst(rst),
    .rsto(Tile_X6Y24_rsto),
    .FrameStrobe(Tile_X6_FrameStrobe),
    .FrameStrobe_O(Tile_X6Y24_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
S_term_custom Tile_X7Y24_S_term_custom (
    .from_SA(Tile_X7Y23_to_SA),
    .from_SB(Tile_X7Y23_to_SB),
    .from_SC(Tile_X7Y23_to_SC),
    .from_SD(Tile_X7Y23_to_SD),
    .from_SF(Tile_X7Y23_to_SF),
    .from_SG(Tile_X7Y23_to_SG),
    .from_SH(Tile_X7Y23_to_SH),
    .from_SI(Tile_X7Y23_to_SI),
    .to_NA(Tile_X7Y24_to_NA),
    .to_NB(Tile_X7Y24_to_NB),
    .to_NC(Tile_X7Y24_to_NC),
    .to_ND(Tile_X7Y24_to_ND),
    .to_NF(Tile_X7Y24_to_NF),
    .to_NG(Tile_X7Y24_to_NG),
    .to_NH(Tile_X7Y24_to_NH),
    .to_NI(Tile_X7Y24_to_NI),
    .UserCLK(UserCLK),
    .UserCLKo(Tile_X7Y24_UserCLKo),
    .rst(rst),
    .rsto(Tile_X7Y24_rsto),
    .FrameStrobe(Tile_X7_FrameStrobe),
    .FrameStrobe_O(Tile_X7Y24_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
S_term_custom Tile_X8Y24_S_term_custom (
    .from_SA(Tile_X8Y23_to_SA),
    .from_SB(Tile_X8Y23_to_SB),
    .from_SC(Tile_X8Y23_to_SC),
    .from_SD(Tile_X8Y23_to_SD),
    .from_SF(Tile_X8Y23_to_SF),
    .from_SG(Tile_X8Y23_to_SG),
    .from_SH(Tile_X8Y23_to_SH),
    .from_SI(Tile_X8Y23_to_SI),
    .to_NA(Tile_X8Y24_to_NA),
    .to_NB(Tile_X8Y24_to_NB),
    .to_NC(Tile_X8Y24_to_NC),
    .to_ND(Tile_X8Y24_to_ND),
    .to_NF(Tile_X8Y24_to_NF),
    .to_NG(Tile_X8Y24_to_NG),
    .to_NH(Tile_X8Y24_to_NH),
    .to_NI(Tile_X8Y24_to_NI),
    .UserCLK(UserCLK),
    .UserCLKo(Tile_X8Y24_UserCLKo),
    .rst(rst),
    .rsto(Tile_X8Y24_rsto),
    .FrameStrobe(Tile_X8_FrameStrobe),
    .FrameStrobe_O(Tile_X8Y24_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
S_term_s1 Tile_X9Y24_S_term_s1 (
    .from_SA_1s(Tile_X9Y23_to_SA_1s),
    .from_SB_1s(Tile_X9Y23_to_SB_1s),
    .from_SC_1s(Tile_X9Y23_to_SC_1s),
    .from_SD_1s(Tile_X9Y23_to_SD_1s),
    .from_SF_1s(Tile_X9Y23_to_SF_1s),
    .from_SG_1s(Tile_X9Y23_to_SG_1s),
    .from_SH_1s(Tile_X9Y23_to_SH_1s),
    .from_SI_1s(Tile_X9Y23_to_SI_1s),
    .to_NA_1s(Tile_X9Y24_to_NA_1s),
    .to_NB_1s(Tile_X9Y24_to_NB_1s),
    .to_NC_1s(Tile_X9Y24_to_NC_1s),
    .to_ND_1s(Tile_X9Y24_to_ND_1s),
    .to_NF_1s(Tile_X9Y24_to_NF_1s),
    .to_NG_1s(Tile_X9Y24_to_NG_1s),
    .to_NH_1s(Tile_X9Y24_to_NH_1s),
    .to_NI_1s(Tile_X9Y24_to_NI_1s),
    .UserCLK(UserCLK),
    .UserCLKo(Tile_X9Y24_UserCLKo),
    .rst(rst),
    .rsto(Tile_X9Y24_rsto),
    .FrameStrobe(Tile_X9_FrameStrobe),
    .FrameStrobe_O(Tile_X9Y24_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
S_term_s1 Tile_X10Y24_S_term_s1 (
    .to_NA_1s(Tile_X10Y24_to_NA_1s),
    .to_NB_1s(Tile_X10Y24_to_NB_1s),
    .to_NC_1s(Tile_X10Y24_to_NC_1s),
    .to_ND_1s(Tile_X10Y24_to_ND_1s),
    .to_NF_1s(Tile_X10Y24_to_NF_1s),
    .to_NG_1s(Tile_X10Y24_to_NG_1s),
    .to_NH_1s(Tile_X10Y24_to_NH_1s),
    .to_NI_1s(Tile_X10Y24_to_NI_1s),
    .UserCLK(UserCLK),
    .UserCLKo(Tile_X10Y24_UserCLKo),
    .rst(rst),
    .rsto(Tile_X10Y24_rsto),
    .FrameStrobe(Tile_X10_FrameStrobe),
    .FrameStrobe_O(Tile_X10Y24_FrameStrobe_O)
);

endmodule