--Template for state register with two shifting directions
-- MixColumns is included and requires 4 clock cycles, 1 for each column
-- S00 first, then S01
--    +---+  +---+  +---+  +---+
--  <-|S00|<-|S01|<-|S02|<-|S03|<-
--    +---+  +---+  +---+  +---+
--    +---+  +---+  +---+  +---+
--  <-|S10|<-|S11|<-|S12|<-|S13|<-
--    +---+  +---+  +---+  +---+
--    +---+  +---+  +---+  +---+
--  <-|S20|<-|S21|<-|S22|<-|S23|<-
--    +---+  +---+  +---+  +---+
--    +---+  +---+  +---+  +---+
--  <-|S30|<-|S31|<-|S32|<-|S33|<-
--    +---+  +---+  +---+  +---+
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity State is
	port(
		clk	: in std_logic;
		selSR: in std_logic;
		selMC: in std_logic;
		inputSer : in std_logic_vector(7 downto 0);
		nReset   : in std_logic;
		input: in std_logic_vector(7 downto 0);
		inMC: in std_logic_vector(31 downto 0);
		output: out std_logic_vector(7 downto 0);
		outMC: out std_logic_vector(31 downto 0)
		);

end entity State;


architecture dfl of State is

	signal inS00ser, inS01ser, inS02ser, inS03ser 	: std_logic_vector(7 downto 0);
	signal inS00par, inS01par, inS02par, inS03par 	: std_logic_vector(7 downto 0);
	signal inS10ser, inS11ser, inS12ser, inS13ser 	: std_logic_vector(7 downto 0);
	signal inS10par, inS11par, inS12par, inS13par 	: std_logic_vector(7 downto 0);
	signal inS20ser, inS21ser, inS22ser, inS23ser 	: std_logic_vector(7 downto 0);
	signal inS20par, inS21par, inS22par, inS23par 	: std_logic_vector(7 downto 0);
	signal inS30ser, inS31ser, inS32ser, inS33ser 	: std_logic_vector(7 downto 0);
	signal inS30par, inS31par, inS32par, inS33par 	: std_logic_vector(7 downto 0);
	
	signal outS00ser, outS01ser, outS02ser, outS03ser 	: std_logic_vector(7 downto 0);
	signal outS00par, outS01par, outS02par, outS03par 	: std_logic_vector(7 downto 0);
	signal outS10ser, outS11ser, outS12ser, outS13ser 	: std_logic_vector(7 downto 0);
	signal outS10par, outS11par, outS12par, outS13par 	: std_logic_vector(7 downto 0);
	signal outS20ser, outS21ser, outS22ser, outS23ser 	: std_logic_vector(7 downto 0);
	signal outS20par, outS21par, outS22par, outS23par 	: std_logic_vector(7 downto 0);
	signal outS30ser, outS31ser, outS32ser, outS33ser 	: std_logic_vector(7 downto 0);
	signal outS30par, outS31par, outS32par, outS33par 	: std_logic_vector(7 downto 0);

component reg is
	generic (NBITS_D0: integer;
		 NBITS_D1: integer);
	port(
		clk	: in std_logic;
		sel	: in std_logic;
		D0	: in std_logic_vector(NBITS_D0 - 1 downto 0);
		D1	: in std_logic_vector(NBITS_D1 - 1 downto 0);
		Q0	: out std_logic_vector(NBITS_D0 -1 downto 0);
		Q1	: out std_logic_vector(NBITS_D1 -1 downto 0)
		);
end component;

	signal outS10ser_MC, outS20ser_MC, outS30ser_MC, input_MC : std_logic_vector(7 downto 0);
	signal nReset_selMC : std_logic;

begin

-----------------------------------------------
--Row 0 
-----------------------------------------------
S00reg: reg
	generic map(NBITS_D0=>8,
				NBITS_D1=>8)
	port map(
		clk => clk,
		sel => selSR,
      	D0 => inS00ser,
  		D1 => inS00par,
      	Q0 => outS00ser,
      	Q1 => outS00par
		);
S01reg: reg
	generic map(NBITS_D0=>8,
				NBITS_D1=>8)
	port map(
		clk => clk,
		sel => selSR,
      	D0 => inS01ser,
		D1 => inS01par,
      	Q0 => outS01ser,
      	Q1 => outS01par
		);
S02reg: reg
	generic map(NBITS_D0=>8,
				NBITS_D1=>8)
	port map(
		clk => clk,
		sel => selSR,
      	D0 => inS02ser,
  		D1 => inS02par,
      	Q0 => outS02ser,
      	Q1 => outS02par
		);
S03reg: reg
	generic map(NBITS_D0=>8,
				NBITS_D1=>8)
	port map(
		clk => clk,
		sel => selSR,
      	D0 => inS03ser,
  		D1 => inS03par,
      	Q0 => outS03ser,
      	Q1 => outS03par
		);
-----------------------------------------------
--Row 1
-----------------------------------------------
S10reg: reg
	generic map(NBITS_D0=>8,
				NBITS_D1=>8)
	port map(
		clk => clk,
		sel => selSR,
      	D0 => inS10ser,
  		D1 => inS10par,
      	Q0 => outS10ser,
      	Q1 => outS10par
		);
S11reg: reg
	generic map(NBITS_D0=>8,
				NBITS_D1=>8)
	port map(
		clk => clk,
		sel => selSR,
      	D0 => inS11ser,
  		D1 => inS11par,
      	Q0 => outS11ser,
      	Q1 => outS11par
		);
S12reg: reg
	generic map(NBITS_D0=>8,
				NBITS_D1=>8)
	port map(
		clk => clk,
		sel => selSR,
      	D0 => inS12ser,
  		D1 => inS12par,
      	Q0 => outS12ser,
      	Q1 => outS12par
		);
S13reg: reg
	generic map(NBITS_D0=>8,
				NBITS_D1=>8)
	port map(
		clk => clk,
		sel => selSR,
      	D0 => inS13ser,
  		D1 => inS13par,
      	Q0 => outS13ser,
      	Q1 => outS13par
		);
-----------------------------------------------
--Row 2
-----------------------------------------------
S20reg: reg
	generic map(NBITS_D0=>8,
				NBITS_D1=>8)
	port map(
		clk => clk,
		sel => selSR,
      	D0 => inS20ser,
  		D1 => inS20par,
      	Q0 => outS20ser,
      	Q1 => outS20par
		);
S21reg: reg
	generic map(NBITS_D0=>8,
				NBITS_D1=>8)
	port map(
		clk => clk,
		sel => selSR,
      	D0 => inS21ser,
  		D1 => inS21par,
      	Q0 => outS21ser,
      	Q1 => outS21par
		);
S22reg: reg
	generic map(NBITS_D0=>8,
				NBITS_D1=>8)
	port map(
		clk => clk,
		sel => selSR,
      	D0 => inS22ser,
  		D1 => inS22par,
      	Q0 => outS22ser,
      	Q1 => outS22par
		);
S23reg: reg
	generic map(NBITS_D0=>8,
				NBITS_D1=>8)
	port map(
		clk => clk,
		sel => selSR,
      	D0 => inS23ser,
  		D1 => inS23par,
      	Q0 => outS23ser,
      	Q1 => outS23par
		);
-----------------------------------------------
--Row 3
-----------------------------------------------
S30reg: reg
	generic map(NBITS_D0=>8,
				NBITS_D1=>8)
	port map(
		clk => clk,
		sel => selSR,
      	D0 => inS30ser,
  		D1 => inS30par,
      	Q0 => outS30ser,
      	Q1 => outS30par
		);
S31reg: reg
	generic map(NBITS_D0=>8,
				NBITS_D1=>8)
	port map(
		clk => clk,
		sel => selSR,
      	D0 => inS31ser,
  		D1 => inS31par,
      	Q0 => outS31ser,
      	Q1 => outS31par
		);
S32reg: reg
	generic map(NBITS_D0=>8,
				NBITS_D1=>8)
	port map(
		clk => clk,
		sel => selSR,
      	D0 => inS32ser,
  		D1 => inS32par,
      	Q0 => outS32ser,
      	Q1 => outS32par
		);
S33reg: reg
	generic map(NBITS_D0=>8,
				NBITS_D1=>8)
	port map(
		clk => clk,
		sel => selSR,
      	D0 => inS33ser,
  		D1 => inS33par,
      	Q0 => outS33ser,
      	Q1 => outS33par
		);

-----------------------------------------------
--8-bit horizontal Wiring, 1 MUX per Row for MC
-----------------------------------------------
--Row 0 
-----------------------------------------------

nReset_selMC <= nReset and selMC;

inS00ser <= outS01ser;
inS01ser <= outS02ser;
inS02ser <= outS03ser;
MUX_inS03ser:  ENTITY work.MUX Generic Map (size => 8) Port Map (S => nReset_selMC, D0 => outS10ser, D1 => inMC(31 downto 24), Q => inS03ser);

-----------------------------------------------
--Row 1
-----------------------------------------------

inS10ser <= outS11ser;
inS11ser <= outS12ser;
inS12ser <= outS13ser;
MUX_inS13ser:  ENTITY work.MUX Generic Map (size => 8) Port Map (S => nReset_selMC, D0 => outS20ser, D1 => inMC(23 downto 16), Q => inS13ser);

-----------------------------------------------
--Row 2
-----------------------------------------------

inS20ser <= outS21ser;
inS21ser <= outS22ser;
inS22ser <= outS23ser;

MUX_inS23ser:  ENTITY work.MUX Generic Map (size => 8) Port Map (S => nReset_selMC, D0 => outS30ser, D1 => inMC(15 downto  8), Q => inS23ser);

-----------------------------------------------
--Row 3 
-----------------------------------------------

inS30ser <= outS31ser;
inS31ser <= outS32ser;
inS32ser <= outS33ser;

MUX_input_MC:  ENTITY work.MUX Generic Map (size => 8) Port Map (S => selMC,  D0 => input,    D1 => inMC(7  downto  0), Q => input_MC);
MUX_inS33ser:  ENTITY work.MUX Generic Map (size => 8) Port Map (S => nReset, D0 => inputSer, D1 => input_MC,           Q => inS33ser);

-----------------------------------------------
--8-bit vertical Wiring
-----------------------------------------------
--Row 0 no shifting
-----------------------------------------------
inS00par <= outS00par;
inS01par <= outS01par;
inS02par <= outS02par;
inS03par <= outS03par;
-----------------------------------------------
--Row 1 left shift by 1 
-----------------------------------------------
inS10par <= outS11par;
inS11par <= outS12par;
inS12par <= outS13par;
inS13par <= outS10par;
-----------------------------------------------
--Row 2 left shift by 2 
-----------------------------------------------
inS20par <= outS22par;
inS21par <= outS23par;
inS22par <= outS20par;
inS23par <= outS21par;
-----------------------------------------------
--Row 3 left shift by 3 
-----------------------------------------------
inS30par <= outS33par;
inS31par <= outS30par;
inS32par <= outS31par;
inS33par <= outS32par;

-----------------------------------------------
--output Wiring 
-----------------------------------------------
outMC <= outS00ser&outS10ser&outS20ser&outS30ser;

output <= outS00ser;

end architecture;
