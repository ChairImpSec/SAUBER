//-----------------------------------------

module top(input wire [22:0] io_in_0t, io_in_0f, io_in_1t, io_in_1f, ctrl_io_in_0t, ctrl_io_in_0f,  output wire [22:0] io_out_0t, io_out_0f, io_out_1t, io_out_1f, io_oeb, ctrl_io_out_0t, ctrl_io_out_0f, ctrl_io_oeb);

    main_SAUBER_Pipeline_d1 generated_module (
        .value_in(io_in_0t[7:0]),

        .start(ctrl_io_in_0t[3:0]),
        .rst(ctrl_io_in_0t[4]),
        .value_out(io_out_0t[19:12]),

    );

//-----------

    assign io_oeb      = 60'b11111111000000000000;
    assign ctrl_io_oeb = 60'b0;

endmodule

module main_SAUBER_Pipeline_d1 (value_in, start, rst, value_out);
    input [7:0] value_in ;
    input [3:0] start ;
    input rst ;
    output [7:0] value_out ;
    wire n9 ;
    wire n10 ;
    wire [3:3] Inc_out ;
    wire [7:0] Sbox_in ;
    wire [3:0] Inc_Reg ;
    wire [3:0] Inc_in ;
    wire \M1.gen_loop_0__M.X ;
    wire \M1.gen_loop_0__M.Y ;
    wire \M1.gen_loop_1__M.X ;
    wire \M1.gen_loop_1__M.Y ;
    wire \M1.gen_loop_2__M.X ;
    wire \M1.gen_loop_2__M.Y ;
    wire \M1.gen_loop_3__M.X ;
    wire \M1.gen_loop_3__M.Y ;
    wire \M1.gen_loop_4__M.X ;
    wire \M1.gen_loop_4__M.Y ;
    wire \M1.gen_loop_5__M.X ;
    wire \M1.gen_loop_5__M.Y ;
    wire \M1.gen_loop_6__M.X ;
    wire \M1.gen_loop_6__M.Y ;
    wire \M1.gen_loop_7__M.X ;
    wire \M1.gen_loop_7__M.Y ;
    wire \SboxInst.T1 ;
    wire \SboxInst.T2 ;
    wire \SboxInst.T3 ;
    wire \SboxInst.T4 ;
    wire \SboxInst.T5 ;
    wire \SboxInst.T6 ;
    wire \SboxInst.T7 ;
    wire \SboxInst.T8 ;
    wire \SboxInst.T9 ;
    wire \SboxInst.T10 ;
    wire \SboxInst.T11 ;
    wire \SboxInst.T12 ;
    wire \SboxInst.T13 ;
    wire \SboxInst.T14 ;
    wire \SboxInst.T15 ;
    wire \SboxInst.T16 ;
    wire \SboxInst.T17 ;
    wire \SboxInst.T18 ;
    wire \SboxInst.T19 ;
    wire \SboxInst.T20 ;
    wire \SboxInst.T21 ;
    wire \SboxInst.T22 ;
    wire \SboxInst.T23 ;
    wire \SboxInst.T24 ;
    wire \SboxInst.T25 ;
    wire \SboxInst.T26 ;
    wire \SboxInst.T27 ;
    wire \SboxInst.M1 ;
    wire \SboxInst.M2 ;
    wire \SboxInst.M3 ;
    wire \SboxInst.M4 ;
    wire \SboxInst.M5 ;
    wire \SboxInst.M6 ;
    wire \SboxInst.M7 ;
    wire \SboxInst.M8 ;
    wire \SboxInst.M9 ;
    wire \SboxInst.M10 ;
    wire \SboxInst.M11 ;
    wire \SboxInst.M12 ;
    wire \SboxInst.M13 ;
    wire \SboxInst.M14 ;
    wire \SboxInst.M15 ;
    wire \SboxInst.M16 ;
    wire \SboxInst.M17 ;
    wire \SboxInst.M18 ;
    wire \SboxInst.M19 ;
    wire \SboxInst.M20 ;
    wire \SboxInst.M21 ;
    wire \SboxInst.M22 ;
    wire \SboxInst.M23 ;
    wire \SboxInst.M24 ;
    wire \SboxInst.M25 ;
    wire \SboxInst.M26 ;
    wire \SboxInst.M27 ;
    wire \SboxInst.M28 ;
    wire \SboxInst.M29 ;
    wire \SboxInst.M30 ;
    wire \SboxInst.M31 ;
    wire \SboxInst.M32 ;
    wire \SboxInst.M33 ;
    wire \SboxInst.M34 ;
    wire \SboxInst.M35 ;
    wire \SboxInst.M36 ;
    wire \SboxInst.M37 ;
    wire \SboxInst.M38 ;
    wire \SboxInst.M39 ;
    wire \SboxInst.M40 ;
    wire \SboxInst.M41 ;
    wire \SboxInst.M42 ;
    wire \SboxInst.M43 ;
    wire \SboxInst.M44 ;
    wire \SboxInst.M45 ;
    wire \SboxInst.M46 ;
    wire \SboxInst.M47 ;
    wire \SboxInst.M48 ;
    wire \SboxInst.M49 ;
    wire \SboxInst.M50 ;
    wire \SboxInst.M51 ;
    wire \SboxInst.M52 ;
    wire \SboxInst.M53 ;
    wire \SboxInst.M54 ;
    wire \SboxInst.M55 ;
    wire \SboxInst.M56 ;
    wire \SboxInst.M57 ;
    wire \SboxInst.M58 ;
    wire \SboxInst.M59 ;
    wire \SboxInst.M60 ;
    wire \SboxInst.M61 ;
    wire \SboxInst.M62 ;
    wire \SboxInst.M63 ;
    wire \SboxInst.L0 ;
    wire \SboxInst.L1 ;
    wire \SboxInst.L2 ;
    wire \SboxInst.L3 ;
    wire \SboxInst.L4 ;
    wire \SboxInst.L5 ;
    wire \SboxInst.L6 ;
    wire \SboxInst.L7 ;
    wire \SboxInst.L8 ;
    wire \SboxInst.L9 ;
    wire \SboxInst.L10 ;
    wire \SboxInst.L11 ;
    wire \SboxInst.L12 ;
    wire \SboxInst.L13 ;
    wire \SboxInst.L14 ;
    wire \SboxInst.L15 ;
    wire \SboxInst.L16 ;
    wire \SboxInst.L17 ;
    wire \SboxInst.L18 ;
    wire \SboxInst.L19 ;
    wire \SboxInst.L20 ;
    wire \SboxInst.L21 ;
    wire \SboxInst.L22 ;
    wire \SboxInst.L23 ;
    wire \SboxInst.L24 ;
    wire \SboxInst.L25 ;
    wire \SboxInst.L26 ;
    wire \SboxInst.L27 ;
    wire \SboxInst.L28 ;
    wire \SboxInst.L29 ;
    wire \M2.gen_loop_0__M.X ;
    wire \M2.gen_loop_0__M.Y ;
    wire \M2.gen_loop_1__M.X ;
    wire \M2.gen_loop_1__M.Y ;
    wire \M2.gen_loop_2__M.X ;
    wire \M2.gen_loop_2__M.Y ;
    wire \M2.gen_loop_3__M.X ;
    wire \M2.gen_loop_3__M.Y ;

    /* cells in depth 0 */
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \M1.gen_loop_0__M.X1.U1 ( .A0_t (value_in[0]), .B0_t (value_out[0]), .Z0_t (\M1.gen_loop_0__M.X ) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \M1.gen_loop_0__M.A.U1 ( .A0_t (Inc_out[3]), .B0_t (\M1.gen_loop_0__M.X ), .Z0_t (\M1.gen_loop_0__M.Y ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \M1.gen_loop_0__M.X2.U1 ( .A0_t (\M1.gen_loop_0__M.Y ), .B0_t (value_in[0]), .Z0_t (Sbox_in[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \M1.gen_loop_1__M.X1.U1 ( .A0_t (value_in[1]), .B0_t (value_out[1]), .Z0_t (\M1.gen_loop_1__M.X ) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \M1.gen_loop_1__M.A.U1 ( .A0_t (Inc_out[3]), .B0_t (\M1.gen_loop_1__M.X ), .Z0_t (\M1.gen_loop_1__M.Y ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \M1.gen_loop_1__M.X2.U1 ( .A0_t (\M1.gen_loop_1__M.Y ), .B0_t (value_in[1]), .Z0_t (Sbox_in[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \M1.gen_loop_2__M.X1.U1 ( .A0_t (value_in[2]), .B0_t (value_out[2]), .Z0_t (\M1.gen_loop_2__M.X ) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \M1.gen_loop_2__M.A.U1 ( .A0_t (Inc_out[3]), .B0_t (\M1.gen_loop_2__M.X ), .Z0_t (\M1.gen_loop_2__M.Y ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \M1.gen_loop_2__M.X2.U1 ( .A0_t (\M1.gen_loop_2__M.Y ), .B0_t (value_in[2]), .Z0_t (Sbox_in[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \M1.gen_loop_3__M.X1.U1 ( .A0_t (value_in[3]), .B0_t (value_out[3]), .Z0_t (\M1.gen_loop_3__M.X ) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \M1.gen_loop_3__M.A.U1 ( .A0_t (Inc_out[3]), .B0_t (\M1.gen_loop_3__M.X ), .Z0_t (\M1.gen_loop_3__M.Y ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \M1.gen_loop_3__M.X2.U1 ( .A0_t (\M1.gen_loop_3__M.Y ), .B0_t (value_in[3]), .Z0_t (Sbox_in[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \M1.gen_loop_4__M.X1.U1 ( .A0_t (value_in[4]), .B0_t (value_out[4]), .Z0_t (\M1.gen_loop_4__M.X ) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \M1.gen_loop_4__M.A.U1 ( .A0_t (Inc_out[3]), .B0_t (\M1.gen_loop_4__M.X ), .Z0_t (\M1.gen_loop_4__M.Y ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \M1.gen_loop_4__M.X2.U1 ( .A0_t (\M1.gen_loop_4__M.Y ), .B0_t (value_in[4]), .Z0_t (Sbox_in[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \M1.gen_loop_5__M.X1.U1 ( .A0_t (value_in[5]), .B0_t (value_out[5]), .Z0_t (\M1.gen_loop_5__M.X ) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \M1.gen_loop_5__M.A.U1 ( .A0_t (Inc_out[3]), .B0_t (\M1.gen_loop_5__M.X ), .Z0_t (\M1.gen_loop_5__M.Y ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \M1.gen_loop_5__M.X2.U1 ( .A0_t (\M1.gen_loop_5__M.Y ), .B0_t (value_in[5]), .Z0_t (Sbox_in[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \M1.gen_loop_6__M.X1.U1 ( .A0_t (value_in[6]), .B0_t (value_out[6]), .Z0_t (\M1.gen_loop_6__M.X ) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \M1.gen_loop_6__M.A.U1 ( .A0_t (Inc_out[3]), .B0_t (\M1.gen_loop_6__M.X ), .Z0_t (\M1.gen_loop_6__M.Y ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \M1.gen_loop_6__M.X2.U1 ( .A0_t (\M1.gen_loop_6__M.Y ), .B0_t (value_in[6]), .Z0_t (Sbox_in[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \M1.gen_loop_7__M.X1.U1 ( .A0_t (value_in[7]), .B0_t (value_out[7]), .Z0_t (\M1.gen_loop_7__M.X ) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \M1.gen_loop_7__M.A.U1 ( .A0_t (Inc_out[3]), .B0_t (\M1.gen_loop_7__M.X ), .Z0_t (\M1.gen_loop_7__M.Y ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \M1.gen_loop_7__M.X2.U1 ( .A0_t (\M1.gen_loop_7__M.Y ), .B0_t (value_in[7]), .Z0_t (Sbox_in[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_T1.U1 ( .A0_t (Sbox_in[7]), .B0_t (Sbox_in[4]), .Z0_t (\SboxInst.T1 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_T2.U1 ( .A0_t (Sbox_in[7]), .B0_t (Sbox_in[2]), .Z0_t (\SboxInst.T2 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_T3.U1 ( .A0_t (Sbox_in[7]), .B0_t (Sbox_in[1]), .Z0_t (\SboxInst.T3 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_T4.U1 ( .A0_t (Sbox_in[4]), .B0_t (Sbox_in[2]), .Z0_t (\SboxInst.T4 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_T5.U1 ( .A0_t (Sbox_in[3]), .B0_t (Sbox_in[1]), .Z0_t (\SboxInst.T5 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_T6.U1 ( .A0_t (\SboxInst.T1 ), .B0_t (\SboxInst.T5 ), .Z0_t (\SboxInst.T6 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_T7.U1 ( .A0_t (Sbox_in[6]), .B0_t (Sbox_in[5]), .Z0_t (\SboxInst.T7 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_T8.U1 ( .A0_t (Sbox_in[0]), .B0_t (\SboxInst.T6 ), .Z0_t (\SboxInst.T8 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_T9.U1 ( .A0_t (Sbox_in[0]), .B0_t (\SboxInst.T7 ), .Z0_t (\SboxInst.T9 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_T10.U1 ( .A0_t (\SboxInst.T6 ), .B0_t (\SboxInst.T7 ), .Z0_t (\SboxInst.T10 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_T11.U1 ( .A0_t (Sbox_in[6]), .B0_t (Sbox_in[2]), .Z0_t (\SboxInst.T11 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_T12.U1 ( .A0_t (Sbox_in[5]), .B0_t (Sbox_in[2]), .Z0_t (\SboxInst.T12 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_T13.U1 ( .A0_t (\SboxInst.T3 ), .B0_t (\SboxInst.T4 ), .Z0_t (\SboxInst.T13 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_T14.U1 ( .A0_t (\SboxInst.T6 ), .B0_t (\SboxInst.T11 ), .Z0_t (\SboxInst.T14 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_T15.U1 ( .A0_t (\SboxInst.T5 ), .B0_t (\SboxInst.T11 ), .Z0_t (\SboxInst.T15 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_T16.U1 ( .A0_t (\SboxInst.T5 ), .B0_t (\SboxInst.T12 ), .Z0_t (\SboxInst.T16 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_T17.U1 ( .A0_t (\SboxInst.T9 ), .B0_t (\SboxInst.T16 ), .Z0_t (\SboxInst.T17 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_T18.U1 ( .A0_t (Sbox_in[4]), .B0_t (Sbox_in[0]), .Z0_t (\SboxInst.T18 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_T19.U1 ( .A0_t (\SboxInst.T7 ), .B0_t (\SboxInst.T18 ), .Z0_t (\SboxInst.T19 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_T20.U1 ( .A0_t (\SboxInst.T1 ), .B0_t (\SboxInst.T19 ), .Z0_t (\SboxInst.T20 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_T21.U1 ( .A0_t (Sbox_in[1]), .B0_t (Sbox_in[0]), .Z0_t (\SboxInst.T21 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_T22.U1 ( .A0_t (\SboxInst.T7 ), .B0_t (\SboxInst.T21 ), .Z0_t (\SboxInst.T22 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_T23.U1 ( .A0_t (\SboxInst.T2 ), .B0_t (\SboxInst.T22 ), .Z0_t (\SboxInst.T23 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_T24.U1 ( .A0_t (\SboxInst.T2 ), .B0_t (\SboxInst.T10 ), .Z0_t (\SboxInst.T24 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_T25.U1 ( .A0_t (\SboxInst.T20 ), .B0_t (\SboxInst.T17 ), .Z0_t (\SboxInst.T25 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_T26.U1 ( .A0_t (\SboxInst.T3 ), .B0_t (\SboxInst.T16 ), .Z0_t (\SboxInst.T26 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_T27.U1 ( .A0_t (\SboxInst.T1 ), .B0_t (\SboxInst.T12 ), .Z0_t (\SboxInst.T27 ) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M1.U1 ( .A0_t (\SboxInst.T13 ), .B0_t (\SboxInst.T6 ), .Z0_t (\SboxInst.M1 ) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M2.U1 ( .A0_t (\SboxInst.T23 ), .B0_t (\SboxInst.T8 ), .Z0_t (\SboxInst.M2 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_M3.U1 ( .A0_t (\SboxInst.T14 ), .B0_t (\SboxInst.M1 ), .Z0_t (\SboxInst.M3 ) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M4.U1 ( .A0_t (\SboxInst.T19 ), .B0_t (Sbox_in[0]), .Z0_t (\SboxInst.M4 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_M5.U1 ( .A0_t (\SboxInst.M4 ), .B0_t (\SboxInst.M1 ), .Z0_t (\SboxInst.M5 ) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M6.U1 ( .A0_t (\SboxInst.T3 ), .B0_t (\SboxInst.T16 ), .Z0_t (\SboxInst.M6 ) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M7.U1 ( .A0_t (\SboxInst.T22 ), .B0_t (\SboxInst.T9 ), .Z0_t (\SboxInst.M7 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_M8.U1 ( .A0_t (\SboxInst.T26 ), .B0_t (\SboxInst.M6 ), .Z0_t (\SboxInst.M8 ) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M9.U1 ( .A0_t (\SboxInst.T20 ), .B0_t (\SboxInst.T17 ), .Z0_t (\SboxInst.M9 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_M10.U1 ( .A0_t (\SboxInst.M9 ), .B0_t (\SboxInst.M6 ), .Z0_t (\SboxInst.M10 ) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M11.U1 ( .A0_t (\SboxInst.T1 ), .B0_t (\SboxInst.T15 ), .Z0_t (\SboxInst.M11 ) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M12.U1 ( .A0_t (\SboxInst.T4 ), .B0_t (\SboxInst.T27 ), .Z0_t (\SboxInst.M12 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_M13.U1 ( .A0_t (\SboxInst.M12 ), .B0_t (\SboxInst.M11 ), .Z0_t (\SboxInst.M13 ) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M14.U1 ( .A0_t (\SboxInst.T2 ), .B0_t (\SboxInst.T10 ), .Z0_t (\SboxInst.M14 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_M15.U1 ( .A0_t (\SboxInst.M14 ), .B0_t (\SboxInst.M11 ), .Z0_t (\SboxInst.M15 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_M16.U1 ( .A0_t (\SboxInst.M3 ), .B0_t (\SboxInst.M2 ), .Z0_t (\SboxInst.M16 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_M17.U1 ( .A0_t (\SboxInst.M5 ), .B0_t (\SboxInst.T24 ), .Z0_t (\SboxInst.M17 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_M18.U1 ( .A0_t (\SboxInst.M8 ), .B0_t (\SboxInst.M7 ), .Z0_t (\SboxInst.M18 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_M19.U1 ( .A0_t (\SboxInst.M10 ), .B0_t (\SboxInst.M15 ), .Z0_t (\SboxInst.M19 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_M20.U1 ( .A0_t (\SboxInst.M16 ), .B0_t (\SboxInst.M13 ), .Z0_t (\SboxInst.M20 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_M21.U1 ( .A0_t (\SboxInst.M17 ), .B0_t (\SboxInst.M15 ), .Z0_t (\SboxInst.M21 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_M22.U1 ( .A0_t (\SboxInst.M18 ), .B0_t (\SboxInst.M13 ), .Z0_t (\SboxInst.M22 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_M23.U1 ( .A0_t (\SboxInst.M19 ), .B0_t (\SboxInst.T25 ), .Z0_t (\SboxInst.M23 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_M24.U1 ( .A0_t (\SboxInst.M22 ), .B0_t (\SboxInst.M23 ), .Z0_t (\SboxInst.M24 ) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M25.U1 ( .A0_t (\SboxInst.M22 ), .B0_t (\SboxInst.M20 ), .Z0_t (\SboxInst.M25 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_M26.U1 ( .A0_t (\SboxInst.M21 ), .B0_t (\SboxInst.M25 ), .Z0_t (\SboxInst.M26 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_M27.U1 ( .A0_t (\SboxInst.M20 ), .B0_t (\SboxInst.M21 ), .Z0_t (\SboxInst.M27 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_M28.U1 ( .A0_t (\SboxInst.M23 ), .B0_t (\SboxInst.M25 ), .Z0_t (\SboxInst.M28 ) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M29.U1 ( .A0_t (\SboxInst.M28 ), .B0_t (\SboxInst.M27 ), .Z0_t (\SboxInst.M29 ) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M30.U1 ( .A0_t (\SboxInst.M26 ), .B0_t (\SboxInst.M24 ), .Z0_t (\SboxInst.M30 ) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M31.U1 ( .A0_t (\SboxInst.M20 ), .B0_t (\SboxInst.M23 ), .Z0_t (\SboxInst.M31 ) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M32.U1 ( .A0_t (\SboxInst.M27 ), .B0_t (\SboxInst.M31 ), .Z0_t (\SboxInst.M32 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_M33.U1 ( .A0_t (\SboxInst.M27 ), .B0_t (\SboxInst.M25 ), .Z0_t (\SboxInst.M33 ) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M34.U1 ( .A0_t (\SboxInst.M21 ), .B0_t (\SboxInst.M22 ), .Z0_t (\SboxInst.M34 ) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M35.U1 ( .A0_t (\SboxInst.M24 ), .B0_t (\SboxInst.M34 ), .Z0_t (\SboxInst.M35 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_M36.U1 ( .A0_t (\SboxInst.M24 ), .B0_t (\SboxInst.M25 ), .Z0_t (\SboxInst.M36 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_M37.U1 ( .A0_t (\SboxInst.M21 ), .B0_t (\SboxInst.M29 ), .Z0_t (\SboxInst.M37 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_M38.U1 ( .A0_t (\SboxInst.M32 ), .B0_t (\SboxInst.M33 ), .Z0_t (\SboxInst.M38 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_M39.U1 ( .A0_t (\SboxInst.M23 ), .B0_t (\SboxInst.M30 ), .Z0_t (\SboxInst.M39 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_M40.U1 ( .A0_t (\SboxInst.M35 ), .B0_t (\SboxInst.M36 ), .Z0_t (\SboxInst.M40 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_M41.U1 ( .A0_t (\SboxInst.M38 ), .B0_t (\SboxInst.M40 ), .Z0_t (\SboxInst.M41 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_M42.U1 ( .A0_t (\SboxInst.M37 ), .B0_t (\SboxInst.M39 ), .Z0_t (\SboxInst.M42 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_M43.U1 ( .A0_t (\SboxInst.M37 ), .B0_t (\SboxInst.M38 ), .Z0_t (\SboxInst.M43 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_M44.U1 ( .A0_t (\SboxInst.M39 ), .B0_t (\SboxInst.M40 ), .Z0_t (\SboxInst.M44 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_M45.U1 ( .A0_t (\SboxInst.M42 ), .B0_t (\SboxInst.M41 ), .Z0_t (\SboxInst.M45 ) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M46.U1 ( .A0_t (\SboxInst.M44 ), .B0_t (\SboxInst.T6 ), .Z0_t (\SboxInst.M46 ) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M47.U1 ( .A0_t (\SboxInst.M40 ), .B0_t (\SboxInst.T8 ), .Z0_t (\SboxInst.M47 ) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M48.U1 ( .A0_t (\SboxInst.M39 ), .B0_t (Sbox_in[0]), .Z0_t (\SboxInst.M48 ) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M49.U1 ( .A0_t (\SboxInst.M43 ), .B0_t (\SboxInst.T16 ), .Z0_t (\SboxInst.M49 ) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M50.U1 ( .A0_t (\SboxInst.M38 ), .B0_t (\SboxInst.T9 ), .Z0_t (\SboxInst.M50 ) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M51.U1 ( .A0_t (\SboxInst.M37 ), .B0_t (\SboxInst.T17 ), .Z0_t (\SboxInst.M51 ) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M52.U1 ( .A0_t (\SboxInst.M42 ), .B0_t (\SboxInst.T15 ), .Z0_t (\SboxInst.M52 ) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M53.U1 ( .A0_t (\SboxInst.M45 ), .B0_t (\SboxInst.T27 ), .Z0_t (\SboxInst.M53 ) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M54.U1 ( .A0_t (\SboxInst.M41 ), .B0_t (\SboxInst.T10 ), .Z0_t (\SboxInst.M54 ) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M55.U1 ( .A0_t (\SboxInst.M44 ), .B0_t (\SboxInst.T13 ), .Z0_t (\SboxInst.M55 ) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M56.U1 ( .A0_t (\SboxInst.M40 ), .B0_t (\SboxInst.T23 ), .Z0_t (\SboxInst.M56 ) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M57.U1 ( .A0_t (\SboxInst.M39 ), .B0_t (\SboxInst.T19 ), .Z0_t (\SboxInst.M57 ) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M58.U1 ( .A0_t (\SboxInst.M43 ), .B0_t (\SboxInst.T3 ), .Z0_t (\SboxInst.M58 ) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M59.U1 ( .A0_t (\SboxInst.M38 ), .B0_t (\SboxInst.T22 ), .Z0_t (\SboxInst.M59 ) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M60.U1 ( .A0_t (\SboxInst.M37 ), .B0_t (\SboxInst.T20 ), .Z0_t (\SboxInst.M60 ) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M61.U1 ( .A0_t (\SboxInst.M42 ), .B0_t (\SboxInst.T1 ), .Z0_t (\SboxInst.M61 ) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M62.U1 ( .A0_t (\SboxInst.M45 ), .B0_t (\SboxInst.T4 ), .Z0_t (\SboxInst.M62 ) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.AND_M63.U1 ( .A0_t (\SboxInst.M41 ), .B0_t (\SboxInst.T2 ), .Z0_t (\SboxInst.M63 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_L0.U1 ( .A0_t (\SboxInst.M61 ), .B0_t (\SboxInst.M62 ), .Z0_t (\SboxInst.L0 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_L1.U1 ( .A0_t (\SboxInst.M50 ), .B0_t (\SboxInst.M56 ), .Z0_t (\SboxInst.L1 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_L2.U1 ( .A0_t (\SboxInst.M46 ), .B0_t (\SboxInst.M48 ), .Z0_t (\SboxInst.L2 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_L3.U1 ( .A0_t (\SboxInst.M47 ), .B0_t (\SboxInst.M55 ), .Z0_t (\SboxInst.L3 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_L4.U1 ( .A0_t (\SboxInst.M54 ), .B0_t (\SboxInst.M58 ), .Z0_t (\SboxInst.L4 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_L5.U1 ( .A0_t (\SboxInst.M49 ), .B0_t (\SboxInst.M61 ), .Z0_t (\SboxInst.L5 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_L6.U1 ( .A0_t (\SboxInst.M62 ), .B0_t (\SboxInst.L5 ), .Z0_t (\SboxInst.L6 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_L7.U1 ( .A0_t (\SboxInst.M46 ), .B0_t (\SboxInst.L3 ), .Z0_t (\SboxInst.L7 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_L8.U1 ( .A0_t (\SboxInst.M51 ), .B0_t (\SboxInst.M59 ), .Z0_t (\SboxInst.L8 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_L9.U1 ( .A0_t (\SboxInst.M52 ), .B0_t (\SboxInst.M53 ), .Z0_t (\SboxInst.L9 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_L10.U1 ( .A0_t (\SboxInst.M53 ), .B0_t (\SboxInst.L4 ), .Z0_t (\SboxInst.L10 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_L11.U1 ( .A0_t (\SboxInst.M60 ), .B0_t (\SboxInst.L2 ), .Z0_t (\SboxInst.L11 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_L12.U1 ( .A0_t (\SboxInst.M48 ), .B0_t (\SboxInst.M51 ), .Z0_t (\SboxInst.L12 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_L13.U1 ( .A0_t (\SboxInst.M50 ), .B0_t (\SboxInst.L0 ), .Z0_t (\SboxInst.L13 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_L14.U1 ( .A0_t (\SboxInst.M52 ), .B0_t (\SboxInst.M61 ), .Z0_t (\SboxInst.L14 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_L15.U1 ( .A0_t (\SboxInst.M55 ), .B0_t (\SboxInst.L1 ), .Z0_t (\SboxInst.L15 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_L16.U1 ( .A0_t (\SboxInst.M56 ), .B0_t (\SboxInst.L0 ), .Z0_t (\SboxInst.L16 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_L17.U1 ( .A0_t (\SboxInst.M57 ), .B0_t (\SboxInst.L1 ), .Z0_t (\SboxInst.L17 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_L18.U1 ( .A0_t (\SboxInst.M58 ), .B0_t (\SboxInst.L8 ), .Z0_t (\SboxInst.L18 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_L19.U1 ( .A0_t (\SboxInst.M63 ), .B0_t (\SboxInst.L4 ), .Z0_t (\SboxInst.L19 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_L20.U1 ( .A0_t (\SboxInst.L0 ), .B0_t (\SboxInst.L1 ), .Z0_t (\SboxInst.L20 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_L21.U1 ( .A0_t (\SboxInst.L1 ), .B0_t (\SboxInst.L7 ), .Z0_t (\SboxInst.L21 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_L22.U1 ( .A0_t (\SboxInst.L3 ), .B0_t (\SboxInst.L12 ), .Z0_t (\SboxInst.L22 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_L23.U1 ( .A0_t (\SboxInst.L18 ), .B0_t (\SboxInst.L2 ), .Z0_t (\SboxInst.L23 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_L24.U1 ( .A0_t (\SboxInst.L15 ), .B0_t (\SboxInst.L9 ), .Z0_t (\SboxInst.L24 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_L25.U1 ( .A0_t (\SboxInst.L6 ), .B0_t (\SboxInst.L10 ), .Z0_t (\SboxInst.L25 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_L26.U1 ( .A0_t (\SboxInst.L7 ), .B0_t (\SboxInst.L9 ), .Z0_t (\SboxInst.L26 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_L27.U1 ( .A0_t (\SboxInst.L8 ), .B0_t (\SboxInst.L10 ), .Z0_t (\SboxInst.L27 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_L28.U1 ( .A0_t (\SboxInst.L11 ), .B0_t (\SboxInst.L14 ), .Z0_t (\SboxInst.L28 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) \SboxInst.XOR_L29.U1 ( .A0_t (\SboxInst.L11 ), .B0_t (\SboxInst.L17 ), .Z0_t (\SboxInst.L29 ) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) \SboxInst.XOR_S0.U1 ( .A0_t (\SboxInst.L6 ), .B0_t (\SboxInst.L24 ), .Z0_t (value_out[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) \SboxInst.XOR_S1.U1 ( .A0_t (\SboxInst.L16 ), .B0_t (\SboxInst.L26 ), .Z0_t (value_out[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) \SboxInst.XOR_S2.U1 ( .A0_t (\SboxInst.L19 ), .B0_t (\SboxInst.L28 ), .Z0_t (value_out[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) \SboxInst.XOR_S3.U1 ( .A0_t (\SboxInst.L6 ), .B0_t (\SboxInst.L21 ), .Z0_t (value_out[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) \SboxInst.XOR_S4.U1 ( .A0_t (\SboxInst.L20 ), .B0_t (\SboxInst.L22 ), .Z0_t (value_out[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) \SboxInst.XOR_S5.U1 ( .A0_t (\SboxInst.L25 ), .B0_t (\SboxInst.L29 ), .Z0_t (value_out[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) \SboxInst.XOR_S6.U1 ( .A0_t (\SboxInst.L13 ), .B0_t (\SboxInst.L27 ), .Z0_t (value_out[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) \SboxInst.XOR_S7.U1 ( .A0_t (\SboxInst.L6 ), .B0_t (\SboxInst.L23 ), .Z0_t (value_out[0]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) \M2.gen_loop_0__M.X1.U1 ( .A0_t (Inc_Reg[0]), .B0_t (start[0]), .Z0_t (\M2.gen_loop_0__M.X ) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) \M2.gen_loop_0__M.A.U1 ( .A0_t (rst), .B0_t (\M2.gen_loop_0__M.X ), .Z0_t (\M2.gen_loop_0__M.Y ) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) \M2.gen_loop_0__M.X2.U1 ( .A0_t (\M2.gen_loop_0__M.Y ), .B0_t (Inc_Reg[0]), .Z0_t (Inc_in[0]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) \M2.gen_loop_1__M.X1.U1 ( .A0_t (Inc_Reg[1]), .B0_t (start[1]), .Z0_t (\M2.gen_loop_1__M.X ) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) \M2.gen_loop_1__M.A.U1 ( .A0_t (rst), .B0_t (\M2.gen_loop_1__M.X ), .Z0_t (\M2.gen_loop_1__M.Y ) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) \M2.gen_loop_1__M.X2.U1 ( .A0_t (\M2.gen_loop_1__M.Y ), .B0_t (Inc_Reg[1]), .Z0_t (Inc_in[1]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) \M2.gen_loop_2__M.X1.U1 ( .A0_t (Inc_Reg[2]), .B0_t (start[2]), .Z0_t (\M2.gen_loop_2__M.X ) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) \M2.gen_loop_2__M.A.U1 ( .A0_t (rst), .B0_t (\M2.gen_loop_2__M.X ), .Z0_t (\M2.gen_loop_2__M.Y ) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) \M2.gen_loop_2__M.X2.U1 ( .A0_t (\M2.gen_loop_2__M.Y ), .B0_t (Inc_Reg[2]), .Z0_t (Inc_in[2]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) \M2.gen_loop_3__M.X1.U1 ( .A0_t (Inc_Reg[3]), .B0_t (start[3]), .Z0_t (\M2.gen_loop_3__M.X ) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) \M2.gen_loop_3__M.A.U1 ( .A0_t (rst), .B0_t (\M2.gen_loop_3__M.X ), .Z0_t (\M2.gen_loop_3__M.Y ) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) \M2.gen_loop_3__M.X2.U1 ( .A0_t (\M2.gen_loop_3__M.Y ), .B0_t (Inc_Reg[3]), .Z0_t (Inc_in[3]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) U10 ( .A0_t (Inc_in[0]), .B0_t (Inc_in[1]), .Z0_t (n9) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b1), .NL(1'b0)) U12 ( .A0_t (Inc_in[1]), .B0_t (Inc_in[0]), .Z0_t (Inc_Reg[1]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1), .NL(1'b0)) U13 ( .A0_t (n9), .B0_t (Inc_in[2]), .Z0_t (Inc_Reg[2]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) U14 ( .A0_t (n9), .B0_t (Inc_in[2]), .Z0_t (n10) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b0)) U15 ( .A0_t (Inc_in[3]), .B0_t (n10), .Z0_t (Inc_out[3]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1), .NL(1'b0)) new_AGEMA_gate_182 ( .A0_t (Inc_in[0]), .B0_t (1'b0), .Z0_t (Inc_Reg[0]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1), .NL(1'b0)) new_AGEMA_gate_183 ( .A0_t (Inc_out[3]), .B0_t (1'b0), .Z0_t (Inc_Reg[3]) ) ;

    /* register cells */
endmodule