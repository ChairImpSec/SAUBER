/* modified netlist. Source: module AES in file /mnt/c/Users/amirm/Desktop/Papers_in_progress/SAUBER/Design for our FPGA/4-AES_EncSerial_PortParallel/4-AGEMA/AES.v */
/* 0 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 1 register stage(s) in total */

module AES_SAUBER_Pipeline_d1 (plaintext_s0_t, key_s0_t, start_t, plaintext_s0_f, plaintext_s1_t, plaintext_s1_f, key_s0_f, key_s1_t, key_s1_f, start_f, ciphertext_s0_t, done_t, ciphertext_s0_f, ciphertext_s1_t, ciphertext_s1_f, done_f);
    input [127:0] plaintext_s0_t ;
    input [127:0] key_s0_t ;
    input start_t ;
    input [127:0] plaintext_s0_f ;
    input [127:0] plaintext_s1_t ;
    input [127:0] plaintext_s1_f ;
    input [127:0] key_s0_f ;
    input [127:0] key_s1_t ;
    input [127:0] key_s1_f ;
    input start_f ;
    output [127:0] ciphertext_s0_t ;
    output done_t ;
    output [127:0] ciphertext_s0_f ;
    output [127:0] ciphertext_s1_t ;
    output [127:0] ciphertext_s1_f ;
    output done_f ;
    wire nReset ;
    wire selMC ;
    wire selXOR ;
    wire enRCon ;
    wire finalStep ;
    wire intFinal ;
    wire intselXOR ;
    wire notFirst ;
    wire n13 ;
    wire ctrl_n15 ;
    wire ctrl_n11 ;
    wire ctrl_n10 ;
    wire ctrl_n9 ;
    wire ctrl_n8 ;
    wire ctrl_n7 ;
    wire ctrl_n6 ;
    wire ctrl_n5 ;
    wire ctrl_n2 ;
    wire ctrl_seq4Out_1_ ;
    wire ctrl_seq4In_1_ ;
    wire ctrl_nRstSeq4 ;
    wire ctrl_n13 ;
    wire ctrl_seq6Out_4_ ;
    wire ctrl_seq6In_1_ ;
    wire ctrl_seq6In_2_ ;
    wire ctrl_seq6In_3_ ;
    wire ctrl_seq6In_4_ ;
    wire ctrl_seq6_SFF_0_MUXInst_Y ;
    wire ctrl_seq6_SFF_0_MUXInst_X ;
    wire ctrl_seq6_SFF_1_MUXInst_Y ;
    wire ctrl_seq6_SFF_1_MUXInst_X ;
    wire ctrl_seq6_SFF_2_MUXInst_Y ;
    wire ctrl_seq6_SFF_2_MUXInst_X ;
    wire ctrl_seq6_SFF_3_MUXInst_Y ;
    wire ctrl_seq6_SFF_3_MUXInst_X ;
    wire ctrl_seq6_SFF_4_MUXInst_Y ;
    wire ctrl_seq6_SFF_4_MUXInst_X ;
    wire ctrl_seq4_SFF_0_MUXInst_Y ;
    wire ctrl_seq4_SFF_0_MUXInst_X ;
    wire ctrl_seq4_SFF_1_MUXInst_Y ;
    wire ctrl_seq4_SFF_1_MUXInst_X ;
    wire MUX_StateIn_mux_inst_0_Y ;
    wire MUX_StateIn_mux_inst_0_X ;
    wire MUX_StateIn_mux_inst_1_Y ;
    wire MUX_StateIn_mux_inst_1_X ;
    wire MUX_StateIn_mux_inst_2_Y ;
    wire MUX_StateIn_mux_inst_2_X ;
    wire MUX_StateIn_mux_inst_3_Y ;
    wire MUX_StateIn_mux_inst_3_X ;
    wire MUX_StateIn_mux_inst_4_Y ;
    wire MUX_StateIn_mux_inst_4_X ;
    wire MUX_StateIn_mux_inst_5_Y ;
    wire MUX_StateIn_mux_inst_5_X ;
    wire MUX_StateIn_mux_inst_6_Y ;
    wire MUX_StateIn_mux_inst_6_X ;
    wire MUX_StateIn_mux_inst_7_Y ;
    wire MUX_StateIn_mux_inst_7_X ;
    wire stateArray_S00reg_gff_1_SFF_0_MUXInst_Y ;
    wire stateArray_S00reg_gff_1_SFF_0_MUXInst_X ;
    wire stateArray_S00reg_gff_1_SFF_1_MUXInst_Y ;
    wire stateArray_S00reg_gff_1_SFF_1_MUXInst_X ;
    wire stateArray_S00reg_gff_1_SFF_2_MUXInst_Y ;
    wire stateArray_S00reg_gff_1_SFF_2_MUXInst_X ;
    wire stateArray_S00reg_gff_1_SFF_3_MUXInst_Y ;
    wire stateArray_S00reg_gff_1_SFF_3_MUXInst_X ;
    wire stateArray_S00reg_gff_1_SFF_4_MUXInst_Y ;
    wire stateArray_S00reg_gff_1_SFF_4_MUXInst_X ;
    wire stateArray_S00reg_gff_1_SFF_5_MUXInst_Y ;
    wire stateArray_S00reg_gff_1_SFF_5_MUXInst_X ;
    wire stateArray_S00reg_gff_1_SFF_6_MUXInst_Y ;
    wire stateArray_S00reg_gff_1_SFF_6_MUXInst_X ;
    wire stateArray_S00reg_gff_1_SFF_7_MUXInst_Y ;
    wire stateArray_S00reg_gff_1_SFF_7_MUXInst_X ;
    wire stateArray_S01reg_gff_1_SFF_0_MUXInst_Y ;
    wire stateArray_S01reg_gff_1_SFF_0_MUXInst_X ;
    wire stateArray_S01reg_gff_1_SFF_1_MUXInst_Y ;
    wire stateArray_S01reg_gff_1_SFF_1_MUXInst_X ;
    wire stateArray_S01reg_gff_1_SFF_2_MUXInst_Y ;
    wire stateArray_S01reg_gff_1_SFF_2_MUXInst_X ;
    wire stateArray_S01reg_gff_1_SFF_3_MUXInst_Y ;
    wire stateArray_S01reg_gff_1_SFF_3_MUXInst_X ;
    wire stateArray_S01reg_gff_1_SFF_4_MUXInst_Y ;
    wire stateArray_S01reg_gff_1_SFF_4_MUXInst_X ;
    wire stateArray_S01reg_gff_1_SFF_5_MUXInst_Y ;
    wire stateArray_S01reg_gff_1_SFF_5_MUXInst_X ;
    wire stateArray_S01reg_gff_1_SFF_6_MUXInst_Y ;
    wire stateArray_S01reg_gff_1_SFF_6_MUXInst_X ;
    wire stateArray_S01reg_gff_1_SFF_7_MUXInst_Y ;
    wire stateArray_S01reg_gff_1_SFF_7_MUXInst_X ;
    wire stateArray_S02reg_gff_1_SFF_0_MUXInst_Y ;
    wire stateArray_S02reg_gff_1_SFF_0_MUXInst_X ;
    wire stateArray_S02reg_gff_1_SFF_1_MUXInst_Y ;
    wire stateArray_S02reg_gff_1_SFF_1_MUXInst_X ;
    wire stateArray_S02reg_gff_1_SFF_2_MUXInst_Y ;
    wire stateArray_S02reg_gff_1_SFF_2_MUXInst_X ;
    wire stateArray_S02reg_gff_1_SFF_3_MUXInst_Y ;
    wire stateArray_S02reg_gff_1_SFF_3_MUXInst_X ;
    wire stateArray_S02reg_gff_1_SFF_4_MUXInst_Y ;
    wire stateArray_S02reg_gff_1_SFF_4_MUXInst_X ;
    wire stateArray_S02reg_gff_1_SFF_5_MUXInst_Y ;
    wire stateArray_S02reg_gff_1_SFF_5_MUXInst_X ;
    wire stateArray_S02reg_gff_1_SFF_6_MUXInst_Y ;
    wire stateArray_S02reg_gff_1_SFF_6_MUXInst_X ;
    wire stateArray_S02reg_gff_1_SFF_7_MUXInst_Y ;
    wire stateArray_S02reg_gff_1_SFF_7_MUXInst_X ;
    wire stateArray_S03reg_gff_1_SFF_0_MUXInst_Y ;
    wire stateArray_S03reg_gff_1_SFF_0_MUXInst_X ;
    wire stateArray_S03reg_gff_1_SFF_1_MUXInst_Y ;
    wire stateArray_S03reg_gff_1_SFF_1_MUXInst_X ;
    wire stateArray_S03reg_gff_1_SFF_2_MUXInst_Y ;
    wire stateArray_S03reg_gff_1_SFF_2_MUXInst_X ;
    wire stateArray_S03reg_gff_1_SFF_3_MUXInst_Y ;
    wire stateArray_S03reg_gff_1_SFF_3_MUXInst_X ;
    wire stateArray_S03reg_gff_1_SFF_4_MUXInst_Y ;
    wire stateArray_S03reg_gff_1_SFF_4_MUXInst_X ;
    wire stateArray_S03reg_gff_1_SFF_5_MUXInst_Y ;
    wire stateArray_S03reg_gff_1_SFF_5_MUXInst_X ;
    wire stateArray_S03reg_gff_1_SFF_6_MUXInst_Y ;
    wire stateArray_S03reg_gff_1_SFF_6_MUXInst_X ;
    wire stateArray_S03reg_gff_1_SFF_7_MUXInst_Y ;
    wire stateArray_S03reg_gff_1_SFF_7_MUXInst_X ;
    wire stateArray_S10reg_gff_1_SFF_0_MUXInst_Y ;
    wire stateArray_S10reg_gff_1_SFF_0_MUXInst_X ;
    wire stateArray_S10reg_gff_1_SFF_1_MUXInst_Y ;
    wire stateArray_S10reg_gff_1_SFF_1_MUXInst_X ;
    wire stateArray_S10reg_gff_1_SFF_2_MUXInst_Y ;
    wire stateArray_S10reg_gff_1_SFF_2_MUXInst_X ;
    wire stateArray_S10reg_gff_1_SFF_3_MUXInst_Y ;
    wire stateArray_S10reg_gff_1_SFF_3_MUXInst_X ;
    wire stateArray_S10reg_gff_1_SFF_4_MUXInst_Y ;
    wire stateArray_S10reg_gff_1_SFF_4_MUXInst_X ;
    wire stateArray_S10reg_gff_1_SFF_5_MUXInst_Y ;
    wire stateArray_S10reg_gff_1_SFF_5_MUXInst_X ;
    wire stateArray_S10reg_gff_1_SFF_6_MUXInst_Y ;
    wire stateArray_S10reg_gff_1_SFF_6_MUXInst_X ;
    wire stateArray_S10reg_gff_1_SFF_7_MUXInst_Y ;
    wire stateArray_S10reg_gff_1_SFF_7_MUXInst_X ;
    wire stateArray_S11reg_gff_1_SFF_0_MUXInst_Y ;
    wire stateArray_S11reg_gff_1_SFF_0_MUXInst_X ;
    wire stateArray_S11reg_gff_1_SFF_1_MUXInst_Y ;
    wire stateArray_S11reg_gff_1_SFF_1_MUXInst_X ;
    wire stateArray_S11reg_gff_1_SFF_2_MUXInst_Y ;
    wire stateArray_S11reg_gff_1_SFF_2_MUXInst_X ;
    wire stateArray_S11reg_gff_1_SFF_3_MUXInst_Y ;
    wire stateArray_S11reg_gff_1_SFF_3_MUXInst_X ;
    wire stateArray_S11reg_gff_1_SFF_4_MUXInst_Y ;
    wire stateArray_S11reg_gff_1_SFF_4_MUXInst_X ;
    wire stateArray_S11reg_gff_1_SFF_5_MUXInst_Y ;
    wire stateArray_S11reg_gff_1_SFF_5_MUXInst_X ;
    wire stateArray_S11reg_gff_1_SFF_6_MUXInst_Y ;
    wire stateArray_S11reg_gff_1_SFF_6_MUXInst_X ;
    wire stateArray_S11reg_gff_1_SFF_7_MUXInst_Y ;
    wire stateArray_S11reg_gff_1_SFF_7_MUXInst_X ;
    wire stateArray_S12reg_gff_1_SFF_0_MUXInst_Y ;
    wire stateArray_S12reg_gff_1_SFF_0_MUXInst_X ;
    wire stateArray_S12reg_gff_1_SFF_1_MUXInst_Y ;
    wire stateArray_S12reg_gff_1_SFF_1_MUXInst_X ;
    wire stateArray_S12reg_gff_1_SFF_2_MUXInst_Y ;
    wire stateArray_S12reg_gff_1_SFF_2_MUXInst_X ;
    wire stateArray_S12reg_gff_1_SFF_3_MUXInst_Y ;
    wire stateArray_S12reg_gff_1_SFF_3_MUXInst_X ;
    wire stateArray_S12reg_gff_1_SFF_4_MUXInst_Y ;
    wire stateArray_S12reg_gff_1_SFF_4_MUXInst_X ;
    wire stateArray_S12reg_gff_1_SFF_5_MUXInst_Y ;
    wire stateArray_S12reg_gff_1_SFF_5_MUXInst_X ;
    wire stateArray_S12reg_gff_1_SFF_6_MUXInst_Y ;
    wire stateArray_S12reg_gff_1_SFF_6_MUXInst_X ;
    wire stateArray_S12reg_gff_1_SFF_7_MUXInst_Y ;
    wire stateArray_S12reg_gff_1_SFF_7_MUXInst_X ;
    wire stateArray_S13reg_gff_1_SFF_0_MUXInst_Y ;
    wire stateArray_S13reg_gff_1_SFF_0_MUXInst_X ;
    wire stateArray_S13reg_gff_1_SFF_1_MUXInst_Y ;
    wire stateArray_S13reg_gff_1_SFF_1_MUXInst_X ;
    wire stateArray_S13reg_gff_1_SFF_2_MUXInst_Y ;
    wire stateArray_S13reg_gff_1_SFF_2_MUXInst_X ;
    wire stateArray_S13reg_gff_1_SFF_3_MUXInst_Y ;
    wire stateArray_S13reg_gff_1_SFF_3_MUXInst_X ;
    wire stateArray_S13reg_gff_1_SFF_4_MUXInst_Y ;
    wire stateArray_S13reg_gff_1_SFF_4_MUXInst_X ;
    wire stateArray_S13reg_gff_1_SFF_5_MUXInst_Y ;
    wire stateArray_S13reg_gff_1_SFF_5_MUXInst_X ;
    wire stateArray_S13reg_gff_1_SFF_6_MUXInst_Y ;
    wire stateArray_S13reg_gff_1_SFF_6_MUXInst_X ;
    wire stateArray_S13reg_gff_1_SFF_7_MUXInst_Y ;
    wire stateArray_S13reg_gff_1_SFF_7_MUXInst_X ;
    wire stateArray_S20reg_gff_1_SFF_0_MUXInst_Y ;
    wire stateArray_S20reg_gff_1_SFF_0_MUXInst_X ;
    wire stateArray_S20reg_gff_1_SFF_1_MUXInst_Y ;
    wire stateArray_S20reg_gff_1_SFF_1_MUXInst_X ;
    wire stateArray_S20reg_gff_1_SFF_2_MUXInst_Y ;
    wire stateArray_S20reg_gff_1_SFF_2_MUXInst_X ;
    wire stateArray_S20reg_gff_1_SFF_3_MUXInst_Y ;
    wire stateArray_S20reg_gff_1_SFF_3_MUXInst_X ;
    wire stateArray_S20reg_gff_1_SFF_4_MUXInst_Y ;
    wire stateArray_S20reg_gff_1_SFF_4_MUXInst_X ;
    wire stateArray_S20reg_gff_1_SFF_5_MUXInst_Y ;
    wire stateArray_S20reg_gff_1_SFF_5_MUXInst_X ;
    wire stateArray_S20reg_gff_1_SFF_6_MUXInst_Y ;
    wire stateArray_S20reg_gff_1_SFF_6_MUXInst_X ;
    wire stateArray_S20reg_gff_1_SFF_7_MUXInst_Y ;
    wire stateArray_S20reg_gff_1_SFF_7_MUXInst_X ;
    wire stateArray_S21reg_gff_1_SFF_0_MUXInst_Y ;
    wire stateArray_S21reg_gff_1_SFF_0_MUXInst_X ;
    wire stateArray_S21reg_gff_1_SFF_1_MUXInst_Y ;
    wire stateArray_S21reg_gff_1_SFF_1_MUXInst_X ;
    wire stateArray_S21reg_gff_1_SFF_2_MUXInst_Y ;
    wire stateArray_S21reg_gff_1_SFF_2_MUXInst_X ;
    wire stateArray_S21reg_gff_1_SFF_3_MUXInst_Y ;
    wire stateArray_S21reg_gff_1_SFF_3_MUXInst_X ;
    wire stateArray_S21reg_gff_1_SFF_4_MUXInst_Y ;
    wire stateArray_S21reg_gff_1_SFF_4_MUXInst_X ;
    wire stateArray_S21reg_gff_1_SFF_5_MUXInst_Y ;
    wire stateArray_S21reg_gff_1_SFF_5_MUXInst_X ;
    wire stateArray_S21reg_gff_1_SFF_6_MUXInst_Y ;
    wire stateArray_S21reg_gff_1_SFF_6_MUXInst_X ;
    wire stateArray_S21reg_gff_1_SFF_7_MUXInst_Y ;
    wire stateArray_S21reg_gff_1_SFF_7_MUXInst_X ;
    wire stateArray_S22reg_gff_1_SFF_0_MUXInst_Y ;
    wire stateArray_S22reg_gff_1_SFF_0_MUXInst_X ;
    wire stateArray_S22reg_gff_1_SFF_1_MUXInst_Y ;
    wire stateArray_S22reg_gff_1_SFF_1_MUXInst_X ;
    wire stateArray_S22reg_gff_1_SFF_2_MUXInst_Y ;
    wire stateArray_S22reg_gff_1_SFF_2_MUXInst_X ;
    wire stateArray_S22reg_gff_1_SFF_3_MUXInst_Y ;
    wire stateArray_S22reg_gff_1_SFF_3_MUXInst_X ;
    wire stateArray_S22reg_gff_1_SFF_4_MUXInst_Y ;
    wire stateArray_S22reg_gff_1_SFF_4_MUXInst_X ;
    wire stateArray_S22reg_gff_1_SFF_5_MUXInst_Y ;
    wire stateArray_S22reg_gff_1_SFF_5_MUXInst_X ;
    wire stateArray_S22reg_gff_1_SFF_6_MUXInst_Y ;
    wire stateArray_S22reg_gff_1_SFF_6_MUXInst_X ;
    wire stateArray_S22reg_gff_1_SFF_7_MUXInst_Y ;
    wire stateArray_S22reg_gff_1_SFF_7_MUXInst_X ;
    wire stateArray_S23reg_gff_1_SFF_0_MUXInst_Y ;
    wire stateArray_S23reg_gff_1_SFF_0_MUXInst_X ;
    wire stateArray_S23reg_gff_1_SFF_1_MUXInst_Y ;
    wire stateArray_S23reg_gff_1_SFF_1_MUXInst_X ;
    wire stateArray_S23reg_gff_1_SFF_2_MUXInst_Y ;
    wire stateArray_S23reg_gff_1_SFF_2_MUXInst_X ;
    wire stateArray_S23reg_gff_1_SFF_3_MUXInst_Y ;
    wire stateArray_S23reg_gff_1_SFF_3_MUXInst_X ;
    wire stateArray_S23reg_gff_1_SFF_4_MUXInst_Y ;
    wire stateArray_S23reg_gff_1_SFF_4_MUXInst_X ;
    wire stateArray_S23reg_gff_1_SFF_5_MUXInst_Y ;
    wire stateArray_S23reg_gff_1_SFF_5_MUXInst_X ;
    wire stateArray_S23reg_gff_1_SFF_6_MUXInst_Y ;
    wire stateArray_S23reg_gff_1_SFF_6_MUXInst_X ;
    wire stateArray_S23reg_gff_1_SFF_7_MUXInst_Y ;
    wire stateArray_S23reg_gff_1_SFF_7_MUXInst_X ;
    wire stateArray_S30reg_gff_1_SFF_0_MUXInst_Y ;
    wire stateArray_S30reg_gff_1_SFF_0_MUXInst_X ;
    wire stateArray_S30reg_gff_1_SFF_1_MUXInst_Y ;
    wire stateArray_S30reg_gff_1_SFF_1_MUXInst_X ;
    wire stateArray_S30reg_gff_1_SFF_2_MUXInst_Y ;
    wire stateArray_S30reg_gff_1_SFF_2_MUXInst_X ;
    wire stateArray_S30reg_gff_1_SFF_3_MUXInst_Y ;
    wire stateArray_S30reg_gff_1_SFF_3_MUXInst_X ;
    wire stateArray_S30reg_gff_1_SFF_4_MUXInst_Y ;
    wire stateArray_S30reg_gff_1_SFF_4_MUXInst_X ;
    wire stateArray_S30reg_gff_1_SFF_5_MUXInst_Y ;
    wire stateArray_S30reg_gff_1_SFF_5_MUXInst_X ;
    wire stateArray_S30reg_gff_1_SFF_6_MUXInst_Y ;
    wire stateArray_S30reg_gff_1_SFF_6_MUXInst_X ;
    wire stateArray_S30reg_gff_1_SFF_7_MUXInst_Y ;
    wire stateArray_S30reg_gff_1_SFF_7_MUXInst_X ;
    wire stateArray_S31reg_gff_1_SFF_0_MUXInst_Y ;
    wire stateArray_S31reg_gff_1_SFF_0_MUXInst_X ;
    wire stateArray_S31reg_gff_1_SFF_1_MUXInst_Y ;
    wire stateArray_S31reg_gff_1_SFF_1_MUXInst_X ;
    wire stateArray_S31reg_gff_1_SFF_2_MUXInst_Y ;
    wire stateArray_S31reg_gff_1_SFF_2_MUXInst_X ;
    wire stateArray_S31reg_gff_1_SFF_3_MUXInst_Y ;
    wire stateArray_S31reg_gff_1_SFF_3_MUXInst_X ;
    wire stateArray_S31reg_gff_1_SFF_4_MUXInst_Y ;
    wire stateArray_S31reg_gff_1_SFF_4_MUXInst_X ;
    wire stateArray_S31reg_gff_1_SFF_5_MUXInst_Y ;
    wire stateArray_S31reg_gff_1_SFF_5_MUXInst_X ;
    wire stateArray_S31reg_gff_1_SFF_6_MUXInst_Y ;
    wire stateArray_S31reg_gff_1_SFF_6_MUXInst_X ;
    wire stateArray_S31reg_gff_1_SFF_7_MUXInst_Y ;
    wire stateArray_S31reg_gff_1_SFF_7_MUXInst_X ;
    wire stateArray_S32reg_gff_1_SFF_0_MUXInst_Y ;
    wire stateArray_S32reg_gff_1_SFF_0_MUXInst_X ;
    wire stateArray_S32reg_gff_1_SFF_1_MUXInst_Y ;
    wire stateArray_S32reg_gff_1_SFF_1_MUXInst_X ;
    wire stateArray_S32reg_gff_1_SFF_2_MUXInst_Y ;
    wire stateArray_S32reg_gff_1_SFF_2_MUXInst_X ;
    wire stateArray_S32reg_gff_1_SFF_3_MUXInst_Y ;
    wire stateArray_S32reg_gff_1_SFF_3_MUXInst_X ;
    wire stateArray_S32reg_gff_1_SFF_4_MUXInst_Y ;
    wire stateArray_S32reg_gff_1_SFF_4_MUXInst_X ;
    wire stateArray_S32reg_gff_1_SFF_5_MUXInst_Y ;
    wire stateArray_S32reg_gff_1_SFF_5_MUXInst_X ;
    wire stateArray_S32reg_gff_1_SFF_6_MUXInst_Y ;
    wire stateArray_S32reg_gff_1_SFF_6_MUXInst_X ;
    wire stateArray_S32reg_gff_1_SFF_7_MUXInst_Y ;
    wire stateArray_S32reg_gff_1_SFF_7_MUXInst_X ;
    wire stateArray_S33reg_gff_1_SFF_0_MUXInst_Y ;
    wire stateArray_S33reg_gff_1_SFF_0_MUXInst_X ;
    wire stateArray_S33reg_gff_1_SFF_1_MUXInst_Y ;
    wire stateArray_S33reg_gff_1_SFF_1_MUXInst_X ;
    wire stateArray_S33reg_gff_1_SFF_2_MUXInst_Y ;
    wire stateArray_S33reg_gff_1_SFF_2_MUXInst_X ;
    wire stateArray_S33reg_gff_1_SFF_3_MUXInst_Y ;
    wire stateArray_S33reg_gff_1_SFF_3_MUXInst_X ;
    wire stateArray_S33reg_gff_1_SFF_4_MUXInst_Y ;
    wire stateArray_S33reg_gff_1_SFF_4_MUXInst_X ;
    wire stateArray_S33reg_gff_1_SFF_5_MUXInst_Y ;
    wire stateArray_S33reg_gff_1_SFF_5_MUXInst_X ;
    wire stateArray_S33reg_gff_1_SFF_6_MUXInst_Y ;
    wire stateArray_S33reg_gff_1_SFF_6_MUXInst_X ;
    wire stateArray_S33reg_gff_1_SFF_7_MUXInst_Y ;
    wire stateArray_S33reg_gff_1_SFF_7_MUXInst_X ;
    wire stateArray_MUX_inS00ser_mux_inst_0_Y ;
    wire stateArray_MUX_inS00ser_mux_inst_0_X ;
    wire stateArray_MUX_inS00ser_mux_inst_1_Y ;
    wire stateArray_MUX_inS00ser_mux_inst_1_X ;
    wire stateArray_MUX_inS00ser_mux_inst_2_Y ;
    wire stateArray_MUX_inS00ser_mux_inst_2_X ;
    wire stateArray_MUX_inS00ser_mux_inst_3_Y ;
    wire stateArray_MUX_inS00ser_mux_inst_3_X ;
    wire stateArray_MUX_inS00ser_mux_inst_4_Y ;
    wire stateArray_MUX_inS00ser_mux_inst_4_X ;
    wire stateArray_MUX_inS00ser_mux_inst_5_Y ;
    wire stateArray_MUX_inS00ser_mux_inst_5_X ;
    wire stateArray_MUX_inS00ser_mux_inst_6_Y ;
    wire stateArray_MUX_inS00ser_mux_inst_6_X ;
    wire stateArray_MUX_inS00ser_mux_inst_7_Y ;
    wire stateArray_MUX_inS00ser_mux_inst_7_X ;
    wire stateArray_MUX_inS01ser_mux_inst_0_Y ;
    wire stateArray_MUX_inS01ser_mux_inst_0_X ;
    wire stateArray_MUX_inS01ser_mux_inst_1_Y ;
    wire stateArray_MUX_inS01ser_mux_inst_1_X ;
    wire stateArray_MUX_inS01ser_mux_inst_2_Y ;
    wire stateArray_MUX_inS01ser_mux_inst_2_X ;
    wire stateArray_MUX_inS01ser_mux_inst_3_Y ;
    wire stateArray_MUX_inS01ser_mux_inst_3_X ;
    wire stateArray_MUX_inS01ser_mux_inst_4_Y ;
    wire stateArray_MUX_inS01ser_mux_inst_4_X ;
    wire stateArray_MUX_inS01ser_mux_inst_5_Y ;
    wire stateArray_MUX_inS01ser_mux_inst_5_X ;
    wire stateArray_MUX_inS01ser_mux_inst_6_Y ;
    wire stateArray_MUX_inS01ser_mux_inst_6_X ;
    wire stateArray_MUX_inS01ser_mux_inst_7_Y ;
    wire stateArray_MUX_inS01ser_mux_inst_7_X ;
    wire stateArray_MUX_inS02ser_mux_inst_0_Y ;
    wire stateArray_MUX_inS02ser_mux_inst_0_X ;
    wire stateArray_MUX_inS02ser_mux_inst_1_Y ;
    wire stateArray_MUX_inS02ser_mux_inst_1_X ;
    wire stateArray_MUX_inS02ser_mux_inst_2_Y ;
    wire stateArray_MUX_inS02ser_mux_inst_2_X ;
    wire stateArray_MUX_inS02ser_mux_inst_3_Y ;
    wire stateArray_MUX_inS02ser_mux_inst_3_X ;
    wire stateArray_MUX_inS02ser_mux_inst_4_Y ;
    wire stateArray_MUX_inS02ser_mux_inst_4_X ;
    wire stateArray_MUX_inS02ser_mux_inst_5_Y ;
    wire stateArray_MUX_inS02ser_mux_inst_5_X ;
    wire stateArray_MUX_inS02ser_mux_inst_6_Y ;
    wire stateArray_MUX_inS02ser_mux_inst_6_X ;
    wire stateArray_MUX_inS02ser_mux_inst_7_Y ;
    wire stateArray_MUX_inS02ser_mux_inst_7_X ;
    wire stateArray_MUX_outS10_MC_mux_inst_0_Y ;
    wire stateArray_MUX_outS10_MC_mux_inst_0_X ;
    wire stateArray_MUX_outS10_MC_mux_inst_1_Y ;
    wire stateArray_MUX_outS10_MC_mux_inst_1_X ;
    wire stateArray_MUX_outS10_MC_mux_inst_2_Y ;
    wire stateArray_MUX_outS10_MC_mux_inst_2_X ;
    wire stateArray_MUX_outS10_MC_mux_inst_3_Y ;
    wire stateArray_MUX_outS10_MC_mux_inst_3_X ;
    wire stateArray_MUX_outS10_MC_mux_inst_4_Y ;
    wire stateArray_MUX_outS10_MC_mux_inst_4_X ;
    wire stateArray_MUX_outS10_MC_mux_inst_5_Y ;
    wire stateArray_MUX_outS10_MC_mux_inst_5_X ;
    wire stateArray_MUX_outS10_MC_mux_inst_6_Y ;
    wire stateArray_MUX_outS10_MC_mux_inst_6_X ;
    wire stateArray_MUX_outS10_MC_mux_inst_7_Y ;
    wire stateArray_MUX_outS10_MC_mux_inst_7_X ;
    wire stateArray_MUX_inS03ser_mux_inst_0_Y ;
    wire stateArray_MUX_inS03ser_mux_inst_0_X ;
    wire stateArray_MUX_inS03ser_mux_inst_1_Y ;
    wire stateArray_MUX_inS03ser_mux_inst_1_X ;
    wire stateArray_MUX_inS03ser_mux_inst_2_Y ;
    wire stateArray_MUX_inS03ser_mux_inst_2_X ;
    wire stateArray_MUX_inS03ser_mux_inst_3_Y ;
    wire stateArray_MUX_inS03ser_mux_inst_3_X ;
    wire stateArray_MUX_inS03ser_mux_inst_4_Y ;
    wire stateArray_MUX_inS03ser_mux_inst_4_X ;
    wire stateArray_MUX_inS03ser_mux_inst_5_Y ;
    wire stateArray_MUX_inS03ser_mux_inst_5_X ;
    wire stateArray_MUX_inS03ser_mux_inst_6_Y ;
    wire stateArray_MUX_inS03ser_mux_inst_6_X ;
    wire stateArray_MUX_inS03ser_mux_inst_7_Y ;
    wire stateArray_MUX_inS03ser_mux_inst_7_X ;
    wire stateArray_MUX_inS10ser_mux_inst_0_Y ;
    wire stateArray_MUX_inS10ser_mux_inst_0_X ;
    wire stateArray_MUX_inS10ser_mux_inst_1_Y ;
    wire stateArray_MUX_inS10ser_mux_inst_1_X ;
    wire stateArray_MUX_inS10ser_mux_inst_2_Y ;
    wire stateArray_MUX_inS10ser_mux_inst_2_X ;
    wire stateArray_MUX_inS10ser_mux_inst_3_Y ;
    wire stateArray_MUX_inS10ser_mux_inst_3_X ;
    wire stateArray_MUX_inS10ser_mux_inst_4_Y ;
    wire stateArray_MUX_inS10ser_mux_inst_4_X ;
    wire stateArray_MUX_inS10ser_mux_inst_5_Y ;
    wire stateArray_MUX_inS10ser_mux_inst_5_X ;
    wire stateArray_MUX_inS10ser_mux_inst_6_Y ;
    wire stateArray_MUX_inS10ser_mux_inst_6_X ;
    wire stateArray_MUX_inS10ser_mux_inst_7_Y ;
    wire stateArray_MUX_inS10ser_mux_inst_7_X ;
    wire stateArray_MUX_inS11ser_mux_inst_0_Y ;
    wire stateArray_MUX_inS11ser_mux_inst_0_X ;
    wire stateArray_MUX_inS11ser_mux_inst_1_Y ;
    wire stateArray_MUX_inS11ser_mux_inst_1_X ;
    wire stateArray_MUX_inS11ser_mux_inst_2_Y ;
    wire stateArray_MUX_inS11ser_mux_inst_2_X ;
    wire stateArray_MUX_inS11ser_mux_inst_3_Y ;
    wire stateArray_MUX_inS11ser_mux_inst_3_X ;
    wire stateArray_MUX_inS11ser_mux_inst_4_Y ;
    wire stateArray_MUX_inS11ser_mux_inst_4_X ;
    wire stateArray_MUX_inS11ser_mux_inst_5_Y ;
    wire stateArray_MUX_inS11ser_mux_inst_5_X ;
    wire stateArray_MUX_inS11ser_mux_inst_6_Y ;
    wire stateArray_MUX_inS11ser_mux_inst_6_X ;
    wire stateArray_MUX_inS11ser_mux_inst_7_Y ;
    wire stateArray_MUX_inS11ser_mux_inst_7_X ;
    wire stateArray_MUX_inS12ser_mux_inst_0_Y ;
    wire stateArray_MUX_inS12ser_mux_inst_0_X ;
    wire stateArray_MUX_inS12ser_mux_inst_1_Y ;
    wire stateArray_MUX_inS12ser_mux_inst_1_X ;
    wire stateArray_MUX_inS12ser_mux_inst_2_Y ;
    wire stateArray_MUX_inS12ser_mux_inst_2_X ;
    wire stateArray_MUX_inS12ser_mux_inst_3_Y ;
    wire stateArray_MUX_inS12ser_mux_inst_3_X ;
    wire stateArray_MUX_inS12ser_mux_inst_4_Y ;
    wire stateArray_MUX_inS12ser_mux_inst_4_X ;
    wire stateArray_MUX_inS12ser_mux_inst_5_Y ;
    wire stateArray_MUX_inS12ser_mux_inst_5_X ;
    wire stateArray_MUX_inS12ser_mux_inst_6_Y ;
    wire stateArray_MUX_inS12ser_mux_inst_6_X ;
    wire stateArray_MUX_inS12ser_mux_inst_7_Y ;
    wire stateArray_MUX_inS12ser_mux_inst_7_X ;
    wire stateArray_MUX_outS20_MC_mux_inst_0_Y ;
    wire stateArray_MUX_outS20_MC_mux_inst_0_X ;
    wire stateArray_MUX_outS20_MC_mux_inst_1_Y ;
    wire stateArray_MUX_outS20_MC_mux_inst_1_X ;
    wire stateArray_MUX_outS20_MC_mux_inst_2_Y ;
    wire stateArray_MUX_outS20_MC_mux_inst_2_X ;
    wire stateArray_MUX_outS20_MC_mux_inst_3_Y ;
    wire stateArray_MUX_outS20_MC_mux_inst_3_X ;
    wire stateArray_MUX_outS20_MC_mux_inst_4_Y ;
    wire stateArray_MUX_outS20_MC_mux_inst_4_X ;
    wire stateArray_MUX_outS20_MC_mux_inst_5_Y ;
    wire stateArray_MUX_outS20_MC_mux_inst_5_X ;
    wire stateArray_MUX_outS20_MC_mux_inst_6_Y ;
    wire stateArray_MUX_outS20_MC_mux_inst_6_X ;
    wire stateArray_MUX_outS20_MC_mux_inst_7_Y ;
    wire stateArray_MUX_outS20_MC_mux_inst_7_X ;
    wire stateArray_MUX_inS13ser_mux_inst_0_Y ;
    wire stateArray_MUX_inS13ser_mux_inst_0_X ;
    wire stateArray_MUX_inS13ser_mux_inst_1_Y ;
    wire stateArray_MUX_inS13ser_mux_inst_1_X ;
    wire stateArray_MUX_inS13ser_mux_inst_2_Y ;
    wire stateArray_MUX_inS13ser_mux_inst_2_X ;
    wire stateArray_MUX_inS13ser_mux_inst_3_Y ;
    wire stateArray_MUX_inS13ser_mux_inst_3_X ;
    wire stateArray_MUX_inS13ser_mux_inst_4_Y ;
    wire stateArray_MUX_inS13ser_mux_inst_4_X ;
    wire stateArray_MUX_inS13ser_mux_inst_5_Y ;
    wire stateArray_MUX_inS13ser_mux_inst_5_X ;
    wire stateArray_MUX_inS13ser_mux_inst_6_Y ;
    wire stateArray_MUX_inS13ser_mux_inst_6_X ;
    wire stateArray_MUX_inS13ser_mux_inst_7_Y ;
    wire stateArray_MUX_inS13ser_mux_inst_7_X ;
    wire stateArray_MUX_inS20ser_mux_inst_0_Y ;
    wire stateArray_MUX_inS20ser_mux_inst_0_X ;
    wire stateArray_MUX_inS20ser_mux_inst_1_Y ;
    wire stateArray_MUX_inS20ser_mux_inst_1_X ;
    wire stateArray_MUX_inS20ser_mux_inst_2_Y ;
    wire stateArray_MUX_inS20ser_mux_inst_2_X ;
    wire stateArray_MUX_inS20ser_mux_inst_3_Y ;
    wire stateArray_MUX_inS20ser_mux_inst_3_X ;
    wire stateArray_MUX_inS20ser_mux_inst_4_Y ;
    wire stateArray_MUX_inS20ser_mux_inst_4_X ;
    wire stateArray_MUX_inS20ser_mux_inst_5_Y ;
    wire stateArray_MUX_inS20ser_mux_inst_5_X ;
    wire stateArray_MUX_inS20ser_mux_inst_6_Y ;
    wire stateArray_MUX_inS20ser_mux_inst_6_X ;
    wire stateArray_MUX_inS20ser_mux_inst_7_Y ;
    wire stateArray_MUX_inS20ser_mux_inst_7_X ;
    wire stateArray_MUX_inS21ser_mux_inst_0_Y ;
    wire stateArray_MUX_inS21ser_mux_inst_0_X ;
    wire stateArray_MUX_inS21ser_mux_inst_1_Y ;
    wire stateArray_MUX_inS21ser_mux_inst_1_X ;
    wire stateArray_MUX_inS21ser_mux_inst_2_Y ;
    wire stateArray_MUX_inS21ser_mux_inst_2_X ;
    wire stateArray_MUX_inS21ser_mux_inst_3_Y ;
    wire stateArray_MUX_inS21ser_mux_inst_3_X ;
    wire stateArray_MUX_inS21ser_mux_inst_4_Y ;
    wire stateArray_MUX_inS21ser_mux_inst_4_X ;
    wire stateArray_MUX_inS21ser_mux_inst_5_Y ;
    wire stateArray_MUX_inS21ser_mux_inst_5_X ;
    wire stateArray_MUX_inS21ser_mux_inst_6_Y ;
    wire stateArray_MUX_inS21ser_mux_inst_6_X ;
    wire stateArray_MUX_inS21ser_mux_inst_7_Y ;
    wire stateArray_MUX_inS21ser_mux_inst_7_X ;
    wire stateArray_MUX_inS22ser_mux_inst_0_Y ;
    wire stateArray_MUX_inS22ser_mux_inst_0_X ;
    wire stateArray_MUX_inS22ser_mux_inst_1_Y ;
    wire stateArray_MUX_inS22ser_mux_inst_1_X ;
    wire stateArray_MUX_inS22ser_mux_inst_2_Y ;
    wire stateArray_MUX_inS22ser_mux_inst_2_X ;
    wire stateArray_MUX_inS22ser_mux_inst_3_Y ;
    wire stateArray_MUX_inS22ser_mux_inst_3_X ;
    wire stateArray_MUX_inS22ser_mux_inst_4_Y ;
    wire stateArray_MUX_inS22ser_mux_inst_4_X ;
    wire stateArray_MUX_inS22ser_mux_inst_5_Y ;
    wire stateArray_MUX_inS22ser_mux_inst_5_X ;
    wire stateArray_MUX_inS22ser_mux_inst_6_Y ;
    wire stateArray_MUX_inS22ser_mux_inst_6_X ;
    wire stateArray_MUX_inS22ser_mux_inst_7_Y ;
    wire stateArray_MUX_inS22ser_mux_inst_7_X ;
    wire stateArray_MUX_outS30_MC_mux_inst_0_Y ;
    wire stateArray_MUX_outS30_MC_mux_inst_0_X ;
    wire stateArray_MUX_outS30_MC_mux_inst_1_Y ;
    wire stateArray_MUX_outS30_MC_mux_inst_1_X ;
    wire stateArray_MUX_outS30_MC_mux_inst_2_Y ;
    wire stateArray_MUX_outS30_MC_mux_inst_2_X ;
    wire stateArray_MUX_outS30_MC_mux_inst_3_Y ;
    wire stateArray_MUX_outS30_MC_mux_inst_3_X ;
    wire stateArray_MUX_outS30_MC_mux_inst_4_Y ;
    wire stateArray_MUX_outS30_MC_mux_inst_4_X ;
    wire stateArray_MUX_outS30_MC_mux_inst_5_Y ;
    wire stateArray_MUX_outS30_MC_mux_inst_5_X ;
    wire stateArray_MUX_outS30_MC_mux_inst_6_Y ;
    wire stateArray_MUX_outS30_MC_mux_inst_6_X ;
    wire stateArray_MUX_outS30_MC_mux_inst_7_Y ;
    wire stateArray_MUX_outS30_MC_mux_inst_7_X ;
    wire stateArray_MUX_inS23ser_mux_inst_0_Y ;
    wire stateArray_MUX_inS23ser_mux_inst_0_X ;
    wire stateArray_MUX_inS23ser_mux_inst_1_Y ;
    wire stateArray_MUX_inS23ser_mux_inst_1_X ;
    wire stateArray_MUX_inS23ser_mux_inst_2_Y ;
    wire stateArray_MUX_inS23ser_mux_inst_2_X ;
    wire stateArray_MUX_inS23ser_mux_inst_3_Y ;
    wire stateArray_MUX_inS23ser_mux_inst_3_X ;
    wire stateArray_MUX_inS23ser_mux_inst_4_Y ;
    wire stateArray_MUX_inS23ser_mux_inst_4_X ;
    wire stateArray_MUX_inS23ser_mux_inst_5_Y ;
    wire stateArray_MUX_inS23ser_mux_inst_5_X ;
    wire stateArray_MUX_inS23ser_mux_inst_6_Y ;
    wire stateArray_MUX_inS23ser_mux_inst_6_X ;
    wire stateArray_MUX_inS23ser_mux_inst_7_Y ;
    wire stateArray_MUX_inS23ser_mux_inst_7_X ;
    wire stateArray_MUX_inS30ser_mux_inst_0_Y ;
    wire stateArray_MUX_inS30ser_mux_inst_0_X ;
    wire stateArray_MUX_inS30ser_mux_inst_1_Y ;
    wire stateArray_MUX_inS30ser_mux_inst_1_X ;
    wire stateArray_MUX_inS30ser_mux_inst_2_Y ;
    wire stateArray_MUX_inS30ser_mux_inst_2_X ;
    wire stateArray_MUX_inS30ser_mux_inst_3_Y ;
    wire stateArray_MUX_inS30ser_mux_inst_3_X ;
    wire stateArray_MUX_inS30ser_mux_inst_4_Y ;
    wire stateArray_MUX_inS30ser_mux_inst_4_X ;
    wire stateArray_MUX_inS30ser_mux_inst_5_Y ;
    wire stateArray_MUX_inS30ser_mux_inst_5_X ;
    wire stateArray_MUX_inS30ser_mux_inst_6_Y ;
    wire stateArray_MUX_inS30ser_mux_inst_6_X ;
    wire stateArray_MUX_inS30ser_mux_inst_7_Y ;
    wire stateArray_MUX_inS30ser_mux_inst_7_X ;
    wire stateArray_MUX_inS31ser_mux_inst_0_Y ;
    wire stateArray_MUX_inS31ser_mux_inst_0_X ;
    wire stateArray_MUX_inS31ser_mux_inst_1_Y ;
    wire stateArray_MUX_inS31ser_mux_inst_1_X ;
    wire stateArray_MUX_inS31ser_mux_inst_2_Y ;
    wire stateArray_MUX_inS31ser_mux_inst_2_X ;
    wire stateArray_MUX_inS31ser_mux_inst_3_Y ;
    wire stateArray_MUX_inS31ser_mux_inst_3_X ;
    wire stateArray_MUX_inS31ser_mux_inst_4_Y ;
    wire stateArray_MUX_inS31ser_mux_inst_4_X ;
    wire stateArray_MUX_inS31ser_mux_inst_5_Y ;
    wire stateArray_MUX_inS31ser_mux_inst_5_X ;
    wire stateArray_MUX_inS31ser_mux_inst_6_Y ;
    wire stateArray_MUX_inS31ser_mux_inst_6_X ;
    wire stateArray_MUX_inS31ser_mux_inst_7_Y ;
    wire stateArray_MUX_inS31ser_mux_inst_7_X ;
    wire stateArray_MUX_inS32ser_mux_inst_0_Y ;
    wire stateArray_MUX_inS32ser_mux_inst_0_X ;
    wire stateArray_MUX_inS32ser_mux_inst_1_Y ;
    wire stateArray_MUX_inS32ser_mux_inst_1_X ;
    wire stateArray_MUX_inS32ser_mux_inst_2_Y ;
    wire stateArray_MUX_inS32ser_mux_inst_2_X ;
    wire stateArray_MUX_inS32ser_mux_inst_3_Y ;
    wire stateArray_MUX_inS32ser_mux_inst_3_X ;
    wire stateArray_MUX_inS32ser_mux_inst_4_Y ;
    wire stateArray_MUX_inS32ser_mux_inst_4_X ;
    wire stateArray_MUX_inS32ser_mux_inst_5_Y ;
    wire stateArray_MUX_inS32ser_mux_inst_5_X ;
    wire stateArray_MUX_inS32ser_mux_inst_6_Y ;
    wire stateArray_MUX_inS32ser_mux_inst_6_X ;
    wire stateArray_MUX_inS32ser_mux_inst_7_Y ;
    wire stateArray_MUX_inS32ser_mux_inst_7_X ;
    wire stateArray_MUX_input_MC_mux_inst_0_Y ;
    wire stateArray_MUX_input_MC_mux_inst_0_X ;
    wire stateArray_MUX_input_MC_mux_inst_1_Y ;
    wire stateArray_MUX_input_MC_mux_inst_1_X ;
    wire stateArray_MUX_input_MC_mux_inst_2_Y ;
    wire stateArray_MUX_input_MC_mux_inst_2_X ;
    wire stateArray_MUX_input_MC_mux_inst_3_Y ;
    wire stateArray_MUX_input_MC_mux_inst_3_X ;
    wire stateArray_MUX_input_MC_mux_inst_4_Y ;
    wire stateArray_MUX_input_MC_mux_inst_4_X ;
    wire stateArray_MUX_input_MC_mux_inst_5_Y ;
    wire stateArray_MUX_input_MC_mux_inst_5_X ;
    wire stateArray_MUX_input_MC_mux_inst_6_Y ;
    wire stateArray_MUX_input_MC_mux_inst_6_X ;
    wire stateArray_MUX_input_MC_mux_inst_7_Y ;
    wire stateArray_MUX_input_MC_mux_inst_7_X ;
    wire stateArray_MUX_inS33ser_mux_inst_0_Y ;
    wire stateArray_MUX_inS33ser_mux_inst_0_X ;
    wire stateArray_MUX_inS33ser_mux_inst_1_Y ;
    wire stateArray_MUX_inS33ser_mux_inst_1_X ;
    wire stateArray_MUX_inS33ser_mux_inst_2_Y ;
    wire stateArray_MUX_inS33ser_mux_inst_2_X ;
    wire stateArray_MUX_inS33ser_mux_inst_3_Y ;
    wire stateArray_MUX_inS33ser_mux_inst_3_X ;
    wire stateArray_MUX_inS33ser_mux_inst_4_Y ;
    wire stateArray_MUX_inS33ser_mux_inst_4_X ;
    wire stateArray_MUX_inS33ser_mux_inst_5_Y ;
    wire stateArray_MUX_inS33ser_mux_inst_5_X ;
    wire stateArray_MUX_inS33ser_mux_inst_6_Y ;
    wire stateArray_MUX_inS33ser_mux_inst_6_X ;
    wire stateArray_MUX_inS33ser_mux_inst_7_Y ;
    wire stateArray_MUX_inS33ser_mux_inst_7_X ;
    wire MUX_StateInMC_mux_inst_0_Y ;
    wire MUX_StateInMC_mux_inst_0_X ;
    wire MUX_StateInMC_mux_inst_1_Y ;
    wire MUX_StateInMC_mux_inst_1_X ;
    wire MUX_StateInMC_mux_inst_2_Y ;
    wire MUX_StateInMC_mux_inst_2_X ;
    wire MUX_StateInMC_mux_inst_3_Y ;
    wire MUX_StateInMC_mux_inst_3_X ;
    wire MUX_StateInMC_mux_inst_4_Y ;
    wire MUX_StateInMC_mux_inst_4_X ;
    wire MUX_StateInMC_mux_inst_5_Y ;
    wire MUX_StateInMC_mux_inst_5_X ;
    wire MUX_StateInMC_mux_inst_6_Y ;
    wire MUX_StateInMC_mux_inst_6_X ;
    wire MUX_StateInMC_mux_inst_7_Y ;
    wire MUX_StateInMC_mux_inst_7_X ;
    wire MUX_StateInMC_mux_inst_8_Y ;
    wire MUX_StateInMC_mux_inst_8_X ;
    wire MUX_StateInMC_mux_inst_9_Y ;
    wire MUX_StateInMC_mux_inst_9_X ;
    wire MUX_StateInMC_mux_inst_10_Y ;
    wire MUX_StateInMC_mux_inst_10_X ;
    wire MUX_StateInMC_mux_inst_11_Y ;
    wire MUX_StateInMC_mux_inst_11_X ;
    wire MUX_StateInMC_mux_inst_12_Y ;
    wire MUX_StateInMC_mux_inst_12_X ;
    wire MUX_StateInMC_mux_inst_13_Y ;
    wire MUX_StateInMC_mux_inst_13_X ;
    wire MUX_StateInMC_mux_inst_14_Y ;
    wire MUX_StateInMC_mux_inst_14_X ;
    wire MUX_StateInMC_mux_inst_15_Y ;
    wire MUX_StateInMC_mux_inst_15_X ;
    wire MUX_StateInMC_mux_inst_16_Y ;
    wire MUX_StateInMC_mux_inst_16_X ;
    wire MUX_StateInMC_mux_inst_17_Y ;
    wire MUX_StateInMC_mux_inst_17_X ;
    wire MUX_StateInMC_mux_inst_18_Y ;
    wire MUX_StateInMC_mux_inst_18_X ;
    wire MUX_StateInMC_mux_inst_19_Y ;
    wire MUX_StateInMC_mux_inst_19_X ;
    wire MUX_StateInMC_mux_inst_20_Y ;
    wire MUX_StateInMC_mux_inst_20_X ;
    wire MUX_StateInMC_mux_inst_21_Y ;
    wire MUX_StateInMC_mux_inst_21_X ;
    wire MUX_StateInMC_mux_inst_22_Y ;
    wire MUX_StateInMC_mux_inst_22_X ;
    wire MUX_StateInMC_mux_inst_23_Y ;
    wire MUX_StateInMC_mux_inst_23_X ;
    wire MUX_StateInMC_mux_inst_24_Y ;
    wire MUX_StateInMC_mux_inst_24_X ;
    wire MUX_StateInMC_mux_inst_25_Y ;
    wire MUX_StateInMC_mux_inst_25_X ;
    wire MUX_StateInMC_mux_inst_26_Y ;
    wire MUX_StateInMC_mux_inst_26_X ;
    wire MUX_StateInMC_mux_inst_27_Y ;
    wire MUX_StateInMC_mux_inst_27_X ;
    wire MUX_StateInMC_mux_inst_28_Y ;
    wire MUX_StateInMC_mux_inst_28_X ;
    wire MUX_StateInMC_mux_inst_29_Y ;
    wire MUX_StateInMC_mux_inst_29_X ;
    wire MUX_StateInMC_mux_inst_30_Y ;
    wire MUX_StateInMC_mux_inst_30_X ;
    wire MUX_StateInMC_mux_inst_31_Y ;
    wire MUX_StateInMC_mux_inst_31_X ;
    wire KeyArray_n40 ;
    wire KeyArray_n39 ;
    wire KeyArray_n38 ;
    wire KeyArray_n37 ;
    wire KeyArray_n36 ;
    wire KeyArray_n35 ;
    wire KeyArray_n34 ;
    wire KeyArray_n33 ;
    wire KeyArray_outS01ser_0_ ;
    wire KeyArray_outS01ser_1_ ;
    wire KeyArray_outS01ser_2_ ;
    wire KeyArray_outS01ser_3_ ;
    wire KeyArray_outS01ser_4_ ;
    wire KeyArray_outS01ser_5_ ;
    wire KeyArray_outS01ser_6_ ;
    wire KeyArray_outS01ser_7_ ;
    wire KeyArray_S00reg_gff_1_SFF_0_n2 ;
    wire KeyArray_S00reg_gff_1_SFF_0_n1 ;
    wire KeyArray_S00reg_gff_1_SFF_0_QD ;
    wire KeyArray_S00reg_gff_1_SFF_0_MUXInst_Y ;
    wire KeyArray_S00reg_gff_1_SFF_0_MUXInst_X ;
    wire KeyArray_S00reg_gff_1_SFF_1_n2 ;
    wire KeyArray_S00reg_gff_1_SFF_1_n1 ;
    wire KeyArray_S00reg_gff_1_SFF_1_QD ;
    wire KeyArray_S00reg_gff_1_SFF_1_MUXInst_Y ;
    wire KeyArray_S00reg_gff_1_SFF_1_MUXInst_X ;
    wire KeyArray_S00reg_gff_1_SFF_2_n2 ;
    wire KeyArray_S00reg_gff_1_SFF_2_n1 ;
    wire KeyArray_S00reg_gff_1_SFF_2_QD ;
    wire KeyArray_S00reg_gff_1_SFF_2_MUXInst_Y ;
    wire KeyArray_S00reg_gff_1_SFF_2_MUXInst_X ;
    wire KeyArray_S00reg_gff_1_SFF_3_n2 ;
    wire KeyArray_S00reg_gff_1_SFF_3_n1 ;
    wire KeyArray_S00reg_gff_1_SFF_3_QD ;
    wire KeyArray_S00reg_gff_1_SFF_3_MUXInst_Y ;
    wire KeyArray_S00reg_gff_1_SFF_3_MUXInst_X ;
    wire KeyArray_S00reg_gff_1_SFF_4_n2 ;
    wire KeyArray_S00reg_gff_1_SFF_4_n1 ;
    wire KeyArray_S00reg_gff_1_SFF_4_QD ;
    wire KeyArray_S00reg_gff_1_SFF_4_MUXInst_Y ;
    wire KeyArray_S00reg_gff_1_SFF_4_MUXInst_X ;
    wire KeyArray_S00reg_gff_1_SFF_5_n2 ;
    wire KeyArray_S00reg_gff_1_SFF_5_n1 ;
    wire KeyArray_S00reg_gff_1_SFF_5_QD ;
    wire KeyArray_S00reg_gff_1_SFF_5_MUXInst_Y ;
    wire KeyArray_S00reg_gff_1_SFF_5_MUXInst_X ;
    wire KeyArray_S00reg_gff_1_SFF_6_n2 ;
    wire KeyArray_S00reg_gff_1_SFF_6_n1 ;
    wire KeyArray_S00reg_gff_1_SFF_6_QD ;
    wire KeyArray_S00reg_gff_1_SFF_6_MUXInst_Y ;
    wire KeyArray_S00reg_gff_1_SFF_6_MUXInst_X ;
    wire KeyArray_S00reg_gff_1_SFF_7_n2 ;
    wire KeyArray_S00reg_gff_1_SFF_7_n1 ;
    wire KeyArray_S00reg_gff_1_SFF_7_QD ;
    wire KeyArray_S00reg_gff_1_SFF_7_MUXInst_Y ;
    wire KeyArray_S00reg_gff_1_SFF_7_MUXInst_X ;
    wire KeyArray_S01reg_gff_1_SFF_0_n2 ;
    wire KeyArray_S01reg_gff_1_SFF_0_n1 ;
    wire KeyArray_S01reg_gff_1_SFF_0_QD ;
    wire KeyArray_S01reg_gff_1_SFF_0_MUXInst_Y ;
    wire KeyArray_S01reg_gff_1_SFF_0_MUXInst_X ;
    wire KeyArray_S01reg_gff_1_SFF_1_n2 ;
    wire KeyArray_S01reg_gff_1_SFF_1_n1 ;
    wire KeyArray_S01reg_gff_1_SFF_1_QD ;
    wire KeyArray_S01reg_gff_1_SFF_1_MUXInst_Y ;
    wire KeyArray_S01reg_gff_1_SFF_1_MUXInst_X ;
    wire KeyArray_S01reg_gff_1_SFF_2_n2 ;
    wire KeyArray_S01reg_gff_1_SFF_2_n1 ;
    wire KeyArray_S01reg_gff_1_SFF_2_QD ;
    wire KeyArray_S01reg_gff_1_SFF_2_MUXInst_Y ;
    wire KeyArray_S01reg_gff_1_SFF_2_MUXInst_X ;
    wire KeyArray_S01reg_gff_1_SFF_3_n2 ;
    wire KeyArray_S01reg_gff_1_SFF_3_n1 ;
    wire KeyArray_S01reg_gff_1_SFF_3_QD ;
    wire KeyArray_S01reg_gff_1_SFF_3_MUXInst_Y ;
    wire KeyArray_S01reg_gff_1_SFF_3_MUXInst_X ;
    wire KeyArray_S01reg_gff_1_SFF_4_n2 ;
    wire KeyArray_S01reg_gff_1_SFF_4_n1 ;
    wire KeyArray_S01reg_gff_1_SFF_4_QD ;
    wire KeyArray_S01reg_gff_1_SFF_4_MUXInst_Y ;
    wire KeyArray_S01reg_gff_1_SFF_4_MUXInst_X ;
    wire KeyArray_S01reg_gff_1_SFF_5_n2 ;
    wire KeyArray_S01reg_gff_1_SFF_5_n1 ;
    wire KeyArray_S01reg_gff_1_SFF_5_QD ;
    wire KeyArray_S01reg_gff_1_SFF_5_MUXInst_Y ;
    wire KeyArray_S01reg_gff_1_SFF_5_MUXInst_X ;
    wire KeyArray_S01reg_gff_1_SFF_6_n2 ;
    wire KeyArray_S01reg_gff_1_SFF_6_n1 ;
    wire KeyArray_S01reg_gff_1_SFF_6_QD ;
    wire KeyArray_S01reg_gff_1_SFF_6_MUXInst_Y ;
    wire KeyArray_S01reg_gff_1_SFF_6_MUXInst_X ;
    wire KeyArray_S01reg_gff_1_SFF_7_n2 ;
    wire KeyArray_S01reg_gff_1_SFF_7_n1 ;
    wire KeyArray_S01reg_gff_1_SFF_7_QD ;
    wire KeyArray_S01reg_gff_1_SFF_7_MUXInst_Y ;
    wire KeyArray_S01reg_gff_1_SFF_7_MUXInst_X ;
    wire KeyArray_S02reg_gff_1_SFF_0_n2 ;
    wire KeyArray_S02reg_gff_1_SFF_0_n1 ;
    wire KeyArray_S02reg_gff_1_SFF_0_QD ;
    wire KeyArray_S02reg_gff_1_SFF_0_MUXInst_Y ;
    wire KeyArray_S02reg_gff_1_SFF_0_MUXInst_X ;
    wire KeyArray_S02reg_gff_1_SFF_1_n2 ;
    wire KeyArray_S02reg_gff_1_SFF_1_n1 ;
    wire KeyArray_S02reg_gff_1_SFF_1_QD ;
    wire KeyArray_S02reg_gff_1_SFF_1_MUXInst_Y ;
    wire KeyArray_S02reg_gff_1_SFF_1_MUXInst_X ;
    wire KeyArray_S02reg_gff_1_SFF_2_n2 ;
    wire KeyArray_S02reg_gff_1_SFF_2_n1 ;
    wire KeyArray_S02reg_gff_1_SFF_2_QD ;
    wire KeyArray_S02reg_gff_1_SFF_2_MUXInst_Y ;
    wire KeyArray_S02reg_gff_1_SFF_2_MUXInst_X ;
    wire KeyArray_S02reg_gff_1_SFF_3_n2 ;
    wire KeyArray_S02reg_gff_1_SFF_3_n1 ;
    wire KeyArray_S02reg_gff_1_SFF_3_QD ;
    wire KeyArray_S02reg_gff_1_SFF_3_MUXInst_Y ;
    wire KeyArray_S02reg_gff_1_SFF_3_MUXInst_X ;
    wire KeyArray_S02reg_gff_1_SFF_4_n2 ;
    wire KeyArray_S02reg_gff_1_SFF_4_n1 ;
    wire KeyArray_S02reg_gff_1_SFF_4_QD ;
    wire KeyArray_S02reg_gff_1_SFF_4_MUXInst_Y ;
    wire KeyArray_S02reg_gff_1_SFF_4_MUXInst_X ;
    wire KeyArray_S02reg_gff_1_SFF_5_n2 ;
    wire KeyArray_S02reg_gff_1_SFF_5_n1 ;
    wire KeyArray_S02reg_gff_1_SFF_5_QD ;
    wire KeyArray_S02reg_gff_1_SFF_5_MUXInst_Y ;
    wire KeyArray_S02reg_gff_1_SFF_5_MUXInst_X ;
    wire KeyArray_S02reg_gff_1_SFF_6_n2 ;
    wire KeyArray_S02reg_gff_1_SFF_6_n1 ;
    wire KeyArray_S02reg_gff_1_SFF_6_QD ;
    wire KeyArray_S02reg_gff_1_SFF_6_MUXInst_Y ;
    wire KeyArray_S02reg_gff_1_SFF_6_MUXInst_X ;
    wire KeyArray_S02reg_gff_1_SFF_7_n2 ;
    wire KeyArray_S02reg_gff_1_SFF_7_n1 ;
    wire KeyArray_S02reg_gff_1_SFF_7_QD ;
    wire KeyArray_S02reg_gff_1_SFF_7_MUXInst_Y ;
    wire KeyArray_S02reg_gff_1_SFF_7_MUXInst_X ;
    wire KeyArray_S03reg_gff_1_SFF_0_n2 ;
    wire KeyArray_S03reg_gff_1_SFF_0_n1 ;
    wire KeyArray_S03reg_gff_1_SFF_0_QD ;
    wire KeyArray_S03reg_gff_1_SFF_0_MUXInst_Y ;
    wire KeyArray_S03reg_gff_1_SFF_0_MUXInst_X ;
    wire KeyArray_S03reg_gff_1_SFF_1_n2 ;
    wire KeyArray_S03reg_gff_1_SFF_1_n1 ;
    wire KeyArray_S03reg_gff_1_SFF_1_QD ;
    wire KeyArray_S03reg_gff_1_SFF_1_MUXInst_Y ;
    wire KeyArray_S03reg_gff_1_SFF_1_MUXInst_X ;
    wire KeyArray_S03reg_gff_1_SFF_2_n2 ;
    wire KeyArray_S03reg_gff_1_SFF_2_n1 ;
    wire KeyArray_S03reg_gff_1_SFF_2_QD ;
    wire KeyArray_S03reg_gff_1_SFF_2_MUXInst_Y ;
    wire KeyArray_S03reg_gff_1_SFF_2_MUXInst_X ;
    wire KeyArray_S03reg_gff_1_SFF_3_n2 ;
    wire KeyArray_S03reg_gff_1_SFF_3_n1 ;
    wire KeyArray_S03reg_gff_1_SFF_3_QD ;
    wire KeyArray_S03reg_gff_1_SFF_3_MUXInst_Y ;
    wire KeyArray_S03reg_gff_1_SFF_3_MUXInst_X ;
    wire KeyArray_S03reg_gff_1_SFF_4_n2 ;
    wire KeyArray_S03reg_gff_1_SFF_4_n1 ;
    wire KeyArray_S03reg_gff_1_SFF_4_QD ;
    wire KeyArray_S03reg_gff_1_SFF_4_MUXInst_Y ;
    wire KeyArray_S03reg_gff_1_SFF_4_MUXInst_X ;
    wire KeyArray_S03reg_gff_1_SFF_5_n2 ;
    wire KeyArray_S03reg_gff_1_SFF_5_n1 ;
    wire KeyArray_S03reg_gff_1_SFF_5_QD ;
    wire KeyArray_S03reg_gff_1_SFF_5_MUXInst_Y ;
    wire KeyArray_S03reg_gff_1_SFF_5_MUXInst_X ;
    wire KeyArray_S03reg_gff_1_SFF_6_n2 ;
    wire KeyArray_S03reg_gff_1_SFF_6_n1 ;
    wire KeyArray_S03reg_gff_1_SFF_6_QD ;
    wire KeyArray_S03reg_gff_1_SFF_6_MUXInst_Y ;
    wire KeyArray_S03reg_gff_1_SFF_6_MUXInst_X ;
    wire KeyArray_S03reg_gff_1_SFF_7_n2 ;
    wire KeyArray_S03reg_gff_1_SFF_7_n1 ;
    wire KeyArray_S03reg_gff_1_SFF_7_QD ;
    wire KeyArray_S03reg_gff_1_SFF_7_MUXInst_Y ;
    wire KeyArray_S03reg_gff_1_SFF_7_MUXInst_X ;
    wire KeyArray_S10reg_gff_1_SFF_0_n2 ;
    wire KeyArray_S10reg_gff_1_SFF_0_n1 ;
    wire KeyArray_S10reg_gff_1_SFF_0_QD ;
    wire KeyArray_S10reg_gff_1_SFF_0_MUXInst_Y ;
    wire KeyArray_S10reg_gff_1_SFF_0_MUXInst_X ;
    wire KeyArray_S10reg_gff_1_SFF_1_n2 ;
    wire KeyArray_S10reg_gff_1_SFF_1_n1 ;
    wire KeyArray_S10reg_gff_1_SFF_1_QD ;
    wire KeyArray_S10reg_gff_1_SFF_1_MUXInst_Y ;
    wire KeyArray_S10reg_gff_1_SFF_1_MUXInst_X ;
    wire KeyArray_S10reg_gff_1_SFF_2_n2 ;
    wire KeyArray_S10reg_gff_1_SFF_2_n1 ;
    wire KeyArray_S10reg_gff_1_SFF_2_QD ;
    wire KeyArray_S10reg_gff_1_SFF_2_MUXInst_Y ;
    wire KeyArray_S10reg_gff_1_SFF_2_MUXInst_X ;
    wire KeyArray_S10reg_gff_1_SFF_3_n2 ;
    wire KeyArray_S10reg_gff_1_SFF_3_n1 ;
    wire KeyArray_S10reg_gff_1_SFF_3_QD ;
    wire KeyArray_S10reg_gff_1_SFF_3_MUXInst_Y ;
    wire KeyArray_S10reg_gff_1_SFF_3_MUXInst_X ;
    wire KeyArray_S10reg_gff_1_SFF_4_n2 ;
    wire KeyArray_S10reg_gff_1_SFF_4_n1 ;
    wire KeyArray_S10reg_gff_1_SFF_4_QD ;
    wire KeyArray_S10reg_gff_1_SFF_4_MUXInst_Y ;
    wire KeyArray_S10reg_gff_1_SFF_4_MUXInst_X ;
    wire KeyArray_S10reg_gff_1_SFF_5_n2 ;
    wire KeyArray_S10reg_gff_1_SFF_5_n1 ;
    wire KeyArray_S10reg_gff_1_SFF_5_QD ;
    wire KeyArray_S10reg_gff_1_SFF_5_MUXInst_Y ;
    wire KeyArray_S10reg_gff_1_SFF_5_MUXInst_X ;
    wire KeyArray_S10reg_gff_1_SFF_6_n2 ;
    wire KeyArray_S10reg_gff_1_SFF_6_n1 ;
    wire KeyArray_S10reg_gff_1_SFF_6_QD ;
    wire KeyArray_S10reg_gff_1_SFF_6_MUXInst_Y ;
    wire KeyArray_S10reg_gff_1_SFF_6_MUXInst_X ;
    wire KeyArray_S10reg_gff_1_SFF_7_n2 ;
    wire KeyArray_S10reg_gff_1_SFF_7_n1 ;
    wire KeyArray_S10reg_gff_1_SFF_7_QD ;
    wire KeyArray_S10reg_gff_1_SFF_7_MUXInst_Y ;
    wire KeyArray_S10reg_gff_1_SFF_7_MUXInst_X ;
    wire KeyArray_S11reg_gff_1_SFF_0_n2 ;
    wire KeyArray_S11reg_gff_1_SFF_0_n1 ;
    wire KeyArray_S11reg_gff_1_SFF_0_QD ;
    wire KeyArray_S11reg_gff_1_SFF_0_MUXInst_Y ;
    wire KeyArray_S11reg_gff_1_SFF_0_MUXInst_X ;
    wire KeyArray_S11reg_gff_1_SFF_1_n2 ;
    wire KeyArray_S11reg_gff_1_SFF_1_n1 ;
    wire KeyArray_S11reg_gff_1_SFF_1_QD ;
    wire KeyArray_S11reg_gff_1_SFF_1_MUXInst_Y ;
    wire KeyArray_S11reg_gff_1_SFF_1_MUXInst_X ;
    wire KeyArray_S11reg_gff_1_SFF_2_n2 ;
    wire KeyArray_S11reg_gff_1_SFF_2_n1 ;
    wire KeyArray_S11reg_gff_1_SFF_2_QD ;
    wire KeyArray_S11reg_gff_1_SFF_2_MUXInst_Y ;
    wire KeyArray_S11reg_gff_1_SFF_2_MUXInst_X ;
    wire KeyArray_S11reg_gff_1_SFF_3_n2 ;
    wire KeyArray_S11reg_gff_1_SFF_3_n1 ;
    wire KeyArray_S11reg_gff_1_SFF_3_QD ;
    wire KeyArray_S11reg_gff_1_SFF_3_MUXInst_Y ;
    wire KeyArray_S11reg_gff_1_SFF_3_MUXInst_X ;
    wire KeyArray_S11reg_gff_1_SFF_4_n2 ;
    wire KeyArray_S11reg_gff_1_SFF_4_n1 ;
    wire KeyArray_S11reg_gff_1_SFF_4_QD ;
    wire KeyArray_S11reg_gff_1_SFF_4_MUXInst_Y ;
    wire KeyArray_S11reg_gff_1_SFF_4_MUXInst_X ;
    wire KeyArray_S11reg_gff_1_SFF_5_n2 ;
    wire KeyArray_S11reg_gff_1_SFF_5_n1 ;
    wire KeyArray_S11reg_gff_1_SFF_5_QD ;
    wire KeyArray_S11reg_gff_1_SFF_5_MUXInst_Y ;
    wire KeyArray_S11reg_gff_1_SFF_5_MUXInst_X ;
    wire KeyArray_S11reg_gff_1_SFF_6_n2 ;
    wire KeyArray_S11reg_gff_1_SFF_6_n1 ;
    wire KeyArray_S11reg_gff_1_SFF_6_QD ;
    wire KeyArray_S11reg_gff_1_SFF_6_MUXInst_Y ;
    wire KeyArray_S11reg_gff_1_SFF_6_MUXInst_X ;
    wire KeyArray_S11reg_gff_1_SFF_7_n2 ;
    wire KeyArray_S11reg_gff_1_SFF_7_n1 ;
    wire KeyArray_S11reg_gff_1_SFF_7_QD ;
    wire KeyArray_S11reg_gff_1_SFF_7_MUXInst_Y ;
    wire KeyArray_S11reg_gff_1_SFF_7_MUXInst_X ;
    wire KeyArray_S12reg_gff_1_SFF_0_n2 ;
    wire KeyArray_S12reg_gff_1_SFF_0_n1 ;
    wire KeyArray_S12reg_gff_1_SFF_0_QD ;
    wire KeyArray_S12reg_gff_1_SFF_0_MUXInst_Y ;
    wire KeyArray_S12reg_gff_1_SFF_0_MUXInst_X ;
    wire KeyArray_S12reg_gff_1_SFF_1_n2 ;
    wire KeyArray_S12reg_gff_1_SFF_1_n1 ;
    wire KeyArray_S12reg_gff_1_SFF_1_QD ;
    wire KeyArray_S12reg_gff_1_SFF_1_MUXInst_Y ;
    wire KeyArray_S12reg_gff_1_SFF_1_MUXInst_X ;
    wire KeyArray_S12reg_gff_1_SFF_2_n2 ;
    wire KeyArray_S12reg_gff_1_SFF_2_n1 ;
    wire KeyArray_S12reg_gff_1_SFF_2_QD ;
    wire KeyArray_S12reg_gff_1_SFF_2_MUXInst_Y ;
    wire KeyArray_S12reg_gff_1_SFF_2_MUXInst_X ;
    wire KeyArray_S12reg_gff_1_SFF_3_n2 ;
    wire KeyArray_S12reg_gff_1_SFF_3_n1 ;
    wire KeyArray_S12reg_gff_1_SFF_3_QD ;
    wire KeyArray_S12reg_gff_1_SFF_3_MUXInst_Y ;
    wire KeyArray_S12reg_gff_1_SFF_3_MUXInst_X ;
    wire KeyArray_S12reg_gff_1_SFF_4_n2 ;
    wire KeyArray_S12reg_gff_1_SFF_4_n1 ;
    wire KeyArray_S12reg_gff_1_SFF_4_QD ;
    wire KeyArray_S12reg_gff_1_SFF_4_MUXInst_Y ;
    wire KeyArray_S12reg_gff_1_SFF_4_MUXInst_X ;
    wire KeyArray_S12reg_gff_1_SFF_5_n2 ;
    wire KeyArray_S12reg_gff_1_SFF_5_n1 ;
    wire KeyArray_S12reg_gff_1_SFF_5_QD ;
    wire KeyArray_S12reg_gff_1_SFF_5_MUXInst_Y ;
    wire KeyArray_S12reg_gff_1_SFF_5_MUXInst_X ;
    wire KeyArray_S12reg_gff_1_SFF_6_n2 ;
    wire KeyArray_S12reg_gff_1_SFF_6_n1 ;
    wire KeyArray_S12reg_gff_1_SFF_6_QD ;
    wire KeyArray_S12reg_gff_1_SFF_6_MUXInst_Y ;
    wire KeyArray_S12reg_gff_1_SFF_6_MUXInst_X ;
    wire KeyArray_S12reg_gff_1_SFF_7_n2 ;
    wire KeyArray_S12reg_gff_1_SFF_7_n1 ;
    wire KeyArray_S12reg_gff_1_SFF_7_QD ;
    wire KeyArray_S12reg_gff_1_SFF_7_MUXInst_Y ;
    wire KeyArray_S12reg_gff_1_SFF_7_MUXInst_X ;
    wire KeyArray_S13reg_gff_1_SFF_0_n2 ;
    wire KeyArray_S13reg_gff_1_SFF_0_n1 ;
    wire KeyArray_S13reg_gff_1_SFF_0_QD ;
    wire KeyArray_S13reg_gff_1_SFF_0_MUXInst_Y ;
    wire KeyArray_S13reg_gff_1_SFF_0_MUXInst_X ;
    wire KeyArray_S13reg_gff_1_SFF_1_n2 ;
    wire KeyArray_S13reg_gff_1_SFF_1_n1 ;
    wire KeyArray_S13reg_gff_1_SFF_1_QD ;
    wire KeyArray_S13reg_gff_1_SFF_1_MUXInst_Y ;
    wire KeyArray_S13reg_gff_1_SFF_1_MUXInst_X ;
    wire KeyArray_S13reg_gff_1_SFF_2_n2 ;
    wire KeyArray_S13reg_gff_1_SFF_2_n1 ;
    wire KeyArray_S13reg_gff_1_SFF_2_QD ;
    wire KeyArray_S13reg_gff_1_SFF_2_MUXInst_Y ;
    wire KeyArray_S13reg_gff_1_SFF_2_MUXInst_X ;
    wire KeyArray_S13reg_gff_1_SFF_3_n2 ;
    wire KeyArray_S13reg_gff_1_SFF_3_n1 ;
    wire KeyArray_S13reg_gff_1_SFF_3_QD ;
    wire KeyArray_S13reg_gff_1_SFF_3_MUXInst_Y ;
    wire KeyArray_S13reg_gff_1_SFF_3_MUXInst_X ;
    wire KeyArray_S13reg_gff_1_SFF_4_n2 ;
    wire KeyArray_S13reg_gff_1_SFF_4_n1 ;
    wire KeyArray_S13reg_gff_1_SFF_4_QD ;
    wire KeyArray_S13reg_gff_1_SFF_4_MUXInst_Y ;
    wire KeyArray_S13reg_gff_1_SFF_4_MUXInst_X ;
    wire KeyArray_S13reg_gff_1_SFF_5_n2 ;
    wire KeyArray_S13reg_gff_1_SFF_5_n1 ;
    wire KeyArray_S13reg_gff_1_SFF_5_QD ;
    wire KeyArray_S13reg_gff_1_SFF_5_MUXInst_Y ;
    wire KeyArray_S13reg_gff_1_SFF_5_MUXInst_X ;
    wire KeyArray_S13reg_gff_1_SFF_6_n2 ;
    wire KeyArray_S13reg_gff_1_SFF_6_n1 ;
    wire KeyArray_S13reg_gff_1_SFF_6_QD ;
    wire KeyArray_S13reg_gff_1_SFF_6_MUXInst_Y ;
    wire KeyArray_S13reg_gff_1_SFF_6_MUXInst_X ;
    wire KeyArray_S13reg_gff_1_SFF_7_n2 ;
    wire KeyArray_S13reg_gff_1_SFF_7_n1 ;
    wire KeyArray_S13reg_gff_1_SFF_7_QD ;
    wire KeyArray_S13reg_gff_1_SFF_7_MUXInst_Y ;
    wire KeyArray_S13reg_gff_1_SFF_7_MUXInst_X ;
    wire KeyArray_S20reg_gff_1_SFF_0_n2 ;
    wire KeyArray_S20reg_gff_1_SFF_0_n1 ;
    wire KeyArray_S20reg_gff_1_SFF_0_QD ;
    wire KeyArray_S20reg_gff_1_SFF_0_MUXInst_Y ;
    wire KeyArray_S20reg_gff_1_SFF_0_MUXInst_X ;
    wire KeyArray_S20reg_gff_1_SFF_1_n2 ;
    wire KeyArray_S20reg_gff_1_SFF_1_n1 ;
    wire KeyArray_S20reg_gff_1_SFF_1_QD ;
    wire KeyArray_S20reg_gff_1_SFF_1_MUXInst_Y ;
    wire KeyArray_S20reg_gff_1_SFF_1_MUXInst_X ;
    wire KeyArray_S20reg_gff_1_SFF_2_n2 ;
    wire KeyArray_S20reg_gff_1_SFF_2_n1 ;
    wire KeyArray_S20reg_gff_1_SFF_2_QD ;
    wire KeyArray_S20reg_gff_1_SFF_2_MUXInst_Y ;
    wire KeyArray_S20reg_gff_1_SFF_2_MUXInst_X ;
    wire KeyArray_S20reg_gff_1_SFF_3_n2 ;
    wire KeyArray_S20reg_gff_1_SFF_3_n1 ;
    wire KeyArray_S20reg_gff_1_SFF_3_QD ;
    wire KeyArray_S20reg_gff_1_SFF_3_MUXInst_Y ;
    wire KeyArray_S20reg_gff_1_SFF_3_MUXInst_X ;
    wire KeyArray_S20reg_gff_1_SFF_4_n2 ;
    wire KeyArray_S20reg_gff_1_SFF_4_n1 ;
    wire KeyArray_S20reg_gff_1_SFF_4_QD ;
    wire KeyArray_S20reg_gff_1_SFF_4_MUXInst_Y ;
    wire KeyArray_S20reg_gff_1_SFF_4_MUXInst_X ;
    wire KeyArray_S20reg_gff_1_SFF_5_n2 ;
    wire KeyArray_S20reg_gff_1_SFF_5_n1 ;
    wire KeyArray_S20reg_gff_1_SFF_5_QD ;
    wire KeyArray_S20reg_gff_1_SFF_5_MUXInst_Y ;
    wire KeyArray_S20reg_gff_1_SFF_5_MUXInst_X ;
    wire KeyArray_S20reg_gff_1_SFF_6_n2 ;
    wire KeyArray_S20reg_gff_1_SFF_6_n1 ;
    wire KeyArray_S20reg_gff_1_SFF_6_QD ;
    wire KeyArray_S20reg_gff_1_SFF_6_MUXInst_Y ;
    wire KeyArray_S20reg_gff_1_SFF_6_MUXInst_X ;
    wire KeyArray_S20reg_gff_1_SFF_7_n2 ;
    wire KeyArray_S20reg_gff_1_SFF_7_n1 ;
    wire KeyArray_S20reg_gff_1_SFF_7_QD ;
    wire KeyArray_S20reg_gff_1_SFF_7_MUXInst_Y ;
    wire KeyArray_S20reg_gff_1_SFF_7_MUXInst_X ;
    wire KeyArray_S21reg_gff_1_SFF_0_n2 ;
    wire KeyArray_S21reg_gff_1_SFF_0_n1 ;
    wire KeyArray_S21reg_gff_1_SFF_0_QD ;
    wire KeyArray_S21reg_gff_1_SFF_0_MUXInst_Y ;
    wire KeyArray_S21reg_gff_1_SFF_0_MUXInst_X ;
    wire KeyArray_S21reg_gff_1_SFF_1_n2 ;
    wire KeyArray_S21reg_gff_1_SFF_1_n1 ;
    wire KeyArray_S21reg_gff_1_SFF_1_QD ;
    wire KeyArray_S21reg_gff_1_SFF_1_MUXInst_Y ;
    wire KeyArray_S21reg_gff_1_SFF_1_MUXInst_X ;
    wire KeyArray_S21reg_gff_1_SFF_2_n2 ;
    wire KeyArray_S21reg_gff_1_SFF_2_n1 ;
    wire KeyArray_S21reg_gff_1_SFF_2_QD ;
    wire KeyArray_S21reg_gff_1_SFF_2_MUXInst_Y ;
    wire KeyArray_S21reg_gff_1_SFF_2_MUXInst_X ;
    wire KeyArray_S21reg_gff_1_SFF_3_n2 ;
    wire KeyArray_S21reg_gff_1_SFF_3_n1 ;
    wire KeyArray_S21reg_gff_1_SFF_3_QD ;
    wire KeyArray_S21reg_gff_1_SFF_3_MUXInst_Y ;
    wire KeyArray_S21reg_gff_1_SFF_3_MUXInst_X ;
    wire KeyArray_S21reg_gff_1_SFF_4_n2 ;
    wire KeyArray_S21reg_gff_1_SFF_4_n1 ;
    wire KeyArray_S21reg_gff_1_SFF_4_QD ;
    wire KeyArray_S21reg_gff_1_SFF_4_MUXInst_Y ;
    wire KeyArray_S21reg_gff_1_SFF_4_MUXInst_X ;
    wire KeyArray_S21reg_gff_1_SFF_5_n2 ;
    wire KeyArray_S21reg_gff_1_SFF_5_n1 ;
    wire KeyArray_S21reg_gff_1_SFF_5_QD ;
    wire KeyArray_S21reg_gff_1_SFF_5_MUXInst_Y ;
    wire KeyArray_S21reg_gff_1_SFF_5_MUXInst_X ;
    wire KeyArray_S21reg_gff_1_SFF_6_n2 ;
    wire KeyArray_S21reg_gff_1_SFF_6_n1 ;
    wire KeyArray_S21reg_gff_1_SFF_6_QD ;
    wire KeyArray_S21reg_gff_1_SFF_6_MUXInst_Y ;
    wire KeyArray_S21reg_gff_1_SFF_6_MUXInst_X ;
    wire KeyArray_S21reg_gff_1_SFF_7_n2 ;
    wire KeyArray_S21reg_gff_1_SFF_7_n1 ;
    wire KeyArray_S21reg_gff_1_SFF_7_QD ;
    wire KeyArray_S21reg_gff_1_SFF_7_MUXInst_Y ;
    wire KeyArray_S21reg_gff_1_SFF_7_MUXInst_X ;
    wire KeyArray_S22reg_gff_1_SFF_0_n2 ;
    wire KeyArray_S22reg_gff_1_SFF_0_n1 ;
    wire KeyArray_S22reg_gff_1_SFF_0_QD ;
    wire KeyArray_S22reg_gff_1_SFF_0_MUXInst_Y ;
    wire KeyArray_S22reg_gff_1_SFF_0_MUXInst_X ;
    wire KeyArray_S22reg_gff_1_SFF_1_n2 ;
    wire KeyArray_S22reg_gff_1_SFF_1_n1 ;
    wire KeyArray_S22reg_gff_1_SFF_1_QD ;
    wire KeyArray_S22reg_gff_1_SFF_1_MUXInst_Y ;
    wire KeyArray_S22reg_gff_1_SFF_1_MUXInst_X ;
    wire KeyArray_S22reg_gff_1_SFF_2_n2 ;
    wire KeyArray_S22reg_gff_1_SFF_2_n1 ;
    wire KeyArray_S22reg_gff_1_SFF_2_QD ;
    wire KeyArray_S22reg_gff_1_SFF_2_MUXInst_Y ;
    wire KeyArray_S22reg_gff_1_SFF_2_MUXInst_X ;
    wire KeyArray_S22reg_gff_1_SFF_3_n2 ;
    wire KeyArray_S22reg_gff_1_SFF_3_n1 ;
    wire KeyArray_S22reg_gff_1_SFF_3_QD ;
    wire KeyArray_S22reg_gff_1_SFF_3_MUXInst_Y ;
    wire KeyArray_S22reg_gff_1_SFF_3_MUXInst_X ;
    wire KeyArray_S22reg_gff_1_SFF_4_n2 ;
    wire KeyArray_S22reg_gff_1_SFF_4_n1 ;
    wire KeyArray_S22reg_gff_1_SFF_4_QD ;
    wire KeyArray_S22reg_gff_1_SFF_4_MUXInst_Y ;
    wire KeyArray_S22reg_gff_1_SFF_4_MUXInst_X ;
    wire KeyArray_S22reg_gff_1_SFF_5_n2 ;
    wire KeyArray_S22reg_gff_1_SFF_5_n1 ;
    wire KeyArray_S22reg_gff_1_SFF_5_QD ;
    wire KeyArray_S22reg_gff_1_SFF_5_MUXInst_Y ;
    wire KeyArray_S22reg_gff_1_SFF_5_MUXInst_X ;
    wire KeyArray_S22reg_gff_1_SFF_6_n2 ;
    wire KeyArray_S22reg_gff_1_SFF_6_n1 ;
    wire KeyArray_S22reg_gff_1_SFF_6_QD ;
    wire KeyArray_S22reg_gff_1_SFF_6_MUXInst_Y ;
    wire KeyArray_S22reg_gff_1_SFF_6_MUXInst_X ;
    wire KeyArray_S22reg_gff_1_SFF_7_n2 ;
    wire KeyArray_S22reg_gff_1_SFF_7_n1 ;
    wire KeyArray_S22reg_gff_1_SFF_7_QD ;
    wire KeyArray_S22reg_gff_1_SFF_7_MUXInst_Y ;
    wire KeyArray_S22reg_gff_1_SFF_7_MUXInst_X ;
    wire KeyArray_S23reg_gff_1_SFF_0_n2 ;
    wire KeyArray_S23reg_gff_1_SFF_0_n1 ;
    wire KeyArray_S23reg_gff_1_SFF_0_QD ;
    wire KeyArray_S23reg_gff_1_SFF_0_MUXInst_Y ;
    wire KeyArray_S23reg_gff_1_SFF_0_MUXInst_X ;
    wire KeyArray_S23reg_gff_1_SFF_1_n2 ;
    wire KeyArray_S23reg_gff_1_SFF_1_n1 ;
    wire KeyArray_S23reg_gff_1_SFF_1_QD ;
    wire KeyArray_S23reg_gff_1_SFF_1_MUXInst_Y ;
    wire KeyArray_S23reg_gff_1_SFF_1_MUXInst_X ;
    wire KeyArray_S23reg_gff_1_SFF_2_n2 ;
    wire KeyArray_S23reg_gff_1_SFF_2_n1 ;
    wire KeyArray_S23reg_gff_1_SFF_2_QD ;
    wire KeyArray_S23reg_gff_1_SFF_2_MUXInst_Y ;
    wire KeyArray_S23reg_gff_1_SFF_2_MUXInst_X ;
    wire KeyArray_S23reg_gff_1_SFF_3_n2 ;
    wire KeyArray_S23reg_gff_1_SFF_3_n1 ;
    wire KeyArray_S23reg_gff_1_SFF_3_QD ;
    wire KeyArray_S23reg_gff_1_SFF_3_MUXInst_Y ;
    wire KeyArray_S23reg_gff_1_SFF_3_MUXInst_X ;
    wire KeyArray_S23reg_gff_1_SFF_4_n2 ;
    wire KeyArray_S23reg_gff_1_SFF_4_n1 ;
    wire KeyArray_S23reg_gff_1_SFF_4_QD ;
    wire KeyArray_S23reg_gff_1_SFF_4_MUXInst_Y ;
    wire KeyArray_S23reg_gff_1_SFF_4_MUXInst_X ;
    wire KeyArray_S23reg_gff_1_SFF_5_n2 ;
    wire KeyArray_S23reg_gff_1_SFF_5_n1 ;
    wire KeyArray_S23reg_gff_1_SFF_5_QD ;
    wire KeyArray_S23reg_gff_1_SFF_5_MUXInst_Y ;
    wire KeyArray_S23reg_gff_1_SFF_5_MUXInst_X ;
    wire KeyArray_S23reg_gff_1_SFF_6_n2 ;
    wire KeyArray_S23reg_gff_1_SFF_6_n1 ;
    wire KeyArray_S23reg_gff_1_SFF_6_QD ;
    wire KeyArray_S23reg_gff_1_SFF_6_MUXInst_Y ;
    wire KeyArray_S23reg_gff_1_SFF_6_MUXInst_X ;
    wire KeyArray_S23reg_gff_1_SFF_7_n2 ;
    wire KeyArray_S23reg_gff_1_SFF_7_n1 ;
    wire KeyArray_S23reg_gff_1_SFF_7_QD ;
    wire KeyArray_S23reg_gff_1_SFF_7_MUXInst_Y ;
    wire KeyArray_S23reg_gff_1_SFF_7_MUXInst_X ;
    wire KeyArray_S30reg_gff_1_SFF_0_n2 ;
    wire KeyArray_S30reg_gff_1_SFF_0_n1 ;
    wire KeyArray_S30reg_gff_1_SFF_0_QD ;
    wire KeyArray_S30reg_gff_1_SFF_0_MUXInst_Y ;
    wire KeyArray_S30reg_gff_1_SFF_0_MUXInst_X ;
    wire KeyArray_S30reg_gff_1_SFF_1_n2 ;
    wire KeyArray_S30reg_gff_1_SFF_1_n1 ;
    wire KeyArray_S30reg_gff_1_SFF_1_QD ;
    wire KeyArray_S30reg_gff_1_SFF_1_MUXInst_Y ;
    wire KeyArray_S30reg_gff_1_SFF_1_MUXInst_X ;
    wire KeyArray_S30reg_gff_1_SFF_2_n2 ;
    wire KeyArray_S30reg_gff_1_SFF_2_n1 ;
    wire KeyArray_S30reg_gff_1_SFF_2_QD ;
    wire KeyArray_S30reg_gff_1_SFF_2_MUXInst_Y ;
    wire KeyArray_S30reg_gff_1_SFF_2_MUXInst_X ;
    wire KeyArray_S30reg_gff_1_SFF_3_n2 ;
    wire KeyArray_S30reg_gff_1_SFF_3_n1 ;
    wire KeyArray_S30reg_gff_1_SFF_3_QD ;
    wire KeyArray_S30reg_gff_1_SFF_3_MUXInst_Y ;
    wire KeyArray_S30reg_gff_1_SFF_3_MUXInst_X ;
    wire KeyArray_S30reg_gff_1_SFF_4_n2 ;
    wire KeyArray_S30reg_gff_1_SFF_4_n1 ;
    wire KeyArray_S30reg_gff_1_SFF_4_QD ;
    wire KeyArray_S30reg_gff_1_SFF_4_MUXInst_Y ;
    wire KeyArray_S30reg_gff_1_SFF_4_MUXInst_X ;
    wire KeyArray_S30reg_gff_1_SFF_5_n2 ;
    wire KeyArray_S30reg_gff_1_SFF_5_n1 ;
    wire KeyArray_S30reg_gff_1_SFF_5_QD ;
    wire KeyArray_S30reg_gff_1_SFF_5_MUXInst_Y ;
    wire KeyArray_S30reg_gff_1_SFF_5_MUXInst_X ;
    wire KeyArray_S30reg_gff_1_SFF_6_n2 ;
    wire KeyArray_S30reg_gff_1_SFF_6_n1 ;
    wire KeyArray_S30reg_gff_1_SFF_6_QD ;
    wire KeyArray_S30reg_gff_1_SFF_6_MUXInst_Y ;
    wire KeyArray_S30reg_gff_1_SFF_6_MUXInst_X ;
    wire KeyArray_S30reg_gff_1_SFF_7_n2 ;
    wire KeyArray_S30reg_gff_1_SFF_7_n1 ;
    wire KeyArray_S30reg_gff_1_SFF_7_QD ;
    wire KeyArray_S30reg_gff_1_SFF_7_MUXInst_Y ;
    wire KeyArray_S30reg_gff_1_SFF_7_MUXInst_X ;
    wire KeyArray_S31reg_gff_1_SFF_0_n2 ;
    wire KeyArray_S31reg_gff_1_SFF_0_n1 ;
    wire KeyArray_S31reg_gff_1_SFF_0_QD ;
    wire KeyArray_S31reg_gff_1_SFF_0_MUXInst_Y ;
    wire KeyArray_S31reg_gff_1_SFF_0_MUXInst_X ;
    wire KeyArray_S31reg_gff_1_SFF_1_n2 ;
    wire KeyArray_S31reg_gff_1_SFF_1_n1 ;
    wire KeyArray_S31reg_gff_1_SFF_1_QD ;
    wire KeyArray_S31reg_gff_1_SFF_1_MUXInst_Y ;
    wire KeyArray_S31reg_gff_1_SFF_1_MUXInst_X ;
    wire KeyArray_S31reg_gff_1_SFF_2_n2 ;
    wire KeyArray_S31reg_gff_1_SFF_2_n1 ;
    wire KeyArray_S31reg_gff_1_SFF_2_QD ;
    wire KeyArray_S31reg_gff_1_SFF_2_MUXInst_Y ;
    wire KeyArray_S31reg_gff_1_SFF_2_MUXInst_X ;
    wire KeyArray_S31reg_gff_1_SFF_3_n2 ;
    wire KeyArray_S31reg_gff_1_SFF_3_n1 ;
    wire KeyArray_S31reg_gff_1_SFF_3_QD ;
    wire KeyArray_S31reg_gff_1_SFF_3_MUXInst_Y ;
    wire KeyArray_S31reg_gff_1_SFF_3_MUXInst_X ;
    wire KeyArray_S31reg_gff_1_SFF_4_n2 ;
    wire KeyArray_S31reg_gff_1_SFF_4_n1 ;
    wire KeyArray_S31reg_gff_1_SFF_4_QD ;
    wire KeyArray_S31reg_gff_1_SFF_4_MUXInst_Y ;
    wire KeyArray_S31reg_gff_1_SFF_4_MUXInst_X ;
    wire KeyArray_S31reg_gff_1_SFF_5_n2 ;
    wire KeyArray_S31reg_gff_1_SFF_5_n1 ;
    wire KeyArray_S31reg_gff_1_SFF_5_QD ;
    wire KeyArray_S31reg_gff_1_SFF_5_MUXInst_Y ;
    wire KeyArray_S31reg_gff_1_SFF_5_MUXInst_X ;
    wire KeyArray_S31reg_gff_1_SFF_6_n2 ;
    wire KeyArray_S31reg_gff_1_SFF_6_n1 ;
    wire KeyArray_S31reg_gff_1_SFF_6_QD ;
    wire KeyArray_S31reg_gff_1_SFF_6_MUXInst_Y ;
    wire KeyArray_S31reg_gff_1_SFF_6_MUXInst_X ;
    wire KeyArray_S31reg_gff_1_SFF_7_n2 ;
    wire KeyArray_S31reg_gff_1_SFF_7_n1 ;
    wire KeyArray_S31reg_gff_1_SFF_7_QD ;
    wire KeyArray_S31reg_gff_1_SFF_7_MUXInst_Y ;
    wire KeyArray_S31reg_gff_1_SFF_7_MUXInst_X ;
    wire KeyArray_S32reg_gff_1_SFF_0_n2 ;
    wire KeyArray_S32reg_gff_1_SFF_0_n1 ;
    wire KeyArray_S32reg_gff_1_SFF_0_QD ;
    wire KeyArray_S32reg_gff_1_SFF_0_MUXInst_Y ;
    wire KeyArray_S32reg_gff_1_SFF_0_MUXInst_X ;
    wire KeyArray_S32reg_gff_1_SFF_1_n2 ;
    wire KeyArray_S32reg_gff_1_SFF_1_n1 ;
    wire KeyArray_S32reg_gff_1_SFF_1_QD ;
    wire KeyArray_S32reg_gff_1_SFF_1_MUXInst_Y ;
    wire KeyArray_S32reg_gff_1_SFF_1_MUXInst_X ;
    wire KeyArray_S32reg_gff_1_SFF_2_n2 ;
    wire KeyArray_S32reg_gff_1_SFF_2_n1 ;
    wire KeyArray_S32reg_gff_1_SFF_2_QD ;
    wire KeyArray_S32reg_gff_1_SFF_2_MUXInst_Y ;
    wire KeyArray_S32reg_gff_1_SFF_2_MUXInst_X ;
    wire KeyArray_S32reg_gff_1_SFF_3_n2 ;
    wire KeyArray_S32reg_gff_1_SFF_3_n1 ;
    wire KeyArray_S32reg_gff_1_SFF_3_QD ;
    wire KeyArray_S32reg_gff_1_SFF_3_MUXInst_Y ;
    wire KeyArray_S32reg_gff_1_SFF_3_MUXInst_X ;
    wire KeyArray_S32reg_gff_1_SFF_4_n2 ;
    wire KeyArray_S32reg_gff_1_SFF_4_n1 ;
    wire KeyArray_S32reg_gff_1_SFF_4_QD ;
    wire KeyArray_S32reg_gff_1_SFF_4_MUXInst_Y ;
    wire KeyArray_S32reg_gff_1_SFF_4_MUXInst_X ;
    wire KeyArray_S32reg_gff_1_SFF_5_n2 ;
    wire KeyArray_S32reg_gff_1_SFF_5_n1 ;
    wire KeyArray_S32reg_gff_1_SFF_5_QD ;
    wire KeyArray_S32reg_gff_1_SFF_5_MUXInst_Y ;
    wire KeyArray_S32reg_gff_1_SFF_5_MUXInst_X ;
    wire KeyArray_S32reg_gff_1_SFF_6_n2 ;
    wire KeyArray_S32reg_gff_1_SFF_6_n1 ;
    wire KeyArray_S32reg_gff_1_SFF_6_QD ;
    wire KeyArray_S32reg_gff_1_SFF_6_MUXInst_Y ;
    wire KeyArray_S32reg_gff_1_SFF_6_MUXInst_X ;
    wire KeyArray_S32reg_gff_1_SFF_7_n2 ;
    wire KeyArray_S32reg_gff_1_SFF_7_n1 ;
    wire KeyArray_S32reg_gff_1_SFF_7_QD ;
    wire KeyArray_S32reg_gff_1_SFF_7_MUXInst_Y ;
    wire KeyArray_S32reg_gff_1_SFF_7_MUXInst_X ;
    wire KeyArray_S33reg_gff_1_SFF_0_n2 ;
    wire KeyArray_S33reg_gff_1_SFF_0_n1 ;
    wire KeyArray_S33reg_gff_1_SFF_0_QD ;
    wire KeyArray_S33reg_gff_1_SFF_0_MUXInst_Y ;
    wire KeyArray_S33reg_gff_1_SFF_0_MUXInst_X ;
    wire KeyArray_S33reg_gff_1_SFF_1_n2 ;
    wire KeyArray_S33reg_gff_1_SFF_1_n1 ;
    wire KeyArray_S33reg_gff_1_SFF_1_QD ;
    wire KeyArray_S33reg_gff_1_SFF_1_MUXInst_Y ;
    wire KeyArray_S33reg_gff_1_SFF_1_MUXInst_X ;
    wire KeyArray_S33reg_gff_1_SFF_2_n2 ;
    wire KeyArray_S33reg_gff_1_SFF_2_n1 ;
    wire KeyArray_S33reg_gff_1_SFF_2_QD ;
    wire KeyArray_S33reg_gff_1_SFF_2_MUXInst_Y ;
    wire KeyArray_S33reg_gff_1_SFF_2_MUXInst_X ;
    wire KeyArray_S33reg_gff_1_SFF_3_n2 ;
    wire KeyArray_S33reg_gff_1_SFF_3_n1 ;
    wire KeyArray_S33reg_gff_1_SFF_3_QD ;
    wire KeyArray_S33reg_gff_1_SFF_3_MUXInst_Y ;
    wire KeyArray_S33reg_gff_1_SFF_3_MUXInst_X ;
    wire KeyArray_S33reg_gff_1_SFF_4_n2 ;
    wire KeyArray_S33reg_gff_1_SFF_4_n1 ;
    wire KeyArray_S33reg_gff_1_SFF_4_QD ;
    wire KeyArray_S33reg_gff_1_SFF_4_MUXInst_Y ;
    wire KeyArray_S33reg_gff_1_SFF_4_MUXInst_X ;
    wire KeyArray_S33reg_gff_1_SFF_5_n2 ;
    wire KeyArray_S33reg_gff_1_SFF_5_n1 ;
    wire KeyArray_S33reg_gff_1_SFF_5_QD ;
    wire KeyArray_S33reg_gff_1_SFF_5_MUXInst_Y ;
    wire KeyArray_S33reg_gff_1_SFF_5_MUXInst_X ;
    wire KeyArray_S33reg_gff_1_SFF_6_n2 ;
    wire KeyArray_S33reg_gff_1_SFF_6_n1 ;
    wire KeyArray_S33reg_gff_1_SFF_6_QD ;
    wire KeyArray_S33reg_gff_1_SFF_6_MUXInst_Y ;
    wire KeyArray_S33reg_gff_1_SFF_6_MUXInst_X ;
    wire KeyArray_S33reg_gff_1_SFF_7_n2 ;
    wire KeyArray_S33reg_gff_1_SFF_7_n1 ;
    wire KeyArray_S33reg_gff_1_SFF_7_QD ;
    wire KeyArray_S33reg_gff_1_SFF_7_MUXInst_Y ;
    wire KeyArray_S33reg_gff_1_SFF_7_MUXInst_X ;
    wire KeyArray_MUX_selXOR_mux_inst_0_Y ;
    wire KeyArray_MUX_selXOR_mux_inst_0_X ;
    wire KeyArray_MUX_selXOR_mux_inst_1_Y ;
    wire KeyArray_MUX_selXOR_mux_inst_1_X ;
    wire KeyArray_MUX_selXOR_mux_inst_2_Y ;
    wire KeyArray_MUX_selXOR_mux_inst_2_X ;
    wire KeyArray_MUX_selXOR_mux_inst_3_Y ;
    wire KeyArray_MUX_selXOR_mux_inst_3_X ;
    wire KeyArray_MUX_selXOR_mux_inst_4_Y ;
    wire KeyArray_MUX_selXOR_mux_inst_4_X ;
    wire KeyArray_MUX_selXOR_mux_inst_5_Y ;
    wire KeyArray_MUX_selXOR_mux_inst_5_X ;
    wire KeyArray_MUX_selXOR_mux_inst_6_Y ;
    wire KeyArray_MUX_selXOR_mux_inst_6_X ;
    wire KeyArray_MUX_selXOR_mux_inst_7_Y ;
    wire KeyArray_MUX_selXOR_mux_inst_7_X ;
    wire KeyArray_MUX_inS00ser_mux_inst_0_Y ;
    wire KeyArray_MUX_inS00ser_mux_inst_0_X ;
    wire KeyArray_MUX_inS00ser_mux_inst_1_Y ;
    wire KeyArray_MUX_inS00ser_mux_inst_1_X ;
    wire KeyArray_MUX_inS00ser_mux_inst_2_Y ;
    wire KeyArray_MUX_inS00ser_mux_inst_2_X ;
    wire KeyArray_MUX_inS00ser_mux_inst_3_Y ;
    wire KeyArray_MUX_inS00ser_mux_inst_3_X ;
    wire KeyArray_MUX_inS00ser_mux_inst_4_Y ;
    wire KeyArray_MUX_inS00ser_mux_inst_4_X ;
    wire KeyArray_MUX_inS00ser_mux_inst_5_Y ;
    wire KeyArray_MUX_inS00ser_mux_inst_5_X ;
    wire KeyArray_MUX_inS00ser_mux_inst_6_Y ;
    wire KeyArray_MUX_inS00ser_mux_inst_6_X ;
    wire KeyArray_MUX_inS00ser_mux_inst_7_Y ;
    wire KeyArray_MUX_inS00ser_mux_inst_7_X ;
    wire KeyArray_MUX_inS01ser_mux_inst_0_Y ;
    wire KeyArray_MUX_inS01ser_mux_inst_0_X ;
    wire KeyArray_MUX_inS01ser_mux_inst_1_Y ;
    wire KeyArray_MUX_inS01ser_mux_inst_1_X ;
    wire KeyArray_MUX_inS01ser_mux_inst_2_Y ;
    wire KeyArray_MUX_inS01ser_mux_inst_2_X ;
    wire KeyArray_MUX_inS01ser_mux_inst_3_Y ;
    wire KeyArray_MUX_inS01ser_mux_inst_3_X ;
    wire KeyArray_MUX_inS01ser_mux_inst_4_Y ;
    wire KeyArray_MUX_inS01ser_mux_inst_4_X ;
    wire KeyArray_MUX_inS01ser_mux_inst_5_Y ;
    wire KeyArray_MUX_inS01ser_mux_inst_5_X ;
    wire KeyArray_MUX_inS01ser_mux_inst_6_Y ;
    wire KeyArray_MUX_inS01ser_mux_inst_6_X ;
    wire KeyArray_MUX_inS01ser_mux_inst_7_Y ;
    wire KeyArray_MUX_inS01ser_mux_inst_7_X ;
    wire KeyArray_MUX_inS02ser_mux_inst_0_Y ;
    wire KeyArray_MUX_inS02ser_mux_inst_0_X ;
    wire KeyArray_MUX_inS02ser_mux_inst_1_Y ;
    wire KeyArray_MUX_inS02ser_mux_inst_1_X ;
    wire KeyArray_MUX_inS02ser_mux_inst_2_Y ;
    wire KeyArray_MUX_inS02ser_mux_inst_2_X ;
    wire KeyArray_MUX_inS02ser_mux_inst_3_Y ;
    wire KeyArray_MUX_inS02ser_mux_inst_3_X ;
    wire KeyArray_MUX_inS02ser_mux_inst_4_Y ;
    wire KeyArray_MUX_inS02ser_mux_inst_4_X ;
    wire KeyArray_MUX_inS02ser_mux_inst_5_Y ;
    wire KeyArray_MUX_inS02ser_mux_inst_5_X ;
    wire KeyArray_MUX_inS02ser_mux_inst_6_Y ;
    wire KeyArray_MUX_inS02ser_mux_inst_6_X ;
    wire KeyArray_MUX_inS02ser_mux_inst_7_Y ;
    wire KeyArray_MUX_inS02ser_mux_inst_7_X ;
    wire KeyArray_MUX_inS03ser_mux_inst_0_Y ;
    wire KeyArray_MUX_inS03ser_mux_inst_0_X ;
    wire KeyArray_MUX_inS03ser_mux_inst_1_Y ;
    wire KeyArray_MUX_inS03ser_mux_inst_1_X ;
    wire KeyArray_MUX_inS03ser_mux_inst_2_Y ;
    wire KeyArray_MUX_inS03ser_mux_inst_2_X ;
    wire KeyArray_MUX_inS03ser_mux_inst_3_Y ;
    wire KeyArray_MUX_inS03ser_mux_inst_3_X ;
    wire KeyArray_MUX_inS03ser_mux_inst_4_Y ;
    wire KeyArray_MUX_inS03ser_mux_inst_4_X ;
    wire KeyArray_MUX_inS03ser_mux_inst_5_Y ;
    wire KeyArray_MUX_inS03ser_mux_inst_5_X ;
    wire KeyArray_MUX_inS03ser_mux_inst_6_Y ;
    wire KeyArray_MUX_inS03ser_mux_inst_6_X ;
    wire KeyArray_MUX_inS03ser_mux_inst_7_Y ;
    wire KeyArray_MUX_inS03ser_mux_inst_7_X ;
    wire KeyArray_MUX_inS10ser_mux_inst_0_Y ;
    wire KeyArray_MUX_inS10ser_mux_inst_0_X ;
    wire KeyArray_MUX_inS10ser_mux_inst_1_Y ;
    wire KeyArray_MUX_inS10ser_mux_inst_1_X ;
    wire KeyArray_MUX_inS10ser_mux_inst_2_Y ;
    wire KeyArray_MUX_inS10ser_mux_inst_2_X ;
    wire KeyArray_MUX_inS10ser_mux_inst_3_Y ;
    wire KeyArray_MUX_inS10ser_mux_inst_3_X ;
    wire KeyArray_MUX_inS10ser_mux_inst_4_Y ;
    wire KeyArray_MUX_inS10ser_mux_inst_4_X ;
    wire KeyArray_MUX_inS10ser_mux_inst_5_Y ;
    wire KeyArray_MUX_inS10ser_mux_inst_5_X ;
    wire KeyArray_MUX_inS10ser_mux_inst_6_Y ;
    wire KeyArray_MUX_inS10ser_mux_inst_6_X ;
    wire KeyArray_MUX_inS10ser_mux_inst_7_Y ;
    wire KeyArray_MUX_inS10ser_mux_inst_7_X ;
    wire KeyArray_MUX_inS11ser_mux_inst_0_Y ;
    wire KeyArray_MUX_inS11ser_mux_inst_0_X ;
    wire KeyArray_MUX_inS11ser_mux_inst_1_Y ;
    wire KeyArray_MUX_inS11ser_mux_inst_1_X ;
    wire KeyArray_MUX_inS11ser_mux_inst_2_Y ;
    wire KeyArray_MUX_inS11ser_mux_inst_2_X ;
    wire KeyArray_MUX_inS11ser_mux_inst_3_Y ;
    wire KeyArray_MUX_inS11ser_mux_inst_3_X ;
    wire KeyArray_MUX_inS11ser_mux_inst_4_Y ;
    wire KeyArray_MUX_inS11ser_mux_inst_4_X ;
    wire KeyArray_MUX_inS11ser_mux_inst_5_Y ;
    wire KeyArray_MUX_inS11ser_mux_inst_5_X ;
    wire KeyArray_MUX_inS11ser_mux_inst_6_Y ;
    wire KeyArray_MUX_inS11ser_mux_inst_6_X ;
    wire KeyArray_MUX_inS11ser_mux_inst_7_Y ;
    wire KeyArray_MUX_inS11ser_mux_inst_7_X ;
    wire KeyArray_MUX_inS12ser_mux_inst_0_Y ;
    wire KeyArray_MUX_inS12ser_mux_inst_0_X ;
    wire KeyArray_MUX_inS12ser_mux_inst_1_Y ;
    wire KeyArray_MUX_inS12ser_mux_inst_1_X ;
    wire KeyArray_MUX_inS12ser_mux_inst_2_Y ;
    wire KeyArray_MUX_inS12ser_mux_inst_2_X ;
    wire KeyArray_MUX_inS12ser_mux_inst_3_Y ;
    wire KeyArray_MUX_inS12ser_mux_inst_3_X ;
    wire KeyArray_MUX_inS12ser_mux_inst_4_Y ;
    wire KeyArray_MUX_inS12ser_mux_inst_4_X ;
    wire KeyArray_MUX_inS12ser_mux_inst_5_Y ;
    wire KeyArray_MUX_inS12ser_mux_inst_5_X ;
    wire KeyArray_MUX_inS12ser_mux_inst_6_Y ;
    wire KeyArray_MUX_inS12ser_mux_inst_6_X ;
    wire KeyArray_MUX_inS12ser_mux_inst_7_Y ;
    wire KeyArray_MUX_inS12ser_mux_inst_7_X ;
    wire KeyArray_MUX_inS13ser_mux_inst_0_Y ;
    wire KeyArray_MUX_inS13ser_mux_inst_0_X ;
    wire KeyArray_MUX_inS13ser_mux_inst_1_Y ;
    wire KeyArray_MUX_inS13ser_mux_inst_1_X ;
    wire KeyArray_MUX_inS13ser_mux_inst_2_Y ;
    wire KeyArray_MUX_inS13ser_mux_inst_2_X ;
    wire KeyArray_MUX_inS13ser_mux_inst_3_Y ;
    wire KeyArray_MUX_inS13ser_mux_inst_3_X ;
    wire KeyArray_MUX_inS13ser_mux_inst_4_Y ;
    wire KeyArray_MUX_inS13ser_mux_inst_4_X ;
    wire KeyArray_MUX_inS13ser_mux_inst_5_Y ;
    wire KeyArray_MUX_inS13ser_mux_inst_5_X ;
    wire KeyArray_MUX_inS13ser_mux_inst_6_Y ;
    wire KeyArray_MUX_inS13ser_mux_inst_6_X ;
    wire KeyArray_MUX_inS13ser_mux_inst_7_Y ;
    wire KeyArray_MUX_inS13ser_mux_inst_7_X ;
    wire KeyArray_MUX_inS20ser_mux_inst_0_Y ;
    wire KeyArray_MUX_inS20ser_mux_inst_0_X ;
    wire KeyArray_MUX_inS20ser_mux_inst_1_Y ;
    wire KeyArray_MUX_inS20ser_mux_inst_1_X ;
    wire KeyArray_MUX_inS20ser_mux_inst_2_Y ;
    wire KeyArray_MUX_inS20ser_mux_inst_2_X ;
    wire KeyArray_MUX_inS20ser_mux_inst_3_Y ;
    wire KeyArray_MUX_inS20ser_mux_inst_3_X ;
    wire KeyArray_MUX_inS20ser_mux_inst_4_Y ;
    wire KeyArray_MUX_inS20ser_mux_inst_4_X ;
    wire KeyArray_MUX_inS20ser_mux_inst_5_Y ;
    wire KeyArray_MUX_inS20ser_mux_inst_5_X ;
    wire KeyArray_MUX_inS20ser_mux_inst_6_Y ;
    wire KeyArray_MUX_inS20ser_mux_inst_6_X ;
    wire KeyArray_MUX_inS20ser_mux_inst_7_Y ;
    wire KeyArray_MUX_inS20ser_mux_inst_7_X ;
    wire KeyArray_MUX_inS21ser_mux_inst_0_Y ;
    wire KeyArray_MUX_inS21ser_mux_inst_0_X ;
    wire KeyArray_MUX_inS21ser_mux_inst_1_Y ;
    wire KeyArray_MUX_inS21ser_mux_inst_1_X ;
    wire KeyArray_MUX_inS21ser_mux_inst_2_Y ;
    wire KeyArray_MUX_inS21ser_mux_inst_2_X ;
    wire KeyArray_MUX_inS21ser_mux_inst_3_Y ;
    wire KeyArray_MUX_inS21ser_mux_inst_3_X ;
    wire KeyArray_MUX_inS21ser_mux_inst_4_Y ;
    wire KeyArray_MUX_inS21ser_mux_inst_4_X ;
    wire KeyArray_MUX_inS21ser_mux_inst_5_Y ;
    wire KeyArray_MUX_inS21ser_mux_inst_5_X ;
    wire KeyArray_MUX_inS21ser_mux_inst_6_Y ;
    wire KeyArray_MUX_inS21ser_mux_inst_6_X ;
    wire KeyArray_MUX_inS21ser_mux_inst_7_Y ;
    wire KeyArray_MUX_inS21ser_mux_inst_7_X ;
    wire KeyArray_MUX_inS22ser_mux_inst_0_Y ;
    wire KeyArray_MUX_inS22ser_mux_inst_0_X ;
    wire KeyArray_MUX_inS22ser_mux_inst_1_Y ;
    wire KeyArray_MUX_inS22ser_mux_inst_1_X ;
    wire KeyArray_MUX_inS22ser_mux_inst_2_Y ;
    wire KeyArray_MUX_inS22ser_mux_inst_2_X ;
    wire KeyArray_MUX_inS22ser_mux_inst_3_Y ;
    wire KeyArray_MUX_inS22ser_mux_inst_3_X ;
    wire KeyArray_MUX_inS22ser_mux_inst_4_Y ;
    wire KeyArray_MUX_inS22ser_mux_inst_4_X ;
    wire KeyArray_MUX_inS22ser_mux_inst_5_Y ;
    wire KeyArray_MUX_inS22ser_mux_inst_5_X ;
    wire KeyArray_MUX_inS22ser_mux_inst_6_Y ;
    wire KeyArray_MUX_inS22ser_mux_inst_6_X ;
    wire KeyArray_MUX_inS22ser_mux_inst_7_Y ;
    wire KeyArray_MUX_inS22ser_mux_inst_7_X ;
    wire KeyArray_MUX_inS23ser_mux_inst_0_Y ;
    wire KeyArray_MUX_inS23ser_mux_inst_0_X ;
    wire KeyArray_MUX_inS23ser_mux_inst_1_Y ;
    wire KeyArray_MUX_inS23ser_mux_inst_1_X ;
    wire KeyArray_MUX_inS23ser_mux_inst_2_Y ;
    wire KeyArray_MUX_inS23ser_mux_inst_2_X ;
    wire KeyArray_MUX_inS23ser_mux_inst_3_Y ;
    wire KeyArray_MUX_inS23ser_mux_inst_3_X ;
    wire KeyArray_MUX_inS23ser_mux_inst_4_Y ;
    wire KeyArray_MUX_inS23ser_mux_inst_4_X ;
    wire KeyArray_MUX_inS23ser_mux_inst_5_Y ;
    wire KeyArray_MUX_inS23ser_mux_inst_5_X ;
    wire KeyArray_MUX_inS23ser_mux_inst_6_Y ;
    wire KeyArray_MUX_inS23ser_mux_inst_6_X ;
    wire KeyArray_MUX_inS23ser_mux_inst_7_Y ;
    wire KeyArray_MUX_inS23ser_mux_inst_7_X ;
    wire KeyArray_MUX_inS30ser_mux_inst_0_Y ;
    wire KeyArray_MUX_inS30ser_mux_inst_0_X ;
    wire KeyArray_MUX_inS30ser_mux_inst_1_Y ;
    wire KeyArray_MUX_inS30ser_mux_inst_1_X ;
    wire KeyArray_MUX_inS30ser_mux_inst_2_Y ;
    wire KeyArray_MUX_inS30ser_mux_inst_2_X ;
    wire KeyArray_MUX_inS30ser_mux_inst_3_Y ;
    wire KeyArray_MUX_inS30ser_mux_inst_3_X ;
    wire KeyArray_MUX_inS30ser_mux_inst_4_Y ;
    wire KeyArray_MUX_inS30ser_mux_inst_4_X ;
    wire KeyArray_MUX_inS30ser_mux_inst_5_Y ;
    wire KeyArray_MUX_inS30ser_mux_inst_5_X ;
    wire KeyArray_MUX_inS30ser_mux_inst_6_Y ;
    wire KeyArray_MUX_inS30ser_mux_inst_6_X ;
    wire KeyArray_MUX_inS30ser_mux_inst_7_Y ;
    wire KeyArray_MUX_inS30ser_mux_inst_7_X ;
    wire KeyArray_MUX_inS31ser_mux_inst_0_Y ;
    wire KeyArray_MUX_inS31ser_mux_inst_0_X ;
    wire KeyArray_MUX_inS31ser_mux_inst_1_Y ;
    wire KeyArray_MUX_inS31ser_mux_inst_1_X ;
    wire KeyArray_MUX_inS31ser_mux_inst_2_Y ;
    wire KeyArray_MUX_inS31ser_mux_inst_2_X ;
    wire KeyArray_MUX_inS31ser_mux_inst_3_Y ;
    wire KeyArray_MUX_inS31ser_mux_inst_3_X ;
    wire KeyArray_MUX_inS31ser_mux_inst_4_Y ;
    wire KeyArray_MUX_inS31ser_mux_inst_4_X ;
    wire KeyArray_MUX_inS31ser_mux_inst_5_Y ;
    wire KeyArray_MUX_inS31ser_mux_inst_5_X ;
    wire KeyArray_MUX_inS31ser_mux_inst_6_Y ;
    wire KeyArray_MUX_inS31ser_mux_inst_6_X ;
    wire KeyArray_MUX_inS31ser_mux_inst_7_Y ;
    wire KeyArray_MUX_inS31ser_mux_inst_7_X ;
    wire KeyArray_MUX_inS32ser_mux_inst_0_Y ;
    wire KeyArray_MUX_inS32ser_mux_inst_0_X ;
    wire KeyArray_MUX_inS32ser_mux_inst_1_Y ;
    wire KeyArray_MUX_inS32ser_mux_inst_1_X ;
    wire KeyArray_MUX_inS32ser_mux_inst_2_Y ;
    wire KeyArray_MUX_inS32ser_mux_inst_2_X ;
    wire KeyArray_MUX_inS32ser_mux_inst_3_Y ;
    wire KeyArray_MUX_inS32ser_mux_inst_3_X ;
    wire KeyArray_MUX_inS32ser_mux_inst_4_Y ;
    wire KeyArray_MUX_inS32ser_mux_inst_4_X ;
    wire KeyArray_MUX_inS32ser_mux_inst_5_Y ;
    wire KeyArray_MUX_inS32ser_mux_inst_5_X ;
    wire KeyArray_MUX_inS32ser_mux_inst_6_Y ;
    wire KeyArray_MUX_inS32ser_mux_inst_6_X ;
    wire KeyArray_MUX_inS32ser_mux_inst_7_Y ;
    wire KeyArray_MUX_inS32ser_mux_inst_7_X ;
    wire KeyArray_MUX_inS33ser_mux_inst_0_Y ;
    wire KeyArray_MUX_inS33ser_mux_inst_0_X ;
    wire KeyArray_MUX_inS33ser_mux_inst_1_Y ;
    wire KeyArray_MUX_inS33ser_mux_inst_1_X ;
    wire KeyArray_MUX_inS33ser_mux_inst_2_Y ;
    wire KeyArray_MUX_inS33ser_mux_inst_2_X ;
    wire KeyArray_MUX_inS33ser_mux_inst_3_Y ;
    wire KeyArray_MUX_inS33ser_mux_inst_3_X ;
    wire KeyArray_MUX_inS33ser_mux_inst_4_Y ;
    wire KeyArray_MUX_inS33ser_mux_inst_4_X ;
    wire KeyArray_MUX_inS33ser_mux_inst_5_Y ;
    wire KeyArray_MUX_inS33ser_mux_inst_5_X ;
    wire KeyArray_MUX_inS33ser_mux_inst_6_Y ;
    wire KeyArray_MUX_inS33ser_mux_inst_6_X ;
    wire KeyArray_MUX_inS33ser_mux_inst_7_Y ;
    wire KeyArray_MUX_inS33ser_mux_inst_7_X ;
    wire MixColumns_line0_n16 ;
    wire MixColumns_line0_n15 ;
    wire MixColumns_line0_n14 ;
    wire MixColumns_line0_n13 ;
    wire MixColumns_line0_n12 ;
    wire MixColumns_line0_n11 ;
    wire MixColumns_line0_n10 ;
    wire MixColumns_line0_n9 ;
    wire MixColumns_line0_n8 ;
    wire MixColumns_line0_n7 ;
    wire MixColumns_line0_n6 ;
    wire MixColumns_line0_n5 ;
    wire MixColumns_line0_n4 ;
    wire MixColumns_line0_n3 ;
    wire MixColumns_line0_n2 ;
    wire MixColumns_line0_n1 ;
    wire MixColumns_line1_n16 ;
    wire MixColumns_line1_n15 ;
    wire MixColumns_line1_n14 ;
    wire MixColumns_line1_n13 ;
    wire MixColumns_line1_n12 ;
    wire MixColumns_line1_n11 ;
    wire MixColumns_line1_n10 ;
    wire MixColumns_line1_n9 ;
    wire MixColumns_line1_n8 ;
    wire MixColumns_line1_n7 ;
    wire MixColumns_line1_n6 ;
    wire MixColumns_line1_n5 ;
    wire MixColumns_line1_n4 ;
    wire MixColumns_line1_n3 ;
    wire MixColumns_line1_n2 ;
    wire MixColumns_line1_n1 ;
    wire MixColumns_line1_S02_1_ ;
    wire MixColumns_line1_S02_3_ ;
    wire MixColumns_line1_S02_4_ ;
    wire MixColumns_line2_n16 ;
    wire MixColumns_line2_n15 ;
    wire MixColumns_line2_n14 ;
    wire MixColumns_line2_n13 ;
    wire MixColumns_line2_n12 ;
    wire MixColumns_line2_n11 ;
    wire MixColumns_line2_n10 ;
    wire MixColumns_line2_n9 ;
    wire MixColumns_line2_n8 ;
    wire MixColumns_line2_n7 ;
    wire MixColumns_line2_n6 ;
    wire MixColumns_line2_n5 ;
    wire MixColumns_line2_n4 ;
    wire MixColumns_line2_n3 ;
    wire MixColumns_line2_n2 ;
    wire MixColumns_line2_n1 ;
    wire MixColumns_line2_S02_1_ ;
    wire MixColumns_line2_S02_3_ ;
    wire MixColumns_line2_S02_4_ ;
    wire MixColumns_line3_n16 ;
    wire MixColumns_line3_n15 ;
    wire MixColumns_line3_n14 ;
    wire MixColumns_line3_n13 ;
    wire MixColumns_line3_n12 ;
    wire MixColumns_line3_n11 ;
    wire MixColumns_line3_n10 ;
    wire MixColumns_line3_n9 ;
    wire MixColumns_line3_n8 ;
    wire MixColumns_line3_n7 ;
    wire MixColumns_line3_n6 ;
    wire MixColumns_line3_n5 ;
    wire MixColumns_line3_n4 ;
    wire MixColumns_line3_n3 ;
    wire MixColumns_line3_n2 ;
    wire MixColumns_line3_n1 ;
    wire MixColumns_line3_S02_1_ ;
    wire MixColumns_line3_S02_3_ ;
    wire MixColumns_line3_S02_4_ ;
    wire MixColumns_line3_timesTHREE_input2_1_ ;
    wire MixColumns_line3_timesTHREE_input2_3_ ;
    wire MixColumns_line3_timesTHREE_input2_4_ ;
    wire calcRCon_n42 ;
    wire calcRCon_n41 ;
    wire calcRCon_n40 ;
    wire calcRCon_n39 ;
    wire calcRCon_n38 ;
    wire calcRCon_n37 ;
    wire calcRCon_n36 ;
    wire calcRCon_n35 ;
    wire calcRCon_n34 ;
    wire calcRCon_n33 ;
    wire calcRCon_n32 ;
    wire calcRCon_n31 ;
    wire calcRCon_n30 ;
    wire calcRCon_n29 ;
    wire calcRCon_n28 ;
    wire calcRCon_n27 ;
    wire calcRCon_n26 ;
    wire calcRCon_n25 ;
    wire calcRCon_n24 ;
    wire calcRCon_n23 ;
    wire calcRCon_n22 ;
    wire calcRCon_n21 ;
    wire calcRCon_n20 ;
    wire calcRCon_n19 ;
    wire calcRCon_n18 ;
    wire calcRCon_n17 ;
    wire calcRCon_n16 ;
    wire calcRCon_n15 ;
    wire calcRCon_n14 ;
    wire calcRCon_n13 ;
    wire calcRCon_n9 ;
    wire calcRCon_n8 ;
    wire calcRCon_n7 ;
    wire calcRCon_s_current_state_0_ ;
    wire calcRCon_s_current_state_1_ ;
    wire calcRCon_s_current_state_2_ ;
    wire calcRCon_s_current_state_3_ ;
    wire calcRCon_s_current_state_4_ ;
    wire calcRCon_s_current_state_5_ ;
    wire calcRCon_s_current_state_6_ ;
    wire calcRCon_s_current_state_7_ ;
    wire MUX_SboxIn_mux_inst_0_Y ;
    wire MUX_SboxIn_mux_inst_0_X ;
    wire MUX_SboxIn_mux_inst_1_Y ;
    wire MUX_SboxIn_mux_inst_1_X ;
    wire MUX_SboxIn_mux_inst_2_Y ;
    wire MUX_SboxIn_mux_inst_2_X ;
    wire MUX_SboxIn_mux_inst_3_Y ;
    wire MUX_SboxIn_mux_inst_3_X ;
    wire MUX_SboxIn_mux_inst_4_Y ;
    wire MUX_SboxIn_mux_inst_4_X ;
    wire MUX_SboxIn_mux_inst_5_Y ;
    wire MUX_SboxIn_mux_inst_5_X ;
    wire MUX_SboxIn_mux_inst_6_Y ;
    wire MUX_SboxIn_mux_inst_6_X ;
    wire MUX_SboxIn_mux_inst_7_Y ;
    wire MUX_SboxIn_mux_inst_7_X ;
    wire Inst_bSbox_L29 ;
    wire Inst_bSbox_L28 ;
    wire Inst_bSbox_L27 ;
    wire Inst_bSbox_L26 ;
    wire Inst_bSbox_L25 ;
    wire Inst_bSbox_L24 ;
    wire Inst_bSbox_L23 ;
    wire Inst_bSbox_L22 ;
    wire Inst_bSbox_L21 ;
    wire Inst_bSbox_L20 ;
    wire Inst_bSbox_L19 ;
    wire Inst_bSbox_L18 ;
    wire Inst_bSbox_L17 ;
    wire Inst_bSbox_L16 ;
    wire Inst_bSbox_L15 ;
    wire Inst_bSbox_L14 ;
    wire Inst_bSbox_L13 ;
    wire Inst_bSbox_L12 ;
    wire Inst_bSbox_L11 ;
    wire Inst_bSbox_L10 ;
    wire Inst_bSbox_L9 ;
    wire Inst_bSbox_L8 ;
    wire Inst_bSbox_L7 ;
    wire Inst_bSbox_L6 ;
    wire Inst_bSbox_L5 ;
    wire Inst_bSbox_L4 ;
    wire Inst_bSbox_L3 ;
    wire Inst_bSbox_L2 ;
    wire Inst_bSbox_L1 ;
    wire Inst_bSbox_L0 ;
    wire Inst_bSbox_M63 ;
    wire Inst_bSbox_M62 ;
    wire Inst_bSbox_M61 ;
    wire Inst_bSbox_M60 ;
    wire Inst_bSbox_M59 ;
    wire Inst_bSbox_M58 ;
    wire Inst_bSbox_M57 ;
    wire Inst_bSbox_M56 ;
    wire Inst_bSbox_M55 ;
    wire Inst_bSbox_M54 ;
    wire Inst_bSbox_M53 ;
    wire Inst_bSbox_M52 ;
    wire Inst_bSbox_M51 ;
    wire Inst_bSbox_M50 ;
    wire Inst_bSbox_M49 ;
    wire Inst_bSbox_M48 ;
    wire Inst_bSbox_M47 ;
    wire Inst_bSbox_M46 ;
    wire Inst_bSbox_M45 ;
    wire Inst_bSbox_M44 ;
    wire Inst_bSbox_M43 ;
    wire Inst_bSbox_M42 ;
    wire Inst_bSbox_M41 ;
    wire Inst_bSbox_M40 ;
    wire Inst_bSbox_M39 ;
    wire Inst_bSbox_M38 ;
    wire Inst_bSbox_M37 ;
    wire Inst_bSbox_M36 ;
    wire Inst_bSbox_M35 ;
    wire Inst_bSbox_M34 ;
    wire Inst_bSbox_M33 ;
    wire Inst_bSbox_M32 ;
    wire Inst_bSbox_M31 ;
    wire Inst_bSbox_M30 ;
    wire Inst_bSbox_M29 ;
    wire Inst_bSbox_M28 ;
    wire Inst_bSbox_M27 ;
    wire Inst_bSbox_M26 ;
    wire Inst_bSbox_M25 ;
    wire Inst_bSbox_M24 ;
    wire Inst_bSbox_M23 ;
    wire Inst_bSbox_M22 ;
    wire Inst_bSbox_M21 ;
    wire Inst_bSbox_M20 ;
    wire Inst_bSbox_M19 ;
    wire Inst_bSbox_M18 ;
    wire Inst_bSbox_M17 ;
    wire Inst_bSbox_M16 ;
    wire Inst_bSbox_M15 ;
    wire Inst_bSbox_M14 ;
    wire Inst_bSbox_M13 ;
    wire Inst_bSbox_M12 ;
    wire Inst_bSbox_M11 ;
    wire Inst_bSbox_M10 ;
    wire Inst_bSbox_M9 ;
    wire Inst_bSbox_M8 ;
    wire Inst_bSbox_M7 ;
    wire Inst_bSbox_M6 ;
    wire Inst_bSbox_M5 ;
    wire Inst_bSbox_M4 ;
    wire Inst_bSbox_M3 ;
    wire Inst_bSbox_M2 ;
    wire Inst_bSbox_M1 ;
    wire Inst_bSbox_T27 ;
    wire Inst_bSbox_T26 ;
    wire Inst_bSbox_T25 ;
    wire Inst_bSbox_T24 ;
    wire Inst_bSbox_T23 ;
    wire Inst_bSbox_T22 ;
    wire Inst_bSbox_T21 ;
    wire Inst_bSbox_T20 ;
    wire Inst_bSbox_T19 ;
    wire Inst_bSbox_T18 ;
    wire Inst_bSbox_T17 ;
    wire Inst_bSbox_T16 ;
    wire Inst_bSbox_T15 ;
    wire Inst_bSbox_T14 ;
    wire Inst_bSbox_T13 ;
    wire Inst_bSbox_T12 ;
    wire Inst_bSbox_T11 ;
    wire Inst_bSbox_T10 ;
    wire Inst_bSbox_T9 ;
    wire Inst_bSbox_T8 ;
    wire Inst_bSbox_T7 ;
    wire Inst_bSbox_T6 ;
    wire Inst_bSbox_T5 ;
    wire Inst_bSbox_T4 ;
    wire Inst_bSbox_T3 ;
    wire Inst_bSbox_T2 ;
    wire Inst_bSbox_T1 ;
    wire [7:0] SboxOut ;
    wire [7:0] StateOutXORroundKey ;
    wire [7:0] StateIn ;
    wire [31:0] StateInMC ;
    wire [31:0] MCout ;
    wire [7:0] keyStateIn ;
    wire [7:0] roundConstant ;
    wire [7:0] keySBIn ;
    wire [7:0] SboxIn ;
    wire [7:0] stateArray_input_MC ;
    wire [7:0] stateArray_outS30ser_MC ;
    wire [7:0] stateArray_outS20ser_MC ;
    wire [7:0] stateArray_outS10ser_MC ;
    wire [7:0] stateArray_inS33ser ;
    wire [7:0] stateArray_inS32ser ;
    wire [7:0] stateArray_inS31ser ;
    wire [7:0] stateArray_inS30ser ;
    wire [7:0] stateArray_inS23ser ;
    wire [7:0] stateArray_inS22ser ;
    wire [7:0] stateArray_inS21ser ;
    wire [7:0] stateArray_inS20ser ;
    wire [7:0] stateArray_inS13ser ;
    wire [7:0] stateArray_inS12ser ;
    wire [7:0] stateArray_inS11ser ;
    wire [7:0] stateArray_inS10ser ;
    wire [7:0] stateArray_inS03ser ;
    wire [7:0] stateArray_inS02ser ;
    wire [7:0] stateArray_inS01ser ;
    wire [7:0] stateArray_inS00ser ;
    wire [7:0] KeyArray_outS01ser_p ;
    wire [7:0] KeyArray_outS01ser_XOR_00 ;
    wire [7:0] KeyArray_outS33ser ;
    wire [7:0] KeyArray_inS33ser ;
    wire [7:0] KeyArray_outS32ser ;
    wire [7:0] KeyArray_inS32ser ;
    wire [7:0] KeyArray_outS31ser ;
    wire [7:0] KeyArray_inS31ser ;
    wire [7:0] KeyArray_outS30ser ;
    wire [7:0] KeyArray_inS30par ;
    wire [7:0] KeyArray_inS30ser ;
    wire [7:0] KeyArray_outS23ser ;
    wire [7:0] KeyArray_inS23ser ;
    wire [7:0] KeyArray_outS22ser ;
    wire [7:0] KeyArray_inS22ser ;
    wire [7:0] KeyArray_outS21ser ;
    wire [7:0] KeyArray_inS21ser ;
    wire [7:0] KeyArray_outS20ser ;
    wire [7:0] KeyArray_inS20ser ;
    wire [7:0] KeyArray_inS13ser ;
    wire [7:0] KeyArray_outS12ser ;
    wire [7:0] KeyArray_inS12ser ;
    wire [7:0] KeyArray_outS11ser ;
    wire [7:0] KeyArray_inS11ser ;
    wire [7:0] KeyArray_outS10ser ;
    wire [7:0] KeyArray_inS10ser ;
    wire [7:0] KeyArray_outS03ser ;
    wire [7:0] KeyArray_inS03ser ;
    wire [7:0] KeyArray_outS02ser ;
    wire [7:0] KeyArray_inS02ser ;
    wire [7:0] KeyArray_inS01ser ;
    wire [7:0] KeyArray_inS00ser ;
    wire [7:0] MixColumns_line0_S13 ;
    wire [4:1] MixColumns_line0_S02 ;
    wire [4:1] MixColumns_line0_timesTHREE_input2 ;
    wire [7:0] MixColumns_line1_S13 ;
    wire [4:1] MixColumns_line1_timesTHREE_input2 ;
    wire [7:0] MixColumns_line2_S13 ;
    wire [4:1] MixColumns_line2_timesTHREE_input2 ;
    wire [7:0] MixColumns_line3_S13 ;
    wire new_AGEMA_signal_3432 ;
    wire new_AGEMA_signal_3433 ;
    wire new_AGEMA_signal_3434 ;
    wire new_AGEMA_signal_3435 ;
    wire new_AGEMA_signal_3436 ;
    wire new_AGEMA_signal_3437 ;
    wire new_AGEMA_signal_3441 ;
    wire new_AGEMA_signal_3442 ;
    wire new_AGEMA_signal_3443 ;
    wire new_AGEMA_signal_3444 ;
    wire new_AGEMA_signal_3445 ;
    wire new_AGEMA_signal_3446 ;
    wire new_AGEMA_signal_3450 ;
    wire new_AGEMA_signal_3451 ;
    wire new_AGEMA_signal_3452 ;
    wire new_AGEMA_signal_3453 ;
    wire new_AGEMA_signal_3454 ;
    wire new_AGEMA_signal_3455 ;
    wire new_AGEMA_signal_3459 ;
    wire new_AGEMA_signal_3460 ;
    wire new_AGEMA_signal_3461 ;
    wire new_AGEMA_signal_3462 ;
    wire new_AGEMA_signal_3463 ;
    wire new_AGEMA_signal_3464 ;
    wire new_AGEMA_signal_3468 ;
    wire new_AGEMA_signal_3469 ;
    wire new_AGEMA_signal_3470 ;
    wire new_AGEMA_signal_3471 ;
    wire new_AGEMA_signal_3472 ;
    wire new_AGEMA_signal_3473 ;
    wire new_AGEMA_signal_3477 ;
    wire new_AGEMA_signal_3478 ;
    wire new_AGEMA_signal_3479 ;
    wire new_AGEMA_signal_3480 ;
    wire new_AGEMA_signal_3481 ;
    wire new_AGEMA_signal_3482 ;
    wire new_AGEMA_signal_3486 ;
    wire new_AGEMA_signal_3487 ;
    wire new_AGEMA_signal_3488 ;
    wire new_AGEMA_signal_3489 ;
    wire new_AGEMA_signal_3490 ;
    wire new_AGEMA_signal_3491 ;
    wire new_AGEMA_signal_3495 ;
    wire new_AGEMA_signal_3496 ;
    wire new_AGEMA_signal_3497 ;
    wire new_AGEMA_signal_3498 ;
    wire new_AGEMA_signal_3499 ;
    wire new_AGEMA_signal_3500 ;
    wire new_AGEMA_signal_3501 ;
    wire new_AGEMA_signal_3502 ;
    wire new_AGEMA_signal_3503 ;
    wire new_AGEMA_signal_3504 ;
    wire new_AGEMA_signal_3505 ;
    wire new_AGEMA_signal_3506 ;
    wire new_AGEMA_signal_3507 ;
    wire new_AGEMA_signal_3508 ;
    wire new_AGEMA_signal_3509 ;
    wire new_AGEMA_signal_3510 ;
    wire new_AGEMA_signal_3511 ;
    wire new_AGEMA_signal_3512 ;
    wire new_AGEMA_signal_3513 ;
    wire new_AGEMA_signal_3514 ;
    wire new_AGEMA_signal_3515 ;
    wire new_AGEMA_signal_3516 ;
    wire new_AGEMA_signal_3517 ;
    wire new_AGEMA_signal_3518 ;
    wire new_AGEMA_signal_3519 ;
    wire new_AGEMA_signal_3520 ;
    wire new_AGEMA_signal_3521 ;
    wire new_AGEMA_signal_3528 ;
    wire new_AGEMA_signal_3529 ;
    wire new_AGEMA_signal_3530 ;
    wire new_AGEMA_signal_3537 ;
    wire new_AGEMA_signal_3538 ;
    wire new_AGEMA_signal_3539 ;
    wire new_AGEMA_signal_3546 ;
    wire new_AGEMA_signal_3547 ;
    wire new_AGEMA_signal_3548 ;
    wire new_AGEMA_signal_3555 ;
    wire new_AGEMA_signal_3556 ;
    wire new_AGEMA_signal_3557 ;
    wire new_AGEMA_signal_3564 ;
    wire new_AGEMA_signal_3565 ;
    wire new_AGEMA_signal_3566 ;
    wire new_AGEMA_signal_3573 ;
    wire new_AGEMA_signal_3574 ;
    wire new_AGEMA_signal_3575 ;
    wire new_AGEMA_signal_3582 ;
    wire new_AGEMA_signal_3583 ;
    wire new_AGEMA_signal_3584 ;
    wire new_AGEMA_signal_3591 ;
    wire new_AGEMA_signal_3592 ;
    wire new_AGEMA_signal_3593 ;
    wire new_AGEMA_signal_3600 ;
    wire new_AGEMA_signal_3601 ;
    wire new_AGEMA_signal_3602 ;
    wire new_AGEMA_signal_3609 ;
    wire new_AGEMA_signal_3610 ;
    wire new_AGEMA_signal_3611 ;
    wire new_AGEMA_signal_3618 ;
    wire new_AGEMA_signal_3619 ;
    wire new_AGEMA_signal_3620 ;
    wire new_AGEMA_signal_3627 ;
    wire new_AGEMA_signal_3628 ;
    wire new_AGEMA_signal_3629 ;
    wire new_AGEMA_signal_3636 ;
    wire new_AGEMA_signal_3637 ;
    wire new_AGEMA_signal_3638 ;
    wire new_AGEMA_signal_3645 ;
    wire new_AGEMA_signal_3646 ;
    wire new_AGEMA_signal_3647 ;
    wire new_AGEMA_signal_3654 ;
    wire new_AGEMA_signal_3655 ;
    wire new_AGEMA_signal_3656 ;
    wire new_AGEMA_signal_3663 ;
    wire new_AGEMA_signal_3664 ;
    wire new_AGEMA_signal_3665 ;
    wire new_AGEMA_signal_3672 ;
    wire new_AGEMA_signal_3673 ;
    wire new_AGEMA_signal_3674 ;
    wire new_AGEMA_signal_3681 ;
    wire new_AGEMA_signal_3682 ;
    wire new_AGEMA_signal_3683 ;
    wire new_AGEMA_signal_3690 ;
    wire new_AGEMA_signal_3691 ;
    wire new_AGEMA_signal_3692 ;
    wire new_AGEMA_signal_3699 ;
    wire new_AGEMA_signal_3700 ;
    wire new_AGEMA_signal_3701 ;
    wire new_AGEMA_signal_3708 ;
    wire new_AGEMA_signal_3709 ;
    wire new_AGEMA_signal_3710 ;
    wire new_AGEMA_signal_3717 ;
    wire new_AGEMA_signal_3718 ;
    wire new_AGEMA_signal_3719 ;
    wire new_AGEMA_signal_3726 ;
    wire new_AGEMA_signal_3727 ;
    wire new_AGEMA_signal_3728 ;
    wire new_AGEMA_signal_3735 ;
    wire new_AGEMA_signal_3736 ;
    wire new_AGEMA_signal_3737 ;
    wire new_AGEMA_signal_3744 ;
    wire new_AGEMA_signal_3745 ;
    wire new_AGEMA_signal_3746 ;
    wire new_AGEMA_signal_3753 ;
    wire new_AGEMA_signal_3754 ;
    wire new_AGEMA_signal_3755 ;
    wire new_AGEMA_signal_3762 ;
    wire new_AGEMA_signal_3763 ;
    wire new_AGEMA_signal_3764 ;
    wire new_AGEMA_signal_3771 ;
    wire new_AGEMA_signal_3772 ;
    wire new_AGEMA_signal_3773 ;
    wire new_AGEMA_signal_3780 ;
    wire new_AGEMA_signal_3781 ;
    wire new_AGEMA_signal_3782 ;
    wire new_AGEMA_signal_3789 ;
    wire new_AGEMA_signal_3790 ;
    wire new_AGEMA_signal_3791 ;
    wire new_AGEMA_signal_3798 ;
    wire new_AGEMA_signal_3799 ;
    wire new_AGEMA_signal_3800 ;
    wire new_AGEMA_signal_3807 ;
    wire new_AGEMA_signal_3808 ;
    wire new_AGEMA_signal_3809 ;
    wire new_AGEMA_signal_3816 ;
    wire new_AGEMA_signal_3817 ;
    wire new_AGEMA_signal_3818 ;
    wire new_AGEMA_signal_3825 ;
    wire new_AGEMA_signal_3826 ;
    wire new_AGEMA_signal_3827 ;
    wire new_AGEMA_signal_3834 ;
    wire new_AGEMA_signal_3835 ;
    wire new_AGEMA_signal_3836 ;
    wire new_AGEMA_signal_3843 ;
    wire new_AGEMA_signal_3844 ;
    wire new_AGEMA_signal_3845 ;
    wire new_AGEMA_signal_3852 ;
    wire new_AGEMA_signal_3853 ;
    wire new_AGEMA_signal_3854 ;
    wire new_AGEMA_signal_3861 ;
    wire new_AGEMA_signal_3862 ;
    wire new_AGEMA_signal_3863 ;
    wire new_AGEMA_signal_3870 ;
    wire new_AGEMA_signal_3871 ;
    wire new_AGEMA_signal_3872 ;
    wire new_AGEMA_signal_3879 ;
    wire new_AGEMA_signal_3880 ;
    wire new_AGEMA_signal_3881 ;
    wire new_AGEMA_signal_3888 ;
    wire new_AGEMA_signal_3889 ;
    wire new_AGEMA_signal_3890 ;
    wire new_AGEMA_signal_3897 ;
    wire new_AGEMA_signal_3898 ;
    wire new_AGEMA_signal_3899 ;
    wire new_AGEMA_signal_3906 ;
    wire new_AGEMA_signal_3907 ;
    wire new_AGEMA_signal_3908 ;
    wire new_AGEMA_signal_3915 ;
    wire new_AGEMA_signal_3916 ;
    wire new_AGEMA_signal_3917 ;
    wire new_AGEMA_signal_3924 ;
    wire new_AGEMA_signal_3925 ;
    wire new_AGEMA_signal_3926 ;
    wire new_AGEMA_signal_3933 ;
    wire new_AGEMA_signal_3934 ;
    wire new_AGEMA_signal_3935 ;
    wire new_AGEMA_signal_3942 ;
    wire new_AGEMA_signal_3943 ;
    wire new_AGEMA_signal_3944 ;
    wire new_AGEMA_signal_3951 ;
    wire new_AGEMA_signal_3952 ;
    wire new_AGEMA_signal_3953 ;
    wire new_AGEMA_signal_3960 ;
    wire new_AGEMA_signal_3961 ;
    wire new_AGEMA_signal_3962 ;
    wire new_AGEMA_signal_3969 ;
    wire new_AGEMA_signal_3970 ;
    wire new_AGEMA_signal_3971 ;
    wire new_AGEMA_signal_3978 ;
    wire new_AGEMA_signal_3979 ;
    wire new_AGEMA_signal_3980 ;
    wire new_AGEMA_signal_3987 ;
    wire new_AGEMA_signal_3988 ;
    wire new_AGEMA_signal_3989 ;
    wire new_AGEMA_signal_3996 ;
    wire new_AGEMA_signal_3997 ;
    wire new_AGEMA_signal_3998 ;
    wire new_AGEMA_signal_4005 ;
    wire new_AGEMA_signal_4006 ;
    wire new_AGEMA_signal_4007 ;
    wire new_AGEMA_signal_4014 ;
    wire new_AGEMA_signal_4015 ;
    wire new_AGEMA_signal_4016 ;
    wire new_AGEMA_signal_4023 ;
    wire new_AGEMA_signal_4024 ;
    wire new_AGEMA_signal_4025 ;
    wire new_AGEMA_signal_4032 ;
    wire new_AGEMA_signal_4033 ;
    wire new_AGEMA_signal_4034 ;
    wire new_AGEMA_signal_4041 ;
    wire new_AGEMA_signal_4042 ;
    wire new_AGEMA_signal_4043 ;
    wire new_AGEMA_signal_4050 ;
    wire new_AGEMA_signal_4051 ;
    wire new_AGEMA_signal_4052 ;
    wire new_AGEMA_signal_4059 ;
    wire new_AGEMA_signal_4060 ;
    wire new_AGEMA_signal_4061 ;
    wire new_AGEMA_signal_4068 ;
    wire new_AGEMA_signal_4069 ;
    wire new_AGEMA_signal_4070 ;
    wire new_AGEMA_signal_4077 ;
    wire new_AGEMA_signal_4078 ;
    wire new_AGEMA_signal_4079 ;
    wire new_AGEMA_signal_4086 ;
    wire new_AGEMA_signal_4087 ;
    wire new_AGEMA_signal_4088 ;
    wire new_AGEMA_signal_4095 ;
    wire new_AGEMA_signal_4096 ;
    wire new_AGEMA_signal_4097 ;
    wire new_AGEMA_signal_4104 ;
    wire new_AGEMA_signal_4105 ;
    wire new_AGEMA_signal_4106 ;
    wire new_AGEMA_signal_4113 ;
    wire new_AGEMA_signal_4114 ;
    wire new_AGEMA_signal_4115 ;
    wire new_AGEMA_signal_4122 ;
    wire new_AGEMA_signal_4123 ;
    wire new_AGEMA_signal_4124 ;
    wire new_AGEMA_signal_4131 ;
    wire new_AGEMA_signal_4132 ;
    wire new_AGEMA_signal_4133 ;
    wire new_AGEMA_signal_4140 ;
    wire new_AGEMA_signal_4141 ;
    wire new_AGEMA_signal_4142 ;
    wire new_AGEMA_signal_4149 ;
    wire new_AGEMA_signal_4150 ;
    wire new_AGEMA_signal_4151 ;
    wire new_AGEMA_signal_4158 ;
    wire new_AGEMA_signal_4159 ;
    wire new_AGEMA_signal_4160 ;
    wire new_AGEMA_signal_4167 ;
    wire new_AGEMA_signal_4168 ;
    wire new_AGEMA_signal_4169 ;
    wire new_AGEMA_signal_4176 ;
    wire new_AGEMA_signal_4177 ;
    wire new_AGEMA_signal_4178 ;
    wire new_AGEMA_signal_4185 ;
    wire new_AGEMA_signal_4186 ;
    wire new_AGEMA_signal_4187 ;
    wire new_AGEMA_signal_4194 ;
    wire new_AGEMA_signal_4195 ;
    wire new_AGEMA_signal_4196 ;
    wire new_AGEMA_signal_4203 ;
    wire new_AGEMA_signal_4204 ;
    wire new_AGEMA_signal_4205 ;
    wire new_AGEMA_signal_4212 ;
    wire new_AGEMA_signal_4213 ;
    wire new_AGEMA_signal_4214 ;
    wire new_AGEMA_signal_4221 ;
    wire new_AGEMA_signal_4222 ;
    wire new_AGEMA_signal_4223 ;
    wire new_AGEMA_signal_4230 ;
    wire new_AGEMA_signal_4231 ;
    wire new_AGEMA_signal_4232 ;
    wire new_AGEMA_signal_4239 ;
    wire new_AGEMA_signal_4240 ;
    wire new_AGEMA_signal_4241 ;
    wire new_AGEMA_signal_4248 ;
    wire new_AGEMA_signal_4249 ;
    wire new_AGEMA_signal_4250 ;
    wire new_AGEMA_signal_4257 ;
    wire new_AGEMA_signal_4258 ;
    wire new_AGEMA_signal_4259 ;
    wire new_AGEMA_signal_4266 ;
    wire new_AGEMA_signal_4267 ;
    wire new_AGEMA_signal_4268 ;
    wire new_AGEMA_signal_4275 ;
    wire new_AGEMA_signal_4276 ;
    wire new_AGEMA_signal_4277 ;
    wire new_AGEMA_signal_4284 ;
    wire new_AGEMA_signal_4285 ;
    wire new_AGEMA_signal_4286 ;
    wire new_AGEMA_signal_4293 ;
    wire new_AGEMA_signal_4294 ;
    wire new_AGEMA_signal_4295 ;
    wire new_AGEMA_signal_4302 ;
    wire new_AGEMA_signal_4303 ;
    wire new_AGEMA_signal_4304 ;
    wire new_AGEMA_signal_4311 ;
    wire new_AGEMA_signal_4312 ;
    wire new_AGEMA_signal_4313 ;
    wire new_AGEMA_signal_4320 ;
    wire new_AGEMA_signal_4321 ;
    wire new_AGEMA_signal_4322 ;
    wire new_AGEMA_signal_4329 ;
    wire new_AGEMA_signal_4330 ;
    wire new_AGEMA_signal_4331 ;
    wire new_AGEMA_signal_4338 ;
    wire new_AGEMA_signal_4339 ;
    wire new_AGEMA_signal_4340 ;
    wire new_AGEMA_signal_4347 ;
    wire new_AGEMA_signal_4348 ;
    wire new_AGEMA_signal_4349 ;
    wire new_AGEMA_signal_4356 ;
    wire new_AGEMA_signal_4357 ;
    wire new_AGEMA_signal_4358 ;
    wire new_AGEMA_signal_4365 ;
    wire new_AGEMA_signal_4366 ;
    wire new_AGEMA_signal_4367 ;
    wire new_AGEMA_signal_4374 ;
    wire new_AGEMA_signal_4375 ;
    wire new_AGEMA_signal_4376 ;
    wire new_AGEMA_signal_4383 ;
    wire new_AGEMA_signal_4384 ;
    wire new_AGEMA_signal_4385 ;
    wire new_AGEMA_signal_4386 ;
    wire new_AGEMA_signal_4387 ;
    wire new_AGEMA_signal_4388 ;
    wire new_AGEMA_signal_4389 ;
    wire new_AGEMA_signal_4390 ;
    wire new_AGEMA_signal_4391 ;
    wire new_AGEMA_signal_4392 ;
    wire new_AGEMA_signal_4393 ;
    wire new_AGEMA_signal_4394 ;
    wire new_AGEMA_signal_4395 ;
    wire new_AGEMA_signal_4396 ;
    wire new_AGEMA_signal_4397 ;
    wire new_AGEMA_signal_4398 ;
    wire new_AGEMA_signal_4399 ;
    wire new_AGEMA_signal_4400 ;
    wire new_AGEMA_signal_4401 ;
    wire new_AGEMA_signal_4402 ;
    wire new_AGEMA_signal_4403 ;
    wire new_AGEMA_signal_4404 ;
    wire new_AGEMA_signal_4405 ;
    wire new_AGEMA_signal_4406 ;
    wire new_AGEMA_signal_4407 ;
    wire new_AGEMA_signal_4408 ;
    wire new_AGEMA_signal_4409 ;
    wire new_AGEMA_signal_4410 ;
    wire new_AGEMA_signal_4411 ;
    wire new_AGEMA_signal_4412 ;
    wire new_AGEMA_signal_4413 ;
    wire new_AGEMA_signal_4414 ;
    wire new_AGEMA_signal_4415 ;
    wire new_AGEMA_signal_4416 ;
    wire new_AGEMA_signal_4417 ;
    wire new_AGEMA_signal_4418 ;
    wire new_AGEMA_signal_4419 ;
    wire new_AGEMA_signal_4420 ;
    wire new_AGEMA_signal_4421 ;
    wire new_AGEMA_signal_4422 ;
    wire new_AGEMA_signal_4423 ;
    wire new_AGEMA_signal_4424 ;
    wire new_AGEMA_signal_4425 ;
    wire new_AGEMA_signal_4426 ;
    wire new_AGEMA_signal_4427 ;
    wire new_AGEMA_signal_4428 ;
    wire new_AGEMA_signal_4429 ;
    wire new_AGEMA_signal_4430 ;
    wire new_AGEMA_signal_4431 ;
    wire new_AGEMA_signal_4432 ;
    wire new_AGEMA_signal_4433 ;
    wire new_AGEMA_signal_4437 ;
    wire new_AGEMA_signal_4438 ;
    wire new_AGEMA_signal_4439 ;
    wire new_AGEMA_signal_4440 ;
    wire new_AGEMA_signal_4441 ;
    wire new_AGEMA_signal_4442 ;
    wire new_AGEMA_signal_4446 ;
    wire new_AGEMA_signal_4447 ;
    wire new_AGEMA_signal_4448 ;
    wire new_AGEMA_signal_4449 ;
    wire new_AGEMA_signal_4450 ;
    wire new_AGEMA_signal_4451 ;
    wire new_AGEMA_signal_4455 ;
    wire new_AGEMA_signal_4456 ;
    wire new_AGEMA_signal_4457 ;
    wire new_AGEMA_signal_4458 ;
    wire new_AGEMA_signal_4459 ;
    wire new_AGEMA_signal_4460 ;
    wire new_AGEMA_signal_4464 ;
    wire new_AGEMA_signal_4465 ;
    wire new_AGEMA_signal_4466 ;
    wire new_AGEMA_signal_4467 ;
    wire new_AGEMA_signal_4468 ;
    wire new_AGEMA_signal_4469 ;
    wire new_AGEMA_signal_4473 ;
    wire new_AGEMA_signal_4474 ;
    wire new_AGEMA_signal_4475 ;
    wire new_AGEMA_signal_4476 ;
    wire new_AGEMA_signal_4477 ;
    wire new_AGEMA_signal_4478 ;
    wire new_AGEMA_signal_4482 ;
    wire new_AGEMA_signal_4483 ;
    wire new_AGEMA_signal_4484 ;
    wire new_AGEMA_signal_4485 ;
    wire new_AGEMA_signal_4486 ;
    wire new_AGEMA_signal_4487 ;
    wire new_AGEMA_signal_4491 ;
    wire new_AGEMA_signal_4492 ;
    wire new_AGEMA_signal_4493 ;
    wire new_AGEMA_signal_4494 ;
    wire new_AGEMA_signal_4495 ;
    wire new_AGEMA_signal_4496 ;
    wire new_AGEMA_signal_4500 ;
    wire new_AGEMA_signal_4501 ;
    wire new_AGEMA_signal_4502 ;
    wire new_AGEMA_signal_4503 ;
    wire new_AGEMA_signal_4504 ;
    wire new_AGEMA_signal_4505 ;
    wire new_AGEMA_signal_4509 ;
    wire new_AGEMA_signal_4510 ;
    wire new_AGEMA_signal_4511 ;
    wire new_AGEMA_signal_4512 ;
    wire new_AGEMA_signal_4513 ;
    wire new_AGEMA_signal_4514 ;
    wire new_AGEMA_signal_4518 ;
    wire new_AGEMA_signal_4519 ;
    wire new_AGEMA_signal_4520 ;
    wire new_AGEMA_signal_4521 ;
    wire new_AGEMA_signal_4522 ;
    wire new_AGEMA_signal_4523 ;
    wire new_AGEMA_signal_4527 ;
    wire new_AGEMA_signal_4528 ;
    wire new_AGEMA_signal_4529 ;
    wire new_AGEMA_signal_4530 ;
    wire new_AGEMA_signal_4531 ;
    wire new_AGEMA_signal_4532 ;
    wire new_AGEMA_signal_4536 ;
    wire new_AGEMA_signal_4537 ;
    wire new_AGEMA_signal_4538 ;
    wire new_AGEMA_signal_4539 ;
    wire new_AGEMA_signal_4540 ;
    wire new_AGEMA_signal_4541 ;
    wire new_AGEMA_signal_4545 ;
    wire new_AGEMA_signal_4546 ;
    wire new_AGEMA_signal_4547 ;
    wire new_AGEMA_signal_4548 ;
    wire new_AGEMA_signal_4549 ;
    wire new_AGEMA_signal_4550 ;
    wire new_AGEMA_signal_4554 ;
    wire new_AGEMA_signal_4555 ;
    wire new_AGEMA_signal_4556 ;
    wire new_AGEMA_signal_4557 ;
    wire new_AGEMA_signal_4558 ;
    wire new_AGEMA_signal_4559 ;
    wire new_AGEMA_signal_4563 ;
    wire new_AGEMA_signal_4564 ;
    wire new_AGEMA_signal_4565 ;
    wire new_AGEMA_signal_4566 ;
    wire new_AGEMA_signal_4567 ;
    wire new_AGEMA_signal_4568 ;
    wire new_AGEMA_signal_4572 ;
    wire new_AGEMA_signal_4573 ;
    wire new_AGEMA_signal_4574 ;
    wire new_AGEMA_signal_4575 ;
    wire new_AGEMA_signal_4576 ;
    wire new_AGEMA_signal_4577 ;
    wire new_AGEMA_signal_4581 ;
    wire new_AGEMA_signal_4582 ;
    wire new_AGEMA_signal_4583 ;
    wire new_AGEMA_signal_4584 ;
    wire new_AGEMA_signal_4585 ;
    wire new_AGEMA_signal_4586 ;
    wire new_AGEMA_signal_4590 ;
    wire new_AGEMA_signal_4591 ;
    wire new_AGEMA_signal_4592 ;
    wire new_AGEMA_signal_4593 ;
    wire new_AGEMA_signal_4594 ;
    wire new_AGEMA_signal_4595 ;
    wire new_AGEMA_signal_4599 ;
    wire new_AGEMA_signal_4600 ;
    wire new_AGEMA_signal_4601 ;
    wire new_AGEMA_signal_4602 ;
    wire new_AGEMA_signal_4603 ;
    wire new_AGEMA_signal_4604 ;
    wire new_AGEMA_signal_4608 ;
    wire new_AGEMA_signal_4609 ;
    wire new_AGEMA_signal_4610 ;
    wire new_AGEMA_signal_4611 ;
    wire new_AGEMA_signal_4612 ;
    wire new_AGEMA_signal_4613 ;
    wire new_AGEMA_signal_4617 ;
    wire new_AGEMA_signal_4618 ;
    wire new_AGEMA_signal_4619 ;
    wire new_AGEMA_signal_4620 ;
    wire new_AGEMA_signal_4621 ;
    wire new_AGEMA_signal_4622 ;
    wire new_AGEMA_signal_4626 ;
    wire new_AGEMA_signal_4627 ;
    wire new_AGEMA_signal_4628 ;
    wire new_AGEMA_signal_4629 ;
    wire new_AGEMA_signal_4630 ;
    wire new_AGEMA_signal_4631 ;
    wire new_AGEMA_signal_4635 ;
    wire new_AGEMA_signal_4636 ;
    wire new_AGEMA_signal_4637 ;
    wire new_AGEMA_signal_4638 ;
    wire new_AGEMA_signal_4639 ;
    wire new_AGEMA_signal_4640 ;
    wire new_AGEMA_signal_4644 ;
    wire new_AGEMA_signal_4645 ;
    wire new_AGEMA_signal_4646 ;
    wire new_AGEMA_signal_4647 ;
    wire new_AGEMA_signal_4648 ;
    wire new_AGEMA_signal_4649 ;
    wire new_AGEMA_signal_4653 ;
    wire new_AGEMA_signal_4654 ;
    wire new_AGEMA_signal_4655 ;
    wire new_AGEMA_signal_4656 ;
    wire new_AGEMA_signal_4657 ;
    wire new_AGEMA_signal_4658 ;
    wire new_AGEMA_signal_4662 ;
    wire new_AGEMA_signal_4663 ;
    wire new_AGEMA_signal_4664 ;
    wire new_AGEMA_signal_4665 ;
    wire new_AGEMA_signal_4666 ;
    wire new_AGEMA_signal_4667 ;
    wire new_AGEMA_signal_4671 ;
    wire new_AGEMA_signal_4672 ;
    wire new_AGEMA_signal_4673 ;
    wire new_AGEMA_signal_4674 ;
    wire new_AGEMA_signal_4675 ;
    wire new_AGEMA_signal_4676 ;
    wire new_AGEMA_signal_4680 ;
    wire new_AGEMA_signal_4681 ;
    wire new_AGEMA_signal_4682 ;
    wire new_AGEMA_signal_4683 ;
    wire new_AGEMA_signal_4684 ;
    wire new_AGEMA_signal_4685 ;
    wire new_AGEMA_signal_4689 ;
    wire new_AGEMA_signal_4690 ;
    wire new_AGEMA_signal_4691 ;
    wire new_AGEMA_signal_4692 ;
    wire new_AGEMA_signal_4693 ;
    wire new_AGEMA_signal_4694 ;
    wire new_AGEMA_signal_4698 ;
    wire new_AGEMA_signal_4699 ;
    wire new_AGEMA_signal_4700 ;
    wire new_AGEMA_signal_4701 ;
    wire new_AGEMA_signal_4702 ;
    wire new_AGEMA_signal_4703 ;
    wire new_AGEMA_signal_4707 ;
    wire new_AGEMA_signal_4708 ;
    wire new_AGEMA_signal_4709 ;
    wire new_AGEMA_signal_4710 ;
    wire new_AGEMA_signal_4711 ;
    wire new_AGEMA_signal_4712 ;
    wire new_AGEMA_signal_4716 ;
    wire new_AGEMA_signal_4717 ;
    wire new_AGEMA_signal_4718 ;
    wire new_AGEMA_signal_4719 ;
    wire new_AGEMA_signal_4720 ;
    wire new_AGEMA_signal_4721 ;
    wire new_AGEMA_signal_4725 ;
    wire new_AGEMA_signal_4726 ;
    wire new_AGEMA_signal_4727 ;
    wire new_AGEMA_signal_4728 ;
    wire new_AGEMA_signal_4729 ;
    wire new_AGEMA_signal_4730 ;
    wire new_AGEMA_signal_4734 ;
    wire new_AGEMA_signal_4735 ;
    wire new_AGEMA_signal_4736 ;
    wire new_AGEMA_signal_4737 ;
    wire new_AGEMA_signal_4738 ;
    wire new_AGEMA_signal_4739 ;
    wire new_AGEMA_signal_4743 ;
    wire new_AGEMA_signal_4744 ;
    wire new_AGEMA_signal_4745 ;
    wire new_AGEMA_signal_4746 ;
    wire new_AGEMA_signal_4747 ;
    wire new_AGEMA_signal_4748 ;
    wire new_AGEMA_signal_4752 ;
    wire new_AGEMA_signal_4753 ;
    wire new_AGEMA_signal_4754 ;
    wire new_AGEMA_signal_4755 ;
    wire new_AGEMA_signal_4756 ;
    wire new_AGEMA_signal_4757 ;
    wire new_AGEMA_signal_4761 ;
    wire new_AGEMA_signal_4762 ;
    wire new_AGEMA_signal_4763 ;
    wire new_AGEMA_signal_4764 ;
    wire new_AGEMA_signal_4765 ;
    wire new_AGEMA_signal_4766 ;
    wire new_AGEMA_signal_4770 ;
    wire new_AGEMA_signal_4771 ;
    wire new_AGEMA_signal_4772 ;
    wire new_AGEMA_signal_4773 ;
    wire new_AGEMA_signal_4774 ;
    wire new_AGEMA_signal_4775 ;
    wire new_AGEMA_signal_4779 ;
    wire new_AGEMA_signal_4780 ;
    wire new_AGEMA_signal_4781 ;
    wire new_AGEMA_signal_4782 ;
    wire new_AGEMA_signal_4783 ;
    wire new_AGEMA_signal_4784 ;
    wire new_AGEMA_signal_4788 ;
    wire new_AGEMA_signal_4789 ;
    wire new_AGEMA_signal_4790 ;
    wire new_AGEMA_signal_4791 ;
    wire new_AGEMA_signal_4792 ;
    wire new_AGEMA_signal_4793 ;
    wire new_AGEMA_signal_4797 ;
    wire new_AGEMA_signal_4798 ;
    wire new_AGEMA_signal_4799 ;
    wire new_AGEMA_signal_4800 ;
    wire new_AGEMA_signal_4801 ;
    wire new_AGEMA_signal_4802 ;
    wire new_AGEMA_signal_4806 ;
    wire new_AGEMA_signal_4807 ;
    wire new_AGEMA_signal_4808 ;
    wire new_AGEMA_signal_4809 ;
    wire new_AGEMA_signal_4810 ;
    wire new_AGEMA_signal_4811 ;
    wire new_AGEMA_signal_4815 ;
    wire new_AGEMA_signal_4816 ;
    wire new_AGEMA_signal_4817 ;
    wire new_AGEMA_signal_4818 ;
    wire new_AGEMA_signal_4819 ;
    wire new_AGEMA_signal_4820 ;
    wire new_AGEMA_signal_4824 ;
    wire new_AGEMA_signal_4825 ;
    wire new_AGEMA_signal_4826 ;
    wire new_AGEMA_signal_4827 ;
    wire new_AGEMA_signal_4828 ;
    wire new_AGEMA_signal_4829 ;
    wire new_AGEMA_signal_4833 ;
    wire new_AGEMA_signal_4834 ;
    wire new_AGEMA_signal_4835 ;
    wire new_AGEMA_signal_4836 ;
    wire new_AGEMA_signal_4837 ;
    wire new_AGEMA_signal_4838 ;
    wire new_AGEMA_signal_4842 ;
    wire new_AGEMA_signal_4843 ;
    wire new_AGEMA_signal_4844 ;
    wire new_AGEMA_signal_4845 ;
    wire new_AGEMA_signal_4846 ;
    wire new_AGEMA_signal_4847 ;
    wire new_AGEMA_signal_4851 ;
    wire new_AGEMA_signal_4852 ;
    wire new_AGEMA_signal_4853 ;
    wire new_AGEMA_signal_4854 ;
    wire new_AGEMA_signal_4855 ;
    wire new_AGEMA_signal_4856 ;
    wire new_AGEMA_signal_4860 ;
    wire new_AGEMA_signal_4861 ;
    wire new_AGEMA_signal_4862 ;
    wire new_AGEMA_signal_4863 ;
    wire new_AGEMA_signal_4864 ;
    wire new_AGEMA_signal_4865 ;
    wire new_AGEMA_signal_4869 ;
    wire new_AGEMA_signal_4870 ;
    wire new_AGEMA_signal_4871 ;
    wire new_AGEMA_signal_4872 ;
    wire new_AGEMA_signal_4873 ;
    wire new_AGEMA_signal_4874 ;
    wire new_AGEMA_signal_4878 ;
    wire new_AGEMA_signal_4879 ;
    wire new_AGEMA_signal_4880 ;
    wire new_AGEMA_signal_4881 ;
    wire new_AGEMA_signal_4882 ;
    wire new_AGEMA_signal_4883 ;
    wire new_AGEMA_signal_4887 ;
    wire new_AGEMA_signal_4888 ;
    wire new_AGEMA_signal_4889 ;
    wire new_AGEMA_signal_4890 ;
    wire new_AGEMA_signal_4891 ;
    wire new_AGEMA_signal_4892 ;
    wire new_AGEMA_signal_4896 ;
    wire new_AGEMA_signal_4897 ;
    wire new_AGEMA_signal_4898 ;
    wire new_AGEMA_signal_4899 ;
    wire new_AGEMA_signal_4900 ;
    wire new_AGEMA_signal_4901 ;
    wire new_AGEMA_signal_4905 ;
    wire new_AGEMA_signal_4906 ;
    wire new_AGEMA_signal_4907 ;
    wire new_AGEMA_signal_4908 ;
    wire new_AGEMA_signal_4909 ;
    wire new_AGEMA_signal_4910 ;
    wire new_AGEMA_signal_4914 ;
    wire new_AGEMA_signal_4915 ;
    wire new_AGEMA_signal_4916 ;
    wire new_AGEMA_signal_4917 ;
    wire new_AGEMA_signal_4918 ;
    wire new_AGEMA_signal_4919 ;
    wire new_AGEMA_signal_4923 ;
    wire new_AGEMA_signal_4924 ;
    wire new_AGEMA_signal_4925 ;
    wire new_AGEMA_signal_4926 ;
    wire new_AGEMA_signal_4927 ;
    wire new_AGEMA_signal_4928 ;
    wire new_AGEMA_signal_4932 ;
    wire new_AGEMA_signal_4933 ;
    wire new_AGEMA_signal_4934 ;
    wire new_AGEMA_signal_4935 ;
    wire new_AGEMA_signal_4936 ;
    wire new_AGEMA_signal_4937 ;
    wire new_AGEMA_signal_4941 ;
    wire new_AGEMA_signal_4942 ;
    wire new_AGEMA_signal_4943 ;
    wire new_AGEMA_signal_4944 ;
    wire new_AGEMA_signal_4945 ;
    wire new_AGEMA_signal_4946 ;
    wire new_AGEMA_signal_4950 ;
    wire new_AGEMA_signal_4951 ;
    wire new_AGEMA_signal_4952 ;
    wire new_AGEMA_signal_4953 ;
    wire new_AGEMA_signal_4954 ;
    wire new_AGEMA_signal_4955 ;
    wire new_AGEMA_signal_4959 ;
    wire new_AGEMA_signal_4960 ;
    wire new_AGEMA_signal_4961 ;
    wire new_AGEMA_signal_4962 ;
    wire new_AGEMA_signal_4963 ;
    wire new_AGEMA_signal_4964 ;
    wire new_AGEMA_signal_4968 ;
    wire new_AGEMA_signal_4969 ;
    wire new_AGEMA_signal_4970 ;
    wire new_AGEMA_signal_4971 ;
    wire new_AGEMA_signal_4972 ;
    wire new_AGEMA_signal_4973 ;
    wire new_AGEMA_signal_4977 ;
    wire new_AGEMA_signal_4978 ;
    wire new_AGEMA_signal_4979 ;
    wire new_AGEMA_signal_4980 ;
    wire new_AGEMA_signal_4981 ;
    wire new_AGEMA_signal_4982 ;
    wire new_AGEMA_signal_4986 ;
    wire new_AGEMA_signal_4987 ;
    wire new_AGEMA_signal_4988 ;
    wire new_AGEMA_signal_4989 ;
    wire new_AGEMA_signal_4990 ;
    wire new_AGEMA_signal_4991 ;
    wire new_AGEMA_signal_4995 ;
    wire new_AGEMA_signal_4996 ;
    wire new_AGEMA_signal_4997 ;
    wire new_AGEMA_signal_4998 ;
    wire new_AGEMA_signal_4999 ;
    wire new_AGEMA_signal_5000 ;
    wire new_AGEMA_signal_5004 ;
    wire new_AGEMA_signal_5005 ;
    wire new_AGEMA_signal_5006 ;
    wire new_AGEMA_signal_5007 ;
    wire new_AGEMA_signal_5008 ;
    wire new_AGEMA_signal_5009 ;
    wire new_AGEMA_signal_5013 ;
    wire new_AGEMA_signal_5014 ;
    wire new_AGEMA_signal_5015 ;
    wire new_AGEMA_signal_5016 ;
    wire new_AGEMA_signal_5017 ;
    wire new_AGEMA_signal_5018 ;
    wire new_AGEMA_signal_5022 ;
    wire new_AGEMA_signal_5023 ;
    wire new_AGEMA_signal_5024 ;
    wire new_AGEMA_signal_5025 ;
    wire new_AGEMA_signal_5026 ;
    wire new_AGEMA_signal_5027 ;
    wire new_AGEMA_signal_5031 ;
    wire new_AGEMA_signal_5032 ;
    wire new_AGEMA_signal_5033 ;
    wire new_AGEMA_signal_5034 ;
    wire new_AGEMA_signal_5035 ;
    wire new_AGEMA_signal_5036 ;
    wire new_AGEMA_signal_5040 ;
    wire new_AGEMA_signal_5041 ;
    wire new_AGEMA_signal_5042 ;
    wire new_AGEMA_signal_5043 ;
    wire new_AGEMA_signal_5044 ;
    wire new_AGEMA_signal_5045 ;
    wire new_AGEMA_signal_5049 ;
    wire new_AGEMA_signal_5050 ;
    wire new_AGEMA_signal_5051 ;
    wire new_AGEMA_signal_5052 ;
    wire new_AGEMA_signal_5053 ;
    wire new_AGEMA_signal_5054 ;
    wire new_AGEMA_signal_5058 ;
    wire new_AGEMA_signal_5059 ;
    wire new_AGEMA_signal_5060 ;
    wire new_AGEMA_signal_5061 ;
    wire new_AGEMA_signal_5062 ;
    wire new_AGEMA_signal_5063 ;
    wire new_AGEMA_signal_5067 ;
    wire new_AGEMA_signal_5068 ;
    wire new_AGEMA_signal_5069 ;
    wire new_AGEMA_signal_5070 ;
    wire new_AGEMA_signal_5071 ;
    wire new_AGEMA_signal_5072 ;
    wire new_AGEMA_signal_5076 ;
    wire new_AGEMA_signal_5077 ;
    wire new_AGEMA_signal_5078 ;
    wire new_AGEMA_signal_5079 ;
    wire new_AGEMA_signal_5080 ;
    wire new_AGEMA_signal_5081 ;
    wire new_AGEMA_signal_5085 ;
    wire new_AGEMA_signal_5086 ;
    wire new_AGEMA_signal_5087 ;
    wire new_AGEMA_signal_5088 ;
    wire new_AGEMA_signal_5089 ;
    wire new_AGEMA_signal_5090 ;
    wire new_AGEMA_signal_5094 ;
    wire new_AGEMA_signal_5095 ;
    wire new_AGEMA_signal_5096 ;
    wire new_AGEMA_signal_5097 ;
    wire new_AGEMA_signal_5098 ;
    wire new_AGEMA_signal_5099 ;
    wire new_AGEMA_signal_5103 ;
    wire new_AGEMA_signal_5104 ;
    wire new_AGEMA_signal_5105 ;
    wire new_AGEMA_signal_5106 ;
    wire new_AGEMA_signal_5107 ;
    wire new_AGEMA_signal_5108 ;
    wire new_AGEMA_signal_5112 ;
    wire new_AGEMA_signal_5113 ;
    wire new_AGEMA_signal_5114 ;
    wire new_AGEMA_signal_5115 ;
    wire new_AGEMA_signal_5116 ;
    wire new_AGEMA_signal_5117 ;
    wire new_AGEMA_signal_5121 ;
    wire new_AGEMA_signal_5122 ;
    wire new_AGEMA_signal_5123 ;
    wire new_AGEMA_signal_5124 ;
    wire new_AGEMA_signal_5125 ;
    wire new_AGEMA_signal_5126 ;
    wire new_AGEMA_signal_5130 ;
    wire new_AGEMA_signal_5131 ;
    wire new_AGEMA_signal_5132 ;
    wire new_AGEMA_signal_5133 ;
    wire new_AGEMA_signal_5134 ;
    wire new_AGEMA_signal_5135 ;
    wire new_AGEMA_signal_5139 ;
    wire new_AGEMA_signal_5140 ;
    wire new_AGEMA_signal_5141 ;
    wire new_AGEMA_signal_5142 ;
    wire new_AGEMA_signal_5143 ;
    wire new_AGEMA_signal_5144 ;
    wire new_AGEMA_signal_5148 ;
    wire new_AGEMA_signal_5149 ;
    wire new_AGEMA_signal_5150 ;
    wire new_AGEMA_signal_5151 ;
    wire new_AGEMA_signal_5152 ;
    wire new_AGEMA_signal_5153 ;
    wire new_AGEMA_signal_5157 ;
    wire new_AGEMA_signal_5158 ;
    wire new_AGEMA_signal_5159 ;
    wire new_AGEMA_signal_5160 ;
    wire new_AGEMA_signal_5161 ;
    wire new_AGEMA_signal_5162 ;
    wire new_AGEMA_signal_5166 ;
    wire new_AGEMA_signal_5167 ;
    wire new_AGEMA_signal_5168 ;
    wire new_AGEMA_signal_5169 ;
    wire new_AGEMA_signal_5170 ;
    wire new_AGEMA_signal_5171 ;
    wire new_AGEMA_signal_5175 ;
    wire new_AGEMA_signal_5176 ;
    wire new_AGEMA_signal_5177 ;
    wire new_AGEMA_signal_5178 ;
    wire new_AGEMA_signal_5179 ;
    wire new_AGEMA_signal_5180 ;
    wire new_AGEMA_signal_5184 ;
    wire new_AGEMA_signal_5185 ;
    wire new_AGEMA_signal_5186 ;
    wire new_AGEMA_signal_5187 ;
    wire new_AGEMA_signal_5188 ;
    wire new_AGEMA_signal_5189 ;
    wire new_AGEMA_signal_5193 ;
    wire new_AGEMA_signal_5194 ;
    wire new_AGEMA_signal_5195 ;
    wire new_AGEMA_signal_5196 ;
    wire new_AGEMA_signal_5197 ;
    wire new_AGEMA_signal_5198 ;
    wire new_AGEMA_signal_5202 ;
    wire new_AGEMA_signal_5203 ;
    wire new_AGEMA_signal_5204 ;
    wire new_AGEMA_signal_5205 ;
    wire new_AGEMA_signal_5206 ;
    wire new_AGEMA_signal_5207 ;
    wire new_AGEMA_signal_5211 ;
    wire new_AGEMA_signal_5212 ;
    wire new_AGEMA_signal_5213 ;
    wire new_AGEMA_signal_5214 ;
    wire new_AGEMA_signal_5215 ;
    wire new_AGEMA_signal_5216 ;
    wire new_AGEMA_signal_5220 ;
    wire new_AGEMA_signal_5221 ;
    wire new_AGEMA_signal_5222 ;
    wire new_AGEMA_signal_5223 ;
    wire new_AGEMA_signal_5224 ;
    wire new_AGEMA_signal_5225 ;
    wire new_AGEMA_signal_5229 ;
    wire new_AGEMA_signal_5230 ;
    wire new_AGEMA_signal_5231 ;
    wire new_AGEMA_signal_5232 ;
    wire new_AGEMA_signal_5233 ;
    wire new_AGEMA_signal_5234 ;
    wire new_AGEMA_signal_5238 ;
    wire new_AGEMA_signal_5239 ;
    wire new_AGEMA_signal_5240 ;
    wire new_AGEMA_signal_5241 ;
    wire new_AGEMA_signal_5242 ;
    wire new_AGEMA_signal_5243 ;
    wire new_AGEMA_signal_5247 ;
    wire new_AGEMA_signal_5248 ;
    wire new_AGEMA_signal_5249 ;
    wire new_AGEMA_signal_5250 ;
    wire new_AGEMA_signal_5251 ;
    wire new_AGEMA_signal_5252 ;
    wire new_AGEMA_signal_5256 ;
    wire new_AGEMA_signal_5257 ;
    wire new_AGEMA_signal_5258 ;
    wire new_AGEMA_signal_5259 ;
    wire new_AGEMA_signal_5260 ;
    wire new_AGEMA_signal_5261 ;
    wire new_AGEMA_signal_5265 ;
    wire new_AGEMA_signal_5266 ;
    wire new_AGEMA_signal_5267 ;
    wire new_AGEMA_signal_5268 ;
    wire new_AGEMA_signal_5269 ;
    wire new_AGEMA_signal_5270 ;
    wire new_AGEMA_signal_5274 ;
    wire new_AGEMA_signal_5275 ;
    wire new_AGEMA_signal_5276 ;
    wire new_AGEMA_signal_5277 ;
    wire new_AGEMA_signal_5278 ;
    wire new_AGEMA_signal_5279 ;
    wire new_AGEMA_signal_5283 ;
    wire new_AGEMA_signal_5284 ;
    wire new_AGEMA_signal_5285 ;
    wire new_AGEMA_signal_5286 ;
    wire new_AGEMA_signal_5287 ;
    wire new_AGEMA_signal_5288 ;
    wire new_AGEMA_signal_5292 ;
    wire new_AGEMA_signal_5293 ;
    wire new_AGEMA_signal_5294 ;
    wire new_AGEMA_signal_5295 ;
    wire new_AGEMA_signal_5296 ;
    wire new_AGEMA_signal_5297 ;
    wire new_AGEMA_signal_5301 ;
    wire new_AGEMA_signal_5302 ;
    wire new_AGEMA_signal_5303 ;
    wire new_AGEMA_signal_5304 ;
    wire new_AGEMA_signal_5305 ;
    wire new_AGEMA_signal_5306 ;
    wire new_AGEMA_signal_5310 ;
    wire new_AGEMA_signal_5311 ;
    wire new_AGEMA_signal_5312 ;
    wire new_AGEMA_signal_5313 ;
    wire new_AGEMA_signal_5314 ;
    wire new_AGEMA_signal_5315 ;
    wire new_AGEMA_signal_5319 ;
    wire new_AGEMA_signal_5320 ;
    wire new_AGEMA_signal_5321 ;
    wire new_AGEMA_signal_5322 ;
    wire new_AGEMA_signal_5323 ;
    wire new_AGEMA_signal_5324 ;
    wire new_AGEMA_signal_5328 ;
    wire new_AGEMA_signal_5329 ;
    wire new_AGEMA_signal_5330 ;
    wire new_AGEMA_signal_5331 ;
    wire new_AGEMA_signal_5332 ;
    wire new_AGEMA_signal_5333 ;
    wire new_AGEMA_signal_5337 ;
    wire new_AGEMA_signal_5338 ;
    wire new_AGEMA_signal_5339 ;
    wire new_AGEMA_signal_5340 ;
    wire new_AGEMA_signal_5341 ;
    wire new_AGEMA_signal_5342 ;
    wire new_AGEMA_signal_5346 ;
    wire new_AGEMA_signal_5347 ;
    wire new_AGEMA_signal_5348 ;
    wire new_AGEMA_signal_5349 ;
    wire new_AGEMA_signal_5350 ;
    wire new_AGEMA_signal_5351 ;
    wire new_AGEMA_signal_5355 ;
    wire new_AGEMA_signal_5356 ;
    wire new_AGEMA_signal_5357 ;
    wire new_AGEMA_signal_5358 ;
    wire new_AGEMA_signal_5359 ;
    wire new_AGEMA_signal_5360 ;
    wire new_AGEMA_signal_5364 ;
    wire new_AGEMA_signal_5365 ;
    wire new_AGEMA_signal_5366 ;
    wire new_AGEMA_signal_5367 ;
    wire new_AGEMA_signal_5368 ;
    wire new_AGEMA_signal_5369 ;
    wire new_AGEMA_signal_5373 ;
    wire new_AGEMA_signal_5374 ;
    wire new_AGEMA_signal_5375 ;
    wire new_AGEMA_signal_5376 ;
    wire new_AGEMA_signal_5377 ;
    wire new_AGEMA_signal_5378 ;
    wire new_AGEMA_signal_5382 ;
    wire new_AGEMA_signal_5383 ;
    wire new_AGEMA_signal_5384 ;
    wire new_AGEMA_signal_5385 ;
    wire new_AGEMA_signal_5386 ;
    wire new_AGEMA_signal_5387 ;
    wire new_AGEMA_signal_5391 ;
    wire new_AGEMA_signal_5392 ;
    wire new_AGEMA_signal_5393 ;
    wire new_AGEMA_signal_5394 ;
    wire new_AGEMA_signal_5395 ;
    wire new_AGEMA_signal_5396 ;
    wire new_AGEMA_signal_5400 ;
    wire new_AGEMA_signal_5401 ;
    wire new_AGEMA_signal_5402 ;
    wire new_AGEMA_signal_5403 ;
    wire new_AGEMA_signal_5404 ;
    wire new_AGEMA_signal_5405 ;
    wire new_AGEMA_signal_5409 ;
    wire new_AGEMA_signal_5410 ;
    wire new_AGEMA_signal_5411 ;
    wire new_AGEMA_signal_5412 ;
    wire new_AGEMA_signal_5413 ;
    wire new_AGEMA_signal_5414 ;
    wire new_AGEMA_signal_5418 ;
    wire new_AGEMA_signal_5419 ;
    wire new_AGEMA_signal_5420 ;
    wire new_AGEMA_signal_5421 ;
    wire new_AGEMA_signal_5422 ;
    wire new_AGEMA_signal_5423 ;
    wire new_AGEMA_signal_5427 ;
    wire new_AGEMA_signal_5428 ;
    wire new_AGEMA_signal_5429 ;
    wire new_AGEMA_signal_5430 ;
    wire new_AGEMA_signal_5431 ;
    wire new_AGEMA_signal_5432 ;
    wire new_AGEMA_signal_5436 ;
    wire new_AGEMA_signal_5437 ;
    wire new_AGEMA_signal_5438 ;
    wire new_AGEMA_signal_5439 ;
    wire new_AGEMA_signal_5440 ;
    wire new_AGEMA_signal_5441 ;
    wire new_AGEMA_signal_5445 ;
    wire new_AGEMA_signal_5446 ;
    wire new_AGEMA_signal_5447 ;
    wire new_AGEMA_signal_5451 ;
    wire new_AGEMA_signal_5452 ;
    wire new_AGEMA_signal_5453 ;
    wire new_AGEMA_signal_5457 ;
    wire new_AGEMA_signal_5458 ;
    wire new_AGEMA_signal_5459 ;
    wire new_AGEMA_signal_5463 ;
    wire new_AGEMA_signal_5464 ;
    wire new_AGEMA_signal_5465 ;
    wire new_AGEMA_signal_5469 ;
    wire new_AGEMA_signal_5470 ;
    wire new_AGEMA_signal_5471 ;
    wire new_AGEMA_signal_5475 ;
    wire new_AGEMA_signal_5476 ;
    wire new_AGEMA_signal_5477 ;
    wire new_AGEMA_signal_5481 ;
    wire new_AGEMA_signal_5482 ;
    wire new_AGEMA_signal_5483 ;
    wire new_AGEMA_signal_5487 ;
    wire new_AGEMA_signal_5488 ;
    wire new_AGEMA_signal_5489 ;
    wire new_AGEMA_signal_5496 ;
    wire new_AGEMA_signal_5497 ;
    wire new_AGEMA_signal_5498 ;
    wire new_AGEMA_signal_5505 ;
    wire new_AGEMA_signal_5506 ;
    wire new_AGEMA_signal_5507 ;
    wire new_AGEMA_signal_5514 ;
    wire new_AGEMA_signal_5515 ;
    wire new_AGEMA_signal_5516 ;
    wire new_AGEMA_signal_5523 ;
    wire new_AGEMA_signal_5524 ;
    wire new_AGEMA_signal_5525 ;
    wire new_AGEMA_signal_5532 ;
    wire new_AGEMA_signal_5533 ;
    wire new_AGEMA_signal_5534 ;
    wire new_AGEMA_signal_5541 ;
    wire new_AGEMA_signal_5542 ;
    wire new_AGEMA_signal_5543 ;
    wire new_AGEMA_signal_5550 ;
    wire new_AGEMA_signal_5551 ;
    wire new_AGEMA_signal_5552 ;
    wire new_AGEMA_signal_5559 ;
    wire new_AGEMA_signal_5560 ;
    wire new_AGEMA_signal_5561 ;
    wire new_AGEMA_signal_5562 ;
    wire new_AGEMA_signal_5563 ;
    wire new_AGEMA_signal_5564 ;
    wire new_AGEMA_signal_5565 ;
    wire new_AGEMA_signal_5566 ;
    wire new_AGEMA_signal_5567 ;
    wire new_AGEMA_signal_5568 ;
    wire new_AGEMA_signal_5569 ;
    wire new_AGEMA_signal_5570 ;
    wire new_AGEMA_signal_5577 ;
    wire new_AGEMA_signal_5578 ;
    wire new_AGEMA_signal_5579 ;
    wire new_AGEMA_signal_5583 ;
    wire new_AGEMA_signal_5584 ;
    wire new_AGEMA_signal_5585 ;
    wire new_AGEMA_signal_5589 ;
    wire new_AGEMA_signal_5590 ;
    wire new_AGEMA_signal_5591 ;
    wire new_AGEMA_signal_5598 ;
    wire new_AGEMA_signal_5599 ;
    wire new_AGEMA_signal_5600 ;
    wire new_AGEMA_signal_5604 ;
    wire new_AGEMA_signal_5605 ;
    wire new_AGEMA_signal_5606 ;
    wire new_AGEMA_signal_5610 ;
    wire new_AGEMA_signal_5611 ;
    wire new_AGEMA_signal_5612 ;
    wire new_AGEMA_signal_5613 ;
    wire new_AGEMA_signal_5614 ;
    wire new_AGEMA_signal_5615 ;
    wire new_AGEMA_signal_5616 ;
    wire new_AGEMA_signal_5617 ;
    wire new_AGEMA_signal_5618 ;
    wire new_AGEMA_signal_5619 ;
    wire new_AGEMA_signal_5620 ;
    wire new_AGEMA_signal_5621 ;
    wire new_AGEMA_signal_5622 ;
    wire new_AGEMA_signal_5623 ;
    wire new_AGEMA_signal_5624 ;
    wire new_AGEMA_signal_5625 ;
    wire new_AGEMA_signal_5626 ;
    wire new_AGEMA_signal_5627 ;
    wire new_AGEMA_signal_5628 ;
    wire new_AGEMA_signal_5629 ;
    wire new_AGEMA_signal_5630 ;
    wire new_AGEMA_signal_5631 ;
    wire new_AGEMA_signal_5632 ;
    wire new_AGEMA_signal_5633 ;
    wire new_AGEMA_signal_5634 ;
    wire new_AGEMA_signal_5635 ;
    wire new_AGEMA_signal_5636 ;
    wire new_AGEMA_signal_5637 ;
    wire new_AGEMA_signal_5638 ;
    wire new_AGEMA_signal_5639 ;
    wire new_AGEMA_signal_5640 ;
    wire new_AGEMA_signal_5641 ;
    wire new_AGEMA_signal_5642 ;
    wire new_AGEMA_signal_5643 ;
    wire new_AGEMA_signal_5644 ;
    wire new_AGEMA_signal_5645 ;
    wire new_AGEMA_signal_5646 ;
    wire new_AGEMA_signal_5647 ;
    wire new_AGEMA_signal_5648 ;
    wire new_AGEMA_signal_5649 ;
    wire new_AGEMA_signal_5650 ;
    wire new_AGEMA_signal_5651 ;
    wire new_AGEMA_signal_5652 ;
    wire new_AGEMA_signal_5653 ;
    wire new_AGEMA_signal_5654 ;
    wire new_AGEMA_signal_5655 ;
    wire new_AGEMA_signal_5656 ;
    wire new_AGEMA_signal_5657 ;
    wire new_AGEMA_signal_5658 ;
    wire new_AGEMA_signal_5659 ;
    wire new_AGEMA_signal_5660 ;
    wire new_AGEMA_signal_5661 ;
    wire new_AGEMA_signal_5662 ;
    wire new_AGEMA_signal_5663 ;
    wire new_AGEMA_signal_5664 ;
    wire new_AGEMA_signal_5665 ;
    wire new_AGEMA_signal_5666 ;
    wire new_AGEMA_signal_5667 ;
    wire new_AGEMA_signal_5668 ;
    wire new_AGEMA_signal_5669 ;
    wire new_AGEMA_signal_5670 ;
    wire new_AGEMA_signal_5671 ;
    wire new_AGEMA_signal_5672 ;
    wire new_AGEMA_signal_5673 ;
    wire new_AGEMA_signal_5674 ;
    wire new_AGEMA_signal_5675 ;
    wire new_AGEMA_signal_5676 ;
    wire new_AGEMA_signal_5677 ;
    wire new_AGEMA_signal_5678 ;
    wire new_AGEMA_signal_5679 ;
    wire new_AGEMA_signal_5680 ;
    wire new_AGEMA_signal_5681 ;
    wire new_AGEMA_signal_5682 ;
    wire new_AGEMA_signal_5683 ;
    wire new_AGEMA_signal_5684 ;
    wire new_AGEMA_signal_5685 ;
    wire new_AGEMA_signal_5686 ;
    wire new_AGEMA_signal_5687 ;
    wire new_AGEMA_signal_5688 ;
    wire new_AGEMA_signal_5689 ;
    wire new_AGEMA_signal_5690 ;
    wire new_AGEMA_signal_5691 ;
    wire new_AGEMA_signal_5692 ;
    wire new_AGEMA_signal_5693 ;
    wire new_AGEMA_signal_5694 ;
    wire new_AGEMA_signal_5695 ;
    wire new_AGEMA_signal_5696 ;
    wire new_AGEMA_signal_5697 ;
    wire new_AGEMA_signal_5698 ;
    wire new_AGEMA_signal_5699 ;
    wire new_AGEMA_signal_5700 ;
    wire new_AGEMA_signal_5701 ;
    wire new_AGEMA_signal_5702 ;
    wire new_AGEMA_signal_5703 ;
    wire new_AGEMA_signal_5704 ;
    wire new_AGEMA_signal_5705 ;
    wire new_AGEMA_signal_5706 ;
    wire new_AGEMA_signal_5707 ;
    wire new_AGEMA_signal_5708 ;
    wire new_AGEMA_signal_5709 ;
    wire new_AGEMA_signal_5710 ;
    wire new_AGEMA_signal_5711 ;
    wire new_AGEMA_signal_5712 ;
    wire new_AGEMA_signal_5713 ;
    wire new_AGEMA_signal_5714 ;
    wire new_AGEMA_signal_5715 ;
    wire new_AGEMA_signal_5716 ;
    wire new_AGEMA_signal_5717 ;
    wire new_AGEMA_signal_5718 ;
    wire new_AGEMA_signal_5719 ;
    wire new_AGEMA_signal_5720 ;
    wire new_AGEMA_signal_5721 ;
    wire new_AGEMA_signal_5722 ;
    wire new_AGEMA_signal_5723 ;
    wire new_AGEMA_signal_5724 ;
    wire new_AGEMA_signal_5725 ;
    wire new_AGEMA_signal_5726 ;
    wire new_AGEMA_signal_5727 ;
    wire new_AGEMA_signal_5728 ;
    wire new_AGEMA_signal_5729 ;
    wire new_AGEMA_signal_5730 ;
    wire new_AGEMA_signal_5731 ;
    wire new_AGEMA_signal_5732 ;
    wire new_AGEMA_signal_5733 ;
    wire new_AGEMA_signal_5734 ;
    wire new_AGEMA_signal_5735 ;
    wire new_AGEMA_signal_5736 ;
    wire new_AGEMA_signal_5737 ;
    wire new_AGEMA_signal_5738 ;
    wire new_AGEMA_signal_5739 ;
    wire new_AGEMA_signal_5740 ;
    wire new_AGEMA_signal_5741 ;
    wire new_AGEMA_signal_5742 ;
    wire new_AGEMA_signal_5743 ;
    wire new_AGEMA_signal_5744 ;
    wire new_AGEMA_signal_5745 ;
    wire new_AGEMA_signal_5746 ;
    wire new_AGEMA_signal_5747 ;
    wire new_AGEMA_signal_5748 ;
    wire new_AGEMA_signal_5749 ;
    wire new_AGEMA_signal_5750 ;
    wire new_AGEMA_signal_5751 ;
    wire new_AGEMA_signal_5752 ;
    wire new_AGEMA_signal_5753 ;
    wire new_AGEMA_signal_5754 ;
    wire new_AGEMA_signal_5755 ;
    wire new_AGEMA_signal_5756 ;
    wire new_AGEMA_signal_5757 ;
    wire new_AGEMA_signal_5758 ;
    wire new_AGEMA_signal_5759 ;
    wire new_AGEMA_signal_5760 ;
    wire new_AGEMA_signal_5761 ;
    wire new_AGEMA_signal_5762 ;
    wire new_AGEMA_signal_5763 ;
    wire new_AGEMA_signal_5764 ;
    wire new_AGEMA_signal_5765 ;
    wire new_AGEMA_signal_5766 ;
    wire new_AGEMA_signal_5767 ;
    wire new_AGEMA_signal_5768 ;
    wire new_AGEMA_signal_5769 ;
    wire new_AGEMA_signal_5770 ;
    wire new_AGEMA_signal_5771 ;
    wire new_AGEMA_signal_5772 ;
    wire new_AGEMA_signal_5773 ;
    wire new_AGEMA_signal_5774 ;
    wire new_AGEMA_signal_5775 ;
    wire new_AGEMA_signal_5776 ;
    wire new_AGEMA_signal_5777 ;
    wire new_AGEMA_signal_5778 ;
    wire new_AGEMA_signal_5779 ;
    wire new_AGEMA_signal_5780 ;
    wire new_AGEMA_signal_5781 ;
    wire new_AGEMA_signal_5782 ;
    wire new_AGEMA_signal_5783 ;
    wire new_AGEMA_signal_5784 ;
    wire new_AGEMA_signal_5785 ;
    wire new_AGEMA_signal_5786 ;
    wire new_AGEMA_signal_5787 ;
    wire new_AGEMA_signal_5788 ;
    wire new_AGEMA_signal_5789 ;
    wire new_AGEMA_signal_5790 ;
    wire new_AGEMA_signal_5791 ;
    wire new_AGEMA_signal_5792 ;
    wire new_AGEMA_signal_5793 ;
    wire new_AGEMA_signal_5794 ;
    wire new_AGEMA_signal_5795 ;
    wire new_AGEMA_signal_5796 ;
    wire new_AGEMA_signal_5797 ;
    wire new_AGEMA_signal_5798 ;
    wire new_AGEMA_signal_5799 ;
    wire new_AGEMA_signal_5800 ;
    wire new_AGEMA_signal_5801 ;
    wire new_AGEMA_signal_5802 ;
    wire new_AGEMA_signal_5803 ;
    wire new_AGEMA_signal_5804 ;
    wire new_AGEMA_signal_5805 ;
    wire new_AGEMA_signal_5806 ;
    wire new_AGEMA_signal_5807 ;
    wire new_AGEMA_signal_5808 ;
    wire new_AGEMA_signal_5809 ;
    wire new_AGEMA_signal_5810 ;
    wire new_AGEMA_signal_5811 ;
    wire new_AGEMA_signal_5812 ;
    wire new_AGEMA_signal_5813 ;
    wire new_AGEMA_signal_5814 ;
    wire new_AGEMA_signal_5815 ;
    wire new_AGEMA_signal_5817 ;
    wire new_AGEMA_signal_5818 ;
    wire new_AGEMA_signal_5819 ;
    wire new_AGEMA_signal_5820 ;
    wire new_AGEMA_signal_5821 ;
    wire new_AGEMA_signal_5822 ;
    wire new_AGEMA_signal_5823 ;
    wire new_AGEMA_signal_5824 ;
    wire new_AGEMA_signal_5825 ;
    wire new_AGEMA_signal_5826 ;
    wire new_AGEMA_signal_5827 ;
    wire new_AGEMA_signal_5828 ;
    wire new_AGEMA_signal_5829 ;
    wire new_AGEMA_signal_5830 ;
    wire new_AGEMA_signal_5831 ;
    wire new_AGEMA_signal_5832 ;
    wire new_AGEMA_signal_5833 ;
    wire new_AGEMA_signal_5834 ;
    wire new_AGEMA_signal_5835 ;
    wire new_AGEMA_signal_5836 ;
    wire new_AGEMA_signal_5837 ;
    wire new_AGEMA_signal_5838 ;
    wire new_AGEMA_signal_5839 ;
    wire new_AGEMA_signal_5840 ;
    wire new_AGEMA_signal_5841 ;
    wire new_AGEMA_signal_5842 ;
    wire new_AGEMA_signal_5843 ;
    wire new_AGEMA_signal_5844 ;
    wire new_AGEMA_signal_5845 ;
    wire new_AGEMA_signal_5846 ;
    wire new_AGEMA_signal_5847 ;
    wire new_AGEMA_signal_5848 ;
    wire new_AGEMA_signal_5849 ;
    wire new_AGEMA_signal_5850 ;
    wire new_AGEMA_signal_5851 ;
    wire new_AGEMA_signal_5852 ;
    wire new_AGEMA_signal_5853 ;
    wire new_AGEMA_signal_5854 ;
    wire new_AGEMA_signal_5855 ;
    wire new_AGEMA_signal_5856 ;
    wire new_AGEMA_signal_5857 ;
    wire new_AGEMA_signal_5858 ;
    wire new_AGEMA_signal_5859 ;
    wire new_AGEMA_signal_5860 ;
    wire new_AGEMA_signal_5861 ;
    wire new_AGEMA_signal_5862 ;
    wire new_AGEMA_signal_5863 ;
    wire new_AGEMA_signal_5864 ;
    wire new_AGEMA_signal_5865 ;
    wire new_AGEMA_signal_5866 ;
    wire new_AGEMA_signal_5867 ;
    wire new_AGEMA_signal_5868 ;
    wire new_AGEMA_signal_5869 ;
    wire new_AGEMA_signal_5870 ;
    wire new_AGEMA_signal_5871 ;
    wire new_AGEMA_signal_5872 ;
    wire new_AGEMA_signal_5873 ;
    wire new_AGEMA_signal_5874 ;
    wire new_AGEMA_signal_5875 ;
    wire new_AGEMA_signal_5876 ;
    wire new_AGEMA_signal_5877 ;
    wire new_AGEMA_signal_5878 ;
    wire new_AGEMA_signal_5879 ;
    wire new_AGEMA_signal_5880 ;
    wire new_AGEMA_signal_5881 ;
    wire new_AGEMA_signal_5882 ;
    wire new_AGEMA_signal_5883 ;
    wire new_AGEMA_signal_5884 ;
    wire new_AGEMA_signal_5885 ;
    wire new_AGEMA_signal_5886 ;
    wire new_AGEMA_signal_5887 ;
    wire new_AGEMA_signal_5888 ;
    wire new_AGEMA_signal_5889 ;
    wire new_AGEMA_signal_5890 ;
    wire new_AGEMA_signal_5891 ;
    wire new_AGEMA_signal_5892 ;
    wire new_AGEMA_signal_5893 ;
    wire new_AGEMA_signal_5894 ;
    wire new_AGEMA_signal_5895 ;
    wire new_AGEMA_signal_5896 ;
    wire new_AGEMA_signal_5897 ;
    wire new_AGEMA_signal_5898 ;
    wire new_AGEMA_signal_5899 ;
    wire new_AGEMA_signal_5900 ;
    wire new_AGEMA_signal_5901 ;
    wire new_AGEMA_signal_5902 ;
    wire new_AGEMA_signal_5903 ;
    wire new_AGEMA_signal_5904 ;
    wire new_AGEMA_signal_5905 ;
    wire new_AGEMA_signal_5906 ;
    wire new_AGEMA_signal_5907 ;
    wire new_AGEMA_signal_5908 ;
    wire new_AGEMA_signal_5909 ;
    wire new_AGEMA_signal_5910 ;
    wire new_AGEMA_signal_5911 ;
    wire new_AGEMA_signal_5912 ;
    wire new_AGEMA_signal_5913 ;
    wire new_AGEMA_signal_5914 ;
    wire new_AGEMA_signal_5915 ;
    wire new_AGEMA_signal_5916 ;
    wire new_AGEMA_signal_5917 ;
    wire new_AGEMA_signal_5918 ;
    wire new_AGEMA_signal_5919 ;
    wire new_AGEMA_signal_5920 ;
    wire new_AGEMA_signal_5921 ;
    wire new_AGEMA_signal_5922 ;
    wire new_AGEMA_signal_5923 ;
    wire new_AGEMA_signal_5924 ;
    wire new_AGEMA_signal_5925 ;
    wire new_AGEMA_signal_5926 ;
    wire new_AGEMA_signal_5927 ;
    wire new_AGEMA_signal_5928 ;
    wire new_AGEMA_signal_5929 ;
    wire new_AGEMA_signal_5930 ;
    wire new_AGEMA_signal_5931 ;
    wire new_AGEMA_signal_5932 ;
    wire new_AGEMA_signal_5933 ;
    wire new_AGEMA_signal_5934 ;
    wire new_AGEMA_signal_5935 ;
    wire new_AGEMA_signal_5936 ;
    wire new_AGEMA_signal_5937 ;
    wire new_AGEMA_signal_5938 ;
    wire new_AGEMA_signal_5939 ;
    wire new_AGEMA_signal_5940 ;
    wire new_AGEMA_signal_5941 ;
    wire new_AGEMA_signal_5942 ;
    wire new_AGEMA_signal_5943 ;
    wire new_AGEMA_signal_5944 ;
    wire new_AGEMA_signal_5945 ;
    wire new_AGEMA_signal_5946 ;
    wire new_AGEMA_signal_5947 ;
    wire new_AGEMA_signal_5948 ;
    wire new_AGEMA_signal_5949 ;
    wire new_AGEMA_signal_5950 ;
    wire new_AGEMA_signal_5951 ;
    wire new_AGEMA_signal_5952 ;
    wire new_AGEMA_signal_5953 ;
    wire new_AGEMA_signal_5954 ;
    wire new_AGEMA_signal_5955 ;
    wire new_AGEMA_signal_5956 ;
    wire new_AGEMA_signal_5957 ;
    wire new_AGEMA_signal_5958 ;
    wire new_AGEMA_signal_5959 ;
    wire new_AGEMA_signal_5960 ;
    wire new_AGEMA_signal_5961 ;
    wire new_AGEMA_signal_5962 ;
    wire new_AGEMA_signal_5963 ;
    wire new_AGEMA_signal_5964 ;
    wire new_AGEMA_signal_5965 ;
    wire new_AGEMA_signal_5966 ;
    wire new_AGEMA_signal_5967 ;
    wire new_AGEMA_signal_5968 ;
    wire new_AGEMA_signal_5969 ;
    wire new_AGEMA_signal_5970 ;
    wire new_AGEMA_signal_5971 ;
    wire new_AGEMA_signal_5972 ;
    wire new_AGEMA_signal_5973 ;
    wire new_AGEMA_signal_5974 ;
    wire new_AGEMA_signal_5975 ;
    wire new_AGEMA_signal_5976 ;
    wire new_AGEMA_signal_5977 ;
    wire new_AGEMA_signal_5978 ;
    wire new_AGEMA_signal_5979 ;
    wire new_AGEMA_signal_5980 ;
    wire new_AGEMA_signal_5981 ;
    wire new_AGEMA_signal_5982 ;
    wire new_AGEMA_signal_5983 ;
    wire new_AGEMA_signal_5984 ;
    wire new_AGEMA_signal_5985 ;
    wire new_AGEMA_signal_5986 ;
    wire new_AGEMA_signal_5987 ;
    wire new_AGEMA_signal_5988 ;
    wire new_AGEMA_signal_5989 ;
    wire new_AGEMA_signal_5990 ;
    wire new_AGEMA_signal_5991 ;
    wire new_AGEMA_signal_5992 ;
    wire new_AGEMA_signal_5993 ;
    wire new_AGEMA_signal_5994 ;
    wire new_AGEMA_signal_5995 ;
    wire new_AGEMA_signal_5996 ;
    wire new_AGEMA_signal_5997 ;
    wire new_AGEMA_signal_5998 ;
    wire new_AGEMA_signal_5999 ;
    wire new_AGEMA_signal_6000 ;
    wire new_AGEMA_signal_6001 ;
    wire new_AGEMA_signal_6002 ;
    wire new_AGEMA_signal_6003 ;
    wire new_AGEMA_signal_6004 ;
    wire new_AGEMA_signal_6005 ;
    wire new_AGEMA_signal_6006 ;
    wire new_AGEMA_signal_6007 ;
    wire new_AGEMA_signal_6008 ;
    wire new_AGEMA_signal_6009 ;
    wire new_AGEMA_signal_6010 ;
    wire new_AGEMA_signal_6011 ;
    wire new_AGEMA_signal_6012 ;
    wire new_AGEMA_signal_6013 ;
    wire new_AGEMA_signal_6014 ;
    wire new_AGEMA_signal_6015 ;
    wire new_AGEMA_signal_6016 ;
    wire new_AGEMA_signal_6017 ;
    wire new_AGEMA_signal_6018 ;
    wire new_AGEMA_signal_6019 ;
    wire new_AGEMA_signal_6020 ;
    wire new_AGEMA_signal_6021 ;
    wire new_AGEMA_signal_6022 ;
    wire new_AGEMA_signal_6023 ;
    wire new_AGEMA_signal_6024 ;
    wire new_AGEMA_signal_6025 ;
    wire new_AGEMA_signal_6026 ;
    wire new_AGEMA_signal_6027 ;
    wire new_AGEMA_signal_6028 ;
    wire new_AGEMA_signal_6029 ;
    wire new_AGEMA_signal_6030 ;
    wire new_AGEMA_signal_6031 ;
    wire new_AGEMA_signal_6032 ;
    wire new_AGEMA_signal_6033 ;
    wire new_AGEMA_signal_6034 ;
    wire new_AGEMA_signal_6035 ;
    wire new_AGEMA_signal_6036 ;
    wire new_AGEMA_signal_6037 ;
    wire new_AGEMA_signal_6038 ;
    wire new_AGEMA_signal_6039 ;
    wire new_AGEMA_signal_6040 ;
    wire new_AGEMA_signal_6041 ;
    wire new_AGEMA_signal_6042 ;
    wire new_AGEMA_signal_6043 ;
    wire new_AGEMA_signal_6044 ;
    wire new_AGEMA_signal_6045 ;
    wire new_AGEMA_signal_6046 ;
    wire new_AGEMA_signal_6047 ;
    wire new_AGEMA_signal_6048 ;
    wire new_AGEMA_signal_6049 ;
    wire new_AGEMA_signal_6050 ;
    wire new_AGEMA_signal_6051 ;
    wire new_AGEMA_signal_6052 ;
    wire new_AGEMA_signal_6053 ;
    wire new_AGEMA_signal_6054 ;
    wire new_AGEMA_signal_6055 ;
    wire new_AGEMA_signal_6056 ;
    wire new_AGEMA_signal_6057 ;
    wire new_AGEMA_signal_6058 ;
    wire new_AGEMA_signal_6059 ;
    wire new_AGEMA_signal_6060 ;
    wire new_AGEMA_signal_6061 ;
    wire new_AGEMA_signal_6062 ;
    wire new_AGEMA_signal_6063 ;
    wire new_AGEMA_signal_6064 ;
    wire new_AGEMA_signal_6065 ;
    wire new_AGEMA_signal_6066 ;
    wire new_AGEMA_signal_6067 ;
    wire new_AGEMA_signal_6068 ;
    wire new_AGEMA_signal_6069 ;
    wire new_AGEMA_signal_6070 ;
    wire new_AGEMA_signal_6071 ;
    wire new_AGEMA_signal_6072 ;
    wire new_AGEMA_signal_6073 ;
    wire new_AGEMA_signal_6074 ;
    wire new_AGEMA_signal_6075 ;
    wire new_AGEMA_signal_6076 ;
    wire new_AGEMA_signal_6077 ;
    wire new_AGEMA_signal_6078 ;
    wire new_AGEMA_signal_6079 ;
    wire new_AGEMA_signal_6080 ;
    wire new_AGEMA_signal_6081 ;
    wire new_AGEMA_signal_6082 ;
    wire new_AGEMA_signal_6083 ;
    wire new_AGEMA_signal_6084 ;
    wire new_AGEMA_signal_6085 ;
    wire new_AGEMA_signal_6086 ;
    wire new_AGEMA_signal_6087 ;
    wire new_AGEMA_signal_6088 ;
    wire new_AGEMA_signal_6089 ;
    wire new_AGEMA_signal_6090 ;
    wire new_AGEMA_signal_6091 ;
    wire new_AGEMA_signal_6092 ;
    wire new_AGEMA_signal_6093 ;
    wire new_AGEMA_signal_6094 ;
    wire new_AGEMA_signal_6095 ;
    wire new_AGEMA_signal_6096 ;
    wire new_AGEMA_signal_6097 ;
    wire new_AGEMA_signal_6098 ;
    wire new_AGEMA_signal_6099 ;
    wire new_AGEMA_signal_6100 ;
    wire new_AGEMA_signal_6101 ;
    wire new_AGEMA_signal_6102 ;
    wire new_AGEMA_signal_6103 ;
    wire new_AGEMA_signal_6104 ;
    wire new_AGEMA_signal_6105 ;
    wire new_AGEMA_signal_6106 ;
    wire new_AGEMA_signal_6107 ;
    wire new_AGEMA_signal_6108 ;
    wire new_AGEMA_signal_6109 ;
    wire new_AGEMA_signal_6110 ;
    wire new_AGEMA_signal_6111 ;
    wire new_AGEMA_signal_6112 ;
    wire new_AGEMA_signal_6113 ;
    wire new_AGEMA_signal_6114 ;
    wire new_AGEMA_signal_6115 ;
    wire new_AGEMA_signal_6116 ;
    wire new_AGEMA_signal_6117 ;
    wire new_AGEMA_signal_6118 ;
    wire new_AGEMA_signal_6119 ;
    wire new_AGEMA_signal_6120 ;
    wire new_AGEMA_signal_6121 ;
    wire new_AGEMA_signal_6122 ;
    wire new_AGEMA_signal_6123 ;
    wire new_AGEMA_signal_6124 ;
    wire new_AGEMA_signal_6125 ;
    wire new_AGEMA_signal_6126 ;
    wire new_AGEMA_signal_6127 ;
    wire new_AGEMA_signal_6128 ;
    wire new_AGEMA_signal_6129 ;
    wire new_AGEMA_signal_6130 ;
    wire new_AGEMA_signal_6131 ;
    wire new_AGEMA_signal_6132 ;
    wire new_AGEMA_signal_6133 ;
    wire new_AGEMA_signal_6134 ;
    wire new_AGEMA_signal_6135 ;
    wire new_AGEMA_signal_6136 ;
    wire new_AGEMA_signal_6137 ;
    wire new_AGEMA_signal_6138 ;
    wire new_AGEMA_signal_6139 ;
    wire new_AGEMA_signal_6140 ;
    wire new_AGEMA_signal_6141 ;
    wire new_AGEMA_signal_6142 ;
    wire new_AGEMA_signal_6143 ;
    wire new_AGEMA_signal_6144 ;
    wire new_AGEMA_signal_6145 ;
    wire new_AGEMA_signal_6146 ;
    wire new_AGEMA_signal_6147 ;
    wire new_AGEMA_signal_6148 ;
    wire new_AGEMA_signal_6149 ;
    wire new_AGEMA_signal_6150 ;
    wire new_AGEMA_signal_6151 ;
    wire new_AGEMA_signal_6152 ;
    wire new_AGEMA_signal_6153 ;
    wire new_AGEMA_signal_6154 ;
    wire new_AGEMA_signal_6155 ;
    wire new_AGEMA_signal_6156 ;
    wire new_AGEMA_signal_6157 ;
    wire new_AGEMA_signal_6158 ;
    wire new_AGEMA_signal_6159 ;
    wire new_AGEMA_signal_6160 ;
    wire new_AGEMA_signal_6161 ;
    wire new_AGEMA_signal_6162 ;
    wire new_AGEMA_signal_6163 ;
    wire new_AGEMA_signal_6164 ;
    wire new_AGEMA_signal_6165 ;
    wire new_AGEMA_signal_6166 ;
    wire new_AGEMA_signal_6167 ;
    wire new_AGEMA_signal_6168 ;
    wire new_AGEMA_signal_6169 ;
    wire new_AGEMA_signal_6170 ;
    wire new_AGEMA_signal_6171 ;
    wire new_AGEMA_signal_6172 ;
    wire new_AGEMA_signal_6173 ;
    wire new_AGEMA_signal_6174 ;
    wire new_AGEMA_signal_6175 ;
    wire new_AGEMA_signal_6176 ;
    wire new_AGEMA_signal_6177 ;
    wire new_AGEMA_signal_6178 ;
    wire new_AGEMA_signal_6179 ;
    wire new_AGEMA_signal_6180 ;
    wire new_AGEMA_signal_6181 ;
    wire new_AGEMA_signal_6182 ;
    wire new_AGEMA_signal_6183 ;
    wire new_AGEMA_signal_6184 ;
    wire new_AGEMA_signal_6185 ;
    wire new_AGEMA_signal_6186 ;
    wire new_AGEMA_signal_6187 ;
    wire new_AGEMA_signal_6188 ;
    wire new_AGEMA_signal_6189 ;
    wire new_AGEMA_signal_6190 ;
    wire new_AGEMA_signal_6191 ;
    wire new_AGEMA_signal_6192 ;
    wire new_AGEMA_signal_6193 ;
    wire new_AGEMA_signal_6194 ;
    wire new_AGEMA_signal_6195 ;
    wire new_AGEMA_signal_6196 ;
    wire new_AGEMA_signal_6197 ;
    wire new_AGEMA_signal_6198 ;
    wire new_AGEMA_signal_6199 ;
    wire new_AGEMA_signal_6200 ;
    wire new_AGEMA_signal_6201 ;
    wire new_AGEMA_signal_6202 ;
    wire new_AGEMA_signal_6203 ;
    wire new_AGEMA_signal_6204 ;
    wire new_AGEMA_signal_6205 ;
    wire new_AGEMA_signal_6206 ;
    wire new_AGEMA_signal_6207 ;
    wire new_AGEMA_signal_6208 ;
    wire new_AGEMA_signal_6209 ;
    wire new_AGEMA_signal_6210 ;
    wire new_AGEMA_signal_6211 ;
    wire new_AGEMA_signal_6212 ;
    wire new_AGEMA_signal_6213 ;
    wire new_AGEMA_signal_6214 ;
    wire new_AGEMA_signal_6215 ;
    wire new_AGEMA_signal_6216 ;
    wire new_AGEMA_signal_6217 ;
    wire new_AGEMA_signal_6218 ;
    wire new_AGEMA_signal_6219 ;
    wire new_AGEMA_signal_6220 ;
    wire new_AGEMA_signal_6221 ;
    wire new_AGEMA_signal_6222 ;
    wire new_AGEMA_signal_6223 ;
    wire new_AGEMA_signal_6224 ;
    wire new_AGEMA_signal_6225 ;
    wire new_AGEMA_signal_6226 ;
    wire new_AGEMA_signal_6227 ;
    wire new_AGEMA_signal_6228 ;
    wire new_AGEMA_signal_6229 ;
    wire new_AGEMA_signal_6230 ;
    wire new_AGEMA_signal_6231 ;
    wire new_AGEMA_signal_6232 ;
    wire new_AGEMA_signal_6233 ;
    wire new_AGEMA_signal_6234 ;
    wire new_AGEMA_signal_6235 ;
    wire new_AGEMA_signal_6236 ;
    wire new_AGEMA_signal_6237 ;
    wire new_AGEMA_signal_6238 ;
    wire new_AGEMA_signal_6239 ;
    wire new_AGEMA_signal_6240 ;
    wire new_AGEMA_signal_6241 ;
    wire new_AGEMA_signal_6242 ;
    wire new_AGEMA_signal_6243 ;
    wire new_AGEMA_signal_6244 ;
    wire new_AGEMA_signal_6245 ;
    wire new_AGEMA_signal_6246 ;
    wire new_AGEMA_signal_6247 ;
    wire new_AGEMA_signal_6248 ;
    wire new_AGEMA_signal_6249 ;
    wire new_AGEMA_signal_6250 ;
    wire new_AGEMA_signal_6251 ;
    wire new_AGEMA_signal_6252 ;
    wire new_AGEMA_signal_6253 ;
    wire new_AGEMA_signal_6254 ;
    wire new_AGEMA_signal_6255 ;
    wire new_AGEMA_signal_6256 ;
    wire new_AGEMA_signal_6257 ;
    wire new_AGEMA_signal_6258 ;
    wire new_AGEMA_signal_6259 ;
    wire new_AGEMA_signal_6260 ;
    wire new_AGEMA_signal_6261 ;
    wire new_AGEMA_signal_6262 ;
    wire new_AGEMA_signal_6263 ;
    wire new_AGEMA_signal_6264 ;
    wire new_AGEMA_signal_6265 ;
    wire new_AGEMA_signal_6266 ;
    wire new_AGEMA_signal_6267 ;
    wire new_AGEMA_signal_6268 ;
    wire new_AGEMA_signal_6269 ;
    wire new_AGEMA_signal_6270 ;
    wire new_AGEMA_signal_6271 ;
    wire new_AGEMA_signal_6272 ;
    wire new_AGEMA_signal_6273 ;
    wire new_AGEMA_signal_6274 ;
    wire new_AGEMA_signal_6275 ;
    wire new_AGEMA_signal_6276 ;
    wire new_AGEMA_signal_6277 ;
    wire new_AGEMA_signal_6278 ;
    wire new_AGEMA_signal_6279 ;
    wire new_AGEMA_signal_6280 ;
    wire new_AGEMA_signal_6281 ;
    wire new_AGEMA_signal_6282 ;
    wire new_AGEMA_signal_6283 ;
    wire new_AGEMA_signal_6284 ;
    wire new_AGEMA_signal_6285 ;
    wire new_AGEMA_signal_6286 ;
    wire new_AGEMA_signal_6287 ;
    wire new_AGEMA_signal_6288 ;
    wire new_AGEMA_signal_6289 ;
    wire new_AGEMA_signal_6290 ;
    wire new_AGEMA_signal_6291 ;
    wire new_AGEMA_signal_6292 ;
    wire new_AGEMA_signal_6293 ;
    wire new_AGEMA_signal_6294 ;
    wire new_AGEMA_signal_6295 ;
    wire new_AGEMA_signal_6296 ;
    wire new_AGEMA_signal_6297 ;
    wire new_AGEMA_signal_6298 ;
    wire new_AGEMA_signal_6299 ;
    wire new_AGEMA_signal_6300 ;
    wire new_AGEMA_signal_6301 ;
    wire new_AGEMA_signal_6302 ;
    wire new_AGEMA_signal_6303 ;
    wire new_AGEMA_signal_6304 ;
    wire new_AGEMA_signal_6305 ;
    wire new_AGEMA_signal_6306 ;
    wire new_AGEMA_signal_6307 ;
    wire new_AGEMA_signal_6308 ;
    wire new_AGEMA_signal_6309 ;
    wire new_AGEMA_signal_6310 ;
    wire new_AGEMA_signal_6311 ;
    wire new_AGEMA_signal_6312 ;
    wire new_AGEMA_signal_6313 ;
    wire new_AGEMA_signal_6314 ;
    wire new_AGEMA_signal_6315 ;
    wire new_AGEMA_signal_6316 ;
    wire new_AGEMA_signal_6317 ;
    wire new_AGEMA_signal_6318 ;
    wire new_AGEMA_signal_6319 ;
    wire new_AGEMA_signal_6320 ;
    wire new_AGEMA_signal_6321 ;
    wire new_AGEMA_signal_6322 ;
    wire new_AGEMA_signal_6323 ;
    wire new_AGEMA_signal_6324 ;
    wire new_AGEMA_signal_6325 ;
    wire new_AGEMA_signal_6326 ;
    wire new_AGEMA_signal_6327 ;
    wire new_AGEMA_signal_6328 ;
    wire new_AGEMA_signal_6329 ;
    wire new_AGEMA_signal_6330 ;
    wire new_AGEMA_signal_6331 ;
    wire new_AGEMA_signal_6332 ;
    wire new_AGEMA_signal_6333 ;
    wire new_AGEMA_signal_6334 ;
    wire new_AGEMA_signal_6335 ;
    wire new_AGEMA_signal_6336 ;
    wire new_AGEMA_signal_6337 ;
    wire new_AGEMA_signal_6338 ;
    wire new_AGEMA_signal_6339 ;
    wire new_AGEMA_signal_6340 ;
    wire new_AGEMA_signal_6341 ;
    wire new_AGEMA_signal_6342 ;
    wire new_AGEMA_signal_6343 ;
    wire new_AGEMA_signal_6344 ;
    wire new_AGEMA_signal_6345 ;
    wire new_AGEMA_signal_6346 ;
    wire new_AGEMA_signal_6347 ;
    wire new_AGEMA_signal_6348 ;
    wire new_AGEMA_signal_6349 ;
    wire new_AGEMA_signal_6350 ;
    wire new_AGEMA_signal_6351 ;
    wire new_AGEMA_signal_6352 ;
    wire new_AGEMA_signal_6353 ;
    wire new_AGEMA_signal_6354 ;
    wire new_AGEMA_signal_6355 ;
    wire new_AGEMA_signal_6356 ;
    wire new_AGEMA_signal_6357 ;
    wire new_AGEMA_signal_6358 ;
    wire new_AGEMA_signal_6359 ;
    wire new_AGEMA_signal_6360 ;
    wire new_AGEMA_signal_6361 ;
    wire new_AGEMA_signal_6362 ;
    wire new_AGEMA_signal_6363 ;
    wire new_AGEMA_signal_6364 ;
    wire new_AGEMA_signal_6365 ;
    wire new_AGEMA_signal_6366 ;
    wire new_AGEMA_signal_6367 ;
    wire new_AGEMA_signal_6368 ;
    wire new_AGEMA_signal_6369 ;
    wire new_AGEMA_signal_6370 ;
    wire new_AGEMA_signal_6371 ;
    wire new_AGEMA_signal_6372 ;
    wire new_AGEMA_signal_6373 ;
    wire new_AGEMA_signal_6374 ;
    wire new_AGEMA_signal_6375 ;
    wire new_AGEMA_signal_6376 ;
    wire new_AGEMA_signal_6377 ;
    wire new_AGEMA_signal_6378 ;
    wire new_AGEMA_signal_6379 ;
    wire new_AGEMA_signal_6380 ;
    wire new_AGEMA_signal_6381 ;
    wire new_AGEMA_signal_6382 ;
    wire new_AGEMA_signal_6383 ;
    wire new_AGEMA_signal_6384 ;
    wire new_AGEMA_signal_6385 ;
    wire new_AGEMA_signal_6386 ;
    wire new_AGEMA_signal_6387 ;
    wire new_AGEMA_signal_6388 ;
    wire new_AGEMA_signal_6389 ;
    wire new_AGEMA_signal_6390 ;
    wire new_AGEMA_signal_6391 ;
    wire new_AGEMA_signal_6392 ;
    wire new_AGEMA_signal_6393 ;
    wire new_AGEMA_signal_6394 ;
    wire new_AGEMA_signal_6395 ;
    wire new_AGEMA_signal_6396 ;
    wire new_AGEMA_signal_6397 ;
    wire new_AGEMA_signal_6398 ;
    wire new_AGEMA_signal_6399 ;
    wire new_AGEMA_signal_6400 ;
    wire new_AGEMA_signal_6401 ;
    wire new_AGEMA_signal_6402 ;
    wire new_AGEMA_signal_6403 ;
    wire new_AGEMA_signal_6404 ;
    wire new_AGEMA_signal_6405 ;
    wire new_AGEMA_signal_6406 ;
    wire new_AGEMA_signal_6407 ;
    wire new_AGEMA_signal_6408 ;
    wire new_AGEMA_signal_6409 ;
    wire new_AGEMA_signal_6410 ;
    wire new_AGEMA_signal_6411 ;
    wire new_AGEMA_signal_6412 ;
    wire new_AGEMA_signal_6413 ;
    wire new_AGEMA_signal_6414 ;
    wire new_AGEMA_signal_6415 ;
    wire new_AGEMA_signal_6416 ;
    wire new_AGEMA_signal_6417 ;
    wire new_AGEMA_signal_6418 ;
    wire new_AGEMA_signal_6419 ;
    wire new_AGEMA_signal_6420 ;
    wire new_AGEMA_signal_6421 ;
    wire new_AGEMA_signal_6422 ;
    wire new_AGEMA_signal_6423 ;
    wire new_AGEMA_signal_6424 ;
    wire new_AGEMA_signal_6425 ;
    wire new_AGEMA_signal_6426 ;
    wire new_AGEMA_signal_6427 ;
    wire new_AGEMA_signal_6428 ;
    wire new_AGEMA_signal_6429 ;
    wire new_AGEMA_signal_6430 ;
    wire new_AGEMA_signal_6431 ;
    wire new_AGEMA_signal_6432 ;
    wire new_AGEMA_signal_6433 ;
    wire new_AGEMA_signal_6434 ;
    wire new_AGEMA_signal_6435 ;
    wire new_AGEMA_signal_6436 ;
    wire new_AGEMA_signal_6437 ;
    wire new_AGEMA_signal_6438 ;
    wire new_AGEMA_signal_6439 ;
    wire new_AGEMA_signal_6440 ;
    wire new_AGEMA_signal_6441 ;
    wire new_AGEMA_signal_6442 ;
    wire new_AGEMA_signal_6443 ;
    wire new_AGEMA_signal_6444 ;
    wire new_AGEMA_signal_6445 ;
    wire new_AGEMA_signal_6446 ;
    wire new_AGEMA_signal_6447 ;
    wire new_AGEMA_signal_6448 ;
    wire new_AGEMA_signal_6449 ;
    wire new_AGEMA_signal_6450 ;
    wire new_AGEMA_signal_6451 ;
    wire new_AGEMA_signal_6452 ;
    wire new_AGEMA_signal_6453 ;
    wire new_AGEMA_signal_6454 ;
    wire new_AGEMA_signal_6455 ;
    wire new_AGEMA_signal_6456 ;
    wire new_AGEMA_signal_6457 ;
    wire new_AGEMA_signal_6458 ;
    wire new_AGEMA_signal_6459 ;
    wire new_AGEMA_signal_6460 ;
    wire new_AGEMA_signal_6461 ;
    wire new_AGEMA_signal_6462 ;
    wire new_AGEMA_signal_6463 ;
    wire new_AGEMA_signal_6464 ;
    wire new_AGEMA_signal_6465 ;
    wire new_AGEMA_signal_6466 ;
    wire new_AGEMA_signal_6467 ;
    wire new_AGEMA_signal_6468 ;
    wire new_AGEMA_signal_6469 ;
    wire new_AGEMA_signal_6470 ;
    wire new_AGEMA_signal_6471 ;
    wire new_AGEMA_signal_6472 ;
    wire new_AGEMA_signal_6473 ;
    wire new_AGEMA_signal_6474 ;
    wire new_AGEMA_signal_6475 ;
    wire new_AGEMA_signal_6476 ;
    wire new_AGEMA_signal_6477 ;
    wire new_AGEMA_signal_6478 ;
    wire new_AGEMA_signal_6479 ;
    wire new_AGEMA_signal_6480 ;
    wire new_AGEMA_signal_6481 ;
    wire new_AGEMA_signal_6482 ;
    wire new_AGEMA_signal_6483 ;
    wire new_AGEMA_signal_6484 ;
    wire new_AGEMA_signal_6485 ;
    wire new_AGEMA_signal_6486 ;
    wire new_AGEMA_signal_6487 ;
    wire new_AGEMA_signal_6488 ;
    wire new_AGEMA_signal_6489 ;
    wire new_AGEMA_signal_6490 ;
    wire new_AGEMA_signal_6491 ;
    wire new_AGEMA_signal_6492 ;
    wire new_AGEMA_signal_6493 ;
    wire new_AGEMA_signal_6494 ;
    wire new_AGEMA_signal_6495 ;
    wire new_AGEMA_signal_6496 ;
    wire new_AGEMA_signal_6497 ;
    wire new_AGEMA_signal_6498 ;
    wire new_AGEMA_signal_6499 ;
    wire new_AGEMA_signal_6500 ;
    wire new_AGEMA_signal_6501 ;
    wire new_AGEMA_signal_6502 ;
    wire new_AGEMA_signal_6503 ;
    wire new_AGEMA_signal_6504 ;
    wire new_AGEMA_signal_6505 ;
    wire new_AGEMA_signal_6506 ;
    wire new_AGEMA_signal_6507 ;
    wire new_AGEMA_signal_6508 ;
    wire new_AGEMA_signal_6509 ;
    wire new_AGEMA_signal_6510 ;
    wire new_AGEMA_signal_6511 ;
    wire new_AGEMA_signal_6512 ;
    wire new_AGEMA_signal_6513 ;
    wire new_AGEMA_signal_6514 ;
    wire new_AGEMA_signal_6515 ;
    wire new_AGEMA_signal_6516 ;
    wire new_AGEMA_signal_6517 ;
    wire new_AGEMA_signal_6518 ;
    wire new_AGEMA_signal_6519 ;
    wire new_AGEMA_signal_6520 ;
    wire new_AGEMA_signal_6521 ;
    wire new_AGEMA_signal_6522 ;
    wire new_AGEMA_signal_6523 ;
    wire new_AGEMA_signal_6524 ;
    wire new_AGEMA_signal_6525 ;
    wire new_AGEMA_signal_6526 ;
    wire new_AGEMA_signal_6527 ;
    wire new_AGEMA_signal_6528 ;
    wire new_AGEMA_signal_6529 ;
    wire new_AGEMA_signal_6530 ;
    wire new_AGEMA_signal_6531 ;
    wire new_AGEMA_signal_6532 ;
    wire new_AGEMA_signal_6533 ;
    wire new_AGEMA_signal_6534 ;
    wire new_AGEMA_signal_6535 ;
    wire new_AGEMA_signal_6536 ;
    wire new_AGEMA_signal_6537 ;
    wire new_AGEMA_signal_6538 ;
    wire new_AGEMA_signal_6539 ;
    wire new_AGEMA_signal_6540 ;
    wire new_AGEMA_signal_6541 ;
    wire new_AGEMA_signal_6542 ;
    wire new_AGEMA_signal_6543 ;
    wire new_AGEMA_signal_6544 ;
    wire new_AGEMA_signal_6545 ;
    wire new_AGEMA_signal_6546 ;
    wire new_AGEMA_signal_6547 ;
    wire new_AGEMA_signal_6548 ;
    wire new_AGEMA_signal_6549 ;
    wire new_AGEMA_signal_6550 ;
    wire new_AGEMA_signal_6551 ;
    wire new_AGEMA_signal_6552 ;
    wire new_AGEMA_signal_6553 ;
    wire new_AGEMA_signal_6554 ;
    wire new_AGEMA_signal_6555 ;
    wire new_AGEMA_signal_6556 ;
    wire new_AGEMA_signal_6557 ;
    wire new_AGEMA_signal_6558 ;
    wire new_AGEMA_signal_6559 ;
    wire new_AGEMA_signal_6560 ;
    wire new_AGEMA_signal_6561 ;
    wire new_AGEMA_signal_6562 ;
    wire new_AGEMA_signal_6563 ;
    wire new_AGEMA_signal_6564 ;
    wire new_AGEMA_signal_6565 ;
    wire new_AGEMA_signal_6566 ;
    wire new_AGEMA_signal_6567 ;
    wire new_AGEMA_signal_6568 ;
    wire new_AGEMA_signal_6569 ;
    wire new_AGEMA_signal_6570 ;
    wire new_AGEMA_signal_6571 ;
    wire new_AGEMA_signal_6572 ;
    wire new_AGEMA_signal_6573 ;
    wire new_AGEMA_signal_6574 ;
    wire new_AGEMA_signal_6575 ;
    wire new_AGEMA_signal_6576 ;
    wire new_AGEMA_signal_6577 ;
    wire new_AGEMA_signal_6578 ;
    wire new_AGEMA_signal_6579 ;
    wire new_AGEMA_signal_6580 ;
    wire new_AGEMA_signal_6581 ;
    wire new_AGEMA_signal_6582 ;
    wire new_AGEMA_signal_6583 ;
    wire new_AGEMA_signal_6584 ;
    wire new_AGEMA_signal_6585 ;
    wire new_AGEMA_signal_6586 ;
    wire new_AGEMA_signal_6587 ;
    wire new_AGEMA_signal_6588 ;
    wire new_AGEMA_signal_6589 ;
    wire new_AGEMA_signal_6590 ;
    wire new_AGEMA_signal_6591 ;
    wire new_AGEMA_signal_6592 ;
    wire new_AGEMA_signal_6593 ;
    wire new_AGEMA_signal_6594 ;
    wire new_AGEMA_signal_6595 ;
    wire new_AGEMA_signal_6596 ;
    wire new_AGEMA_signal_6597 ;
    wire new_AGEMA_signal_6598 ;
    wire new_AGEMA_signal_6599 ;
    wire new_AGEMA_signal_6600 ;
    wire new_AGEMA_signal_6601 ;
    wire new_AGEMA_signal_6602 ;
    wire new_AGEMA_signal_6603 ;
    wire new_AGEMA_signal_6604 ;
    wire new_AGEMA_signal_6605 ;
    wire new_AGEMA_signal_6606 ;
    wire new_AGEMA_signal_6607 ;
    wire new_AGEMA_signal_6608 ;
    wire new_AGEMA_signal_6609 ;
    wire new_AGEMA_signal_6610 ;
    wire new_AGEMA_signal_6611 ;
    wire new_AGEMA_signal_6612 ;
    wire new_AGEMA_signal_6613 ;
    wire new_AGEMA_signal_6614 ;
    wire new_AGEMA_signal_6615 ;
    wire new_AGEMA_signal_6616 ;
    wire new_AGEMA_signal_6617 ;
    wire new_AGEMA_signal_6618 ;
    wire new_AGEMA_signal_6619 ;
    wire new_AGEMA_signal_6620 ;
    wire new_AGEMA_signal_6621 ;
    wire new_AGEMA_signal_6622 ;
    wire new_AGEMA_signal_6623 ;
    wire new_AGEMA_signal_6624 ;
    wire new_AGEMA_signal_6625 ;
    wire new_AGEMA_signal_6626 ;
    wire new_AGEMA_signal_6627 ;
    wire new_AGEMA_signal_6628 ;
    wire new_AGEMA_signal_6629 ;
    wire new_AGEMA_signal_6630 ;
    wire new_AGEMA_signal_6631 ;
    wire new_AGEMA_signal_6632 ;
    wire new_AGEMA_signal_6633 ;
    wire new_AGEMA_signal_6634 ;
    wire new_AGEMA_signal_6635 ;
    wire new_AGEMA_signal_6636 ;
    wire new_AGEMA_signal_6637 ;
    wire new_AGEMA_signal_6638 ;
    wire new_AGEMA_signal_6639 ;
    wire new_AGEMA_signal_6640 ;
    wire new_AGEMA_signal_6641 ;
    wire new_AGEMA_signal_6642 ;
    wire new_AGEMA_signal_6643 ;
    wire new_AGEMA_signal_6644 ;
    wire new_AGEMA_signal_6645 ;
    wire new_AGEMA_signal_6646 ;
    wire new_AGEMA_signal_6647 ;
    wire new_AGEMA_signal_6648 ;
    wire new_AGEMA_signal_6649 ;
    wire new_AGEMA_signal_6650 ;
    wire new_AGEMA_signal_6651 ;
    wire new_AGEMA_signal_6652 ;
    wire new_AGEMA_signal_6653 ;
    wire new_AGEMA_signal_6654 ;
    wire new_AGEMA_signal_6655 ;
    wire new_AGEMA_signal_6656 ;
    wire new_AGEMA_signal_6657 ;
    wire new_AGEMA_signal_6658 ;
    wire new_AGEMA_signal_6659 ;
    wire new_AGEMA_signal_6660 ;
    wire new_AGEMA_signal_6661 ;
    wire new_AGEMA_signal_6662 ;
    wire new_AGEMA_signal_6663 ;
    wire new_AGEMA_signal_6664 ;
    wire new_AGEMA_signal_6665 ;
    wire new_AGEMA_signal_6666 ;
    wire new_AGEMA_signal_6667 ;
    wire new_AGEMA_signal_6668 ;
    wire new_AGEMA_signal_6669 ;
    wire new_AGEMA_signal_6670 ;
    wire new_AGEMA_signal_6671 ;
    wire new_AGEMA_signal_6672 ;
    wire new_AGEMA_signal_6673 ;
    wire new_AGEMA_signal_6674 ;
    wire new_AGEMA_signal_6675 ;
    wire new_AGEMA_signal_6676 ;
    wire new_AGEMA_signal_6677 ;
    wire new_AGEMA_signal_6678 ;
    wire new_AGEMA_signal_6679 ;
    wire new_AGEMA_signal_6680 ;
    wire new_AGEMA_signal_6681 ;
    wire new_AGEMA_signal_6682 ;
    wire new_AGEMA_signal_6683 ;
    wire new_AGEMA_signal_6684 ;
    wire new_AGEMA_signal_6685 ;
    wire new_AGEMA_signal_6686 ;
    wire new_AGEMA_signal_6687 ;
    wire new_AGEMA_signal_6688 ;
    wire new_AGEMA_signal_6689 ;
    wire new_AGEMA_signal_6690 ;
    wire new_AGEMA_signal_6691 ;
    wire new_AGEMA_signal_6692 ;
    wire new_AGEMA_signal_6693 ;
    wire new_AGEMA_signal_6694 ;
    wire new_AGEMA_signal_6695 ;
    wire new_AGEMA_signal_6696 ;
    wire new_AGEMA_signal_6697 ;
    wire new_AGEMA_signal_6698 ;
    wire new_AGEMA_signal_6699 ;
    wire new_AGEMA_signal_6700 ;
    wire new_AGEMA_signal_6701 ;
    wire new_AGEMA_signal_6702 ;
    wire new_AGEMA_signal_6703 ;
    wire new_AGEMA_signal_6704 ;
    wire new_AGEMA_signal_6705 ;
    wire new_AGEMA_signal_6706 ;
    wire new_AGEMA_signal_6707 ;
    wire new_AGEMA_signal_6708 ;
    wire new_AGEMA_signal_6709 ;
    wire new_AGEMA_signal_6710 ;
    wire new_AGEMA_signal_6711 ;
    wire new_AGEMA_signal_6712 ;
    wire new_AGEMA_signal_6713 ;
    wire new_AGEMA_signal_6714 ;
    wire new_AGEMA_signal_6715 ;
    wire new_AGEMA_signal_6716 ;
    wire new_AGEMA_signal_6717 ;
    wire new_AGEMA_signal_6718 ;
    wire new_AGEMA_signal_6719 ;
    wire new_AGEMA_signal_6720 ;
    wire new_AGEMA_signal_6721 ;
    wire new_AGEMA_signal_6722 ;
    wire new_AGEMA_signal_6723 ;
    wire new_AGEMA_signal_6724 ;
    wire new_AGEMA_signal_6725 ;
    wire new_AGEMA_signal_6726 ;
    wire new_AGEMA_signal_6727 ;
    wire new_AGEMA_signal_6728 ;
    wire new_AGEMA_signal_6729 ;
    wire new_AGEMA_signal_6730 ;
    wire new_AGEMA_signal_6731 ;
    wire new_AGEMA_signal_6732 ;
    wire new_AGEMA_signal_6733 ;
    wire new_AGEMA_signal_6734 ;
    wire new_AGEMA_signal_6735 ;
    wire new_AGEMA_signal_6736 ;
    wire new_AGEMA_signal_6737 ;
    wire new_AGEMA_signal_6738 ;
    wire new_AGEMA_signal_6739 ;
    wire new_AGEMA_signal_6740 ;
    wire new_AGEMA_signal_6741 ;
    wire new_AGEMA_signal_6742 ;
    wire new_AGEMA_signal_6743 ;
    wire new_AGEMA_signal_6744 ;
    wire new_AGEMA_signal_6745 ;
    wire new_AGEMA_signal_6746 ;
    wire new_AGEMA_signal_6747 ;
    wire new_AGEMA_signal_6748 ;
    wire new_AGEMA_signal_6749 ;
    wire new_AGEMA_signal_6750 ;
    wire new_AGEMA_signal_6751 ;
    wire new_AGEMA_signal_6752 ;
    wire new_AGEMA_signal_6753 ;
    wire new_AGEMA_signal_6754 ;
    wire new_AGEMA_signal_6755 ;
    wire new_AGEMA_signal_6756 ;
    wire new_AGEMA_signal_6757 ;
    wire new_AGEMA_signal_6758 ;
    wire new_AGEMA_signal_6759 ;
    wire new_AGEMA_signal_6760 ;
    wire new_AGEMA_signal_6761 ;
    wire new_AGEMA_signal_6762 ;
    wire new_AGEMA_signal_6763 ;
    wire new_AGEMA_signal_6764 ;
    wire new_AGEMA_signal_6765 ;
    wire new_AGEMA_signal_6766 ;
    wire new_AGEMA_signal_6767 ;
    wire new_AGEMA_signal_6768 ;
    wire new_AGEMA_signal_6769 ;
    wire new_AGEMA_signal_6770 ;
    wire new_AGEMA_signal_6771 ;
    wire new_AGEMA_signal_6772 ;
    wire new_AGEMA_signal_6773 ;
    wire new_AGEMA_signal_6774 ;
    wire new_AGEMA_signal_6775 ;
    wire new_AGEMA_signal_6776 ;
    wire new_AGEMA_signal_6777 ;
    wire new_AGEMA_signal_6778 ;
    wire new_AGEMA_signal_6779 ;
    wire new_AGEMA_signal_6780 ;
    wire new_AGEMA_signal_6781 ;
    wire new_AGEMA_signal_6782 ;
    wire new_AGEMA_signal_6783 ;
    wire new_AGEMA_signal_6784 ;
    wire new_AGEMA_signal_6785 ;
    wire new_AGEMA_signal_6786 ;
    wire new_AGEMA_signal_6787 ;
    wire new_AGEMA_signal_6788 ;
    wire new_AGEMA_signal_6789 ;
    wire new_AGEMA_signal_6790 ;
    wire new_AGEMA_signal_6791 ;
    wire new_AGEMA_signal_6792 ;
    wire new_AGEMA_signal_6793 ;
    wire new_AGEMA_signal_6794 ;
    wire new_AGEMA_signal_6795 ;
    wire new_AGEMA_signal_6796 ;
    wire new_AGEMA_signal_6797 ;
    wire new_AGEMA_signal_6798 ;
    wire new_AGEMA_signal_6799 ;
    wire new_AGEMA_signal_6800 ;
    wire new_AGEMA_signal_6801 ;
    wire new_AGEMA_signal_6802 ;
    wire new_AGEMA_signal_6803 ;
    wire new_AGEMA_signal_6804 ;
    wire new_AGEMA_signal_6805 ;
    wire new_AGEMA_signal_6806 ;
    wire new_AGEMA_signal_6807 ;
    wire new_AGEMA_signal_6808 ;
    wire new_AGEMA_signal_6809 ;
    wire new_AGEMA_signal_6810 ;
    wire new_AGEMA_signal_6811 ;
    wire new_AGEMA_signal_6812 ;
    wire new_AGEMA_signal_6813 ;
    wire new_AGEMA_signal_6814 ;
    wire new_AGEMA_signal_6815 ;
    wire new_AGEMA_signal_6816 ;
    wire new_AGEMA_signal_6817 ;
    wire new_AGEMA_signal_6818 ;
    wire new_AGEMA_signal_6819 ;
    wire new_AGEMA_signal_6820 ;
    wire new_AGEMA_signal_6821 ;
    wire new_AGEMA_signal_6822 ;
    wire new_AGEMA_signal_6823 ;
    wire new_AGEMA_signal_6824 ;
    wire new_AGEMA_signal_6825 ;
    wire new_AGEMA_signal_6826 ;
    wire new_AGEMA_signal_6827 ;
    wire new_AGEMA_signal_6828 ;
    wire new_AGEMA_signal_6829 ;
    wire new_AGEMA_signal_6830 ;
    wire new_AGEMA_signal_6831 ;
    wire new_AGEMA_signal_6832 ;
    wire new_AGEMA_signal_6833 ;
    wire new_AGEMA_signal_6834 ;
    wire new_AGEMA_signal_6835 ;
    wire new_AGEMA_signal_6836 ;
    wire new_AGEMA_signal_6837 ;
    wire new_AGEMA_signal_6838 ;
    wire new_AGEMA_signal_6839 ;
    wire new_AGEMA_signal_6840 ;
    wire new_AGEMA_signal_6841 ;
    wire new_AGEMA_signal_6842 ;
    wire new_AGEMA_signal_6843 ;
    wire new_AGEMA_signal_6844 ;
    wire new_AGEMA_signal_6845 ;
    wire new_AGEMA_signal_6846 ;
    wire new_AGEMA_signal_6847 ;
    wire new_AGEMA_signal_6848 ;
    wire new_AGEMA_signal_6849 ;
    wire new_AGEMA_signal_6850 ;
    wire new_AGEMA_signal_6851 ;
    wire new_AGEMA_signal_6852 ;
    wire new_AGEMA_signal_6853 ;
    wire new_AGEMA_signal_6854 ;
    wire new_AGEMA_signal_6855 ;
    wire new_AGEMA_signal_6856 ;
    wire new_AGEMA_signal_6857 ;
    wire new_AGEMA_signal_6858 ;
    wire new_AGEMA_signal_6859 ;
    wire new_AGEMA_signal_6860 ;
    wire new_AGEMA_signal_6861 ;
    wire new_AGEMA_signal_6862 ;
    wire new_AGEMA_signal_6863 ;
    wire new_AGEMA_signal_6864 ;
    wire new_AGEMA_signal_6865 ;
    wire new_AGEMA_signal_6866 ;
    wire new_AGEMA_signal_6867 ;
    wire new_AGEMA_signal_6868 ;
    wire new_AGEMA_signal_6869 ;
    wire new_AGEMA_signal_6870 ;
    wire new_AGEMA_signal_6871 ;
    wire new_AGEMA_signal_6872 ;
    wire new_AGEMA_signal_6873 ;
    wire new_AGEMA_signal_6874 ;
    wire new_AGEMA_signal_6875 ;
    wire new_AGEMA_signal_6876 ;
    wire new_AGEMA_signal_6877 ;
    wire new_AGEMA_signal_6878 ;
    wire new_AGEMA_signal_6879 ;
    wire new_AGEMA_signal_6880 ;
    wire new_AGEMA_signal_6881 ;
    wire new_AGEMA_signal_6882 ;
    wire new_AGEMA_signal_6883 ;
    wire new_AGEMA_signal_6884 ;
    wire new_AGEMA_signal_6885 ;
    wire new_AGEMA_signal_6886 ;
    wire new_AGEMA_signal_6887 ;
    wire new_AGEMA_signal_6888 ;
    wire new_AGEMA_signal_6889 ;
    wire new_AGEMA_signal_6890 ;
    wire new_AGEMA_signal_6891 ;
    wire new_AGEMA_signal_6892 ;
    wire new_AGEMA_signal_6893 ;
    wire new_AGEMA_signal_6894 ;
    wire new_AGEMA_signal_6895 ;
    wire new_AGEMA_signal_6896 ;
    wire new_AGEMA_signal_6897 ;
    wire new_AGEMA_signal_6898 ;
    wire new_AGEMA_signal_6899 ;
    wire new_AGEMA_signal_6900 ;
    wire new_AGEMA_signal_6901 ;
    wire new_AGEMA_signal_6902 ;
    wire new_AGEMA_signal_6903 ;
    wire new_AGEMA_signal_6904 ;
    wire new_AGEMA_signal_6905 ;
    wire new_AGEMA_signal_6906 ;
    wire new_AGEMA_signal_6907 ;
    wire new_AGEMA_signal_6908 ;
    wire new_AGEMA_signal_6909 ;
    wire new_AGEMA_signal_6910 ;
    wire new_AGEMA_signal_6911 ;
    wire new_AGEMA_signal_6912 ;
    wire new_AGEMA_signal_6913 ;
    wire new_AGEMA_signal_6914 ;
    wire new_AGEMA_signal_6915 ;
    wire new_AGEMA_signal_6916 ;
    wire new_AGEMA_signal_6917 ;
    wire new_AGEMA_signal_6918 ;
    wire new_AGEMA_signal_6919 ;
    wire new_AGEMA_signal_6920 ;
    wire new_AGEMA_signal_6921 ;
    wire new_AGEMA_signal_6922 ;
    wire new_AGEMA_signal_6923 ;
    wire new_AGEMA_signal_6924 ;
    wire new_AGEMA_signal_6925 ;
    wire new_AGEMA_signal_6926 ;
    wire new_AGEMA_signal_6927 ;
    wire new_AGEMA_signal_6928 ;
    wire new_AGEMA_signal_6929 ;
    wire new_AGEMA_signal_6930 ;
    wire new_AGEMA_signal_6931 ;
    wire new_AGEMA_signal_6932 ;
    wire new_AGEMA_signal_6933 ;
    wire new_AGEMA_signal_6934 ;
    wire new_AGEMA_signal_6935 ;
    wire new_AGEMA_signal_6936 ;
    wire new_AGEMA_signal_6937 ;
    wire new_AGEMA_signal_6938 ;
    wire new_AGEMA_signal_6939 ;
    wire new_AGEMA_signal_6940 ;
    wire new_AGEMA_signal_6941 ;
    wire new_AGEMA_signal_6942 ;
    wire new_AGEMA_signal_6943 ;
    wire new_AGEMA_signal_6944 ;
    wire new_AGEMA_signal_6945 ;
    wire new_AGEMA_signal_6946 ;
    wire new_AGEMA_signal_6947 ;
    wire new_AGEMA_signal_6948 ;
    wire new_AGEMA_signal_6949 ;
    wire new_AGEMA_signal_6950 ;
    wire new_AGEMA_signal_6951 ;
    wire new_AGEMA_signal_6952 ;
    wire new_AGEMA_signal_6953 ;
    wire new_AGEMA_signal_6954 ;
    wire new_AGEMA_signal_6955 ;
    wire new_AGEMA_signal_6956 ;
    wire new_AGEMA_signal_6957 ;
    wire new_AGEMA_signal_6958 ;
    wire new_AGEMA_signal_6959 ;
    wire new_AGEMA_signal_6960 ;
    wire new_AGEMA_signal_6961 ;
    wire new_AGEMA_signal_6962 ;
    wire new_AGEMA_signal_6963 ;
    wire new_AGEMA_signal_6964 ;
    wire new_AGEMA_signal_6965 ;
    wire new_AGEMA_signal_6966 ;
    wire new_AGEMA_signal_6967 ;
    wire new_AGEMA_signal_6968 ;
    wire new_AGEMA_signal_6969 ;
    wire new_AGEMA_signal_6970 ;
    wire new_AGEMA_signal_6971 ;
    wire new_AGEMA_signal_6972 ;
    wire new_AGEMA_signal_6973 ;
    wire new_AGEMA_signal_6974 ;
    wire new_AGEMA_signal_6975 ;
    wire new_AGEMA_signal_6976 ;
    wire new_AGEMA_signal_6977 ;
    wire new_AGEMA_signal_6978 ;
    wire new_AGEMA_signal_6979 ;
    wire new_AGEMA_signal_6980 ;
    wire new_AGEMA_signal_6981 ;
    wire new_AGEMA_signal_6982 ;
    wire new_AGEMA_signal_6983 ;
    wire new_AGEMA_signal_6984 ;
    wire new_AGEMA_signal_6985 ;
    wire new_AGEMA_signal_6986 ;
    wire new_AGEMA_signal_6987 ;
    wire new_AGEMA_signal_6988 ;
    wire new_AGEMA_signal_6989 ;
    wire new_AGEMA_signal_6990 ;
    wire new_AGEMA_signal_6991 ;
    wire new_AGEMA_signal_6992 ;
    wire new_AGEMA_signal_6993 ;
    wire new_AGEMA_signal_6994 ;
    wire new_AGEMA_signal_6995 ;
    wire new_AGEMA_signal_6996 ;
    wire new_AGEMA_signal_6997 ;
    wire new_AGEMA_signal_6998 ;
    wire new_AGEMA_signal_6999 ;
    wire new_AGEMA_signal_7000 ;
    wire new_AGEMA_signal_7001 ;
    wire new_AGEMA_signal_7002 ;
    wire new_AGEMA_signal_7003 ;
    wire new_AGEMA_signal_7004 ;
    wire new_AGEMA_signal_7005 ;
    wire new_AGEMA_signal_7006 ;
    wire new_AGEMA_signal_7007 ;
    wire new_AGEMA_signal_7008 ;
    wire new_AGEMA_signal_7009 ;
    wire new_AGEMA_signal_7010 ;
    wire new_AGEMA_signal_7011 ;
    wire new_AGEMA_signal_7012 ;
    wire new_AGEMA_signal_7013 ;
    wire new_AGEMA_signal_7014 ;
    wire new_AGEMA_signal_7015 ;
    wire new_AGEMA_signal_7016 ;
    wire new_AGEMA_signal_7017 ;
    wire new_AGEMA_signal_7018 ;
    wire new_AGEMA_signal_7019 ;
    wire new_AGEMA_signal_7020 ;
    wire new_AGEMA_signal_7021 ;
    wire new_AGEMA_signal_7022 ;
    wire new_AGEMA_signal_7023 ;
    wire new_AGEMA_signal_7024 ;
    wire new_AGEMA_signal_7025 ;
    wire new_AGEMA_signal_7026 ;
    wire new_AGEMA_signal_7027 ;
    wire new_AGEMA_signal_7028 ;
    wire new_AGEMA_signal_7029 ;
    wire new_AGEMA_signal_7030 ;
    wire new_AGEMA_signal_7031 ;
    wire new_AGEMA_signal_7032 ;
    wire new_AGEMA_signal_7033 ;
    wire new_AGEMA_signal_7034 ;
    wire new_AGEMA_signal_7035 ;
    wire new_AGEMA_signal_7036 ;
    wire new_AGEMA_signal_7037 ;
    wire new_AGEMA_signal_7038 ;
    wire new_AGEMA_signal_7039 ;
    wire new_AGEMA_signal_7040 ;
    wire new_AGEMA_signal_7041 ;
    wire new_AGEMA_signal_7042 ;
    wire new_AGEMA_signal_7043 ;
    wire new_AGEMA_signal_7044 ;
    wire new_AGEMA_signal_7045 ;
    wire new_AGEMA_signal_7046 ;
    wire new_AGEMA_signal_7047 ;
    wire new_AGEMA_signal_7048 ;
    wire new_AGEMA_signal_7049 ;
    wire new_AGEMA_signal_7050 ;
    wire new_AGEMA_signal_7051 ;
    wire new_AGEMA_signal_7052 ;
    wire new_AGEMA_signal_7053 ;
    wire new_AGEMA_signal_7054 ;
    wire new_AGEMA_signal_7055 ;
    wire new_AGEMA_signal_7056 ;
    wire new_AGEMA_signal_7057 ;
    wire new_AGEMA_signal_7058 ;
    wire new_AGEMA_signal_7059 ;
    wire new_AGEMA_signal_7060 ;
    wire new_AGEMA_signal_7061 ;
    wire new_AGEMA_signal_7062 ;
    wire new_AGEMA_signal_7063 ;
    wire new_AGEMA_signal_7064 ;
    wire new_AGEMA_signal_7065 ;
    wire new_AGEMA_signal_7066 ;
    wire new_AGEMA_signal_7067 ;
    wire new_AGEMA_signal_7068 ;
    wire new_AGEMA_signal_7069 ;
    wire new_AGEMA_signal_7070 ;
    wire new_AGEMA_signal_7071 ;
    wire new_AGEMA_signal_7072 ;
    wire new_AGEMA_signal_7073 ;
    wire new_AGEMA_signal_7074 ;
    wire new_AGEMA_signal_7075 ;
    wire new_AGEMA_signal_7076 ;
    wire new_AGEMA_signal_7077 ;
    wire new_AGEMA_signal_7078 ;
    wire new_AGEMA_signal_7079 ;
    wire new_AGEMA_signal_7080 ;
    wire new_AGEMA_signal_7081 ;
    wire new_AGEMA_signal_7082 ;
    wire new_AGEMA_signal_7083 ;
    wire new_AGEMA_signal_7084 ;
    wire new_AGEMA_signal_7085 ;
    wire new_AGEMA_signal_7086 ;
    wire new_AGEMA_signal_7087 ;
    wire new_AGEMA_signal_7088 ;
    wire new_AGEMA_signal_7089 ;
    wire new_AGEMA_signal_7090 ;
    wire new_AGEMA_signal_7091 ;
    wire new_AGEMA_signal_7092 ;
    wire new_AGEMA_signal_7093 ;
    wire new_AGEMA_signal_7094 ;
    wire new_AGEMA_signal_7095 ;
    wire new_AGEMA_signal_7096 ;
    wire new_AGEMA_signal_7097 ;
    wire new_AGEMA_signal_7098 ;
    wire new_AGEMA_signal_7099 ;
    wire new_AGEMA_signal_7100 ;
    wire new_AGEMA_signal_7101 ;
    wire new_AGEMA_signal_7102 ;
    wire new_AGEMA_signal_7103 ;
    wire new_AGEMA_signal_7104 ;
    wire new_AGEMA_signal_7105 ;
    wire new_AGEMA_signal_7106 ;
    wire new_AGEMA_signal_7107 ;
    wire new_AGEMA_signal_7108 ;
    wire new_AGEMA_signal_7109 ;
    wire new_AGEMA_signal_7110 ;
    wire new_AGEMA_signal_7111 ;
    wire new_AGEMA_signal_7112 ;
    wire new_AGEMA_signal_7113 ;
    wire new_AGEMA_signal_7114 ;
    wire new_AGEMA_signal_7115 ;
    wire new_AGEMA_signal_7116 ;
    wire new_AGEMA_signal_7117 ;
    wire new_AGEMA_signal_7118 ;
    wire new_AGEMA_signal_7119 ;
    wire new_AGEMA_signal_7120 ;
    wire new_AGEMA_signal_7121 ;
    wire new_AGEMA_signal_7122 ;
    wire new_AGEMA_signal_7123 ;
    wire new_AGEMA_signal_7124 ;
    wire new_AGEMA_signal_7125 ;
    wire new_AGEMA_signal_7126 ;
    wire new_AGEMA_signal_7127 ;
    wire new_AGEMA_signal_7128 ;
    wire new_AGEMA_signal_7129 ;
    wire new_AGEMA_signal_7130 ;
    wire new_AGEMA_signal_7131 ;
    wire new_AGEMA_signal_7132 ;
    wire new_AGEMA_signal_7133 ;
    wire new_AGEMA_signal_7134 ;
    wire new_AGEMA_signal_7135 ;
    wire new_AGEMA_signal_7136 ;
    wire new_AGEMA_signal_7137 ;
    wire new_AGEMA_signal_7138 ;
    wire new_AGEMA_signal_7139 ;
    wire new_AGEMA_signal_7140 ;
    wire new_AGEMA_signal_7141 ;
    wire new_AGEMA_signal_7142 ;
    wire new_AGEMA_signal_7143 ;
    wire new_AGEMA_signal_7144 ;
    wire new_AGEMA_signal_7145 ;
    wire new_AGEMA_signal_7146 ;
    wire new_AGEMA_signal_7147 ;
    wire new_AGEMA_signal_7148 ;
    wire new_AGEMA_signal_7149 ;
    wire new_AGEMA_signal_7150 ;
    wire new_AGEMA_signal_7151 ;
    wire new_AGEMA_signal_7152 ;
    wire new_AGEMA_signal_7153 ;
    wire new_AGEMA_signal_7154 ;
    wire new_AGEMA_signal_7155 ;
    wire new_AGEMA_signal_7156 ;
    wire new_AGEMA_signal_7157 ;
    wire new_AGEMA_signal_7158 ;
    wire new_AGEMA_signal_7159 ;
    wire new_AGEMA_signal_7160 ;
    wire new_AGEMA_signal_7161 ;
    wire new_AGEMA_signal_7162 ;
    wire new_AGEMA_signal_7163 ;
    wire new_AGEMA_signal_7164 ;
    wire new_AGEMA_signal_7165 ;
    wire new_AGEMA_signal_7166 ;
    wire new_AGEMA_signal_7167 ;
    wire new_AGEMA_signal_7168 ;
    wire new_AGEMA_signal_7169 ;
    wire new_AGEMA_signal_7170 ;
    wire new_AGEMA_signal_7171 ;
    wire new_AGEMA_signal_7172 ;
    wire new_AGEMA_signal_7173 ;
    wire new_AGEMA_signal_7174 ;
    wire new_AGEMA_signal_7175 ;
    wire new_AGEMA_signal_7176 ;
    wire new_AGEMA_signal_7177 ;
    wire new_AGEMA_signal_7178 ;
    wire new_AGEMA_signal_7179 ;
    wire new_AGEMA_signal_7180 ;
    wire new_AGEMA_signal_7181 ;
    wire new_AGEMA_signal_7182 ;
    wire new_AGEMA_signal_7183 ;
    wire new_AGEMA_signal_7184 ;
    wire new_AGEMA_signal_7185 ;
    wire new_AGEMA_signal_7186 ;
    wire new_AGEMA_signal_7187 ;
    wire new_AGEMA_signal_7188 ;
    wire new_AGEMA_signal_7189 ;
    wire new_AGEMA_signal_7190 ;
    wire new_AGEMA_signal_7191 ;
    wire new_AGEMA_signal_7192 ;
    wire new_AGEMA_signal_7193 ;
    wire new_AGEMA_signal_7194 ;
    wire new_AGEMA_signal_7195 ;
    wire new_AGEMA_signal_7196 ;
    wire new_AGEMA_signal_7197 ;
    wire new_AGEMA_signal_7198 ;
    wire new_AGEMA_signal_7199 ;
    wire new_AGEMA_signal_7200 ;
    wire new_AGEMA_signal_7201 ;
    wire new_AGEMA_signal_7202 ;
    wire new_AGEMA_signal_7203 ;
    wire new_AGEMA_signal_7204 ;
    wire new_AGEMA_signal_7205 ;
    wire new_AGEMA_signal_7206 ;
    wire new_AGEMA_signal_7207 ;
    wire new_AGEMA_signal_7208 ;
    wire new_AGEMA_signal_7209 ;
    wire new_AGEMA_signal_7210 ;
    wire new_AGEMA_signal_7211 ;
    wire new_AGEMA_signal_7212 ;
    wire new_AGEMA_signal_7213 ;
    wire new_AGEMA_signal_7214 ;
    wire new_AGEMA_signal_7215 ;
    wire new_AGEMA_signal_7216 ;
    wire new_AGEMA_signal_7217 ;
    wire new_AGEMA_signal_7218 ;
    wire new_AGEMA_signal_7219 ;
    wire new_AGEMA_signal_7220 ;
    wire new_AGEMA_signal_7221 ;
    wire new_AGEMA_signal_7222 ;
    wire new_AGEMA_signal_7223 ;
    wire new_AGEMA_signal_7224 ;
    wire new_AGEMA_signal_7225 ;
    wire new_AGEMA_signal_7226 ;
    wire new_AGEMA_signal_7227 ;
    wire new_AGEMA_signal_7228 ;
    wire new_AGEMA_signal_7229 ;
    wire new_AGEMA_signal_7230 ;
    wire new_AGEMA_signal_7231 ;
    wire new_AGEMA_signal_7232 ;
    wire new_AGEMA_signal_7233 ;
    wire new_AGEMA_signal_7234 ;
    wire new_AGEMA_signal_7235 ;
    wire new_AGEMA_signal_7236 ;
    wire new_AGEMA_signal_7237 ;
    wire new_AGEMA_signal_7238 ;
    wire new_AGEMA_signal_7239 ;
    wire new_AGEMA_signal_7240 ;
    wire new_AGEMA_signal_7241 ;
    wire new_AGEMA_signal_7242 ;
    wire new_AGEMA_signal_7243 ;
    wire new_AGEMA_signal_7244 ;
    wire new_AGEMA_signal_7245 ;
    wire new_AGEMA_signal_7246 ;
    wire new_AGEMA_signal_7247 ;
    wire new_AGEMA_signal_7248 ;
    wire new_AGEMA_signal_7249 ;
    wire new_AGEMA_signal_7250 ;
    wire new_AGEMA_signal_7251 ;
    wire new_AGEMA_signal_7252 ;
    wire new_AGEMA_signal_7253 ;
    wire new_AGEMA_signal_7254 ;
    wire new_AGEMA_signal_7255 ;
    wire new_AGEMA_signal_7256 ;
    wire new_AGEMA_signal_7257 ;
    wire new_AGEMA_signal_7258 ;
    wire new_AGEMA_signal_7259 ;
    wire new_AGEMA_signal_7260 ;
    wire new_AGEMA_signal_7261 ;
    wire new_AGEMA_signal_7262 ;
    wire new_AGEMA_signal_7263 ;
    wire new_AGEMA_signal_7264 ;
    wire new_AGEMA_signal_7265 ;
    wire new_AGEMA_signal_7266 ;
    wire new_AGEMA_signal_7267 ;
    wire new_AGEMA_signal_7268 ;
    wire new_AGEMA_signal_7269 ;
    wire new_AGEMA_signal_7270 ;
    wire new_AGEMA_signal_7271 ;
    wire new_AGEMA_signal_7272 ;
    wire new_AGEMA_signal_7273 ;
    wire new_AGEMA_signal_7274 ;
    wire new_AGEMA_signal_7275 ;
    wire new_AGEMA_signal_7276 ;
    wire new_AGEMA_signal_7277 ;
    wire new_AGEMA_signal_7278 ;
    wire new_AGEMA_signal_7279 ;
    wire new_AGEMA_signal_7280 ;
    wire new_AGEMA_signal_7281 ;
    wire new_AGEMA_signal_7282 ;
    wire new_AGEMA_signal_7283 ;
    wire new_AGEMA_signal_7284 ;
    wire new_AGEMA_signal_7285 ;
    wire new_AGEMA_signal_7286 ;
    wire new_AGEMA_signal_7287 ;
    wire new_AGEMA_signal_7288 ;
    wire new_AGEMA_signal_7289 ;
    wire new_AGEMA_signal_7290 ;
    wire new_AGEMA_signal_7291 ;
    wire new_AGEMA_signal_7292 ;
    wire new_AGEMA_signal_7293 ;
    wire new_AGEMA_signal_7294 ;
    wire new_AGEMA_signal_7295 ;
    wire new_AGEMA_signal_7296 ;
    wire new_AGEMA_signal_7297 ;
    wire new_AGEMA_signal_7298 ;
    wire new_AGEMA_signal_7299 ;
    wire new_AGEMA_signal_7300 ;
    wire new_AGEMA_signal_7301 ;
    wire new_AGEMA_signal_7302 ;
    wire new_AGEMA_signal_7303 ;
    wire new_AGEMA_signal_7304 ;
    wire new_AGEMA_signal_7305 ;
    wire new_AGEMA_signal_7306 ;
    wire new_AGEMA_signal_7307 ;
    wire new_AGEMA_signal_7308 ;
    wire new_AGEMA_signal_7309 ;
    wire new_AGEMA_signal_7310 ;
    wire new_AGEMA_signal_7311 ;
    wire new_AGEMA_signal_7312 ;
    wire new_AGEMA_signal_7313 ;
    wire new_AGEMA_signal_7314 ;
    wire new_AGEMA_signal_7315 ;
    wire new_AGEMA_signal_7316 ;
    wire new_AGEMA_signal_7317 ;
    wire new_AGEMA_signal_7318 ;
    wire new_AGEMA_signal_7319 ;
    wire new_AGEMA_signal_7320 ;
    wire new_AGEMA_signal_7321 ;
    wire new_AGEMA_signal_7322 ;
    wire new_AGEMA_signal_7323 ;
    wire new_AGEMA_signal_7324 ;
    wire new_AGEMA_signal_7325 ;
    wire new_AGEMA_signal_7326 ;
    wire new_AGEMA_signal_7327 ;
    wire new_AGEMA_signal_7328 ;
    wire new_AGEMA_signal_7329 ;
    wire new_AGEMA_signal_7330 ;
    wire new_AGEMA_signal_7331 ;
    wire new_AGEMA_signal_7332 ;
    wire new_AGEMA_signal_7333 ;
    wire new_AGEMA_signal_7334 ;
    wire new_AGEMA_signal_7335 ;
    wire new_AGEMA_signal_7336 ;
    wire new_AGEMA_signal_7337 ;
    wire new_AGEMA_signal_7338 ;
    wire new_AGEMA_signal_7339 ;
    wire new_AGEMA_signal_7340 ;
    wire new_AGEMA_signal_7341 ;
    wire new_AGEMA_signal_7342 ;
    wire new_AGEMA_signal_7343 ;
    wire new_AGEMA_signal_7344 ;
    wire new_AGEMA_signal_7345 ;
    wire new_AGEMA_signal_7346 ;
    wire new_AGEMA_signal_7347 ;
    wire new_AGEMA_signal_7348 ;
    wire new_AGEMA_signal_7349 ;
    wire new_AGEMA_signal_7350 ;
    wire new_AGEMA_signal_7351 ;
    wire new_AGEMA_signal_7352 ;
    wire new_AGEMA_signal_7353 ;
    wire new_AGEMA_signal_7354 ;
    wire new_AGEMA_signal_7355 ;
    wire new_AGEMA_signal_7356 ;
    wire new_AGEMA_signal_7357 ;
    wire new_AGEMA_signal_7358 ;
    wire new_AGEMA_signal_7359 ;
    wire new_AGEMA_signal_7360 ;
    wire new_AGEMA_signal_7361 ;
    wire new_AGEMA_signal_7362 ;
    wire new_AGEMA_signal_7363 ;
    wire new_AGEMA_signal_7364 ;
    wire new_AGEMA_signal_7365 ;
    wire new_AGEMA_signal_7366 ;
    wire new_AGEMA_signal_7367 ;
    wire new_AGEMA_signal_7368 ;
    wire new_AGEMA_signal_7369 ;
    wire new_AGEMA_signal_7370 ;
    wire new_AGEMA_signal_7371 ;
    wire new_AGEMA_signal_7372 ;
    wire new_AGEMA_signal_7373 ;
    wire new_AGEMA_signal_7374 ;
    wire new_AGEMA_signal_7375 ;
    wire new_AGEMA_signal_7376 ;
    wire new_AGEMA_signal_7377 ;
    wire new_AGEMA_signal_7378 ;
    wire new_AGEMA_signal_7379 ;
    wire new_AGEMA_signal_7380 ;
    wire new_AGEMA_signal_7381 ;
    wire new_AGEMA_signal_7382 ;
    wire new_AGEMA_signal_7383 ;
    wire new_AGEMA_signal_7384 ;
    wire new_AGEMA_signal_7385 ;
    wire new_AGEMA_signal_7386 ;
    wire new_AGEMA_signal_7387 ;
    wire new_AGEMA_signal_7388 ;
    wire new_AGEMA_signal_7389 ;
    wire new_AGEMA_signal_7390 ;
    wire new_AGEMA_signal_7391 ;
    wire new_AGEMA_signal_7392 ;
    wire new_AGEMA_signal_7393 ;
    wire new_AGEMA_signal_7394 ;
    wire new_AGEMA_signal_7395 ;
    wire new_AGEMA_signal_7396 ;
    wire new_AGEMA_signal_7397 ;
    wire new_AGEMA_signal_7398 ;
    wire new_AGEMA_signal_7399 ;
    wire new_AGEMA_signal_7400 ;
    wire new_AGEMA_signal_7401 ;
    wire new_AGEMA_signal_7402 ;
    wire new_AGEMA_signal_7403 ;
    wire new_AGEMA_signal_7404 ;
    wire new_AGEMA_signal_7405 ;
    wire new_AGEMA_signal_7406 ;
    wire new_AGEMA_signal_7407 ;
    wire new_AGEMA_signal_7408 ;
    wire new_AGEMA_signal_7409 ;
    wire new_AGEMA_signal_7410 ;
    wire new_AGEMA_signal_7411 ;
    wire new_AGEMA_signal_7412 ;
    wire new_AGEMA_signal_7413 ;
    wire new_AGEMA_signal_7414 ;
    wire new_AGEMA_signal_7415 ;
    wire new_AGEMA_signal_7416 ;
    wire new_AGEMA_signal_7417 ;
    wire new_AGEMA_signal_7418 ;
    wire new_AGEMA_signal_7419 ;
    wire new_AGEMA_signal_7420 ;
    wire new_AGEMA_signal_7421 ;
    wire new_AGEMA_signal_7422 ;
    wire new_AGEMA_signal_7423 ;
    wire new_AGEMA_signal_7424 ;
    wire new_AGEMA_signal_7425 ;
    wire new_AGEMA_signal_7426 ;
    wire new_AGEMA_signal_7427 ;
    wire new_AGEMA_signal_7428 ;
    wire new_AGEMA_signal_7429 ;
    wire new_AGEMA_signal_7430 ;
    wire new_AGEMA_signal_7431 ;
    wire new_AGEMA_signal_7432 ;
    wire new_AGEMA_signal_7433 ;
    wire new_AGEMA_signal_7434 ;
    wire new_AGEMA_signal_7435 ;
    wire new_AGEMA_signal_7436 ;
    wire new_AGEMA_signal_7437 ;
    wire new_AGEMA_signal_7438 ;
    wire new_AGEMA_signal_7439 ;
    wire new_AGEMA_signal_7440 ;
    wire new_AGEMA_signal_7441 ;
    wire new_AGEMA_signal_7442 ;
    wire new_AGEMA_signal_7443 ;
    wire new_AGEMA_signal_7444 ;
    wire new_AGEMA_signal_7445 ;
    wire new_AGEMA_signal_7446 ;
    wire new_AGEMA_signal_7447 ;
    wire new_AGEMA_signal_7448 ;
    wire new_AGEMA_signal_7449 ;
    wire new_AGEMA_signal_7450 ;
    wire new_AGEMA_signal_7451 ;
    wire new_AGEMA_signal_7452 ;
    wire new_AGEMA_signal_7453 ;
    wire new_AGEMA_signal_7454 ;
    wire new_AGEMA_signal_7455 ;
    wire new_AGEMA_signal_7456 ;
    wire new_AGEMA_signal_7457 ;
    wire new_AGEMA_signal_7458 ;
    wire new_AGEMA_signal_7459 ;
    wire new_AGEMA_signal_7460 ;
    wire new_AGEMA_signal_7461 ;
    wire new_AGEMA_signal_7462 ;
    wire new_AGEMA_signal_7463 ;
    wire new_AGEMA_signal_7464 ;
    wire new_AGEMA_signal_7465 ;
    wire new_AGEMA_signal_7466 ;
    wire new_AGEMA_signal_7467 ;
    wire new_AGEMA_signal_7468 ;
    wire new_AGEMA_signal_7469 ;
    wire new_AGEMA_signal_7470 ;
    wire new_AGEMA_signal_7471 ;
    wire new_AGEMA_signal_7472 ;
    wire new_AGEMA_signal_7473 ;
    wire new_AGEMA_signal_7474 ;
    wire new_AGEMA_signal_7475 ;
    wire new_AGEMA_signal_7476 ;
    wire new_AGEMA_signal_7477 ;
    wire new_AGEMA_signal_7478 ;
    wire new_AGEMA_signal_7479 ;
    wire new_AGEMA_signal_7480 ;
    wire new_AGEMA_signal_7481 ;
    wire new_AGEMA_signal_7482 ;
    wire new_AGEMA_signal_7483 ;
    wire new_AGEMA_signal_7484 ;
    wire new_AGEMA_signal_7485 ;
    wire new_AGEMA_signal_7486 ;
    wire new_AGEMA_signal_7487 ;
    wire new_AGEMA_signal_7488 ;
    wire new_AGEMA_signal_7489 ;
    wire new_AGEMA_signal_7490 ;
    wire new_AGEMA_signal_7491 ;
    wire new_AGEMA_signal_7492 ;
    wire new_AGEMA_signal_7493 ;
    wire new_AGEMA_signal_7494 ;
    wire new_AGEMA_signal_7495 ;
    wire new_AGEMA_signal_7496 ;
    wire new_AGEMA_signal_7497 ;
    wire new_AGEMA_signal_7498 ;
    wire new_AGEMA_signal_7499 ;
    wire new_AGEMA_signal_7500 ;
    wire new_AGEMA_signal_7501 ;
    wire new_AGEMA_signal_7502 ;
    wire new_AGEMA_signal_7503 ;
    wire new_AGEMA_signal_7504 ;
    wire new_AGEMA_signal_7505 ;
    wire new_AGEMA_signal_7506 ;
    wire new_AGEMA_signal_7507 ;
    wire new_AGEMA_signal_7508 ;
    wire new_AGEMA_signal_7509 ;
    wire new_AGEMA_signal_7510 ;
    wire new_AGEMA_signal_7511 ;
    wire new_AGEMA_signal_7512 ;
    wire new_AGEMA_signal_7513 ;
    wire new_AGEMA_signal_7514 ;
    wire new_AGEMA_signal_7515 ;
    wire new_AGEMA_signal_7516 ;
    wire new_AGEMA_signal_7517 ;
    wire new_AGEMA_signal_7518 ;
    wire new_AGEMA_signal_7519 ;
    wire new_AGEMA_signal_7520 ;
    wire new_AGEMA_signal_7521 ;
    wire new_AGEMA_signal_7522 ;
    wire new_AGEMA_signal_7523 ;
    wire new_AGEMA_signal_7524 ;
    wire new_AGEMA_signal_7525 ;
    wire new_AGEMA_signal_7526 ;
    wire new_AGEMA_signal_7527 ;
    wire new_AGEMA_signal_7528 ;
    wire new_AGEMA_signal_7529 ;
    wire new_AGEMA_signal_7530 ;
    wire new_AGEMA_signal_7531 ;
    wire new_AGEMA_signal_7532 ;
    wire new_AGEMA_signal_7533 ;
    wire new_AGEMA_signal_7534 ;
    wire new_AGEMA_signal_7535 ;
    wire new_AGEMA_signal_7536 ;
    wire new_AGEMA_signal_7537 ;
    wire new_AGEMA_signal_7538 ;
    wire new_AGEMA_signal_7539 ;
    wire new_AGEMA_signal_7540 ;
    wire new_AGEMA_signal_7541 ;
    wire new_AGEMA_signal_7542 ;
    wire new_AGEMA_signal_7543 ;
    wire new_AGEMA_signal_7544 ;
    wire new_AGEMA_signal_7545 ;
    wire new_AGEMA_signal_7546 ;
    wire new_AGEMA_signal_7547 ;
    wire new_AGEMA_signal_7548 ;
    wire new_AGEMA_signal_7549 ;
    wire new_AGEMA_signal_7550 ;
    wire new_AGEMA_signal_7551 ;
    wire new_AGEMA_signal_7552 ;
    wire new_AGEMA_signal_7553 ;
    wire new_AGEMA_signal_7554 ;
    wire new_AGEMA_signal_7555 ;
    wire new_AGEMA_signal_7556 ;
    wire new_AGEMA_signal_7557 ;
    wire new_AGEMA_signal_7558 ;
    wire new_AGEMA_signal_7559 ;
    wire new_AGEMA_signal_7560 ;
    wire new_AGEMA_signal_7561 ;
    wire new_AGEMA_signal_7562 ;
    wire new_AGEMA_signal_7563 ;
    wire new_AGEMA_signal_7564 ;
    wire new_AGEMA_signal_7565 ;
    wire new_AGEMA_signal_7566 ;
    wire new_AGEMA_signal_7567 ;
    wire new_AGEMA_signal_7568 ;
    wire new_AGEMA_signal_7569 ;
    wire new_AGEMA_signal_7570 ;
    wire new_AGEMA_signal_7571 ;
    wire new_AGEMA_signal_7572 ;
    wire new_AGEMA_signal_7573 ;
    wire new_AGEMA_signal_7574 ;
    wire new_AGEMA_signal_7575 ;
    wire new_AGEMA_signal_7576 ;
    wire new_AGEMA_signal_7577 ;
    wire new_AGEMA_signal_7578 ;
    wire new_AGEMA_signal_7579 ;
    wire new_AGEMA_signal_7580 ;
    wire new_AGEMA_signal_7581 ;
    wire new_AGEMA_signal_7582 ;
    wire new_AGEMA_signal_7583 ;
    wire new_AGEMA_signal_7584 ;
    wire new_AGEMA_signal_7585 ;
    wire new_AGEMA_signal_7586 ;
    wire new_AGEMA_signal_7587 ;
    wire new_AGEMA_signal_7588 ;
    wire new_AGEMA_signal_7589 ;
    wire new_AGEMA_signal_7590 ;
    wire new_AGEMA_signal_7591 ;
    wire new_AGEMA_signal_7592 ;
    wire new_AGEMA_signal_7593 ;
    wire new_AGEMA_signal_7594 ;
    wire new_AGEMA_signal_7595 ;
    wire new_AGEMA_signal_7596 ;
    wire new_AGEMA_signal_7597 ;
    wire new_AGEMA_signal_7598 ;
    wire new_AGEMA_signal_7599 ;
    wire new_AGEMA_signal_7600 ;
    wire new_AGEMA_signal_7601 ;
    wire new_AGEMA_signal_7602 ;
    wire new_AGEMA_signal_7603 ;
    wire new_AGEMA_signal_7604 ;
    wire new_AGEMA_signal_7605 ;
    wire new_AGEMA_signal_7606 ;
    wire new_AGEMA_signal_7607 ;
    wire new_AGEMA_signal_7608 ;
    wire new_AGEMA_signal_7609 ;
    wire new_AGEMA_signal_7610 ;
    wire new_AGEMA_signal_7611 ;
    wire new_AGEMA_signal_7612 ;
    wire new_AGEMA_signal_7613 ;
    wire new_AGEMA_signal_7614 ;
    wire new_AGEMA_signal_7615 ;
    wire new_AGEMA_signal_7616 ;
    wire new_AGEMA_signal_7617 ;
    wire new_AGEMA_signal_7618 ;
    wire new_AGEMA_signal_7619 ;
    wire new_AGEMA_signal_7620 ;
    wire new_AGEMA_signal_7621 ;
    wire new_AGEMA_signal_7622 ;
    wire new_AGEMA_signal_7623 ;
    wire new_AGEMA_signal_7624 ;
    wire new_AGEMA_signal_7625 ;
    wire new_AGEMA_signal_7626 ;
    wire new_AGEMA_signal_7627 ;
    wire new_AGEMA_signal_7628 ;
    wire new_AGEMA_signal_7629 ;
    wire new_AGEMA_signal_7630 ;
    wire new_AGEMA_signal_7631 ;
    wire new_AGEMA_signal_7632 ;
    wire new_AGEMA_signal_7633 ;
    wire new_AGEMA_signal_7634 ;
    wire new_AGEMA_signal_7635 ;
    wire new_AGEMA_signal_7636 ;
    wire new_AGEMA_signal_7637 ;
    wire new_AGEMA_signal_7638 ;
    wire new_AGEMA_signal_7639 ;
    wire new_AGEMA_signal_7640 ;
    wire new_AGEMA_signal_7641 ;
    wire new_AGEMA_signal_7642 ;
    wire new_AGEMA_signal_7643 ;
    wire new_AGEMA_signal_7644 ;
    wire new_AGEMA_signal_7645 ;
    wire new_AGEMA_signal_7646 ;
    wire new_AGEMA_signal_7647 ;
    wire new_AGEMA_signal_7648 ;
    wire new_AGEMA_signal_7649 ;
    wire new_AGEMA_signal_7650 ;
    wire new_AGEMA_signal_7651 ;
    wire new_AGEMA_signal_7652 ;
    wire new_AGEMA_signal_7653 ;
    wire new_AGEMA_signal_7654 ;
    wire new_AGEMA_signal_7655 ;
    wire new_AGEMA_signal_7656 ;
    wire new_AGEMA_signal_7657 ;
    wire new_AGEMA_signal_7658 ;
    wire new_AGEMA_signal_7659 ;
    wire new_AGEMA_signal_7660 ;
    wire new_AGEMA_signal_7661 ;
    wire new_AGEMA_signal_7662 ;
    wire new_AGEMA_signal_7663 ;
    wire new_AGEMA_signal_7664 ;
    wire new_AGEMA_signal_7665 ;
    wire new_AGEMA_signal_7666 ;
    wire new_AGEMA_signal_7667 ;
    wire new_AGEMA_signal_7668 ;
    wire new_AGEMA_signal_7669 ;
    wire new_AGEMA_signal_7670 ;
    wire new_AGEMA_signal_7671 ;
    wire new_AGEMA_signal_7672 ;
    wire new_AGEMA_signal_7673 ;
    wire new_AGEMA_signal_7674 ;
    wire new_AGEMA_signal_7675 ;
    wire new_AGEMA_signal_7676 ;
    wire new_AGEMA_signal_7677 ;
    wire new_AGEMA_signal_7678 ;
    wire new_AGEMA_signal_7679 ;
    wire new_AGEMA_signal_7680 ;
    wire new_AGEMA_signal_7681 ;
    wire new_AGEMA_signal_7682 ;
    wire new_AGEMA_signal_7683 ;
    wire new_AGEMA_signal_7684 ;
    wire new_AGEMA_signal_7685 ;
    wire new_AGEMA_signal_7686 ;
    wire new_AGEMA_signal_7687 ;
    wire new_AGEMA_signal_7688 ;
    wire new_AGEMA_signal_7689 ;
    wire new_AGEMA_signal_7690 ;
    wire new_AGEMA_signal_7691 ;
    wire new_AGEMA_signal_7692 ;
    wire new_AGEMA_signal_7693 ;
    wire new_AGEMA_signal_7694 ;
    wire new_AGEMA_signal_7695 ;
    wire new_AGEMA_signal_7696 ;
    wire new_AGEMA_signal_7697 ;
    wire new_AGEMA_signal_7698 ;
    wire new_AGEMA_signal_7699 ;
    wire new_AGEMA_signal_7700 ;
    wire new_AGEMA_signal_7701 ;
    wire new_AGEMA_signal_7702 ;
    wire new_AGEMA_signal_7703 ;
    wire new_AGEMA_signal_7704 ;
    wire new_AGEMA_signal_7705 ;
    wire new_AGEMA_signal_7706 ;
    wire new_AGEMA_signal_7707 ;
    wire new_AGEMA_signal_7708 ;
    wire new_AGEMA_signal_7709 ;
    wire new_AGEMA_signal_7710 ;
    wire new_AGEMA_signal_7711 ;
    wire new_AGEMA_signal_7712 ;
    wire new_AGEMA_signal_7713 ;
    wire new_AGEMA_signal_7714 ;
    wire new_AGEMA_signal_7715 ;
    wire new_AGEMA_signal_7716 ;
    wire new_AGEMA_signal_7717 ;
    wire new_AGEMA_signal_7718 ;
    wire new_AGEMA_signal_7719 ;
    wire new_AGEMA_signal_7720 ;
    wire new_AGEMA_signal_7721 ;
    wire new_AGEMA_signal_7722 ;
    wire new_AGEMA_signal_7723 ;
    wire new_AGEMA_signal_7724 ;
    wire new_AGEMA_signal_7725 ;
    wire new_AGEMA_signal_7726 ;
    wire new_AGEMA_signal_7727 ;
    wire new_AGEMA_signal_7728 ;
    wire new_AGEMA_signal_7729 ;
    wire new_AGEMA_signal_7730 ;
    wire new_AGEMA_signal_7731 ;
    wire new_AGEMA_signal_7732 ;
    wire new_AGEMA_signal_7733 ;
    wire new_AGEMA_signal_7734 ;
    wire new_AGEMA_signal_7735 ;
    wire new_AGEMA_signal_7736 ;
    wire new_AGEMA_signal_7737 ;
    wire new_AGEMA_signal_7738 ;
    wire new_AGEMA_signal_7739 ;
    wire new_AGEMA_signal_7740 ;
    wire new_AGEMA_signal_7741 ;
    wire new_AGEMA_signal_7742 ;
    wire new_AGEMA_signal_7743 ;
    wire new_AGEMA_signal_7744 ;
    wire new_AGEMA_signal_7745 ;
    wire new_AGEMA_signal_7746 ;
    wire new_AGEMA_signal_7747 ;
    wire new_AGEMA_signal_7748 ;
    wire new_AGEMA_signal_7749 ;
    wire new_AGEMA_signal_7750 ;
    wire new_AGEMA_signal_7751 ;
    wire new_AGEMA_signal_7752 ;
    wire new_AGEMA_signal_7753 ;
    wire new_AGEMA_signal_7754 ;
    wire new_AGEMA_signal_7755 ;
    wire new_AGEMA_signal_7756 ;
    wire new_AGEMA_signal_7757 ;
    wire new_AGEMA_signal_7758 ;
    wire new_AGEMA_signal_7759 ;
    wire new_AGEMA_signal_7760 ;
    wire new_AGEMA_signal_7761 ;
    wire new_AGEMA_signal_7762 ;
    wire new_AGEMA_signal_7763 ;
    wire new_AGEMA_signal_7764 ;
    wire new_AGEMA_signal_7765 ;
    wire new_AGEMA_signal_7766 ;
    wire new_AGEMA_signal_7767 ;
    wire new_AGEMA_signal_7768 ;
    wire new_AGEMA_signal_7769 ;
    wire new_AGEMA_signal_7770 ;
    wire new_AGEMA_signal_7771 ;
    wire new_AGEMA_signal_7772 ;
    wire new_AGEMA_signal_7773 ;
    wire new_AGEMA_signal_7774 ;
    wire new_AGEMA_signal_7775 ;
    wire new_AGEMA_signal_7776 ;
    wire new_AGEMA_signal_7777 ;
    wire new_AGEMA_signal_7778 ;
    wire new_AGEMA_signal_7779 ;
    wire new_AGEMA_signal_7780 ;
    wire new_AGEMA_signal_7781 ;
    wire new_AGEMA_signal_7782 ;
    wire new_AGEMA_signal_7783 ;
    wire new_AGEMA_signal_7784 ;
    wire new_AGEMA_signal_7785 ;
    wire new_AGEMA_signal_7786 ;
    wire new_AGEMA_signal_7787 ;
    wire new_AGEMA_signal_7788 ;
    wire new_AGEMA_signal_7789 ;
    wire new_AGEMA_signal_7790 ;
    wire new_AGEMA_signal_7791 ;
    wire new_AGEMA_signal_7792 ;
    wire new_AGEMA_signal_7793 ;
    wire new_AGEMA_signal_7794 ;
    wire new_AGEMA_signal_7795 ;
    wire new_AGEMA_signal_7796 ;
    wire new_AGEMA_signal_7797 ;
    wire new_AGEMA_signal_7798 ;
    wire new_AGEMA_signal_7799 ;
    wire new_AGEMA_signal_7800 ;
    wire new_AGEMA_signal_7801 ;
    wire new_AGEMA_signal_7802 ;
    wire new_AGEMA_signal_7803 ;
    wire new_AGEMA_signal_7804 ;
    wire new_AGEMA_signal_7805 ;
    wire new_AGEMA_signal_7806 ;
    wire new_AGEMA_signal_7807 ;
    wire new_AGEMA_signal_7808 ;
    wire new_AGEMA_signal_7809 ;
    wire new_AGEMA_signal_7810 ;
    wire new_AGEMA_signal_7811 ;
    wire new_AGEMA_signal_7812 ;
    wire new_AGEMA_signal_7813 ;
    wire new_AGEMA_signal_7814 ;
    wire new_AGEMA_signal_7815 ;
    wire new_AGEMA_signal_7816 ;
    wire new_AGEMA_signal_7817 ;
    wire new_AGEMA_signal_7818 ;
    wire new_AGEMA_signal_7819 ;
    wire new_AGEMA_signal_7820 ;
    wire new_AGEMA_signal_7821 ;
    wire new_AGEMA_signal_7822 ;
    wire new_AGEMA_signal_7823 ;
    wire new_AGEMA_signal_7824 ;
    wire new_AGEMA_signal_7825 ;
    wire new_AGEMA_signal_7826 ;
    wire new_AGEMA_signal_7827 ;
    wire new_AGEMA_signal_7828 ;
    wire new_AGEMA_signal_7829 ;
    wire new_AGEMA_signal_7830 ;
    wire new_AGEMA_signal_7831 ;
    wire new_AGEMA_signal_7832 ;
    wire new_AGEMA_signal_7833 ;
    wire new_AGEMA_signal_7834 ;
    wire new_AGEMA_signal_7835 ;
    wire new_AGEMA_signal_7836 ;
    wire new_AGEMA_signal_7837 ;
    wire new_AGEMA_signal_7838 ;
    wire new_AGEMA_signal_7839 ;
    wire new_AGEMA_signal_7840 ;
    wire new_AGEMA_signal_7841 ;
    wire new_AGEMA_signal_7842 ;
    wire new_AGEMA_signal_7843 ;
    wire new_AGEMA_signal_7844 ;
    wire new_AGEMA_signal_7845 ;
    wire new_AGEMA_signal_7846 ;
    wire new_AGEMA_signal_7847 ;
    wire new_AGEMA_signal_7848 ;
    wire new_AGEMA_signal_7849 ;
    wire new_AGEMA_signal_7850 ;
    wire new_AGEMA_signal_7851 ;
    wire new_AGEMA_signal_7852 ;
    wire new_AGEMA_signal_7853 ;
    wire new_AGEMA_signal_7854 ;
    wire new_AGEMA_signal_7855 ;
    wire new_AGEMA_signal_7856 ;
    wire new_AGEMA_signal_7857 ;
    wire new_AGEMA_signal_7858 ;
    wire new_AGEMA_signal_7859 ;
    wire new_AGEMA_signal_7860 ;
    wire new_AGEMA_signal_7861 ;
    wire new_AGEMA_signal_7862 ;
    wire new_AGEMA_signal_7863 ;
    wire new_AGEMA_signal_7864 ;
    wire new_AGEMA_signal_7865 ;
    wire new_AGEMA_signal_7866 ;
    wire new_AGEMA_signal_7867 ;
    wire new_AGEMA_signal_7868 ;
    wire new_AGEMA_signal_7869 ;
    wire new_AGEMA_signal_7870 ;
    wire new_AGEMA_signal_7871 ;
    wire new_AGEMA_signal_7872 ;
    wire new_AGEMA_signal_7873 ;
    wire new_AGEMA_signal_7874 ;
    wire new_AGEMA_signal_7875 ;
    wire new_AGEMA_signal_7876 ;
    wire new_AGEMA_signal_7877 ;
    wire new_AGEMA_signal_7878 ;
    wire new_AGEMA_signal_7879 ;
    wire new_AGEMA_signal_7880 ;
    wire new_AGEMA_signal_7881 ;
    wire new_AGEMA_signal_7882 ;
    wire new_AGEMA_signal_7883 ;
    wire new_AGEMA_signal_7884 ;
    wire new_AGEMA_signal_7885 ;
    wire new_AGEMA_signal_7886 ;
    wire new_AGEMA_signal_7887 ;
    wire new_AGEMA_signal_7888 ;
    wire new_AGEMA_signal_7889 ;
    wire new_AGEMA_signal_7890 ;
    wire new_AGEMA_signal_7891 ;
    wire new_AGEMA_signal_7892 ;
    wire new_AGEMA_signal_7893 ;
    wire new_AGEMA_signal_7894 ;
    wire new_AGEMA_signal_7895 ;
    wire new_AGEMA_signal_7896 ;
    wire new_AGEMA_signal_7897 ;
    wire new_AGEMA_signal_7898 ;
    wire new_AGEMA_signal_7899 ;
    wire new_AGEMA_signal_7900 ;
    wire new_AGEMA_signal_7901 ;
    wire new_AGEMA_signal_7902 ;
    wire new_AGEMA_signal_7903 ;
    wire new_AGEMA_signal_7904 ;
    wire new_AGEMA_signal_7905 ;
    wire new_AGEMA_signal_7906 ;
    wire new_AGEMA_signal_7907 ;
    wire new_AGEMA_signal_7908 ;
    wire new_AGEMA_signal_7909 ;
    wire new_AGEMA_signal_7910 ;
    wire new_AGEMA_signal_7911 ;
    wire new_AGEMA_signal_7912 ;
    wire new_AGEMA_signal_7913 ;
    wire new_AGEMA_signal_7914 ;
    wire new_AGEMA_signal_7915 ;
    wire new_AGEMA_signal_7916 ;
    wire new_AGEMA_signal_7917 ;
    wire new_AGEMA_signal_7918 ;
    wire new_AGEMA_signal_7919 ;
    wire new_AGEMA_signal_7920 ;
    wire new_AGEMA_signal_7921 ;
    wire new_AGEMA_signal_7922 ;
    wire new_AGEMA_signal_7923 ;
    wire new_AGEMA_signal_7924 ;
    wire new_AGEMA_signal_7925 ;
    wire new_AGEMA_signal_7926 ;
    wire new_AGEMA_signal_7927 ;
    wire new_AGEMA_signal_7928 ;
    wire new_AGEMA_signal_7929 ;
    wire new_AGEMA_signal_7930 ;
    wire new_AGEMA_signal_7931 ;
    wire new_AGEMA_signal_7932 ;
    wire new_AGEMA_signal_7933 ;
    wire new_AGEMA_signal_7934 ;
    wire new_AGEMA_signal_7935 ;
    wire new_AGEMA_signal_7936 ;
    wire new_AGEMA_signal_7937 ;
    wire new_AGEMA_signal_7938 ;
    wire new_AGEMA_signal_7939 ;
    wire new_AGEMA_signal_7940 ;
    wire new_AGEMA_signal_7941 ;
    wire new_AGEMA_signal_7942 ;
    wire new_AGEMA_signal_7943 ;
    wire new_AGEMA_signal_7944 ;
    wire new_AGEMA_signal_7945 ;
    wire new_AGEMA_signal_7946 ;
    wire new_AGEMA_signal_7947 ;
    wire new_AGEMA_signal_7948 ;
    wire new_AGEMA_signal_7949 ;
    wire new_AGEMA_signal_7950 ;
    wire new_AGEMA_signal_7951 ;
    wire new_AGEMA_signal_7952 ;
    wire new_AGEMA_signal_7953 ;
    wire new_AGEMA_signal_7954 ;
    wire new_AGEMA_signal_7955 ;
    wire new_AGEMA_signal_7956 ;
    wire new_AGEMA_signal_7957 ;
    wire new_AGEMA_signal_7958 ;
    wire new_AGEMA_signal_7959 ;
    wire new_AGEMA_signal_7960 ;
    wire new_AGEMA_signal_7961 ;
    wire new_AGEMA_signal_7962 ;
    wire new_AGEMA_signal_7963 ;
    wire new_AGEMA_signal_7964 ;
    wire new_AGEMA_signal_7965 ;
    wire new_AGEMA_signal_7966 ;
    wire new_AGEMA_signal_7967 ;
    wire new_AGEMA_signal_7968 ;
    wire new_AGEMA_signal_7969 ;
    wire new_AGEMA_signal_7970 ;
    wire new_AGEMA_signal_7971 ;
    wire new_AGEMA_signal_7972 ;
    wire new_AGEMA_signal_7973 ;
    wire new_AGEMA_signal_7974 ;
    wire new_AGEMA_signal_7975 ;
    wire new_AGEMA_signal_7976 ;
    wire new_AGEMA_signal_7977 ;
    wire new_AGEMA_signal_7978 ;
    wire new_AGEMA_signal_7979 ;
    wire new_AGEMA_signal_7980 ;
    wire new_AGEMA_signal_7981 ;
    wire new_AGEMA_signal_7982 ;
    wire new_AGEMA_signal_7983 ;
    wire new_AGEMA_signal_7984 ;
    wire new_AGEMA_signal_7985 ;
    wire new_AGEMA_signal_7986 ;
    wire new_AGEMA_signal_7987 ;
    wire new_AGEMA_signal_7988 ;
    wire new_AGEMA_signal_7989 ;
    wire new_AGEMA_signal_7990 ;
    wire new_AGEMA_signal_7991 ;
    wire new_AGEMA_signal_7992 ;
    wire new_AGEMA_signal_7993 ;
    wire new_AGEMA_signal_7994 ;
    wire new_AGEMA_signal_7995 ;
    wire new_AGEMA_signal_7996 ;
    wire new_AGEMA_signal_7997 ;
    wire new_AGEMA_signal_7998 ;
    wire new_AGEMA_signal_7999 ;
    wire new_AGEMA_signal_8000 ;
    wire new_AGEMA_signal_8001 ;
    wire new_AGEMA_signal_8002 ;
    wire new_AGEMA_signal_8003 ;
    wire new_AGEMA_signal_8004 ;
    wire new_AGEMA_signal_8005 ;
    wire new_AGEMA_signal_8006 ;
    wire new_AGEMA_signal_8007 ;
    wire new_AGEMA_signal_8008 ;
    wire new_AGEMA_signal_8009 ;
    wire new_AGEMA_signal_8010 ;
    wire new_AGEMA_signal_8011 ;
    wire new_AGEMA_signal_8012 ;
    wire new_AGEMA_signal_8013 ;
    wire new_AGEMA_signal_8014 ;
    wire new_AGEMA_signal_8015 ;
    wire new_AGEMA_signal_8016 ;
    wire new_AGEMA_signal_8017 ;
    wire new_AGEMA_signal_8018 ;
    wire new_AGEMA_signal_8019 ;
    wire new_AGEMA_signal_8020 ;
    wire new_AGEMA_signal_8021 ;
    wire new_AGEMA_signal_8022 ;
    wire new_AGEMA_signal_8023 ;
    wire new_AGEMA_signal_8024 ;
    wire new_AGEMA_signal_8025 ;
    wire new_AGEMA_signal_8026 ;
    wire new_AGEMA_signal_8027 ;
    wire new_AGEMA_signal_8028 ;
    wire new_AGEMA_signal_8029 ;
    wire new_AGEMA_signal_8030 ;
    wire new_AGEMA_signal_8031 ;
    wire new_AGEMA_signal_8032 ;
    wire new_AGEMA_signal_8033 ;
    wire new_AGEMA_signal_8034 ;
    wire new_AGEMA_signal_8035 ;
    wire new_AGEMA_signal_8036 ;
    wire new_AGEMA_signal_8037 ;
    wire new_AGEMA_signal_8038 ;
    wire new_AGEMA_signal_8039 ;
    wire new_AGEMA_signal_8040 ;
    wire new_AGEMA_signal_8041 ;
    wire new_AGEMA_signal_8042 ;
    wire new_AGEMA_signal_8043 ;
    wire new_AGEMA_signal_8044 ;
    wire new_AGEMA_signal_8045 ;
    wire new_AGEMA_signal_8046 ;
    wire new_AGEMA_signal_8047 ;
    wire new_AGEMA_signal_8048 ;
    wire new_AGEMA_signal_8049 ;
    wire new_AGEMA_signal_8050 ;
    wire new_AGEMA_signal_8051 ;
    wire new_AGEMA_signal_8052 ;
    wire new_AGEMA_signal_8053 ;
    wire new_AGEMA_signal_8054 ;
    wire new_AGEMA_signal_8055 ;
    wire new_AGEMA_signal_8056 ;
    wire new_AGEMA_signal_8057 ;
    wire new_AGEMA_signal_8058 ;
    wire new_AGEMA_signal_8059 ;
    wire new_AGEMA_signal_8060 ;
    wire new_AGEMA_signal_8061 ;
    wire new_AGEMA_signal_8062 ;
    wire new_AGEMA_signal_8063 ;
    wire new_AGEMA_signal_8064 ;
    wire new_AGEMA_signal_8065 ;
    wire new_AGEMA_signal_8066 ;
    wire new_AGEMA_signal_8067 ;
    wire new_AGEMA_signal_8068 ;
    wire new_AGEMA_signal_8069 ;
    wire new_AGEMA_signal_8070 ;
    wire new_AGEMA_signal_8071 ;
    wire new_AGEMA_signal_8072 ;
    wire new_AGEMA_signal_8073 ;
    wire new_AGEMA_signal_8074 ;
    wire new_AGEMA_signal_8075 ;
    wire new_AGEMA_signal_8076 ;
    wire new_AGEMA_signal_8077 ;
    wire new_AGEMA_signal_8078 ;
    wire new_AGEMA_signal_8079 ;
    wire new_AGEMA_signal_8080 ;
    wire new_AGEMA_signal_8081 ;
    wire new_AGEMA_signal_8082 ;
    wire new_AGEMA_signal_8083 ;
    wire new_AGEMA_signal_8084 ;
    wire new_AGEMA_signal_8085 ;
    wire new_AGEMA_signal_8086 ;
    wire new_AGEMA_signal_8087 ;
    wire new_AGEMA_signal_8088 ;
    wire new_AGEMA_signal_8089 ;
    wire new_AGEMA_signal_8090 ;
    wire new_AGEMA_signal_8091 ;
    wire new_AGEMA_signal_8092 ;
    wire new_AGEMA_signal_8093 ;
    wire new_AGEMA_signal_8094 ;
    wire new_AGEMA_signal_8095 ;
    wire new_AGEMA_signal_8096 ;
    wire new_AGEMA_signal_8097 ;
    wire new_AGEMA_signal_8098 ;
    wire new_AGEMA_signal_8099 ;
    wire new_AGEMA_signal_8100 ;
    wire new_AGEMA_signal_8101 ;
    wire new_AGEMA_signal_8102 ;
    wire new_AGEMA_signal_8103 ;
    wire new_AGEMA_signal_8104 ;
    wire new_AGEMA_signal_8105 ;
    wire new_AGEMA_signal_8106 ;
    wire new_AGEMA_signal_8107 ;
    wire new_AGEMA_signal_8108 ;
    wire new_AGEMA_signal_8109 ;
    wire new_AGEMA_signal_8110 ;
    wire new_AGEMA_signal_8111 ;
    wire new_AGEMA_signal_8112 ;
    wire new_AGEMA_signal_8113 ;
    wire new_AGEMA_signal_8114 ;
    wire new_AGEMA_signal_8115 ;
    wire new_AGEMA_signal_8116 ;
    wire new_AGEMA_signal_8117 ;
    wire new_AGEMA_signal_8118 ;
    wire new_AGEMA_signal_8119 ;
    wire new_AGEMA_signal_8120 ;
    wire new_AGEMA_signal_8121 ;
    wire new_AGEMA_signal_8122 ;
    wire new_AGEMA_signal_8123 ;
    wire new_AGEMA_signal_8124 ;
    wire new_AGEMA_signal_8125 ;
    wire new_AGEMA_signal_8126 ;
    wire new_AGEMA_signal_8127 ;
    wire new_AGEMA_signal_8128 ;
    wire new_AGEMA_signal_8129 ;
    wire new_AGEMA_signal_8130 ;
    wire new_AGEMA_signal_8131 ;
    wire new_AGEMA_signal_8132 ;
    wire new_AGEMA_signal_8133 ;
    wire new_AGEMA_signal_8134 ;
    wire new_AGEMA_signal_8135 ;
    wire new_AGEMA_signal_8136 ;
    wire new_AGEMA_signal_8137 ;
    wire new_AGEMA_signal_8138 ;
    wire new_AGEMA_signal_8139 ;
    wire new_AGEMA_signal_8140 ;
    wire new_AGEMA_signal_8141 ;
    wire new_AGEMA_signal_8142 ;
    wire new_AGEMA_signal_8143 ;
    wire new_AGEMA_signal_8144 ;
    wire new_AGEMA_signal_8145 ;
    wire new_AGEMA_signal_8146 ;
    wire new_AGEMA_signal_8147 ;
    wire new_AGEMA_signal_8148 ;
    wire new_AGEMA_signal_8149 ;
    wire new_AGEMA_signal_8150 ;
    wire new_AGEMA_signal_8151 ;
    wire new_AGEMA_signal_8152 ;
    wire new_AGEMA_signal_8153 ;
    wire new_AGEMA_signal_8154 ;
    wire new_AGEMA_signal_8155 ;
    wire new_AGEMA_signal_8156 ;
    wire new_AGEMA_signal_8157 ;
    wire new_AGEMA_signal_8158 ;
    wire new_AGEMA_signal_8159 ;
    wire new_AGEMA_signal_8160 ;
    wire new_AGEMA_signal_8161 ;
    wire new_AGEMA_signal_8162 ;
    wire new_AGEMA_signal_8163 ;
    wire new_AGEMA_signal_8164 ;
    wire new_AGEMA_signal_8165 ;
    wire new_AGEMA_signal_8166 ;
    wire new_AGEMA_signal_8167 ;
    wire new_AGEMA_signal_8168 ;
    wire new_AGEMA_signal_8169 ;
    wire new_AGEMA_signal_8170 ;
    wire new_AGEMA_signal_8171 ;
    wire new_AGEMA_signal_8172 ;
    wire new_AGEMA_signal_8173 ;
    wire new_AGEMA_signal_8174 ;
    wire new_AGEMA_signal_8175 ;
    wire new_AGEMA_signal_8176 ;
    wire new_AGEMA_signal_8177 ;
    wire new_AGEMA_signal_8178 ;
    wire new_AGEMA_signal_8179 ;
    wire new_AGEMA_signal_8180 ;
    wire new_AGEMA_signal_8181 ;
    wire new_AGEMA_signal_8182 ;
    wire new_AGEMA_signal_8183 ;
    wire new_AGEMA_signal_8184 ;
    wire new_AGEMA_signal_8185 ;
    wire new_AGEMA_signal_8186 ;
    wire new_AGEMA_signal_8187 ;
    wire new_AGEMA_signal_8188 ;
    wire new_AGEMA_signal_8189 ;
    wire new_AGEMA_signal_8190 ;
    wire new_AGEMA_signal_8191 ;
    wire new_AGEMA_signal_8192 ;
    wire new_AGEMA_signal_8193 ;
    wire new_AGEMA_signal_8194 ;
    wire new_AGEMA_signal_8195 ;
    wire new_AGEMA_signal_8196 ;
    wire new_AGEMA_signal_8197 ;
    wire new_AGEMA_signal_8198 ;
    wire new_AGEMA_signal_8199 ;
    wire new_AGEMA_signal_8200 ;
    wire new_AGEMA_signal_8201 ;
    wire new_AGEMA_signal_8202 ;
    wire new_AGEMA_signal_8203 ;
    wire new_AGEMA_signal_8204 ;
    wire new_AGEMA_signal_8205 ;
    wire new_AGEMA_signal_8206 ;
    wire new_AGEMA_signal_8207 ;
    wire new_AGEMA_signal_8208 ;
    wire new_AGEMA_signal_8209 ;
    wire new_AGEMA_signal_8210 ;
    wire new_AGEMA_signal_8211 ;
    wire new_AGEMA_signal_8212 ;
    wire new_AGEMA_signal_8213 ;
    wire new_AGEMA_signal_8214 ;
    wire new_AGEMA_signal_8215 ;
    wire new_AGEMA_signal_8216 ;
    wire new_AGEMA_signal_8217 ;
    wire new_AGEMA_signal_8218 ;
    wire new_AGEMA_signal_8219 ;
    wire new_AGEMA_signal_8220 ;
    wire new_AGEMA_signal_8221 ;
    wire new_AGEMA_signal_8222 ;
    wire new_AGEMA_signal_8223 ;
    wire new_AGEMA_signal_8224 ;
    wire new_AGEMA_signal_8225 ;
    wire new_AGEMA_signal_8226 ;
    wire new_AGEMA_signal_8227 ;
    wire new_AGEMA_signal_8228 ;
    wire new_AGEMA_signal_8229 ;
    wire new_AGEMA_signal_8230 ;
    wire new_AGEMA_signal_8231 ;
    wire new_AGEMA_signal_8232 ;
    wire new_AGEMA_signal_8233 ;
    wire new_AGEMA_signal_8234 ;
    wire new_AGEMA_signal_8235 ;
    wire new_AGEMA_signal_8236 ;
    wire new_AGEMA_signal_8237 ;
    wire new_AGEMA_signal_8238 ;
    wire new_AGEMA_signal_8239 ;
    wire new_AGEMA_signal_8240 ;
    wire new_AGEMA_signal_8241 ;
    wire new_AGEMA_signal_8242 ;
    wire new_AGEMA_signal_8243 ;
    wire new_AGEMA_signal_8244 ;
    wire new_AGEMA_signal_8245 ;
    wire new_AGEMA_signal_8246 ;
    wire new_AGEMA_signal_8247 ;
    wire new_AGEMA_signal_8248 ;
    wire new_AGEMA_signal_8249 ;
    wire new_AGEMA_signal_8250 ;
    wire new_AGEMA_signal_8251 ;
    wire new_AGEMA_signal_8252 ;
    wire new_AGEMA_signal_8253 ;
    wire new_AGEMA_signal_8254 ;
    wire new_AGEMA_signal_8255 ;
    wire new_AGEMA_signal_8256 ;
    wire new_AGEMA_signal_8257 ;
    wire new_AGEMA_signal_8258 ;
    wire new_AGEMA_signal_8259 ;
    wire new_AGEMA_signal_8260 ;
    wire new_AGEMA_signal_8261 ;
    wire new_AGEMA_signal_8262 ;
    wire new_AGEMA_signal_8263 ;
    wire new_AGEMA_signal_8264 ;
    wire new_AGEMA_signal_8265 ;
    wire new_AGEMA_signal_8266 ;
    wire new_AGEMA_signal_8267 ;
    wire new_AGEMA_signal_8268 ;
    wire new_AGEMA_signal_8269 ;
    wire new_AGEMA_signal_8270 ;
    wire new_AGEMA_signal_8271 ;
    wire new_AGEMA_signal_8272 ;
    wire new_AGEMA_signal_8273 ;
    wire new_AGEMA_signal_8274 ;
    wire new_AGEMA_signal_8275 ;
    wire new_AGEMA_signal_8276 ;
    wire new_AGEMA_signal_8277 ;
    wire new_AGEMA_signal_8278 ;
    wire new_AGEMA_signal_8279 ;
    wire new_AGEMA_signal_8280 ;
    wire new_AGEMA_signal_8281 ;
    wire new_AGEMA_signal_8282 ;
    wire new_AGEMA_signal_8283 ;
    wire new_AGEMA_signal_8284 ;
    wire new_AGEMA_signal_8285 ;
    wire new_AGEMA_signal_8286 ;
    wire new_AGEMA_signal_8287 ;
    wire new_AGEMA_signal_8288 ;
    wire new_AGEMA_signal_8289 ;
    wire new_AGEMA_signal_8290 ;
    wire new_AGEMA_signal_8291 ;
    wire new_AGEMA_signal_8292 ;
    wire new_AGEMA_signal_8293 ;
    wire new_AGEMA_signal_8294 ;
    wire new_AGEMA_signal_8295 ;
    wire new_AGEMA_signal_8296 ;
    wire new_AGEMA_signal_8297 ;
    wire new_AGEMA_signal_8298 ;
    wire new_AGEMA_signal_8299 ;
    wire new_AGEMA_signal_8300 ;
    wire new_AGEMA_signal_8301 ;
    wire new_AGEMA_signal_8302 ;
    wire new_AGEMA_signal_8303 ;
    wire new_AGEMA_signal_8304 ;
    wire new_AGEMA_signal_8305 ;
    wire new_AGEMA_signal_8306 ;
    wire new_AGEMA_signal_8307 ;
    wire new_AGEMA_signal_8308 ;
    wire new_AGEMA_signal_8309 ;
    wire new_AGEMA_signal_8310 ;
    wire new_AGEMA_signal_8311 ;
    wire new_AGEMA_signal_8312 ;
    wire new_AGEMA_signal_8313 ;
    wire new_AGEMA_signal_8314 ;
    wire new_AGEMA_signal_8315 ;
    wire new_AGEMA_signal_8316 ;
    wire new_AGEMA_signal_8317 ;
    wire new_AGEMA_signal_8318 ;
    wire new_AGEMA_signal_8319 ;
    wire new_AGEMA_signal_8320 ;
    wire new_AGEMA_signal_8321 ;
    wire new_AGEMA_signal_8322 ;
    wire new_AGEMA_signal_8323 ;
    wire new_AGEMA_signal_8324 ;
    wire new_AGEMA_signal_8325 ;
    wire new_AGEMA_signal_8326 ;
    wire new_AGEMA_signal_8327 ;
    wire new_AGEMA_signal_8328 ;
    wire new_AGEMA_signal_8329 ;
    wire new_AGEMA_signal_8330 ;
    wire new_AGEMA_signal_8331 ;
    wire new_AGEMA_signal_8332 ;
    wire new_AGEMA_signal_8333 ;
    wire new_AGEMA_signal_8334 ;
    wire new_AGEMA_signal_8335 ;
    wire new_AGEMA_signal_8336 ;
    wire new_AGEMA_signal_8337 ;
    wire new_AGEMA_signal_8338 ;
    wire new_AGEMA_signal_8339 ;
    wire new_AGEMA_signal_8340 ;
    wire new_AGEMA_signal_8341 ;
    wire new_AGEMA_signal_8342 ;
    wire new_AGEMA_signal_8343 ;
    wire new_AGEMA_signal_8344 ;
    wire new_AGEMA_signal_8345 ;
    wire new_AGEMA_signal_8346 ;
    wire new_AGEMA_signal_8347 ;
    wire new_AGEMA_signal_8348 ;
    wire new_AGEMA_signal_8349 ;
    wire new_AGEMA_signal_8350 ;
    wire new_AGEMA_signal_8351 ;
    wire new_AGEMA_signal_8352 ;
    wire new_AGEMA_signal_8353 ;
    wire new_AGEMA_signal_8354 ;
    wire new_AGEMA_signal_8355 ;
    wire new_AGEMA_signal_8356 ;
    wire new_AGEMA_signal_8357 ;
    wire new_AGEMA_signal_8358 ;
    wire new_AGEMA_signal_8359 ;
    wire new_AGEMA_signal_8360 ;
    wire new_AGEMA_signal_8361 ;
    wire new_AGEMA_signal_8362 ;
    wire new_AGEMA_signal_8363 ;
    wire new_AGEMA_signal_8364 ;
    wire new_AGEMA_signal_8365 ;
    wire new_AGEMA_signal_8366 ;
    wire new_AGEMA_signal_8367 ;
    wire new_AGEMA_signal_8368 ;
    wire new_AGEMA_signal_8369 ;
    wire new_AGEMA_signal_8370 ;
    wire new_AGEMA_signal_8371 ;
    wire new_AGEMA_signal_8372 ;
    wire new_AGEMA_signal_8373 ;
    wire new_AGEMA_signal_8374 ;
    wire new_AGEMA_signal_8375 ;
    wire new_AGEMA_signal_8376 ;
    wire new_AGEMA_signal_8377 ;
    wire new_AGEMA_signal_8378 ;
    wire new_AGEMA_signal_8379 ;
    wire new_AGEMA_signal_8380 ;
    wire new_AGEMA_signal_8381 ;
    wire new_AGEMA_signal_8382 ;
    wire new_AGEMA_signal_8383 ;
    wire new_AGEMA_signal_8384 ;
    wire new_AGEMA_signal_8385 ;
    wire new_AGEMA_signal_8386 ;
    wire new_AGEMA_signal_8387 ;
    wire new_AGEMA_signal_8388 ;
    wire new_AGEMA_signal_8389 ;
    wire new_AGEMA_signal_8390 ;
    wire new_AGEMA_signal_8391 ;
    wire new_AGEMA_signal_8392 ;
    wire new_AGEMA_signal_8393 ;
    wire new_AGEMA_signal_8394 ;
    wire new_AGEMA_signal_8395 ;
    wire new_AGEMA_signal_8396 ;
    wire new_AGEMA_signal_8397 ;
    wire new_AGEMA_signal_8398 ;
    wire new_AGEMA_signal_8399 ;
    wire new_AGEMA_signal_8400 ;
    wire new_AGEMA_signal_8401 ;
    wire new_AGEMA_signal_8402 ;
    wire new_AGEMA_signal_8403 ;
    wire new_AGEMA_signal_8404 ;
    wire new_AGEMA_signal_8405 ;
    wire new_AGEMA_signal_8406 ;
    wire new_AGEMA_signal_8407 ;
    wire new_AGEMA_signal_8408 ;
    wire new_AGEMA_signal_8409 ;
    wire new_AGEMA_signal_8410 ;
    wire new_AGEMA_signal_8411 ;
    wire new_AGEMA_signal_8412 ;
    wire new_AGEMA_signal_8413 ;
    wire new_AGEMA_signal_8414 ;
    wire new_AGEMA_signal_8415 ;
    wire new_AGEMA_signal_8416 ;
    wire new_AGEMA_signal_8417 ;
    wire new_AGEMA_signal_8418 ;
    wire new_AGEMA_signal_8419 ;
    wire new_AGEMA_signal_8420 ;
    wire new_AGEMA_signal_8421 ;
    wire new_AGEMA_signal_8422 ;
    wire new_AGEMA_signal_8423 ;
    wire new_AGEMA_signal_8424 ;
    wire new_AGEMA_signal_8425 ;
    wire new_AGEMA_signal_8426 ;
    wire new_AGEMA_signal_8427 ;
    wire new_AGEMA_signal_8428 ;
    wire new_AGEMA_signal_8429 ;
    wire new_AGEMA_signal_8430 ;
    wire new_AGEMA_signal_8431 ;
    wire new_AGEMA_signal_8432 ;
    wire new_AGEMA_signal_8433 ;
    wire new_AGEMA_signal_8434 ;
    wire new_AGEMA_signal_8435 ;
    wire new_AGEMA_signal_8436 ;
    wire new_AGEMA_signal_8437 ;
    wire new_AGEMA_signal_8438 ;
    wire new_AGEMA_signal_8439 ;
    wire new_AGEMA_signal_8440 ;
    wire new_AGEMA_signal_8441 ;
    wire new_AGEMA_signal_8442 ;
    wire new_AGEMA_signal_8443 ;
    wire new_AGEMA_signal_8444 ;
    wire new_AGEMA_signal_8445 ;
    wire new_AGEMA_signal_8446 ;
    wire new_AGEMA_signal_8447 ;
    wire new_AGEMA_signal_8448 ;
    wire new_AGEMA_signal_8449 ;
    wire new_AGEMA_signal_8450 ;
    wire new_AGEMA_signal_8451 ;
    wire new_AGEMA_signal_8452 ;
    wire new_AGEMA_signal_8453 ;
    wire new_AGEMA_signal_8454 ;
    wire new_AGEMA_signal_8455 ;
    wire new_AGEMA_signal_8456 ;
    wire new_AGEMA_signal_8457 ;
    wire new_AGEMA_signal_8458 ;
    wire new_AGEMA_signal_8459 ;
    wire new_AGEMA_signal_8460 ;
    wire new_AGEMA_signal_8461 ;
    wire new_AGEMA_signal_8462 ;
    wire new_AGEMA_signal_8463 ;
    wire new_AGEMA_signal_8464 ;
    wire new_AGEMA_signal_8465 ;
    wire new_AGEMA_signal_8466 ;
    wire new_AGEMA_signal_8467 ;
    wire new_AGEMA_signal_8468 ;
    wire new_AGEMA_signal_8469 ;
    wire new_AGEMA_signal_8470 ;
    wire new_AGEMA_signal_8471 ;
    wire new_AGEMA_signal_8472 ;
    wire new_AGEMA_signal_8473 ;
    wire new_AGEMA_signal_8474 ;
    wire new_AGEMA_signal_8475 ;
    wire new_AGEMA_signal_8476 ;
    wire new_AGEMA_signal_8477 ;
    wire new_AGEMA_signal_8478 ;
    wire new_AGEMA_signal_8479 ;
    wire new_AGEMA_signal_8480 ;
    wire new_AGEMA_signal_8481 ;
    wire new_AGEMA_signal_8482 ;
    wire new_AGEMA_signal_8483 ;
    wire new_AGEMA_signal_8484 ;
    wire new_AGEMA_signal_8485 ;
    wire new_AGEMA_signal_8486 ;
    wire new_AGEMA_signal_8487 ;
    wire new_AGEMA_signal_8488 ;
    wire new_AGEMA_signal_8489 ;
    wire new_AGEMA_signal_8490 ;
    wire new_AGEMA_signal_8491 ;
    wire new_AGEMA_signal_8492 ;
    wire new_AGEMA_signal_8493 ;
    wire new_AGEMA_signal_8494 ;
    wire new_AGEMA_signal_8495 ;
    wire new_AGEMA_signal_8496 ;
    wire new_AGEMA_signal_8497 ;
    wire new_AGEMA_signal_8498 ;
    wire new_AGEMA_signal_8499 ;
    wire new_AGEMA_signal_8500 ;
    wire new_AGEMA_signal_8501 ;
    wire new_AGEMA_signal_8502 ;
    wire new_AGEMA_signal_8503 ;
    wire new_AGEMA_signal_8504 ;
    wire new_AGEMA_signal_8505 ;
    wire new_AGEMA_signal_8506 ;
    wire new_AGEMA_signal_8507 ;
    wire new_AGEMA_signal_8508 ;
    wire new_AGEMA_signal_8509 ;
    wire new_AGEMA_signal_8510 ;
    wire new_AGEMA_signal_8511 ;
    wire new_AGEMA_signal_8512 ;
    wire new_AGEMA_signal_8513 ;
    wire new_AGEMA_signal_8514 ;
    wire new_AGEMA_signal_8515 ;
    wire new_AGEMA_signal_8516 ;
    wire new_AGEMA_signal_8517 ;
    wire new_AGEMA_signal_8518 ;
    wire new_AGEMA_signal_8519 ;
    wire new_AGEMA_signal_8520 ;
    wire new_AGEMA_signal_8521 ;
    wire new_AGEMA_signal_8522 ;
    wire new_AGEMA_signal_8523 ;
    wire new_AGEMA_signal_8524 ;
    wire new_AGEMA_signal_8525 ;
    wire new_AGEMA_signal_8526 ;
    wire new_AGEMA_signal_8527 ;
    wire new_AGEMA_signal_8528 ;
    wire new_AGEMA_signal_8529 ;
    wire new_AGEMA_signal_8530 ;
    wire new_AGEMA_signal_8531 ;
    wire new_AGEMA_signal_8532 ;
    wire new_AGEMA_signal_8533 ;
    wire new_AGEMA_signal_8534 ;
    wire new_AGEMA_signal_8535 ;
    wire new_AGEMA_signal_8536 ;
    wire new_AGEMA_signal_8537 ;
    wire new_AGEMA_signal_8538 ;
    wire new_AGEMA_signal_8539 ;
    wire new_AGEMA_signal_8540 ;
    wire new_AGEMA_signal_8541 ;
    wire new_AGEMA_signal_8542 ;
    wire new_AGEMA_signal_8543 ;
    wire new_AGEMA_signal_8544 ;
    wire new_AGEMA_signal_8545 ;
    wire new_AGEMA_signal_8546 ;
    wire new_AGEMA_signal_8547 ;
    wire new_AGEMA_signal_8548 ;
    wire new_AGEMA_signal_8549 ;
    wire new_AGEMA_signal_8550 ;
    wire new_AGEMA_signal_8551 ;
    wire new_AGEMA_signal_8552 ;
    wire new_AGEMA_signal_8553 ;
    wire new_AGEMA_signal_8554 ;
    wire new_AGEMA_signal_8555 ;
    wire new_AGEMA_signal_8556 ;
    wire new_AGEMA_signal_8557 ;
    wire new_AGEMA_signal_8558 ;
    wire new_AGEMA_signal_8559 ;
    wire new_AGEMA_signal_8560 ;
    wire new_AGEMA_signal_8561 ;
    wire new_AGEMA_signal_8562 ;
    wire new_AGEMA_signal_8563 ;
    wire new_AGEMA_signal_8564 ;
    wire new_AGEMA_signal_8565 ;
    wire new_AGEMA_signal_8566 ;
    wire new_AGEMA_signal_8567 ;
    wire new_AGEMA_signal_8568 ;
    wire new_AGEMA_signal_8569 ;
    wire new_AGEMA_signal_8570 ;
    wire new_AGEMA_signal_8571 ;
    wire new_AGEMA_signal_8572 ;
    wire new_AGEMA_signal_8573 ;
    wire new_AGEMA_signal_8574 ;
    wire new_AGEMA_signal_8575 ;
    wire new_AGEMA_signal_8576 ;
    wire new_AGEMA_signal_8577 ;
    wire new_AGEMA_signal_8578 ;
    wire new_AGEMA_signal_8579 ;
    wire new_AGEMA_signal_8580 ;
    wire new_AGEMA_signal_8581 ;
    wire new_AGEMA_signal_8582 ;
    wire new_AGEMA_signal_8583 ;
    wire new_AGEMA_signal_8584 ;
    wire new_AGEMA_signal_8585 ;
    wire new_AGEMA_signal_8586 ;
    wire new_AGEMA_signal_8587 ;
    wire new_AGEMA_signal_8588 ;
    wire new_AGEMA_signal_8589 ;
    wire new_AGEMA_signal_8590 ;
    wire new_AGEMA_signal_8591 ;
    wire new_AGEMA_signal_8592 ;
    wire new_AGEMA_signal_8593 ;
    wire new_AGEMA_signal_8594 ;
    wire new_AGEMA_signal_8595 ;
    wire new_AGEMA_signal_8596 ;
    wire new_AGEMA_signal_8597 ;
    wire new_AGEMA_signal_8598 ;
    wire new_AGEMA_signal_8599 ;
    wire new_AGEMA_signal_8600 ;
    wire new_AGEMA_signal_8601 ;
    wire new_AGEMA_signal_8602 ;
    wire new_AGEMA_signal_8603 ;
    wire new_AGEMA_signal_8604 ;
    wire new_AGEMA_signal_8605 ;
    wire new_AGEMA_signal_8606 ;
    wire new_AGEMA_signal_8607 ;
    wire new_AGEMA_signal_8608 ;
    wire new_AGEMA_signal_8609 ;
    wire new_AGEMA_signal_8610 ;
    wire new_AGEMA_signal_8611 ;
    wire new_AGEMA_signal_8612 ;
    wire new_AGEMA_signal_8613 ;
    wire new_AGEMA_signal_8614 ;
    wire new_AGEMA_signal_8615 ;
    wire new_AGEMA_signal_8616 ;
    wire new_AGEMA_signal_8617 ;
    wire new_AGEMA_signal_8618 ;
    wire new_AGEMA_signal_8619 ;
    wire new_AGEMA_signal_8620 ;
    wire new_AGEMA_signal_8621 ;
    wire new_AGEMA_signal_8622 ;
    wire new_AGEMA_signal_8623 ;
    wire new_AGEMA_signal_8624 ;
    wire new_AGEMA_signal_8625 ;
    wire new_AGEMA_signal_8626 ;
    wire new_AGEMA_signal_8627 ;
    wire new_AGEMA_signal_8628 ;
    wire new_AGEMA_signal_8629 ;
    wire new_AGEMA_signal_8630 ;
    wire new_AGEMA_signal_8631 ;
    wire new_AGEMA_signal_8632 ;
    wire new_AGEMA_signal_8633 ;
    wire new_AGEMA_signal_8634 ;
    wire new_AGEMA_signal_8635 ;
    wire new_AGEMA_signal_8636 ;
    wire new_AGEMA_signal_8637 ;
    wire new_AGEMA_signal_8638 ;
    wire new_AGEMA_signal_8639 ;
    wire new_AGEMA_signal_8640 ;
    wire new_AGEMA_signal_8641 ;
    wire new_AGEMA_signal_8642 ;
    wire new_AGEMA_signal_8643 ;
    wire new_AGEMA_signal_8644 ;
    wire new_AGEMA_signal_8645 ;
    wire new_AGEMA_signal_8646 ;
    wire new_AGEMA_signal_8647 ;
    wire new_AGEMA_signal_8648 ;
    wire new_AGEMA_signal_8649 ;
    wire new_AGEMA_signal_8650 ;
    wire new_AGEMA_signal_8651 ;
    wire new_AGEMA_signal_8652 ;
    wire new_AGEMA_signal_8653 ;
    wire new_AGEMA_signal_8654 ;
    wire new_AGEMA_signal_8655 ;
    wire new_AGEMA_signal_8656 ;
    wire new_AGEMA_signal_8657 ;
    wire new_AGEMA_signal_8658 ;
    wire new_AGEMA_signal_8659 ;
    wire new_AGEMA_signal_8660 ;
    wire new_AGEMA_signal_8661 ;
    wire new_AGEMA_signal_8662 ;
    wire new_AGEMA_signal_8663 ;
    wire new_AGEMA_signal_8664 ;
    wire new_AGEMA_signal_8665 ;
    wire new_AGEMA_signal_8666 ;
    wire new_AGEMA_signal_8667 ;
    wire new_AGEMA_signal_8668 ;
    wire new_AGEMA_signal_8669 ;
    wire new_AGEMA_signal_8670 ;
    wire new_AGEMA_signal_8671 ;
    wire new_AGEMA_signal_8672 ;
    wire new_AGEMA_signal_8673 ;
    wire new_AGEMA_signal_8674 ;
    wire new_AGEMA_signal_8675 ;
    wire new_AGEMA_signal_8676 ;
    wire new_AGEMA_signal_8677 ;
    wire new_AGEMA_signal_8678 ;
    wire new_AGEMA_signal_8679 ;
    wire new_AGEMA_signal_8680 ;
    wire new_AGEMA_signal_8681 ;
    wire new_AGEMA_signal_8682 ;
    wire new_AGEMA_signal_8683 ;
    wire new_AGEMA_signal_8684 ;
    wire new_AGEMA_signal_8685 ;
    wire new_AGEMA_signal_8686 ;
    wire new_AGEMA_signal_8687 ;
    wire new_AGEMA_signal_8688 ;
    wire new_AGEMA_signal_8689 ;
    wire new_AGEMA_signal_8690 ;
    wire new_AGEMA_signal_8691 ;
    wire new_AGEMA_signal_8692 ;
    wire new_AGEMA_signal_8693 ;
    wire new_AGEMA_signal_8694 ;
    wire new_AGEMA_signal_8695 ;
    wire new_AGEMA_signal_8696 ;
    wire new_AGEMA_signal_8697 ;
    wire new_AGEMA_signal_8698 ;
    wire new_AGEMA_signal_8699 ;
    wire new_AGEMA_signal_8700 ;
    wire new_AGEMA_signal_8701 ;
    wire new_AGEMA_signal_8702 ;
    wire new_AGEMA_signal_8703 ;
    wire new_AGEMA_signal_8704 ;
    wire new_AGEMA_signal_8705 ;
    wire new_AGEMA_signal_8706 ;
    wire new_AGEMA_signal_8707 ;
    wire new_AGEMA_signal_8708 ;
    wire new_AGEMA_signal_8709 ;
    wire new_AGEMA_signal_8710 ;
    wire new_AGEMA_signal_8711 ;
    wire new_AGEMA_signal_8712 ;
    wire new_AGEMA_signal_8713 ;
    wire new_AGEMA_signal_8714 ;
    wire new_AGEMA_signal_8715 ;
    wire new_AGEMA_signal_8716 ;
    wire new_AGEMA_signal_8717 ;
    wire new_AGEMA_signal_8718 ;
    wire new_AGEMA_signal_8719 ;
    wire new_AGEMA_signal_8720 ;
    wire new_AGEMA_signal_8721 ;
    wire new_AGEMA_signal_8722 ;
    wire new_AGEMA_signal_8723 ;
    wire new_AGEMA_signal_8724 ;
    wire new_AGEMA_signal_8725 ;
    wire new_AGEMA_signal_8726 ;
    wire new_AGEMA_signal_8727 ;
    wire new_AGEMA_signal_8728 ;
    wire new_AGEMA_signal_8729 ;
    wire new_AGEMA_signal_8730 ;
    wire new_AGEMA_signal_8731 ;
    wire new_AGEMA_signal_8732 ;
    wire new_AGEMA_signal_8733 ;
    wire new_AGEMA_signal_8734 ;
    wire new_AGEMA_signal_8735 ;
    wire new_AGEMA_signal_8736 ;
    wire new_AGEMA_signal_8737 ;
    wire new_AGEMA_signal_8738 ;
    wire new_AGEMA_signal_8739 ;
    wire new_AGEMA_signal_8740 ;
    wire new_AGEMA_signal_8741 ;
    wire new_AGEMA_signal_8742 ;
    wire new_AGEMA_signal_8743 ;
    wire new_AGEMA_signal_8744 ;
    wire new_AGEMA_signal_8745 ;
    wire new_AGEMA_signal_8746 ;
    wire new_AGEMA_signal_8747 ;
    wire new_AGEMA_signal_8748 ;
    wire new_AGEMA_signal_8749 ;
    wire new_AGEMA_signal_8750 ;
    wire new_AGEMA_signal_8751 ;
    wire new_AGEMA_signal_8752 ;
    wire new_AGEMA_signal_8753 ;
    wire new_AGEMA_signal_8754 ;
    wire new_AGEMA_signal_8755 ;
    wire new_AGEMA_signal_8756 ;
    wire new_AGEMA_signal_8757 ;
    wire new_AGEMA_signal_8758 ;
    wire new_AGEMA_signal_8759 ;
    wire new_AGEMA_signal_8760 ;
    wire new_AGEMA_signal_8761 ;
    wire new_AGEMA_signal_8762 ;
    wire new_AGEMA_signal_8763 ;
    wire new_AGEMA_signal_8764 ;
    wire new_AGEMA_signal_8765 ;
    wire new_AGEMA_signal_8766 ;
    wire new_AGEMA_signal_8767 ;
    wire new_AGEMA_signal_8768 ;
    wire new_AGEMA_signal_8769 ;
    wire new_AGEMA_signal_8770 ;
    wire new_AGEMA_signal_8771 ;
    wire new_AGEMA_signal_8772 ;
    wire new_AGEMA_signal_8773 ;
    wire new_AGEMA_signal_8774 ;
    wire new_AGEMA_signal_8775 ;
    wire new_AGEMA_signal_8776 ;
    wire new_AGEMA_signal_8777 ;
    wire new_AGEMA_signal_8778 ;
    wire new_AGEMA_signal_8779 ;
    wire new_AGEMA_signal_8780 ;
    wire new_AGEMA_signal_8781 ;
    wire new_AGEMA_signal_8782 ;
    wire new_AGEMA_signal_8783 ;
    wire new_AGEMA_signal_8784 ;
    wire new_AGEMA_signal_8785 ;
    wire new_AGEMA_signal_8786 ;
    wire new_AGEMA_signal_8787 ;
    wire new_AGEMA_signal_8788 ;
    wire new_AGEMA_signal_8789 ;
    wire new_AGEMA_signal_8790 ;
    wire new_AGEMA_signal_8791 ;
    wire new_AGEMA_signal_8792 ;
    wire new_AGEMA_signal_8793 ;
    wire new_AGEMA_signal_8794 ;
    wire new_AGEMA_signal_8795 ;
    wire new_AGEMA_signal_8796 ;
    wire new_AGEMA_signal_8797 ;
    wire new_AGEMA_signal_8798 ;
    wire new_AGEMA_signal_8799 ;
    wire new_AGEMA_signal_8800 ;
    wire new_AGEMA_signal_8801 ;
    wire new_AGEMA_signal_8802 ;
    wire new_AGEMA_signal_8803 ;
    wire new_AGEMA_signal_8804 ;
    wire new_AGEMA_signal_8805 ;
    wire new_AGEMA_signal_8806 ;
    wire new_AGEMA_signal_8807 ;
    wire new_AGEMA_signal_8808 ;
    wire new_AGEMA_signal_8809 ;
    wire new_AGEMA_signal_8810 ;
    wire new_AGEMA_signal_8811 ;
    wire new_AGEMA_signal_8812 ;
    wire new_AGEMA_signal_8813 ;
    wire new_AGEMA_signal_8814 ;
    wire new_AGEMA_signal_8815 ;
    wire new_AGEMA_signal_8816 ;
    wire new_AGEMA_signal_8817 ;
    wire new_AGEMA_signal_8818 ;
    wire new_AGEMA_signal_8819 ;
    wire new_AGEMA_signal_8820 ;
    wire new_AGEMA_signal_8821 ;
    wire new_AGEMA_signal_8822 ;
    wire new_AGEMA_signal_8823 ;
    wire new_AGEMA_signal_8824 ;
    wire new_AGEMA_signal_8825 ;
    wire new_AGEMA_signal_8826 ;
    wire new_AGEMA_signal_8827 ;
    wire new_AGEMA_signal_8828 ;
    wire new_AGEMA_signal_8829 ;
    wire new_AGEMA_signal_8830 ;
    wire new_AGEMA_signal_8831 ;
    wire new_AGEMA_signal_8832 ;
    wire new_AGEMA_signal_8833 ;
    wire new_AGEMA_signal_8834 ;
    wire new_AGEMA_signal_8835 ;
    wire new_AGEMA_signal_8836 ;
    wire new_AGEMA_signal_8837 ;
    wire new_AGEMA_signal_8838 ;
    wire new_AGEMA_signal_8839 ;
    wire new_AGEMA_signal_8840 ;
    wire new_AGEMA_signal_8841 ;
    wire new_AGEMA_signal_8842 ;
    wire new_AGEMA_signal_8843 ;
    wire new_AGEMA_signal_8844 ;
    wire new_AGEMA_signal_8845 ;
    wire new_AGEMA_signal_8846 ;
    wire new_AGEMA_signal_8847 ;
    wire new_AGEMA_signal_8848 ;
    wire new_AGEMA_signal_8849 ;
    wire new_AGEMA_signal_8850 ;
    wire new_AGEMA_signal_8851 ;
    wire new_AGEMA_signal_8852 ;
    wire new_AGEMA_signal_8853 ;
    wire new_AGEMA_signal_8854 ;
    wire new_AGEMA_signal_8855 ;
    wire new_AGEMA_signal_8856 ;
    wire new_AGEMA_signal_8857 ;
    wire new_AGEMA_signal_8858 ;
    wire new_AGEMA_signal_8859 ;
    wire new_AGEMA_signal_8860 ;
    wire new_AGEMA_signal_8861 ;
    wire new_AGEMA_signal_8862 ;
    wire new_AGEMA_signal_8863 ;
    wire new_AGEMA_signal_8864 ;
    wire new_AGEMA_signal_8865 ;
    wire new_AGEMA_signal_8866 ;
    wire new_AGEMA_signal_8867 ;
    wire new_AGEMA_signal_8868 ;
    wire new_AGEMA_signal_8869 ;
    wire new_AGEMA_signal_8870 ;
    wire new_AGEMA_signal_8871 ;
    wire new_AGEMA_signal_8872 ;
    wire new_AGEMA_signal_8873 ;
    wire new_AGEMA_signal_8874 ;
    wire new_AGEMA_signal_8875 ;
    wire new_AGEMA_signal_8876 ;
    wire new_AGEMA_signal_8877 ;
    wire new_AGEMA_signal_8878 ;
    wire new_AGEMA_signal_8879 ;
    wire new_AGEMA_signal_8880 ;
    wire new_AGEMA_signal_8881 ;
    wire new_AGEMA_signal_8882 ;
    wire new_AGEMA_signal_8883 ;
    wire new_AGEMA_signal_8884 ;
    wire new_AGEMA_signal_8885 ;
    wire new_AGEMA_signal_8886 ;
    wire new_AGEMA_signal_8887 ;
    wire new_AGEMA_signal_8888 ;
    wire new_AGEMA_signal_8889 ;
    wire new_AGEMA_signal_8890 ;
    wire new_AGEMA_signal_8891 ;
    wire new_AGEMA_signal_8892 ;
    wire new_AGEMA_signal_8893 ;
    wire new_AGEMA_signal_8894 ;
    wire new_AGEMA_signal_8895 ;
    wire new_AGEMA_signal_8896 ;
    wire new_AGEMA_signal_8897 ;
    wire new_AGEMA_signal_8898 ;
    wire new_AGEMA_signal_8899 ;
    wire new_AGEMA_signal_8900 ;
    wire new_AGEMA_signal_8901 ;
    wire new_AGEMA_signal_8902 ;
    wire new_AGEMA_signal_8903 ;
    wire new_AGEMA_signal_8904 ;
    wire new_AGEMA_signal_8905 ;
    wire new_AGEMA_signal_8906 ;
    wire new_AGEMA_signal_8907 ;
    wire new_AGEMA_signal_8908 ;
    wire new_AGEMA_signal_8909 ;
    wire new_AGEMA_signal_8910 ;
    wire new_AGEMA_signal_8911 ;
    wire new_AGEMA_signal_8912 ;
    wire new_AGEMA_signal_8913 ;
    wire new_AGEMA_signal_8914 ;
    wire new_AGEMA_signal_8915 ;
    wire new_AGEMA_signal_8916 ;
    wire new_AGEMA_signal_8917 ;
    wire new_AGEMA_signal_8918 ;
    wire new_AGEMA_signal_8919 ;
    wire new_AGEMA_signal_8920 ;
    wire new_AGEMA_signal_8921 ;
    wire new_AGEMA_signal_8922 ;
    wire new_AGEMA_signal_8923 ;
    wire new_AGEMA_signal_8924 ;
    wire new_AGEMA_signal_8925 ;
    wire new_AGEMA_signal_8926 ;
    wire new_AGEMA_signal_8927 ;
    wire new_AGEMA_signal_8928 ;
    wire new_AGEMA_signal_8929 ;
    wire new_AGEMA_signal_8930 ;
    wire new_AGEMA_signal_8931 ;
    wire new_AGEMA_signal_8932 ;
    wire new_AGEMA_signal_8933 ;
    wire new_AGEMA_signal_8934 ;
    wire new_AGEMA_signal_8935 ;
    wire new_AGEMA_signal_8936 ;
    wire new_AGEMA_signal_8937 ;
    wire new_AGEMA_signal_8938 ;
    wire new_AGEMA_signal_8939 ;
    wire new_AGEMA_signal_8940 ;
    wire new_AGEMA_signal_8941 ;
    wire new_AGEMA_signal_8942 ;
    wire new_AGEMA_signal_8943 ;
    wire new_AGEMA_signal_8944 ;
    wire new_AGEMA_signal_8945 ;
    wire new_AGEMA_signal_8946 ;
    wire new_AGEMA_signal_8947 ;
    wire new_AGEMA_signal_8948 ;
    wire new_AGEMA_signal_8949 ;
    wire new_AGEMA_signal_8950 ;
    wire new_AGEMA_signal_8951 ;
    wire new_AGEMA_signal_8952 ;
    wire new_AGEMA_signal_8953 ;
    wire new_AGEMA_signal_8954 ;
    wire new_AGEMA_signal_8955 ;
    wire new_AGEMA_signal_8956 ;
    wire new_AGEMA_signal_8957 ;
    wire new_AGEMA_signal_8958 ;
    wire new_AGEMA_signal_8959 ;
    wire new_AGEMA_signal_8960 ;
    wire new_AGEMA_signal_8961 ;
    wire new_AGEMA_signal_8962 ;
    wire new_AGEMA_signal_8963 ;
    wire new_AGEMA_signal_8964 ;
    wire new_AGEMA_signal_8965 ;
    wire new_AGEMA_signal_8966 ;
    wire new_AGEMA_signal_8967 ;
    wire new_AGEMA_signal_8968 ;
    wire new_AGEMA_signal_8969 ;
    wire new_AGEMA_signal_8970 ;
    wire new_AGEMA_signal_8971 ;
    wire new_AGEMA_signal_8972 ;
    wire new_AGEMA_signal_8973 ;
    wire new_AGEMA_signal_8974 ;
    wire new_AGEMA_signal_8975 ;
    wire new_AGEMA_signal_8976 ;
    wire new_AGEMA_signal_8977 ;
    wire new_AGEMA_signal_8978 ;
    wire new_AGEMA_signal_8979 ;
    wire new_AGEMA_signal_8980 ;
    wire new_AGEMA_signal_8981 ;
    wire new_AGEMA_signal_8982 ;
    wire new_AGEMA_signal_8983 ;
    wire new_AGEMA_signal_8984 ;
    wire new_AGEMA_signal_8985 ;
    wire new_AGEMA_signal_8986 ;
    wire new_AGEMA_signal_8987 ;
    wire new_AGEMA_signal_8988 ;
    wire new_AGEMA_signal_8989 ;
    wire new_AGEMA_signal_8990 ;
    wire new_AGEMA_signal_8991 ;
    wire new_AGEMA_signal_8992 ;
    wire new_AGEMA_signal_8993 ;
    wire new_AGEMA_signal_8994 ;
    wire new_AGEMA_signal_8995 ;
    wire new_AGEMA_signal_8996 ;
    wire new_AGEMA_signal_8997 ;
    wire new_AGEMA_signal_8998 ;
    wire new_AGEMA_signal_8999 ;
    wire new_AGEMA_signal_9000 ;
    wire new_AGEMA_signal_9001 ;
    wire new_AGEMA_signal_9002 ;
    wire new_AGEMA_signal_9003 ;
    wire new_AGEMA_signal_9004 ;
    wire new_AGEMA_signal_9005 ;
    wire new_AGEMA_signal_9006 ;
    wire new_AGEMA_signal_9007 ;
    wire new_AGEMA_signal_9008 ;
    wire new_AGEMA_signal_9009 ;
    wire new_AGEMA_signal_9010 ;
    wire new_AGEMA_signal_9011 ;
    wire new_AGEMA_signal_9012 ;
    wire new_AGEMA_signal_9013 ;
    wire new_AGEMA_signal_9014 ;
    wire new_AGEMA_signal_9015 ;
    wire new_AGEMA_signal_9016 ;
    wire new_AGEMA_signal_9017 ;
    wire new_AGEMA_signal_9018 ;
    wire new_AGEMA_signal_9019 ;
    wire new_AGEMA_signal_9020 ;
    wire new_AGEMA_signal_9021 ;
    wire new_AGEMA_signal_9022 ;
    wire new_AGEMA_signal_9023 ;
    wire new_AGEMA_signal_9024 ;
    wire new_AGEMA_signal_9025 ;
    wire new_AGEMA_signal_9026 ;
    wire new_AGEMA_signal_9027 ;
    wire new_AGEMA_signal_9028 ;
    wire new_AGEMA_signal_9029 ;
    wire new_AGEMA_signal_9030 ;
    wire new_AGEMA_signal_9031 ;
    wire new_AGEMA_signal_9032 ;
    wire new_AGEMA_signal_9033 ;
    wire new_AGEMA_signal_9034 ;
    wire new_AGEMA_signal_9035 ;
    wire new_AGEMA_signal_9036 ;
    wire new_AGEMA_signal_9037 ;
    wire new_AGEMA_signal_9038 ;
    wire new_AGEMA_signal_9039 ;
    wire new_AGEMA_signal_9040 ;
    wire new_AGEMA_signal_9041 ;
    wire new_AGEMA_signal_9042 ;
    wire new_AGEMA_signal_9043 ;
    wire new_AGEMA_signal_9044 ;
    wire new_AGEMA_signal_9045 ;
    wire new_AGEMA_signal_9046 ;
    wire new_AGEMA_signal_9047 ;
    wire new_AGEMA_signal_9048 ;
    wire new_AGEMA_signal_9049 ;
    wire new_AGEMA_signal_9050 ;
    wire new_AGEMA_signal_9051 ;
    wire new_AGEMA_signal_9052 ;
    wire new_AGEMA_signal_9053 ;
    wire new_AGEMA_signal_9054 ;
    wire new_AGEMA_signal_9055 ;
    wire new_AGEMA_signal_9056 ;
    wire new_AGEMA_signal_9057 ;
    wire new_AGEMA_signal_9058 ;
    wire new_AGEMA_signal_9059 ;
    wire new_AGEMA_signal_9060 ;
    wire new_AGEMA_signal_9061 ;
    wire new_AGEMA_signal_9062 ;
    wire new_AGEMA_signal_9063 ;
    wire new_AGEMA_signal_9064 ;
    wire new_AGEMA_signal_9065 ;
    wire new_AGEMA_signal_9066 ;
    wire new_AGEMA_signal_9067 ;
    wire new_AGEMA_signal_9068 ;
    wire new_AGEMA_signal_9069 ;
    wire new_AGEMA_signal_9070 ;
    wire new_AGEMA_signal_9071 ;
    wire new_AGEMA_signal_9072 ;
    wire new_AGEMA_signal_9073 ;
    wire new_AGEMA_signal_9074 ;
    wire new_AGEMA_signal_9075 ;
    wire new_AGEMA_signal_9076 ;
    wire new_AGEMA_signal_9077 ;
    wire new_AGEMA_signal_9078 ;
    wire new_AGEMA_signal_9079 ;
    wire new_AGEMA_signal_9080 ;
    wire new_AGEMA_signal_9081 ;
    wire new_AGEMA_signal_9082 ;
    wire new_AGEMA_signal_9083 ;
    wire new_AGEMA_signal_9084 ;
    wire new_AGEMA_signal_9085 ;
    wire new_AGEMA_signal_9086 ;
    wire new_AGEMA_signal_9087 ;
    wire new_AGEMA_signal_9088 ;
    wire new_AGEMA_signal_9089 ;
    wire new_AGEMA_signal_9090 ;
    wire new_AGEMA_signal_9091 ;
    wire new_AGEMA_signal_9092 ;
    wire new_AGEMA_signal_9093 ;
    wire new_AGEMA_signal_9094 ;
    wire new_AGEMA_signal_9095 ;
    wire new_AGEMA_signal_9096 ;
    wire new_AGEMA_signal_9097 ;
    wire new_AGEMA_signal_9098 ;
    wire new_AGEMA_signal_9099 ;
    wire new_AGEMA_signal_9100 ;
    wire new_AGEMA_signal_9101 ;
    wire new_AGEMA_signal_9102 ;
    wire new_AGEMA_signal_9103 ;
    wire new_AGEMA_signal_9104 ;
    wire new_AGEMA_signal_9105 ;
    wire new_AGEMA_signal_9106 ;
    wire new_AGEMA_signal_9107 ;
    wire new_AGEMA_signal_9108 ;
    wire new_AGEMA_signal_9109 ;
    wire new_AGEMA_signal_9110 ;
    wire new_AGEMA_signal_9111 ;
    wire new_AGEMA_signal_9112 ;
    wire new_AGEMA_signal_9113 ;
    wire new_AGEMA_signal_9114 ;
    wire new_AGEMA_signal_9115 ;
    wire new_AGEMA_signal_9116 ;
    wire new_AGEMA_signal_9117 ;
    wire new_AGEMA_signal_9118 ;
    wire new_AGEMA_signal_9119 ;
    wire new_AGEMA_signal_9120 ;
    wire new_AGEMA_signal_9121 ;
    wire new_AGEMA_signal_9122 ;
    wire new_AGEMA_signal_9123 ;
    wire new_AGEMA_signal_9124 ;
    wire new_AGEMA_signal_9125 ;
    wire new_AGEMA_signal_9126 ;
    wire new_AGEMA_signal_9127 ;
    wire new_AGEMA_signal_9128 ;
    wire new_AGEMA_signal_9129 ;
    wire new_AGEMA_signal_9130 ;
    wire new_AGEMA_signal_9131 ;
    wire new_AGEMA_signal_9132 ;
    wire new_AGEMA_signal_9133 ;
    wire new_AGEMA_signal_9134 ;
    wire new_AGEMA_signal_9135 ;
    wire new_AGEMA_signal_9136 ;
    wire new_AGEMA_signal_9137 ;
    wire new_AGEMA_signal_9138 ;
    wire new_AGEMA_signal_9139 ;
    wire new_AGEMA_signal_9140 ;
    wire new_AGEMA_signal_9141 ;
    wire new_AGEMA_signal_9142 ;
    wire new_AGEMA_signal_9143 ;
    wire new_AGEMA_signal_9144 ;
    wire new_AGEMA_signal_9145 ;
    wire new_AGEMA_signal_9146 ;
    wire new_AGEMA_signal_9147 ;
    wire new_AGEMA_signal_9148 ;
    wire new_AGEMA_signal_9149 ;
    wire new_AGEMA_signal_9150 ;
    wire new_AGEMA_signal_9151 ;
    wire new_AGEMA_signal_9152 ;
    wire new_AGEMA_signal_9153 ;
    wire new_AGEMA_signal_9154 ;
    wire new_AGEMA_signal_9155 ;
    wire new_AGEMA_signal_9156 ;
    wire new_AGEMA_signal_9157 ;
    wire new_AGEMA_signal_9158 ;
    wire new_AGEMA_signal_9159 ;
    wire new_AGEMA_signal_9160 ;
    wire new_AGEMA_signal_9161 ;
    wire new_AGEMA_signal_9162 ;
    wire new_AGEMA_signal_9163 ;
    wire new_AGEMA_signal_9164 ;
    wire new_AGEMA_signal_9165 ;
    wire new_AGEMA_signal_9166 ;
    wire new_AGEMA_signal_9167 ;
    wire new_AGEMA_signal_9168 ;
    wire new_AGEMA_signal_9169 ;
    wire new_AGEMA_signal_9170 ;
    wire new_AGEMA_signal_9171 ;
    wire new_AGEMA_signal_9172 ;
    wire new_AGEMA_signal_9173 ;
    wire new_AGEMA_signal_9174 ;
    wire new_AGEMA_signal_9175 ;
    wire new_AGEMA_signal_9176 ;
    wire new_AGEMA_signal_9177 ;
    wire new_AGEMA_signal_9178 ;
    wire new_AGEMA_signal_9179 ;
    wire new_AGEMA_signal_9180 ;
    wire new_AGEMA_signal_9181 ;
    wire new_AGEMA_signal_9182 ;
    wire new_AGEMA_signal_9183 ;
    wire new_AGEMA_signal_9184 ;
    wire new_AGEMA_signal_9185 ;
    wire new_AGEMA_signal_9186 ;
    wire new_AGEMA_signal_9187 ;
    wire new_AGEMA_signal_9188 ;
    wire new_AGEMA_signal_9189 ;
    wire new_AGEMA_signal_9190 ;
    wire new_AGEMA_signal_9191 ;
    wire new_AGEMA_signal_9192 ;
    wire new_AGEMA_signal_9193 ;
    wire new_AGEMA_signal_9194 ;
    wire new_AGEMA_signal_9195 ;
    wire new_AGEMA_signal_9196 ;
    wire new_AGEMA_signal_9197 ;
    wire new_AGEMA_signal_9198 ;
    wire new_AGEMA_signal_9199 ;
    wire new_AGEMA_signal_9200 ;
    wire new_AGEMA_signal_9201 ;
    wire new_AGEMA_signal_9202 ;
    wire new_AGEMA_signal_9203 ;
    wire new_AGEMA_signal_9204 ;
    wire new_AGEMA_signal_9205 ;
    wire new_AGEMA_signal_9206 ;
    wire new_AGEMA_signal_9207 ;
    wire new_AGEMA_signal_9208 ;
    wire new_AGEMA_signal_9209 ;
    wire new_AGEMA_signal_9210 ;
    wire new_AGEMA_signal_9211 ;
    wire new_AGEMA_signal_9212 ;
    wire new_AGEMA_signal_9213 ;
    wire new_AGEMA_signal_9214 ;
    wire new_AGEMA_signal_9215 ;
    wire new_AGEMA_signal_9216 ;
    wire new_AGEMA_signal_9217 ;
    wire new_AGEMA_signal_9218 ;
    wire new_AGEMA_signal_9219 ;
    wire new_AGEMA_signal_9220 ;
    wire new_AGEMA_signal_9221 ;
    wire new_AGEMA_signal_9222 ;
    wire new_AGEMA_signal_9223 ;
    wire new_AGEMA_signal_9224 ;
    wire new_AGEMA_signal_9225 ;
    wire new_AGEMA_signal_9226 ;
    wire new_AGEMA_signal_9227 ;
    wire new_AGEMA_signal_9228 ;
    wire new_AGEMA_signal_9229 ;
    wire new_AGEMA_signal_9230 ;
    wire new_AGEMA_signal_9231 ;
    wire new_AGEMA_signal_9232 ;
    wire new_AGEMA_signal_9233 ;
    wire new_AGEMA_signal_9234 ;
    wire new_AGEMA_signal_9235 ;
    wire new_AGEMA_signal_9236 ;
    wire new_AGEMA_signal_9237 ;
    wire new_AGEMA_signal_9238 ;
    wire new_AGEMA_signal_9239 ;
    wire new_AGEMA_signal_9240 ;
    wire new_AGEMA_signal_9241 ;
    wire new_AGEMA_signal_9242 ;
    wire new_AGEMA_signal_9243 ;
    wire new_AGEMA_signal_9244 ;
    wire new_AGEMA_signal_9245 ;
    wire new_AGEMA_signal_9246 ;
    wire new_AGEMA_signal_9247 ;
    wire new_AGEMA_signal_9248 ;
    wire new_AGEMA_signal_9249 ;
    wire new_AGEMA_signal_9250 ;
    wire new_AGEMA_signal_9251 ;
    wire new_AGEMA_signal_9252 ;
    wire new_AGEMA_signal_9253 ;
    wire new_AGEMA_signal_9254 ;
    wire new_AGEMA_signal_9255 ;
    wire new_AGEMA_signal_9256 ;
    wire new_AGEMA_signal_9257 ;
    wire new_AGEMA_signal_9258 ;
    wire new_AGEMA_signal_9259 ;
    wire new_AGEMA_signal_9260 ;
    wire new_AGEMA_signal_9261 ;
    wire new_AGEMA_signal_9262 ;
    wire new_AGEMA_signal_9263 ;
    wire new_AGEMA_signal_9264 ;
    wire new_AGEMA_signal_9265 ;
    wire new_AGEMA_signal_9266 ;
    wire new_AGEMA_signal_9267 ;
    wire new_AGEMA_signal_9268 ;
    wire new_AGEMA_signal_9269 ;
    wire new_AGEMA_signal_9270 ;
    wire new_AGEMA_signal_9271 ;
    wire new_AGEMA_signal_9272 ;
    wire new_AGEMA_signal_9273 ;
    wire new_AGEMA_signal_9274 ;
    wire new_AGEMA_signal_9275 ;
    wire new_AGEMA_signal_9276 ;
    wire new_AGEMA_signal_9277 ;
    wire new_AGEMA_signal_9278 ;
    wire new_AGEMA_signal_9279 ;
    wire new_AGEMA_signal_9280 ;
    wire new_AGEMA_signal_9281 ;
    wire new_AGEMA_signal_9282 ;
    wire new_AGEMA_signal_9283 ;
    wire new_AGEMA_signal_9284 ;
    wire new_AGEMA_signal_9285 ;
    wire new_AGEMA_signal_9286 ;
    wire new_AGEMA_signal_9287 ;
    wire new_AGEMA_signal_9288 ;
    wire new_AGEMA_signal_9289 ;
    wire new_AGEMA_signal_9290 ;
    wire new_AGEMA_signal_9291 ;
    wire new_AGEMA_signal_9292 ;
    wire new_AGEMA_signal_9293 ;
    wire new_AGEMA_signal_9294 ;
    wire new_AGEMA_signal_9295 ;
    wire new_AGEMA_signal_9296 ;
    wire new_AGEMA_signal_9297 ;
    wire new_AGEMA_signal_9298 ;
    wire new_AGEMA_signal_9299 ;
    wire new_AGEMA_signal_9300 ;
    wire new_AGEMA_signal_9301 ;
    wire new_AGEMA_signal_9302 ;
    wire new_AGEMA_signal_9304 ;
    wire new_AGEMA_signal_9305 ;
    wire new_AGEMA_signal_9306 ;
    wire new_AGEMA_signal_9307 ;
    wire new_AGEMA_signal_9308 ;
    wire new_AGEMA_signal_9309 ;
    wire new_AGEMA_signal_9310 ;
    wire new_AGEMA_signal_9311 ;
    wire new_AGEMA_signal_9312 ;
    wire new_AGEMA_signal_9313 ;
    wire new_AGEMA_signal_9314 ;
    wire new_AGEMA_signal_9315 ;
    wire new_AGEMA_signal_9316 ;
    wire new_AGEMA_signal_9317 ;
    wire new_AGEMA_signal_9318 ;
    wire new_AGEMA_signal_9319 ;
    wire new_AGEMA_signal_9320 ;
    wire new_AGEMA_signal_9321 ;
    wire new_AGEMA_signal_9322 ;
    wire new_AGEMA_signal_9323 ;
    wire new_AGEMA_signal_9324 ;
    wire new_AGEMA_signal_9325 ;
    wire new_AGEMA_signal_9326 ;
    wire new_AGEMA_signal_9327 ;
    wire new_AGEMA_signal_9328 ;
    wire new_AGEMA_signal_9329 ;
    wire new_AGEMA_signal_9330 ;
    wire new_AGEMA_signal_9331 ;
    wire new_AGEMA_signal_9332 ;
    wire new_AGEMA_signal_9333 ;
    wire new_AGEMA_signal_9334 ;
    wire new_AGEMA_signal_9335 ;
    wire new_AGEMA_signal_9336 ;
    wire new_AGEMA_signal_9337 ;
    wire new_AGEMA_signal_9338 ;
    wire new_AGEMA_signal_9339 ;
    wire new_AGEMA_signal_9340 ;
    wire new_AGEMA_signal_9341 ;
    wire new_AGEMA_signal_9342 ;
    wire new_AGEMA_signal_9343 ;
    wire new_AGEMA_signal_9344 ;
    wire new_AGEMA_signal_9345 ;
    wire new_AGEMA_signal_9346 ;
    wire new_AGEMA_signal_9347 ;
    wire new_AGEMA_signal_9348 ;
    wire new_AGEMA_signal_9349 ;
    wire new_AGEMA_signal_9350 ;
    wire new_AGEMA_signal_9351 ;
    wire new_AGEMA_signal_9352 ;
    wire new_AGEMA_signal_9353 ;
    wire new_AGEMA_signal_9354 ;
    wire new_AGEMA_signal_9355 ;
    wire new_AGEMA_signal_9356 ;
    wire new_AGEMA_signal_9357 ;
    wire new_AGEMA_signal_9358 ;
    wire new_AGEMA_signal_9359 ;
    wire new_AGEMA_signal_9360 ;
    wire new_AGEMA_signal_9361 ;
    wire new_AGEMA_signal_9362 ;
    wire new_AGEMA_signal_9363 ;
    wire new_AGEMA_signal_9364 ;
    wire new_AGEMA_signal_9365 ;
    wire new_AGEMA_signal_9366 ;
    wire new_AGEMA_signal_9367 ;
    wire new_AGEMA_signal_9368 ;
    wire new_AGEMA_signal_9369 ;
    wire new_AGEMA_signal_9370 ;
    wire new_AGEMA_signal_9371 ;
    wire new_AGEMA_signal_9372 ;
    wire new_AGEMA_signal_9373 ;
    wire new_AGEMA_signal_9374 ;
    wire new_AGEMA_signal_9375 ;
    wire new_AGEMA_signal_9376 ;
    wire new_AGEMA_signal_9377 ;
    wire new_AGEMA_signal_9378 ;
    wire new_AGEMA_signal_9379 ;
    wire new_AGEMA_signal_9380 ;
    wire new_AGEMA_signal_9381 ;
    wire new_AGEMA_signal_9382 ;
    wire new_AGEMA_signal_9383 ;
    wire new_AGEMA_signal_9384 ;
    wire new_AGEMA_signal_9385 ;
    wire new_AGEMA_signal_9386 ;
    wire new_AGEMA_signal_9387 ;
    wire new_AGEMA_signal_9388 ;
    wire new_AGEMA_signal_9389 ;
    wire new_AGEMA_signal_9390 ;
    wire new_AGEMA_signal_9391 ;
    wire new_AGEMA_signal_9392 ;
    wire new_AGEMA_signal_9393 ;
    wire new_AGEMA_signal_9394 ;
    wire new_AGEMA_signal_9395 ;
    wire new_AGEMA_signal_9396 ;
    wire new_AGEMA_signal_9397 ;
    wire new_AGEMA_signal_9398 ;
    wire new_AGEMA_signal_9399 ;
    wire new_AGEMA_signal_9400 ;
    wire new_AGEMA_signal_9401 ;
    wire new_AGEMA_signal_9402 ;
    wire new_AGEMA_signal_9403 ;
    wire new_AGEMA_signal_9404 ;
    wire new_AGEMA_signal_9405 ;
    wire new_AGEMA_signal_9406 ;
    wire new_AGEMA_signal_9407 ;
    wire new_AGEMA_signal_9408 ;
    wire new_AGEMA_signal_9409 ;
    wire new_AGEMA_signal_9410 ;
    wire new_AGEMA_signal_9411 ;
    wire new_AGEMA_signal_9412 ;
    wire new_AGEMA_signal_9413 ;
    wire new_AGEMA_signal_9414 ;
    wire new_AGEMA_signal_9415 ;
    wire new_AGEMA_signal_9416 ;
    wire new_AGEMA_signal_9417 ;
    wire new_AGEMA_signal_9418 ;
    wire new_AGEMA_signal_9419 ;
    wire new_AGEMA_signal_9420 ;
    wire new_AGEMA_signal_9421 ;
    wire new_AGEMA_signal_9422 ;
    wire new_AGEMA_signal_9423 ;
    wire new_AGEMA_signal_9424 ;
    wire new_AGEMA_signal_9425 ;
    wire new_AGEMA_signal_9426 ;
    wire new_AGEMA_signal_9427 ;
    wire new_AGEMA_signal_9428 ;
    wire new_AGEMA_signal_9429 ;
    wire new_AGEMA_signal_9430 ;
    wire new_AGEMA_signal_9431 ;
    wire new_AGEMA_signal_9432 ;
    wire new_AGEMA_signal_9433 ;
    wire new_AGEMA_signal_9434 ;
    wire new_AGEMA_signal_9435 ;
    wire new_AGEMA_signal_9436 ;
    wire new_AGEMA_signal_9437 ;
    wire new_AGEMA_signal_9438 ;
    wire new_AGEMA_signal_9439 ;
    wire new_AGEMA_signal_9440 ;
    wire new_AGEMA_signal_9441 ;
    wire new_AGEMA_signal_9442 ;
    wire new_AGEMA_signal_9443 ;
    wire new_AGEMA_signal_9444 ;
    wire new_AGEMA_signal_9445 ;
    wire new_AGEMA_signal_9446 ;
    wire new_AGEMA_signal_9447 ;
    wire new_AGEMA_signal_9448 ;
    wire new_AGEMA_signal_9449 ;
    wire new_AGEMA_signal_9450 ;
    wire new_AGEMA_signal_9451 ;
    wire new_AGEMA_signal_9452 ;
    wire new_AGEMA_signal_9453 ;
    wire new_AGEMA_signal_9454 ;
    wire new_AGEMA_signal_9455 ;
    wire new_AGEMA_signal_9456 ;
    wire new_AGEMA_signal_9457 ;
    wire new_AGEMA_signal_9458 ;
    wire new_AGEMA_signal_9459 ;
    wire new_AGEMA_signal_9460 ;
    wire new_AGEMA_signal_9461 ;
    wire new_AGEMA_signal_9462 ;
    wire new_AGEMA_signal_9463 ;
    wire new_AGEMA_signal_9464 ;
    wire new_AGEMA_signal_9465 ;
    wire new_AGEMA_signal_9466 ;
    wire new_AGEMA_signal_9467 ;
    wire new_AGEMA_signal_9468 ;
    wire new_AGEMA_signal_9469 ;
    wire new_AGEMA_signal_9470 ;
    wire new_AGEMA_signal_9471 ;
    wire new_AGEMA_signal_9472 ;
    wire new_AGEMA_signal_9473 ;
    wire new_AGEMA_signal_9474 ;
    wire new_AGEMA_signal_9475 ;
    wire new_AGEMA_signal_9476 ;
    wire new_AGEMA_signal_9477 ;
    wire new_AGEMA_signal_9478 ;
    wire new_AGEMA_signal_9479 ;
    wire new_AGEMA_signal_9480 ;
    wire new_AGEMA_signal_9481 ;
    wire new_AGEMA_signal_9482 ;
    wire new_AGEMA_signal_9483 ;
    wire new_AGEMA_signal_9484 ;
    wire new_AGEMA_signal_9485 ;
    wire new_AGEMA_signal_9486 ;
    wire new_AGEMA_signal_9487 ;
    wire new_AGEMA_signal_9488 ;
    wire new_AGEMA_signal_9489 ;
    wire new_AGEMA_signal_9490 ;
    wire new_AGEMA_signal_9491 ;
    wire new_AGEMA_signal_9492 ;
    wire new_AGEMA_signal_9493 ;
    wire new_AGEMA_signal_9494 ;
    wire new_AGEMA_signal_9495 ;
    wire new_AGEMA_signal_9496 ;
    wire new_AGEMA_signal_9497 ;
    wire new_AGEMA_signal_9498 ;
    wire new_AGEMA_signal_9499 ;
    wire new_AGEMA_signal_9500 ;
    wire new_AGEMA_signal_9501 ;
    wire new_AGEMA_signal_9502 ;
    wire new_AGEMA_signal_9503 ;
    wire new_AGEMA_signal_9504 ;
    wire new_AGEMA_signal_9505 ;
    wire new_AGEMA_signal_9506 ;
    wire new_AGEMA_signal_9507 ;
    wire new_AGEMA_signal_9508 ;
    wire new_AGEMA_signal_9509 ;
    wire new_AGEMA_signal_9510 ;
    wire new_AGEMA_signal_9511 ;
    wire new_AGEMA_signal_9512 ;
    wire new_AGEMA_signal_9513 ;
    wire new_AGEMA_signal_9514 ;
    wire new_AGEMA_signal_9515 ;
    wire new_AGEMA_signal_9516 ;
    wire new_AGEMA_signal_9517 ;
    wire new_AGEMA_signal_9518 ;
    wire new_AGEMA_signal_9519 ;
    wire new_AGEMA_signal_9520 ;
    wire new_AGEMA_signal_9521 ;
    wire new_AGEMA_signal_9522 ;
    wire new_AGEMA_signal_9523 ;
    wire new_AGEMA_signal_9524 ;
    wire new_AGEMA_signal_9525 ;
    wire new_AGEMA_signal_9526 ;
    wire new_AGEMA_signal_9527 ;
    wire new_AGEMA_signal_9528 ;
    wire new_AGEMA_signal_9529 ;
    wire new_AGEMA_signal_9530 ;
    wire new_AGEMA_signal_9531 ;
    wire new_AGEMA_signal_9532 ;
    wire new_AGEMA_signal_9533 ;
    wire new_AGEMA_signal_9534 ;
    wire new_AGEMA_signal_9535 ;
    wire new_AGEMA_signal_9536 ;
    wire new_AGEMA_signal_9537 ;
    wire new_AGEMA_signal_9538 ;
    wire new_AGEMA_signal_9539 ;
    wire new_AGEMA_signal_9540 ;
    wire new_AGEMA_signal_9541 ;
    wire new_AGEMA_signal_9542 ;
    wire new_AGEMA_signal_9543 ;
    wire new_AGEMA_signal_9544 ;
    wire new_AGEMA_signal_9545 ;
    wire new_AGEMA_signal_9546 ;
    wire new_AGEMA_signal_9547 ;
    wire new_AGEMA_signal_9548 ;
    wire new_AGEMA_signal_9549 ;
    wire new_AGEMA_signal_9550 ;
    wire new_AGEMA_signal_9551 ;
    wire new_AGEMA_signal_9552 ;
    wire new_AGEMA_signal_9553 ;
    wire new_AGEMA_signal_9554 ;
    wire new_AGEMA_signal_9555 ;
    wire new_AGEMA_signal_9556 ;
    wire new_AGEMA_signal_9557 ;
    wire new_AGEMA_signal_9558 ;
    wire new_AGEMA_signal_9559 ;
    wire new_AGEMA_signal_9560 ;
    wire new_AGEMA_signal_9561 ;
    wire new_AGEMA_signal_9562 ;
    wire new_AGEMA_signal_9563 ;
    wire new_AGEMA_signal_9564 ;
    wire new_AGEMA_signal_9565 ;
    wire new_AGEMA_signal_9566 ;
    wire new_AGEMA_signal_9567 ;
    wire new_AGEMA_signal_9568 ;
    wire new_AGEMA_signal_9569 ;
    wire new_AGEMA_signal_9570 ;
    wire new_AGEMA_signal_9571 ;
    wire new_AGEMA_signal_9572 ;
    wire new_AGEMA_signal_9573 ;
    wire new_AGEMA_signal_9574 ;
    wire new_AGEMA_signal_9575 ;
    wire new_AGEMA_signal_9576 ;
    wire new_AGEMA_signal_9577 ;
    wire new_AGEMA_signal_9578 ;
    wire new_AGEMA_signal_9579 ;
    wire new_AGEMA_signal_9580 ;
    wire new_AGEMA_signal_9581 ;
    wire new_AGEMA_signal_9582 ;
    wire new_AGEMA_signal_9583 ;
    wire new_AGEMA_signal_9584 ;
    wire new_AGEMA_signal_9585 ;
    wire new_AGEMA_signal_9586 ;
    wire new_AGEMA_signal_9587 ;
    wire new_AGEMA_signal_9588 ;
    wire new_AGEMA_signal_9589 ;
    wire new_AGEMA_signal_9590 ;
    wire new_AGEMA_signal_9591 ;
    wire new_AGEMA_signal_9592 ;
    wire new_AGEMA_signal_9593 ;
    wire new_AGEMA_signal_9594 ;
    wire new_AGEMA_signal_9595 ;
    wire new_AGEMA_signal_9596 ;
    wire new_AGEMA_signal_9597 ;
    wire new_AGEMA_signal_9598 ;
    wire new_AGEMA_signal_9599 ;
    wire new_AGEMA_signal_9600 ;
    wire new_AGEMA_signal_9601 ;
    wire new_AGEMA_signal_9602 ;
    wire new_AGEMA_signal_9603 ;
    wire new_AGEMA_signal_9604 ;
    wire new_AGEMA_signal_9605 ;
    wire new_AGEMA_signal_9606 ;
    wire new_AGEMA_signal_9607 ;
    wire new_AGEMA_signal_9608 ;
    wire new_AGEMA_signal_9609 ;
    wire new_AGEMA_signal_9610 ;
    wire new_AGEMA_signal_9611 ;
    wire new_AGEMA_signal_9612 ;
    wire new_AGEMA_signal_9613 ;
    wire new_AGEMA_signal_9614 ;
    wire new_AGEMA_signal_9615 ;
    wire new_AGEMA_signal_9616 ;
    wire new_AGEMA_signal_9617 ;
    wire new_AGEMA_signal_9618 ;
    wire new_AGEMA_signal_9619 ;
    wire new_AGEMA_signal_9620 ;
    wire new_AGEMA_signal_9621 ;
    wire new_AGEMA_signal_9622 ;
    wire new_AGEMA_signal_9623 ;
    wire new_AGEMA_signal_9624 ;
    wire new_AGEMA_signal_9625 ;
    wire new_AGEMA_signal_9626 ;
    wire new_AGEMA_signal_9627 ;
    wire new_AGEMA_signal_9628 ;
    wire new_AGEMA_signal_9629 ;
    wire new_AGEMA_signal_9630 ;
    wire new_AGEMA_signal_9631 ;
    wire new_AGEMA_signal_9632 ;
    wire new_AGEMA_signal_9633 ;
    wire new_AGEMA_signal_9634 ;
    wire new_AGEMA_signal_9635 ;
    wire new_AGEMA_signal_9636 ;
    wire new_AGEMA_signal_9637 ;
    wire new_AGEMA_signal_9638 ;
    wire new_AGEMA_signal_9639 ;
    wire new_AGEMA_signal_9640 ;
    wire new_AGEMA_signal_9641 ;
    wire new_AGEMA_signal_9642 ;
    wire new_AGEMA_signal_9643 ;
    wire new_AGEMA_signal_9644 ;
    wire new_AGEMA_signal_9645 ;
    wire new_AGEMA_signal_9646 ;
    wire new_AGEMA_signal_9647 ;
    wire new_AGEMA_signal_9648 ;
    wire new_AGEMA_signal_9649 ;
    wire new_AGEMA_signal_9650 ;
    wire new_AGEMA_signal_9651 ;
    wire new_AGEMA_signal_9652 ;
    wire new_AGEMA_signal_9653 ;
    wire new_AGEMA_signal_9654 ;
    wire new_AGEMA_signal_9655 ;
    wire new_AGEMA_signal_9656 ;
    wire new_AGEMA_signal_9657 ;
    wire new_AGEMA_signal_9658 ;
    wire new_AGEMA_signal_9659 ;
    wire new_AGEMA_signal_9660 ;
    wire new_AGEMA_signal_9661 ;
    wire new_AGEMA_signal_9662 ;
    wire new_AGEMA_signal_9663 ;
    wire new_AGEMA_signal_9664 ;
    wire new_AGEMA_signal_9665 ;
    wire new_AGEMA_signal_9666 ;
    wire new_AGEMA_signal_9667 ;
    wire new_AGEMA_signal_9668 ;
    wire new_AGEMA_signal_9669 ;
    wire new_AGEMA_signal_9670 ;
    wire new_AGEMA_signal_9671 ;
    wire new_AGEMA_signal_9672 ;
    wire new_AGEMA_signal_9673 ;
    wire new_AGEMA_signal_9674 ;
    wire new_AGEMA_signal_9675 ;
    wire new_AGEMA_signal_9676 ;
    wire new_AGEMA_signal_9677 ;
    wire new_AGEMA_signal_9678 ;
    wire new_AGEMA_signal_9679 ;
    wire new_AGEMA_signal_9680 ;
    wire new_AGEMA_signal_9681 ;
    wire new_AGEMA_signal_9682 ;
    wire new_AGEMA_signal_9683 ;
    wire new_AGEMA_signal_9684 ;
    wire new_AGEMA_signal_9685 ;
    wire new_AGEMA_signal_9686 ;
    wire new_AGEMA_signal_9687 ;
    wire new_AGEMA_signal_9688 ;
    wire new_AGEMA_signal_9689 ;
    wire new_AGEMA_signal_9690 ;
    wire new_AGEMA_signal_9691 ;
    wire new_AGEMA_signal_9692 ;
    wire new_AGEMA_signal_9693 ;
    wire new_AGEMA_signal_9694 ;
    wire new_AGEMA_signal_9695 ;
    wire new_AGEMA_signal_9696 ;
    wire new_AGEMA_signal_9697 ;
    wire new_AGEMA_signal_9698 ;
    wire new_AGEMA_signal_9699 ;
    wire new_AGEMA_signal_9700 ;
    wire new_AGEMA_signal_9701 ;
    wire new_AGEMA_signal_9702 ;
    wire new_AGEMA_signal_9703 ;
    wire new_AGEMA_signal_9704 ;
    wire new_AGEMA_signal_9705 ;
    wire new_AGEMA_signal_9706 ;
    wire new_AGEMA_signal_9707 ;
    wire new_AGEMA_signal_9708 ;
    wire new_AGEMA_signal_9709 ;
    wire new_AGEMA_signal_9710 ;
    wire new_AGEMA_signal_9711 ;
    wire new_AGEMA_signal_9712 ;
    wire new_AGEMA_signal_9713 ;
    wire new_AGEMA_signal_9714 ;
    wire new_AGEMA_signal_9715 ;
    wire new_AGEMA_signal_9716 ;
    wire new_AGEMA_signal_9717 ;
    wire new_AGEMA_signal_9718 ;
    wire new_AGEMA_signal_9719 ;
    wire new_AGEMA_signal_9720 ;
    wire new_AGEMA_signal_9721 ;
    wire new_AGEMA_signal_9722 ;
    wire new_AGEMA_signal_9723 ;
    wire new_AGEMA_signal_9724 ;
    wire new_AGEMA_signal_9725 ;
    wire new_AGEMA_signal_9726 ;
    wire new_AGEMA_signal_9727 ;
    wire new_AGEMA_signal_9728 ;
    wire new_AGEMA_signal_9729 ;
    wire new_AGEMA_signal_9730 ;
    wire new_AGEMA_signal_9731 ;
    wire new_AGEMA_signal_9732 ;
    wire new_AGEMA_signal_9733 ;
    wire new_AGEMA_signal_9734 ;
    wire new_AGEMA_signal_9735 ;
    wire new_AGEMA_signal_9736 ;
    wire new_AGEMA_signal_9737 ;
    wire new_AGEMA_signal_9738 ;
    wire new_AGEMA_signal_9739 ;
    wire new_AGEMA_signal_9740 ;
    wire new_AGEMA_signal_9741 ;
    wire new_AGEMA_signal_9742 ;
    wire new_AGEMA_signal_9743 ;
    wire new_AGEMA_signal_9744 ;
    wire new_AGEMA_signal_9745 ;
    wire new_AGEMA_signal_9746 ;
    wire new_AGEMA_signal_9747 ;
    wire new_AGEMA_signal_9748 ;
    wire new_AGEMA_signal_9749 ;
    wire new_AGEMA_signal_9750 ;
    wire new_AGEMA_signal_9751 ;
    wire new_AGEMA_signal_9752 ;
    wire new_AGEMA_signal_9753 ;
    wire new_AGEMA_signal_9754 ;
    wire new_AGEMA_signal_9755 ;
    wire new_AGEMA_signal_9756 ;
    wire new_AGEMA_signal_9757 ;
    wire new_AGEMA_signal_9758 ;
    wire new_AGEMA_signal_9759 ;
    wire new_AGEMA_signal_9760 ;
    wire new_AGEMA_signal_9761 ;
    wire new_AGEMA_signal_9762 ;
    wire new_AGEMA_signal_9763 ;
    wire new_AGEMA_signal_9764 ;
    wire new_AGEMA_signal_9765 ;
    wire new_AGEMA_signal_9766 ;
    wire new_AGEMA_signal_9767 ;
    wire new_AGEMA_signal_9768 ;
    wire new_AGEMA_signal_9769 ;
    wire new_AGEMA_signal_9770 ;
    wire new_AGEMA_signal_9771 ;
    wire new_AGEMA_signal_9772 ;
    wire new_AGEMA_signal_9773 ;
    wire new_AGEMA_signal_9774 ;
    wire new_AGEMA_signal_9775 ;
    wire new_AGEMA_signal_9776 ;
    wire new_AGEMA_signal_9777 ;
    wire new_AGEMA_signal_9778 ;
    wire new_AGEMA_signal_9779 ;
    wire new_AGEMA_signal_9780 ;
    wire new_AGEMA_signal_9781 ;
    wire new_AGEMA_signal_9782 ;
    wire new_AGEMA_signal_9783 ;
    wire new_AGEMA_signal_9784 ;
    wire new_AGEMA_signal_9785 ;
    wire new_AGEMA_signal_9786 ;
    wire new_AGEMA_signal_9787 ;
    wire new_AGEMA_signal_9788 ;
    wire new_AGEMA_signal_9789 ;
    wire new_AGEMA_signal_9790 ;
    wire new_AGEMA_signal_9791 ;
    wire new_AGEMA_signal_9792 ;
    wire new_AGEMA_signal_9793 ;
    wire new_AGEMA_signal_9794 ;
    wire new_AGEMA_signal_9795 ;
    wire new_AGEMA_signal_9796 ;
    wire new_AGEMA_signal_9797 ;
    wire new_AGEMA_signal_9798 ;
    wire new_AGEMA_signal_9799 ;
    wire new_AGEMA_signal_9800 ;
    wire new_AGEMA_signal_9801 ;
    wire new_AGEMA_signal_9802 ;
    wire new_AGEMA_signal_9803 ;
    wire new_AGEMA_signal_9804 ;
    wire new_AGEMA_signal_9805 ;
    wire new_AGEMA_signal_9806 ;
    wire new_AGEMA_signal_9807 ;
    wire new_AGEMA_signal_9808 ;
    wire new_AGEMA_signal_9809 ;
    wire new_AGEMA_signal_9810 ;
    wire new_AGEMA_signal_9811 ;
    wire new_AGEMA_signal_9812 ;
    wire new_AGEMA_signal_9813 ;
    wire new_AGEMA_signal_9814 ;
    wire new_AGEMA_signal_9815 ;
    wire new_AGEMA_signal_9816 ;
    wire new_AGEMA_signal_9817 ;
    wire new_AGEMA_signal_9818 ;
    wire new_AGEMA_signal_9819 ;
    wire new_AGEMA_signal_9820 ;
    wire new_AGEMA_signal_9821 ;
    wire new_AGEMA_signal_9822 ;
    wire new_AGEMA_signal_9823 ;
    wire new_AGEMA_signal_9824 ;
    wire new_AGEMA_signal_9825 ;
    wire new_AGEMA_signal_9826 ;
    wire new_AGEMA_signal_9827 ;
    wire new_AGEMA_signal_9828 ;
    wire new_AGEMA_signal_9829 ;
    wire new_AGEMA_signal_9830 ;
    wire new_AGEMA_signal_9831 ;
    wire new_AGEMA_signal_9832 ;
    wire new_AGEMA_signal_9833 ;
    wire new_AGEMA_signal_9834 ;
    wire new_AGEMA_signal_9835 ;
    wire new_AGEMA_signal_9836 ;
    wire new_AGEMA_signal_9837 ;
    wire new_AGEMA_signal_9838 ;
    wire new_AGEMA_signal_9839 ;
    wire new_AGEMA_signal_9840 ;
    wire new_AGEMA_signal_9841 ;
    wire new_AGEMA_signal_9842 ;
    wire new_AGEMA_signal_9843 ;
    wire new_AGEMA_signal_9844 ;
    wire new_AGEMA_signal_9845 ;
    wire new_AGEMA_signal_9846 ;
    wire new_AGEMA_signal_9847 ;
    wire new_AGEMA_signal_9848 ;
    wire new_AGEMA_signal_9849 ;
    wire new_AGEMA_signal_9850 ;
    wire new_AGEMA_signal_9851 ;
    wire new_AGEMA_signal_9852 ;
    wire new_AGEMA_signal_9853 ;
    wire new_AGEMA_signal_9854 ;
    wire new_AGEMA_signal_9855 ;
    wire new_AGEMA_signal_9856 ;
    wire new_AGEMA_signal_9857 ;
    wire new_AGEMA_signal_9858 ;
    wire new_AGEMA_signal_9859 ;
    wire new_AGEMA_signal_9860 ;
    wire new_AGEMA_signal_9861 ;
    wire new_AGEMA_signal_9862 ;
    wire new_AGEMA_signal_9863 ;
    wire new_AGEMA_signal_9864 ;
    wire new_AGEMA_signal_9865 ;
    wire new_AGEMA_signal_9866 ;
    wire new_AGEMA_signal_9867 ;
    wire new_AGEMA_signal_9868 ;
    wire new_AGEMA_signal_9869 ;
    wire new_AGEMA_signal_9870 ;
    wire new_AGEMA_signal_9871 ;
    wire new_AGEMA_signal_9872 ;
    wire new_AGEMA_signal_9873 ;
    wire new_AGEMA_signal_9874 ;
    wire new_AGEMA_signal_9875 ;
    wire new_AGEMA_signal_9876 ;
    wire new_AGEMA_signal_9877 ;
    wire new_AGEMA_signal_9878 ;
    wire new_AGEMA_signal_9879 ;
    wire new_AGEMA_signal_9880 ;
    wire new_AGEMA_signal_9881 ;
    wire new_AGEMA_signal_9882 ;
    wire new_AGEMA_signal_9883 ;
    wire new_AGEMA_signal_9884 ;
    wire new_AGEMA_signal_9885 ;
    wire new_AGEMA_signal_9886 ;
    wire new_AGEMA_signal_9887 ;
    wire new_AGEMA_signal_9888 ;
    wire new_AGEMA_signal_9889 ;
    wire new_AGEMA_signal_9890 ;
    wire new_AGEMA_signal_9891 ;
    wire new_AGEMA_signal_9892 ;
    wire new_AGEMA_signal_9893 ;
    wire new_AGEMA_signal_9894 ;
    wire new_AGEMA_signal_9895 ;
    wire new_AGEMA_signal_9896 ;
    wire new_AGEMA_signal_9897 ;
    wire new_AGEMA_signal_9898 ;
    wire new_AGEMA_signal_9899 ;
    wire new_AGEMA_signal_9900 ;
    wire new_AGEMA_signal_9901 ;
    wire new_AGEMA_signal_9902 ;
    wire new_AGEMA_signal_9903 ;
    wire new_AGEMA_signal_9904 ;
    wire new_AGEMA_signal_9905 ;
    wire new_AGEMA_signal_9906 ;
    wire new_AGEMA_signal_9907 ;
    wire new_AGEMA_signal_9908 ;
    wire new_AGEMA_signal_9909 ;
    wire new_AGEMA_signal_9910 ;
    wire new_AGEMA_signal_9911 ;
    wire new_AGEMA_signal_9912 ;
    wire new_AGEMA_signal_9913 ;
    wire new_AGEMA_signal_9914 ;
    wire new_AGEMA_signal_9915 ;
    wire new_AGEMA_signal_9916 ;
    wire new_AGEMA_signal_9917 ;
    wire new_AGEMA_signal_9918 ;
    wire new_AGEMA_signal_9919 ;
    wire new_AGEMA_signal_9920 ;
    wire new_AGEMA_signal_9921 ;
    wire new_AGEMA_signal_9922 ;
    wire new_AGEMA_signal_9923 ;
    wire new_AGEMA_signal_9924 ;
    wire new_AGEMA_signal_9925 ;
    wire new_AGEMA_signal_9926 ;
    wire new_AGEMA_signal_9927 ;
    wire new_AGEMA_signal_9928 ;
    wire new_AGEMA_signal_9929 ;
    wire new_AGEMA_signal_9930 ;
    wire new_AGEMA_signal_9931 ;
    wire new_AGEMA_signal_9932 ;
    wire new_AGEMA_signal_9933 ;
    wire new_AGEMA_signal_9934 ;
    wire new_AGEMA_signal_9935 ;
    wire new_AGEMA_signal_9936 ;
    wire new_AGEMA_signal_9937 ;
    wire new_AGEMA_signal_9938 ;
    wire new_AGEMA_signal_9939 ;
    wire new_AGEMA_signal_9940 ;
    wire new_AGEMA_signal_9941 ;
    wire new_AGEMA_signal_9942 ;
    wire new_AGEMA_signal_9943 ;
    wire new_AGEMA_signal_9944 ;
    wire new_AGEMA_signal_9945 ;
    wire new_AGEMA_signal_9946 ;
    wire new_AGEMA_signal_9947 ;
    wire new_AGEMA_signal_9948 ;
    wire new_AGEMA_signal_9949 ;
    wire new_AGEMA_signal_9950 ;
    wire new_AGEMA_signal_9951 ;
    wire new_AGEMA_signal_9952 ;
    wire new_AGEMA_signal_9953 ;
    wire new_AGEMA_signal_9954 ;
    wire new_AGEMA_signal_9955 ;
    wire new_AGEMA_signal_9956 ;
    wire new_AGEMA_signal_9957 ;
    wire new_AGEMA_signal_9958 ;
    wire new_AGEMA_signal_9959 ;
    wire new_AGEMA_signal_9960 ;
    wire new_AGEMA_signal_9961 ;
    wire new_AGEMA_signal_9962 ;
    wire new_AGEMA_signal_9963 ;
    wire new_AGEMA_signal_9964 ;
    wire new_AGEMA_signal_9965 ;
    wire new_AGEMA_signal_9966 ;
    wire new_AGEMA_signal_9967 ;
    wire new_AGEMA_signal_9968 ;
    wire new_AGEMA_signal_9969 ;
    wire new_AGEMA_signal_9970 ;
    wire new_AGEMA_signal_9971 ;
    wire new_AGEMA_signal_9972 ;
    wire new_AGEMA_signal_9973 ;
    wire new_AGEMA_signal_9974 ;
    wire new_AGEMA_signal_9975 ;
    wire new_AGEMA_signal_9976 ;
    wire new_AGEMA_signal_9977 ;
    wire new_AGEMA_signal_9978 ;
    wire new_AGEMA_signal_9979 ;
    wire new_AGEMA_signal_9980 ;
    wire new_AGEMA_signal_9981 ;
    wire new_AGEMA_signal_9982 ;
    wire new_AGEMA_signal_9983 ;
    wire new_AGEMA_signal_9984 ;
    wire new_AGEMA_signal_9985 ;
    wire new_AGEMA_signal_9986 ;
    wire new_AGEMA_signal_9987 ;
    wire new_AGEMA_signal_9988 ;
    wire new_AGEMA_signal_9989 ;
    wire new_AGEMA_signal_9990 ;
    wire new_AGEMA_signal_9991 ;
    wire new_AGEMA_signal_9992 ;
    wire new_AGEMA_signal_9993 ;
    wire new_AGEMA_signal_9994 ;
    wire new_AGEMA_signal_9995 ;
    wire new_AGEMA_signal_9996 ;
    wire new_AGEMA_signal_9997 ;
    wire new_AGEMA_signal_9998 ;
    wire new_AGEMA_signal_9999 ;
    wire new_AGEMA_signal_10000 ;
    wire new_AGEMA_signal_10001 ;
    wire new_AGEMA_signal_10002 ;
    wire new_AGEMA_signal_10003 ;
    wire new_AGEMA_signal_10004 ;
    wire new_AGEMA_signal_10005 ;
    wire new_AGEMA_signal_10006 ;
    wire new_AGEMA_signal_10007 ;
    wire new_AGEMA_signal_10008 ;
    wire new_AGEMA_signal_10009 ;
    wire new_AGEMA_signal_10010 ;
    wire new_AGEMA_signal_10011 ;
    wire new_AGEMA_signal_10012 ;
    wire new_AGEMA_signal_10013 ;
    wire new_AGEMA_signal_10014 ;
    wire new_AGEMA_signal_10015 ;
    wire new_AGEMA_signal_10016 ;
    wire new_AGEMA_signal_10017 ;
    wire new_AGEMA_signal_10018 ;
    wire new_AGEMA_signal_10019 ;
    wire new_AGEMA_signal_10020 ;
    wire new_AGEMA_signal_10021 ;
    wire new_AGEMA_signal_10022 ;
    wire new_AGEMA_signal_10023 ;
    wire new_AGEMA_signal_10024 ;
    wire new_AGEMA_signal_10025 ;
    wire new_AGEMA_signal_10026 ;
    wire new_AGEMA_signal_10027 ;
    wire new_AGEMA_signal_10028 ;
    wire new_AGEMA_signal_10029 ;
    wire new_AGEMA_signal_10030 ;
    wire new_AGEMA_signal_10031 ;
    wire new_AGEMA_signal_10032 ;
    wire new_AGEMA_signal_10033 ;
    wire new_AGEMA_signal_10034 ;
    wire new_AGEMA_signal_10035 ;
    wire new_AGEMA_signal_10036 ;
    wire new_AGEMA_signal_10037 ;
    wire new_AGEMA_signal_10038 ;
    wire new_AGEMA_signal_10039 ;
    wire new_AGEMA_signal_10040 ;
    wire new_AGEMA_signal_10041 ;
    wire new_AGEMA_signal_10042 ;
    wire new_AGEMA_signal_10043 ;
    wire new_AGEMA_signal_10044 ;
    wire new_AGEMA_signal_10045 ;
    wire new_AGEMA_signal_10046 ;
    wire new_AGEMA_signal_10047 ;
    wire new_AGEMA_signal_10048 ;
    wire new_AGEMA_signal_10049 ;
    wire new_AGEMA_signal_10050 ;
    wire new_AGEMA_signal_10051 ;
    wire new_AGEMA_signal_10052 ;
    wire new_AGEMA_signal_10053 ;
    wire new_AGEMA_signal_10054 ;
    wire new_AGEMA_signal_10055 ;
    wire new_AGEMA_signal_10056 ;
    wire new_AGEMA_signal_10057 ;
    wire new_AGEMA_signal_10058 ;
    wire new_AGEMA_signal_10059 ;
    wire new_AGEMA_signal_10060 ;
    wire new_AGEMA_signal_10061 ;
    wire new_AGEMA_signal_10062 ;
    wire new_AGEMA_signal_10063 ;
    wire new_AGEMA_signal_10064 ;
    wire new_AGEMA_signal_10065 ;
    wire new_AGEMA_signal_10066 ;
    wire new_AGEMA_signal_10067 ;
    wire new_AGEMA_signal_10068 ;
    wire new_AGEMA_signal_10069 ;
    wire new_AGEMA_signal_10070 ;
    wire new_AGEMA_signal_10071 ;
    wire new_AGEMA_signal_10072 ;
    wire new_AGEMA_signal_10073 ;
    wire new_AGEMA_signal_10074 ;
    wire new_AGEMA_signal_10075 ;
    wire new_AGEMA_signal_10076 ;
    wire new_AGEMA_signal_10077 ;
    wire new_AGEMA_signal_10078 ;
    wire new_AGEMA_signal_10079 ;
    wire new_AGEMA_signal_10080 ;
    wire new_AGEMA_signal_10081 ;
    wire new_AGEMA_signal_10082 ;
    wire new_AGEMA_signal_10083 ;
    wire new_AGEMA_signal_10084 ;
    wire new_AGEMA_signal_10085 ;
    wire new_AGEMA_signal_10086 ;
    wire new_AGEMA_signal_10087 ;
    wire new_AGEMA_signal_10088 ;
    wire new_AGEMA_signal_10089 ;
    wire new_AGEMA_signal_10090 ;
    wire new_AGEMA_signal_10091 ;
    wire new_AGEMA_signal_10092 ;
    wire new_AGEMA_signal_10093 ;
    wire new_AGEMA_signal_10094 ;
    wire new_AGEMA_signal_10095 ;
    wire new_AGEMA_signal_10096 ;
    wire new_AGEMA_signal_10097 ;
    wire new_AGEMA_signal_10098 ;
    wire new_AGEMA_signal_10099 ;
    wire new_AGEMA_signal_10100 ;
    wire new_AGEMA_signal_10101 ;
    wire new_AGEMA_signal_10102 ;
    wire new_AGEMA_signal_10103 ;
    wire new_AGEMA_signal_10104 ;
    wire new_AGEMA_signal_10105 ;
    wire new_AGEMA_signal_10106 ;
    wire new_AGEMA_signal_10107 ;
    wire new_AGEMA_signal_10108 ;
    wire new_AGEMA_signal_10109 ;
    wire new_AGEMA_signal_10110 ;
    wire new_AGEMA_signal_10111 ;
    wire new_AGEMA_signal_10112 ;
    wire new_AGEMA_signal_10113 ;
    wire new_AGEMA_signal_10114 ;
    wire new_AGEMA_signal_10115 ;
    wire new_AGEMA_signal_10116 ;
    wire new_AGEMA_signal_10117 ;
    wire new_AGEMA_signal_10118 ;
    wire new_AGEMA_signal_10119 ;
    wire new_AGEMA_signal_10120 ;
    wire new_AGEMA_signal_10121 ;
    wire new_AGEMA_signal_10122 ;
    wire new_AGEMA_signal_10123 ;
    wire new_AGEMA_signal_10124 ;
    wire new_AGEMA_signal_10125 ;
    wire new_AGEMA_signal_10126 ;
    wire new_AGEMA_signal_10127 ;
    wire new_AGEMA_signal_10128 ;
    wire new_AGEMA_signal_10129 ;
    wire new_AGEMA_signal_10130 ;
    wire new_AGEMA_signal_10131 ;
    wire new_AGEMA_signal_10132 ;
    wire new_AGEMA_signal_10133 ;
    wire new_AGEMA_signal_10134 ;
    wire new_AGEMA_signal_10135 ;
    wire new_AGEMA_signal_10136 ;
    wire new_AGEMA_signal_10137 ;
    wire new_AGEMA_signal_10138 ;
    wire new_AGEMA_signal_10139 ;
    wire new_AGEMA_signal_10140 ;
    wire new_AGEMA_signal_10141 ;
    wire new_AGEMA_signal_10142 ;
    wire new_AGEMA_signal_10143 ;
    wire new_AGEMA_signal_10144 ;
    wire new_AGEMA_signal_10145 ;
    wire new_AGEMA_signal_10146 ;
    wire new_AGEMA_signal_10147 ;
    wire new_AGEMA_signal_10148 ;
    wire new_AGEMA_signal_10149 ;
    wire new_AGEMA_signal_10150 ;
    wire new_AGEMA_signal_10151 ;
    wire new_AGEMA_signal_10152 ;
    wire new_AGEMA_signal_10153 ;
    wire new_AGEMA_signal_10154 ;
    wire new_AGEMA_signal_10155 ;
    wire new_AGEMA_signal_10156 ;
    wire new_AGEMA_signal_10157 ;
    wire new_AGEMA_signal_10158 ;
    wire new_AGEMA_signal_10159 ;
    wire new_AGEMA_signal_10160 ;
    wire new_AGEMA_signal_10161 ;
    wire new_AGEMA_signal_10162 ;
    wire new_AGEMA_signal_10163 ;
    wire new_AGEMA_signal_10164 ;
    wire new_AGEMA_signal_10165 ;
    wire new_AGEMA_signal_10166 ;
    wire new_AGEMA_signal_10167 ;
    wire new_AGEMA_signal_10168 ;
    wire new_AGEMA_signal_10169 ;
    wire new_AGEMA_signal_10170 ;
    wire new_AGEMA_signal_10171 ;
    wire new_AGEMA_signal_10172 ;
    wire new_AGEMA_signal_10173 ;
    wire new_AGEMA_signal_10174 ;
    wire new_AGEMA_signal_10175 ;
    wire new_AGEMA_signal_10176 ;
    wire new_AGEMA_signal_10177 ;
    wire new_AGEMA_signal_10178 ;
    wire new_AGEMA_signal_10179 ;
    wire new_AGEMA_signal_10180 ;
    wire new_AGEMA_signal_10181 ;
    wire new_AGEMA_signal_10182 ;
    wire new_AGEMA_signal_10183 ;
    wire new_AGEMA_signal_10184 ;
    wire new_AGEMA_signal_10185 ;
    wire new_AGEMA_signal_10186 ;
    wire new_AGEMA_signal_10187 ;
    wire new_AGEMA_signal_10188 ;
    wire new_AGEMA_signal_10189 ;
    wire new_AGEMA_signal_10190 ;
    wire new_AGEMA_signal_10191 ;
    wire new_AGEMA_signal_10192 ;
    wire new_AGEMA_signal_10193 ;
    wire new_AGEMA_signal_10194 ;
    wire new_AGEMA_signal_10195 ;
    wire new_AGEMA_signal_10196 ;
    wire new_AGEMA_signal_10197 ;
    wire new_AGEMA_signal_10198 ;
    wire new_AGEMA_signal_10199 ;
    wire new_AGEMA_signal_10200 ;
    wire new_AGEMA_signal_10201 ;
    wire new_AGEMA_signal_10202 ;
    wire new_AGEMA_signal_10203 ;
    wire new_AGEMA_signal_10204 ;
    wire new_AGEMA_signal_10205 ;
    wire new_AGEMA_signal_10206 ;
    wire new_AGEMA_signal_10207 ;
    wire new_AGEMA_signal_10208 ;
    wire new_AGEMA_signal_10209 ;
    wire new_AGEMA_signal_10210 ;
    wire new_AGEMA_signal_10211 ;
    wire new_AGEMA_signal_10215 ;
    wire new_AGEMA_signal_10216 ;
    wire new_AGEMA_signal_10217 ;
    wire new_AGEMA_signal_10221 ;
    wire new_AGEMA_signal_10222 ;
    wire new_AGEMA_signal_10223 ;
    wire new_AGEMA_signal_10227 ;
    wire new_AGEMA_signal_10228 ;
    wire new_AGEMA_signal_10229 ;
    wire new_AGEMA_signal_10233 ;
    wire new_AGEMA_signal_10234 ;
    wire new_AGEMA_signal_10235 ;
    wire new_AGEMA_signal_10239 ;
    wire new_AGEMA_signal_10240 ;
    wire new_AGEMA_signal_10241 ;
    wire new_AGEMA_signal_10245 ;
    wire new_AGEMA_signal_10246 ;
    wire new_AGEMA_signal_10247 ;
    wire new_AGEMA_signal_10251 ;
    wire new_AGEMA_signal_10252 ;
    wire new_AGEMA_signal_10253 ;
    wire new_AGEMA_signal_10257 ;
    wire new_AGEMA_signal_10258 ;
    wire new_AGEMA_signal_10259 ;
    wire new_AGEMA_signal_10260 ;
    wire new_AGEMA_signal_10261 ;
    wire new_AGEMA_signal_10262 ;
    wire new_AGEMA_signal_10263 ;
    wire new_AGEMA_signal_10264 ;
    wire new_AGEMA_signal_10265 ;
    wire new_AGEMA_signal_10266 ;
    wire new_AGEMA_signal_10267 ;
    wire new_AGEMA_signal_10268 ;
    wire new_AGEMA_signal_10269 ;
    wire new_AGEMA_signal_10270 ;
    wire new_AGEMA_signal_10271 ;
    wire new_AGEMA_signal_10272 ;
    wire new_AGEMA_signal_10273 ;
    wire new_AGEMA_signal_10274 ;
    wire new_AGEMA_signal_10275 ;
    wire new_AGEMA_signal_10276 ;
    wire new_AGEMA_signal_10277 ;
    wire new_AGEMA_signal_10278 ;
    wire new_AGEMA_signal_10279 ;
    wire new_AGEMA_signal_10280 ;
    wire new_AGEMA_signal_10281 ;
    wire new_AGEMA_signal_10282 ;
    wire new_AGEMA_signal_10283 ;
    wire new_AGEMA_signal_10284 ;
    wire new_AGEMA_signal_10285 ;
    wire new_AGEMA_signal_10286 ;
    wire new_AGEMA_signal_10287 ;
    wire new_AGEMA_signal_10288 ;
    wire new_AGEMA_signal_10289 ;
    wire new_AGEMA_signal_10290 ;
    wire new_AGEMA_signal_10291 ;
    wire new_AGEMA_signal_10292 ;
    wire new_AGEMA_signal_10293 ;
    wire new_AGEMA_signal_10294 ;
    wire new_AGEMA_signal_10295 ;
    wire new_AGEMA_signal_10296 ;
    wire new_AGEMA_signal_10297 ;
    wire new_AGEMA_signal_10298 ;
    wire new_AGEMA_signal_10299 ;
    wire new_AGEMA_signal_10300 ;
    wire new_AGEMA_signal_10301 ;
    wire new_AGEMA_signal_10302 ;
    wire new_AGEMA_signal_10303 ;
    wire new_AGEMA_signal_10304 ;
    wire new_AGEMA_signal_10305 ;
    wire new_AGEMA_signal_10306 ;
    wire new_AGEMA_signal_10307 ;
    wire new_AGEMA_signal_10308 ;
    wire new_AGEMA_signal_10309 ;
    wire new_AGEMA_signal_10310 ;
    wire new_AGEMA_signal_10311 ;
    wire new_AGEMA_signal_10312 ;
    wire new_AGEMA_signal_10313 ;
    wire new_AGEMA_signal_10314 ;
    wire new_AGEMA_signal_10315 ;
    wire new_AGEMA_signal_10316 ;
    wire new_AGEMA_signal_10317 ;
    wire new_AGEMA_signal_10318 ;
    wire new_AGEMA_signal_10319 ;
    wire new_AGEMA_signal_10320 ;
    wire new_AGEMA_signal_10321 ;
    wire new_AGEMA_signal_10322 ;
    wire new_AGEMA_signal_10323 ;
    wire new_AGEMA_signal_10324 ;
    wire new_AGEMA_signal_10325 ;
    wire new_AGEMA_signal_10326 ;
    wire new_AGEMA_signal_10327 ;
    wire new_AGEMA_signal_10328 ;
    wire new_AGEMA_signal_10329 ;
    wire new_AGEMA_signal_10330 ;
    wire new_AGEMA_signal_10331 ;
    wire new_AGEMA_signal_10332 ;
    wire new_AGEMA_signal_10333 ;
    wire new_AGEMA_signal_10334 ;
    wire new_AGEMA_signal_10335 ;
    wire new_AGEMA_signal_10336 ;
    wire new_AGEMA_signal_10337 ;
    wire new_AGEMA_signal_10338 ;
    wire new_AGEMA_signal_10339 ;
    wire new_AGEMA_signal_10340 ;
    wire new_AGEMA_signal_10341 ;
    wire new_AGEMA_signal_10342 ;
    wire new_AGEMA_signal_10343 ;
    wire new_AGEMA_signal_10344 ;
    wire new_AGEMA_signal_10345 ;
    wire new_AGEMA_signal_10346 ;
    wire new_AGEMA_signal_10347 ;
    wire new_AGEMA_signal_10348 ;
    wire new_AGEMA_signal_10349 ;
    wire new_AGEMA_signal_10350 ;
    wire new_AGEMA_signal_10351 ;
    wire new_AGEMA_signal_10352 ;
    wire new_AGEMA_signal_10353 ;
    wire new_AGEMA_signal_10354 ;
    wire new_AGEMA_signal_10355 ;
    wire new_AGEMA_signal_10356 ;
    wire new_AGEMA_signal_10357 ;
    wire new_AGEMA_signal_10358 ;
    wire new_AGEMA_signal_10359 ;
    wire new_AGEMA_signal_10360 ;
    wire new_AGEMA_signal_10361 ;
    wire new_AGEMA_signal_10362 ;
    wire new_AGEMA_signal_10363 ;
    wire new_AGEMA_signal_10364 ;
    wire new_AGEMA_signal_10365 ;
    wire new_AGEMA_signal_10366 ;
    wire new_AGEMA_signal_10367 ;
    wire new_AGEMA_signal_10368 ;
    wire new_AGEMA_signal_10369 ;
    wire new_AGEMA_signal_10370 ;
    wire new_AGEMA_signal_10371 ;
    wire new_AGEMA_signal_10372 ;
    wire new_AGEMA_signal_10373 ;
    wire new_AGEMA_signal_10374 ;
    wire new_AGEMA_signal_10375 ;
    wire new_AGEMA_signal_10376 ;
    wire new_AGEMA_signal_10377 ;
    wire new_AGEMA_signal_10378 ;
    wire new_AGEMA_signal_10379 ;
    wire new_AGEMA_signal_10380 ;
    wire new_AGEMA_signal_10381 ;
    wire new_AGEMA_signal_10382 ;
    wire new_AGEMA_signal_10383 ;
    wire new_AGEMA_signal_10384 ;
    wire new_AGEMA_signal_10385 ;
    wire new_AGEMA_signal_10386 ;
    wire new_AGEMA_signal_10387 ;
    wire new_AGEMA_signal_10388 ;
    wire new_AGEMA_signal_10389 ;
    wire new_AGEMA_signal_10390 ;
    wire new_AGEMA_signal_10391 ;
    wire new_AGEMA_signal_10392 ;
    wire new_AGEMA_signal_10393 ;
    wire new_AGEMA_signal_10394 ;
    wire new_AGEMA_signal_10395 ;
    wire new_AGEMA_signal_10396 ;
    wire new_AGEMA_signal_10397 ;
    wire new_AGEMA_signal_10398 ;
    wire new_AGEMA_signal_10399 ;
    wire new_AGEMA_signal_10400 ;
    wire new_AGEMA_signal_10401 ;
    wire new_AGEMA_signal_10402 ;
    wire new_AGEMA_signal_10403 ;
    wire new_AGEMA_signal_10404 ;
    wire new_AGEMA_signal_10405 ;
    wire new_AGEMA_signal_10406 ;
    wire new_AGEMA_signal_10407 ;
    wire new_AGEMA_signal_10408 ;
    wire new_AGEMA_signal_10409 ;
    wire new_AGEMA_signal_10410 ;
    wire new_AGEMA_signal_10411 ;
    wire new_AGEMA_signal_10412 ;
    wire new_AGEMA_signal_10413 ;
    wire new_AGEMA_signal_10414 ;
    wire new_AGEMA_signal_10415 ;
    wire new_AGEMA_signal_10416 ;
    wire new_AGEMA_signal_10417 ;
    wire new_AGEMA_signal_10418 ;
    wire new_AGEMA_signal_10419 ;
    wire new_AGEMA_signal_10420 ;
    wire new_AGEMA_signal_10421 ;
    wire new_AGEMA_signal_10422 ;
    wire new_AGEMA_signal_10423 ;
    wire new_AGEMA_signal_10424 ;
    wire new_AGEMA_signal_10425 ;
    wire new_AGEMA_signal_10426 ;
    wire new_AGEMA_signal_10427 ;
    wire new_AGEMA_signal_10428 ;
    wire new_AGEMA_signal_10429 ;
    wire new_AGEMA_signal_10430 ;
    wire new_AGEMA_signal_10431 ;
    wire new_AGEMA_signal_10432 ;
    wire new_AGEMA_signal_10433 ;
    wire new_AGEMA_signal_10434 ;
    wire new_AGEMA_signal_10435 ;
    wire new_AGEMA_signal_10436 ;
    wire new_AGEMA_signal_10437 ;
    wire new_AGEMA_signal_10438 ;
    wire new_AGEMA_signal_10439 ;
    wire new_AGEMA_signal_10440 ;
    wire new_AGEMA_signal_10441 ;
    wire new_AGEMA_signal_10442 ;
    wire new_AGEMA_signal_10443 ;
    wire new_AGEMA_signal_10444 ;
    wire new_AGEMA_signal_10445 ;
    wire new_AGEMA_signal_10446 ;
    wire new_AGEMA_signal_10447 ;
    wire new_AGEMA_signal_10448 ;
    wire new_AGEMA_signal_10449 ;
    wire new_AGEMA_signal_10450 ;
    wire new_AGEMA_signal_10451 ;
    wire new_AGEMA_signal_10452 ;
    wire new_AGEMA_signal_10453 ;
    wire new_AGEMA_signal_10454 ;
    wire new_AGEMA_signal_10455 ;
    wire new_AGEMA_signal_10456 ;
    wire new_AGEMA_signal_10457 ;
    wire new_AGEMA_signal_10458 ;
    wire new_AGEMA_signal_10459 ;
    wire new_AGEMA_signal_10460 ;
    wire new_AGEMA_signal_10461 ;
    wire new_AGEMA_signal_10462 ;
    wire new_AGEMA_signal_10463 ;
    wire new_AGEMA_signal_10464 ;
    wire new_AGEMA_signal_10465 ;
    wire new_AGEMA_signal_10466 ;
    wire new_AGEMA_signal_10467 ;
    wire new_AGEMA_signal_10468 ;
    wire new_AGEMA_signal_10469 ;
    wire new_AGEMA_signal_10470 ;
    wire new_AGEMA_signal_10471 ;
    wire new_AGEMA_signal_10472 ;
    wire new_AGEMA_signal_10473 ;
    wire new_AGEMA_signal_10474 ;
    wire new_AGEMA_signal_10475 ;
    wire new_AGEMA_signal_10476 ;
    wire new_AGEMA_signal_10477 ;
    wire new_AGEMA_signal_10478 ;
    wire new_AGEMA_signal_10479 ;
    wire new_AGEMA_signal_10480 ;
    wire new_AGEMA_signal_10481 ;
    wire new_AGEMA_signal_10482 ;
    wire new_AGEMA_signal_10483 ;
    wire new_AGEMA_signal_10484 ;
    wire new_AGEMA_signal_10485 ;
    wire new_AGEMA_signal_10486 ;
    wire new_AGEMA_signal_10487 ;
    wire new_AGEMA_signal_10488 ;
    wire new_AGEMA_signal_10489 ;
    wire new_AGEMA_signal_10490 ;
    wire new_AGEMA_signal_10491 ;
    wire new_AGEMA_signal_10492 ;
    wire new_AGEMA_signal_10493 ;
    wire new_AGEMA_signal_10494 ;
    wire new_AGEMA_signal_10495 ;
    wire new_AGEMA_signal_10496 ;
    wire new_AGEMA_signal_10497 ;
    wire new_AGEMA_signal_10498 ;
    wire new_AGEMA_signal_10499 ;
    wire new_AGEMA_signal_10500 ;
    wire new_AGEMA_signal_10501 ;
    wire new_AGEMA_signal_10502 ;
    wire new_AGEMA_signal_10503 ;
    wire new_AGEMA_signal_10504 ;
    wire new_AGEMA_signal_10505 ;
    wire new_AGEMA_signal_10506 ;
    wire new_AGEMA_signal_10507 ;
    wire new_AGEMA_signal_10508 ;
    wire new_AGEMA_signal_10509 ;
    wire new_AGEMA_signal_10510 ;
    wire new_AGEMA_signal_10511 ;
    wire new_AGEMA_signal_10512 ;
    wire new_AGEMA_signal_10513 ;
    wire new_AGEMA_signal_10514 ;
    wire new_AGEMA_signal_10515 ;
    wire new_AGEMA_signal_10516 ;
    wire new_AGEMA_signal_10517 ;
    wire new_AGEMA_signal_10518 ;
    wire new_AGEMA_signal_10519 ;
    wire new_AGEMA_signal_10520 ;
    wire new_AGEMA_signal_10521 ;
    wire new_AGEMA_signal_10522 ;
    wire new_AGEMA_signal_10523 ;
    wire new_AGEMA_signal_10524 ;
    wire new_AGEMA_signal_10525 ;
    wire new_AGEMA_signal_10526 ;
    wire new_AGEMA_signal_10527 ;
    wire new_AGEMA_signal_10528 ;
    wire new_AGEMA_signal_10529 ;
    wire new_AGEMA_signal_10530 ;
    wire new_AGEMA_signal_10531 ;
    wire new_AGEMA_signal_10532 ;
    wire new_AGEMA_signal_10533 ;
    wire new_AGEMA_signal_10534 ;
    wire new_AGEMA_signal_10535 ;
    wire new_AGEMA_signal_10536 ;
    wire new_AGEMA_signal_10537 ;
    wire new_AGEMA_signal_10538 ;
    wire new_AGEMA_signal_10539 ;
    wire new_AGEMA_signal_10540 ;
    wire new_AGEMA_signal_10541 ;
    wire new_AGEMA_signal_10542 ;
    wire new_AGEMA_signal_10543 ;
    wire new_AGEMA_signal_10544 ;
    wire new_AGEMA_signal_10545 ;
    wire new_AGEMA_signal_10546 ;
    wire new_AGEMA_signal_10547 ;
    wire new_AGEMA_signal_10548 ;
    wire new_AGEMA_signal_10549 ;
    wire new_AGEMA_signal_10553 ;
    wire new_AGEMA_signal_10554 ;
    wire new_AGEMA_signal_10555 ;
    wire new_AGEMA_signal_10559 ;
    wire new_AGEMA_signal_10560 ;
    wire new_AGEMA_signal_10561 ;
    wire new_AGEMA_signal_10565 ;
    wire new_AGEMA_signal_10566 ;
    wire new_AGEMA_signal_10567 ;
    wire new_AGEMA_signal_10571 ;
    wire new_AGEMA_signal_10572 ;
    wire new_AGEMA_signal_10573 ;
    wire new_AGEMA_signal_10577 ;
    wire new_AGEMA_signal_10578 ;
    wire new_AGEMA_signal_10579 ;
    wire new_AGEMA_signal_10580 ;
    wire new_AGEMA_signal_10581 ;
    wire new_AGEMA_signal_10582 ;
    wire new_AGEMA_signal_10583 ;
    wire new_AGEMA_signal_10584 ;
    wire new_AGEMA_signal_10585 ;
    wire new_AGEMA_signal_10586 ;
    wire new_AGEMA_signal_10587 ;
    wire new_AGEMA_signal_10588 ;
    wire new_AGEMA_signal_10592 ;
    wire new_AGEMA_signal_10593 ;
    wire new_AGEMA_signal_10594 ;
    wire new_AGEMA_signal_10598 ;
    wire new_AGEMA_signal_10599 ;
    wire new_AGEMA_signal_10600 ;
    wire new_AGEMA_signal_10604 ;
    wire new_AGEMA_signal_10605 ;
    wire new_AGEMA_signal_10606 ;
    wire new_AGEMA_signal_10610 ;
    wire new_AGEMA_signal_10611 ;
    wire new_AGEMA_signal_10612 ;
    wire new_AGEMA_signal_10616 ;
    wire new_AGEMA_signal_10617 ;
    wire new_AGEMA_signal_10618 ;
    wire new_AGEMA_signal_10619 ;
    wire new_AGEMA_signal_10620 ;
    wire new_AGEMA_signal_10621 ;
    wire new_AGEMA_signal_10622 ;
    wire new_AGEMA_signal_10623 ;
    wire new_AGEMA_signal_10624 ;
    wire new_AGEMA_signal_10625 ;
    wire new_AGEMA_signal_10626 ;
    wire new_AGEMA_signal_10627 ;
    wire new_AGEMA_signal_10631 ;
    wire new_AGEMA_signal_10632 ;
    wire new_AGEMA_signal_10633 ;
    wire new_AGEMA_signal_10637 ;
    wire new_AGEMA_signal_10638 ;
    wire new_AGEMA_signal_10639 ;
    wire new_AGEMA_signal_10643 ;
    wire new_AGEMA_signal_10644 ;
    wire new_AGEMA_signal_10645 ;
    wire new_AGEMA_signal_10649 ;
    wire new_AGEMA_signal_10650 ;
    wire new_AGEMA_signal_10651 ;
    wire new_AGEMA_signal_10655 ;
    wire new_AGEMA_signal_10656 ;
    wire new_AGEMA_signal_10657 ;
    wire new_AGEMA_signal_10658 ;
    wire new_AGEMA_signal_10659 ;
    wire new_AGEMA_signal_10660 ;
    wire new_AGEMA_signal_10661 ;
    wire new_AGEMA_signal_10662 ;
    wire new_AGEMA_signal_10663 ;
    wire new_AGEMA_signal_10664 ;
    wire new_AGEMA_signal_10665 ;
    wire new_AGEMA_signal_10666 ;
    wire new_AGEMA_signal_10667 ;
    wire new_AGEMA_signal_10668 ;
    wire new_AGEMA_signal_10669 ;
    wire new_AGEMA_signal_10670 ;
    wire new_AGEMA_signal_10671 ;
    wire new_AGEMA_signal_10672 ;
    wire new_AGEMA_signal_10673 ;
    wire new_AGEMA_signal_10674 ;
    wire new_AGEMA_signal_10675 ;
    wire new_AGEMA_signal_10676 ;
    wire new_AGEMA_signal_10677 ;
    wire new_AGEMA_signal_10678 ;
    wire new_AGEMA_signal_10679 ;
    wire new_AGEMA_signal_10680 ;
    wire new_AGEMA_signal_10681 ;
    wire new_AGEMA_signal_10682 ;
    wire new_AGEMA_signal_10683 ;
    wire new_AGEMA_signal_10684 ;
    wire new_AGEMA_signal_10685 ;
    wire new_AGEMA_signal_10686 ;
    wire new_AGEMA_signal_10687 ;
    wire new_AGEMA_signal_10688 ;
    wire new_AGEMA_signal_10689 ;
    wire new_AGEMA_signal_10690 ;
    wire new_AGEMA_signal_10691 ;
    wire new_AGEMA_signal_10692 ;
    wire new_AGEMA_signal_10693 ;
    wire new_AGEMA_signal_10694 ;
    wire new_AGEMA_signal_10695 ;
    wire new_AGEMA_signal_10696 ;
    wire new_AGEMA_signal_10700 ;
    wire new_AGEMA_signal_10701 ;
    wire new_AGEMA_signal_10702 ;
    wire new_AGEMA_signal_10703 ;
    wire new_AGEMA_signal_10704 ;
    wire new_AGEMA_signal_10705 ;
    wire new_AGEMA_signal_10709 ;
    wire new_AGEMA_signal_10710 ;
    wire new_AGEMA_signal_10711 ;
    wire new_AGEMA_signal_10715 ;
    wire new_AGEMA_signal_10716 ;
    wire new_AGEMA_signal_10717 ;
    wire new_AGEMA_signal_10718 ;
    wire new_AGEMA_signal_10719 ;
    wire new_AGEMA_signal_10720 ;
    wire new_AGEMA_signal_10721 ;
    wire new_AGEMA_signal_10722 ;
    wire new_AGEMA_signal_10723 ;
    wire new_AGEMA_signal_10724 ;
    wire new_AGEMA_signal_10725 ;
    wire new_AGEMA_signal_10726 ;
    wire new_AGEMA_signal_10727 ;
    wire new_AGEMA_signal_10728 ;
    wire new_AGEMA_signal_10729 ;
    wire new_AGEMA_signal_10733 ;
    wire new_AGEMA_signal_10734 ;
    wire new_AGEMA_signal_10735 ;
    wire new_AGEMA_signal_10736 ;
    wire new_AGEMA_signal_10737 ;
    wire new_AGEMA_signal_10738 ;
    wire new_AGEMA_signal_10742 ;
    wire new_AGEMA_signal_10743 ;
    wire new_AGEMA_signal_10744 ;
    wire new_AGEMA_signal_10748 ;
    wire new_AGEMA_signal_10749 ;
    wire new_AGEMA_signal_10750 ;
    wire new_AGEMA_signal_10751 ;
    wire new_AGEMA_signal_10752 ;
    wire new_AGEMA_signal_10753 ;
    wire new_AGEMA_signal_10754 ;
    wire new_AGEMA_signal_10755 ;
    wire new_AGEMA_signal_10756 ;
    wire new_AGEMA_signal_10757 ;
    wire new_AGEMA_signal_10758 ;
    wire new_AGEMA_signal_10759 ;
    wire new_AGEMA_signal_10760 ;
    wire new_AGEMA_signal_10761 ;
    wire new_AGEMA_signal_10762 ;
    wire new_AGEMA_signal_10766 ;
    wire new_AGEMA_signal_10767 ;
    wire new_AGEMA_signal_10768 ;
    wire new_AGEMA_signal_10769 ;
    wire new_AGEMA_signal_10770 ;
    wire new_AGEMA_signal_10771 ;
    wire new_AGEMA_signal_10775 ;
    wire new_AGEMA_signal_10776 ;
    wire new_AGEMA_signal_10777 ;
    wire new_AGEMA_signal_10781 ;
    wire new_AGEMA_signal_10782 ;
    wire new_AGEMA_signal_10783 ;
    wire new_AGEMA_signal_10784 ;
    wire new_AGEMA_signal_10785 ;
    wire new_AGEMA_signal_10786 ;
    wire new_AGEMA_signal_10787 ;
    wire new_AGEMA_signal_10788 ;
    wire new_AGEMA_signal_10789 ;
    wire new_AGEMA_signal_10790 ;
    wire new_AGEMA_signal_10791 ;
    wire new_AGEMA_signal_10792 ;
    wire new_AGEMA_signal_10793 ;
    wire new_AGEMA_signal_10794 ;
    wire new_AGEMA_signal_10795 ;
    wire new_AGEMA_signal_10796 ;
    wire new_AGEMA_signal_10797 ;
    wire new_AGEMA_signal_10798 ;
    wire new_AGEMA_signal_10799 ;
    wire new_AGEMA_signal_10800 ;
    wire new_AGEMA_signal_10801 ;
    wire new_AGEMA_signal_10802 ;
    wire new_AGEMA_signal_10803 ;
    wire new_AGEMA_signal_10804 ;
    wire new_AGEMA_signal_10805 ;
    wire new_AGEMA_signal_10806 ;
    wire new_AGEMA_signal_10807 ;
    wire new_AGEMA_signal_10808 ;
    wire new_AGEMA_signal_10809 ;
    wire new_AGEMA_signal_10810 ;
    wire new_AGEMA_signal_10811 ;
    wire new_AGEMA_signal_10812 ;
    wire new_AGEMA_signal_10813 ;
    wire new_AGEMA_signal_10814 ;
    wire new_AGEMA_signal_10815 ;
    wire new_AGEMA_signal_10816 ;
    wire new_AGEMA_signal_10817 ;
    wire new_AGEMA_signal_10818 ;
    wire new_AGEMA_signal_10819 ;
    wire new_AGEMA_signal_10820 ;
    wire new_AGEMA_signal_10821 ;
    wire new_AGEMA_signal_10822 ;
    wire new_AGEMA_signal_10823 ;
    wire new_AGEMA_signal_10824 ;
    wire new_AGEMA_signal_10825 ;
    wire new_AGEMA_signal_10826 ;
    wire new_AGEMA_signal_10827 ;
    wire new_AGEMA_signal_10828 ;
    wire new_AGEMA_signal_10829 ;
    wire new_AGEMA_signal_10830 ;
    wire new_AGEMA_signal_10831 ;
    wire new_AGEMA_signal_10832 ;
    wire new_AGEMA_signal_10833 ;
    wire new_AGEMA_signal_10834 ;
    wire new_AGEMA_signal_10835 ;
    wire new_AGEMA_signal_10836 ;
    wire new_AGEMA_signal_10837 ;
    wire new_AGEMA_signal_10838 ;
    wire new_AGEMA_signal_10839 ;
    wire new_AGEMA_signal_10840 ;
    wire new_AGEMA_signal_10841 ;
    wire new_AGEMA_signal_10842 ;
    wire new_AGEMA_signal_10843 ;
    wire new_AGEMA_signal_10844 ;
    wire new_AGEMA_signal_10845 ;
    wire new_AGEMA_signal_10846 ;
    wire new_AGEMA_signal_10847 ;
    wire new_AGEMA_signal_10848 ;
    wire new_AGEMA_signal_10849 ;
    wire new_AGEMA_signal_10850 ;
    wire new_AGEMA_signal_10851 ;
    wire new_AGEMA_signal_10852 ;
    wire new_AGEMA_signal_10853 ;
    wire new_AGEMA_signal_10854 ;
    wire new_AGEMA_signal_10855 ;
    wire new_AGEMA_signal_10856 ;
    wire new_AGEMA_signal_10857 ;
    wire new_AGEMA_signal_10858 ;
    wire new_AGEMA_signal_10859 ;
    wire new_AGEMA_signal_10860 ;
    wire new_AGEMA_signal_10861 ;
    wire new_AGEMA_signal_10862 ;
    wire new_AGEMA_signal_10863 ;
    wire new_AGEMA_signal_10864 ;
    wire new_AGEMA_signal_10865 ;
    wire new_AGEMA_signal_10866 ;
    wire new_AGEMA_signal_10867 ;
    wire new_AGEMA_signal_10868 ;
    wire new_AGEMA_signal_10869 ;
    wire new_AGEMA_signal_10870 ;
    wire new_AGEMA_signal_10871 ;
    wire new_AGEMA_signal_10872 ;
    wire new_AGEMA_signal_10873 ;
    wire new_AGEMA_signal_10874 ;
    wire new_AGEMA_signal_10875 ;
    wire new_AGEMA_signal_10876 ;
    wire new_AGEMA_signal_10877 ;
    wire new_AGEMA_signal_10878 ;
    wire new_AGEMA_signal_10879 ;
    wire new_AGEMA_signal_10880 ;
    wire new_AGEMA_signal_10881 ;
    wire new_AGEMA_signal_10882 ;
    wire new_AGEMA_signal_10883 ;
    wire new_AGEMA_signal_10884 ;
    wire new_AGEMA_signal_10885 ;
    wire new_AGEMA_signal_10886 ;
    wire new_AGEMA_signal_10887 ;
    wire new_AGEMA_signal_10888 ;
    wire new_AGEMA_signal_10889 ;
    wire new_AGEMA_signal_10890 ;
    wire new_AGEMA_signal_10891 ;
    wire new_AGEMA_signal_10892 ;
    wire new_AGEMA_signal_10893 ;
    wire new_AGEMA_signal_10894 ;
    wire new_AGEMA_signal_10895 ;
    wire new_AGEMA_signal_10896 ;
    wire new_AGEMA_signal_10897 ;
    wire new_AGEMA_signal_10898 ;
    wire new_AGEMA_signal_10899 ;
    wire new_AGEMA_signal_10900 ;
    wire new_AGEMA_signal_10901 ;
    wire new_AGEMA_signal_10902 ;
    wire new_AGEMA_signal_10903 ;
    wire new_AGEMA_signal_10904 ;
    wire new_AGEMA_signal_10905 ;
    wire new_AGEMA_signal_10906 ;
    wire new_AGEMA_signal_10907 ;
    wire new_AGEMA_signal_10908 ;
    wire new_AGEMA_signal_10909 ;
    wire new_AGEMA_signal_10910 ;
    wire new_AGEMA_signal_10911 ;
    wire new_AGEMA_signal_10912 ;
    wire new_AGEMA_signal_10913 ;
    wire new_AGEMA_signal_10914 ;
    wire new_AGEMA_signal_10915 ;
    wire new_AGEMA_signal_10916 ;
    wire new_AGEMA_signal_10917 ;
    wire new_AGEMA_signal_10918 ;
    wire new_AGEMA_signal_10919 ;
    wire new_AGEMA_signal_10920 ;
    wire new_AGEMA_signal_10921 ;
    wire new_AGEMA_signal_10922 ;
    wire new_AGEMA_signal_10923 ;
    wire new_AGEMA_signal_10924 ;
    wire new_AGEMA_signal_10925 ;
    wire new_AGEMA_signal_10926 ;
    wire new_AGEMA_signal_10927 ;
    wire new_AGEMA_signal_10928 ;
    wire new_AGEMA_signal_10929 ;
    wire new_AGEMA_signal_10930 ;
    wire new_AGEMA_signal_10931 ;
    wire new_AGEMA_signal_10932 ;
    wire new_AGEMA_signal_10933 ;
    wire new_AGEMA_signal_10934 ;
    wire new_AGEMA_signal_10935 ;
    wire new_AGEMA_signal_10936 ;
    wire new_AGEMA_signal_10937 ;
    wire new_AGEMA_signal_10938 ;
    wire new_AGEMA_signal_10939 ;
    wire new_AGEMA_signal_10940 ;
    wire new_AGEMA_signal_10941 ;
    wire new_AGEMA_signal_10942 ;
    wire new_AGEMA_signal_10943 ;
    wire new_AGEMA_signal_10944 ;
    wire new_AGEMA_signal_10945 ;
    wire new_AGEMA_signal_10946 ;
    wire new_AGEMA_signal_10947 ;
    wire new_AGEMA_signal_10948 ;
    wire new_AGEMA_signal_10949 ;
    wire new_AGEMA_signal_10950 ;
    wire new_AGEMA_signal_10951 ;
    wire new_AGEMA_signal_10952 ;
    wire new_AGEMA_signal_10953 ;
    wire new_AGEMA_signal_10954 ;
    wire new_AGEMA_signal_10955 ;
    wire new_AGEMA_signal_10956 ;
    wire new_AGEMA_signal_10957 ;
    wire new_AGEMA_signal_10958 ;
    wire new_AGEMA_signal_10959 ;
    wire new_AGEMA_signal_10960 ;
    wire new_AGEMA_signal_10961 ;
    wire new_AGEMA_signal_10962 ;
    wire new_AGEMA_signal_10963 ;
    wire new_AGEMA_signal_10964 ;
    wire new_AGEMA_signal_10965 ;
    wire new_AGEMA_signal_10966 ;
    wire new_AGEMA_signal_10967 ;
    wire new_AGEMA_signal_10968 ;
    wire new_AGEMA_signal_10969 ;
    wire new_AGEMA_signal_10970 ;
    wire new_AGEMA_signal_10971 ;
    wire new_AGEMA_signal_10972 ;
    wire new_AGEMA_signal_10973 ;
    wire new_AGEMA_signal_10974 ;
    wire new_AGEMA_signal_10975 ;
    wire new_AGEMA_signal_10976 ;
    wire new_AGEMA_signal_10977 ;
    wire new_AGEMA_signal_10978 ;
    wire new_AGEMA_signal_10979 ;
    wire new_AGEMA_signal_10980 ;
    wire new_AGEMA_signal_10981 ;
    wire new_AGEMA_signal_10982 ;
    wire new_AGEMA_signal_10983 ;
    wire new_AGEMA_signal_10984 ;
    wire new_AGEMA_signal_10985 ;
    wire new_AGEMA_signal_10986 ;
    wire new_AGEMA_signal_10987 ;
    wire new_AGEMA_signal_10988 ;
    wire new_AGEMA_signal_10989 ;
    wire new_AGEMA_signal_10990 ;
    wire new_AGEMA_signal_10991 ;
    wire new_AGEMA_signal_10992 ;
    wire new_AGEMA_signal_10993 ;
    wire new_AGEMA_signal_10994 ;
    wire new_AGEMA_signal_10995 ;
    wire new_AGEMA_signal_10996 ;
    wire new_AGEMA_signal_10997 ;
    wire new_AGEMA_signal_10998 ;
    wire new_AGEMA_signal_10999 ;
    wire new_AGEMA_signal_11000 ;
    wire new_AGEMA_signal_11001 ;
    wire new_AGEMA_signal_11002 ;
    wire new_AGEMA_signal_11003 ;
    wire new_AGEMA_signal_11004 ;
    wire new_AGEMA_signal_11005 ;
    wire new_AGEMA_signal_11006 ;
    wire new_AGEMA_signal_11007 ;
    wire new_AGEMA_signal_11008 ;
    wire new_AGEMA_signal_11009 ;
    wire new_AGEMA_signal_11010 ;
    wire new_AGEMA_signal_11011 ;
    wire new_AGEMA_signal_11012 ;
    wire new_AGEMA_signal_11013 ;
    wire new_AGEMA_signal_11014 ;
    wire new_AGEMA_signal_11015 ;
    wire new_AGEMA_signal_11016 ;
    wire new_AGEMA_signal_11017 ;
    wire new_AGEMA_signal_11018 ;
    wire new_AGEMA_signal_11019 ;
    wire new_AGEMA_signal_11020 ;
    wire new_AGEMA_signal_11021 ;
    wire new_AGEMA_signal_11022 ;
    wire new_AGEMA_signal_11023 ;
    wire new_AGEMA_signal_11024 ;
    wire new_AGEMA_signal_11025 ;
    wire new_AGEMA_signal_11026 ;
    wire new_AGEMA_signal_11027 ;
    wire new_AGEMA_signal_11028 ;
    wire new_AGEMA_signal_11029 ;
    wire new_AGEMA_signal_11030 ;
    wire new_AGEMA_signal_11031 ;
    wire new_AGEMA_signal_11032 ;
    wire new_AGEMA_signal_11033 ;
    wire new_AGEMA_signal_11034 ;
    wire new_AGEMA_signal_11035 ;
    wire new_AGEMA_signal_11036 ;
    wire new_AGEMA_signal_11037 ;
    wire new_AGEMA_signal_11038 ;
    wire new_AGEMA_signal_11039 ;
    wire new_AGEMA_signal_11040 ;
    wire new_AGEMA_signal_11041 ;
    wire new_AGEMA_signal_11042 ;
    wire new_AGEMA_signal_11043 ;
    wire new_AGEMA_signal_11044 ;
    wire new_AGEMA_signal_11045 ;
    wire new_AGEMA_signal_11046 ;
    wire new_AGEMA_signal_11047 ;
    wire new_AGEMA_signal_11048 ;
    wire new_AGEMA_signal_11049 ;
    wire new_AGEMA_signal_11050 ;
    wire new_AGEMA_signal_11051 ;
    wire new_AGEMA_signal_11052 ;
    wire new_AGEMA_signal_11053 ;
    wire new_AGEMA_signal_11054 ;
    wire new_AGEMA_signal_11055 ;
    wire new_AGEMA_signal_11056 ;
    wire new_AGEMA_signal_11057 ;
    wire new_AGEMA_signal_11058 ;
    wire new_AGEMA_signal_11059 ;
    wire new_AGEMA_signal_11060 ;
    wire new_AGEMA_signal_11061 ;
    wire new_AGEMA_signal_11062 ;
    wire new_AGEMA_signal_11063 ;
    wire new_AGEMA_signal_11064 ;
    wire new_AGEMA_signal_11065 ;
    wire new_AGEMA_signal_11066 ;
    wire new_AGEMA_signal_11067 ;
    wire new_AGEMA_signal_11068 ;
    wire new_AGEMA_signal_11069 ;
    wire new_AGEMA_signal_11070 ;
    wire new_AGEMA_signal_11071 ;
    wire new_AGEMA_signal_11072 ;
    wire new_AGEMA_signal_11073 ;
    wire new_AGEMA_signal_11074 ;
    wire new_AGEMA_signal_11075 ;
    wire new_AGEMA_signal_11076 ;
    wire new_AGEMA_signal_11077 ;
    wire new_AGEMA_signal_11078 ;
    wire new_AGEMA_signal_11079 ;
    wire new_AGEMA_signal_11080 ;
    wire new_AGEMA_signal_11081 ;
    wire new_AGEMA_signal_11082 ;
    wire new_AGEMA_signal_11083 ;
    wire new_AGEMA_signal_11084 ;
    wire new_AGEMA_signal_11085 ;
    wire new_AGEMA_signal_11086 ;
    wire new_AGEMA_signal_11087 ;
    wire new_AGEMA_signal_11088 ;
    wire new_AGEMA_signal_11089 ;
    wire new_AGEMA_signal_11090 ;
    wire new_AGEMA_signal_11091 ;
    wire new_AGEMA_signal_11092 ;
    wire new_AGEMA_signal_11093 ;
    wire new_AGEMA_signal_11094 ;
    wire new_AGEMA_signal_11095 ;
    wire new_AGEMA_signal_11096 ;
    wire new_AGEMA_signal_11097 ;
    wire new_AGEMA_signal_11098 ;
    wire new_AGEMA_signal_11099 ;
    wire new_AGEMA_signal_11100 ;
    wire new_AGEMA_signal_11101 ;
    wire new_AGEMA_signal_11102 ;
    wire new_AGEMA_signal_11103 ;
    wire new_AGEMA_signal_11104 ;
    wire new_AGEMA_signal_11105 ;
    wire new_AGEMA_signal_11106 ;
    wire new_AGEMA_signal_11107 ;
    wire new_AGEMA_signal_11108 ;
    wire new_AGEMA_signal_11109 ;
    wire new_AGEMA_signal_11110 ;
    wire new_AGEMA_signal_11111 ;
    wire new_AGEMA_signal_11112 ;
    wire new_AGEMA_signal_11113 ;
    wire new_AGEMA_signal_11114 ;
    wire new_AGEMA_signal_11115 ;
    wire new_AGEMA_signal_11116 ;
    wire new_AGEMA_signal_11117 ;
    wire new_AGEMA_signal_11118 ;
    wire new_AGEMA_signal_11119 ;
    wire new_AGEMA_signal_11120 ;
    wire new_AGEMA_signal_11121 ;
    wire new_AGEMA_signal_11122 ;
    wire new_AGEMA_signal_11123 ;
    wire new_AGEMA_signal_11124 ;
    wire new_AGEMA_signal_11125 ;
    wire new_AGEMA_signal_11126 ;
    wire new_AGEMA_signal_11127 ;
    wire new_AGEMA_signal_11128 ;
    wire new_AGEMA_signal_11129 ;
    wire new_AGEMA_signal_11130 ;
    wire new_AGEMA_signal_11131 ;
    wire new_AGEMA_signal_11132 ;
    wire new_AGEMA_signal_11133 ;
    wire new_AGEMA_signal_11134 ;
    wire new_AGEMA_signal_11135 ;
    wire new_AGEMA_signal_11136 ;
    wire new_AGEMA_signal_11137 ;
    wire new_AGEMA_signal_11138 ;
    wire new_AGEMA_signal_11139 ;
    wire new_AGEMA_signal_11140 ;
    wire new_AGEMA_signal_11141 ;
    wire new_AGEMA_signal_11142 ;
    wire new_AGEMA_signal_11143 ;
    wire new_AGEMA_signal_11144 ;
    wire new_AGEMA_signal_11145 ;
    wire new_AGEMA_signal_11146 ;
    wire new_AGEMA_signal_11147 ;
    wire new_AGEMA_signal_11148 ;
    wire new_AGEMA_signal_11149 ;
    wire new_AGEMA_signal_11150 ;
    wire new_AGEMA_signal_11151 ;
    wire new_AGEMA_signal_11152 ;
    wire new_AGEMA_signal_11153 ;
    wire new_AGEMA_signal_11154 ;
    wire new_AGEMA_signal_11155 ;
    wire new_AGEMA_signal_11156 ;
    wire new_AGEMA_signal_11157 ;
    wire new_AGEMA_signal_11158 ;
    wire new_AGEMA_signal_11159 ;
    wire new_AGEMA_signal_11160 ;
    wire new_AGEMA_signal_11161 ;
    wire new_AGEMA_signal_11162 ;
    wire new_AGEMA_signal_11163 ;
    wire new_AGEMA_signal_11164 ;
    wire new_AGEMA_signal_11165 ;
    wire new_AGEMA_signal_11166 ;
    wire new_AGEMA_signal_11167 ;
    wire new_AGEMA_signal_11168 ;
    wire new_AGEMA_signal_11169 ;
    wire new_AGEMA_signal_11170 ;
    wire new_AGEMA_signal_11171 ;
    wire new_AGEMA_signal_11172 ;
    wire new_AGEMA_signal_11173 ;
    wire new_AGEMA_signal_11174 ;
    wire new_AGEMA_signal_11175 ;
    wire new_AGEMA_signal_11176 ;
    wire new_AGEMA_signal_11177 ;
    wire new_AGEMA_signal_11178 ;
    wire new_AGEMA_signal_11179 ;
    wire new_AGEMA_signal_11180 ;
    wire new_AGEMA_signal_11181 ;
    wire new_AGEMA_signal_11182 ;
    wire new_AGEMA_signal_11183 ;
    wire new_AGEMA_signal_11184 ;
    wire new_AGEMA_signal_11185 ;
    wire new_AGEMA_signal_11186 ;
    wire new_AGEMA_signal_11187 ;
    wire new_AGEMA_signal_11188 ;
    wire new_AGEMA_signal_11189 ;
    wire new_AGEMA_signal_11190 ;
    wire new_AGEMA_signal_11191 ;
    wire new_AGEMA_signal_11192 ;
    wire new_AGEMA_signal_11193 ;
    wire new_AGEMA_signal_11194 ;
    wire new_AGEMA_signal_11195 ;
    wire new_AGEMA_signal_11196 ;
    wire new_AGEMA_signal_11197 ;
    wire new_AGEMA_signal_11198 ;
    wire new_AGEMA_signal_11199 ;
    wire new_AGEMA_signal_11200 ;
    wire new_AGEMA_signal_11201 ;
    wire new_AGEMA_signal_11202 ;
    wire new_AGEMA_signal_11203 ;
    wire new_AGEMA_signal_11204 ;
    wire new_AGEMA_signal_11205 ;
    wire new_AGEMA_signal_11206 ;
    wire new_AGEMA_signal_11207 ;
    wire new_AGEMA_signal_11208 ;
    wire new_AGEMA_signal_11209 ;
    wire new_AGEMA_signal_11210 ;
    wire new_AGEMA_signal_11211 ;
    wire new_AGEMA_signal_11212 ;
    wire new_AGEMA_signal_11213 ;
    wire new_AGEMA_signal_11214 ;
    wire new_AGEMA_signal_11215 ;
    wire new_AGEMA_signal_11216 ;
    wire new_AGEMA_signal_11217 ;
    wire new_AGEMA_signal_11218 ;
    wire new_AGEMA_signal_11219 ;
    wire new_AGEMA_signal_11220 ;
    wire new_AGEMA_signal_11221 ;
    wire new_AGEMA_signal_11222 ;
    wire new_AGEMA_signal_11223 ;
    wire new_AGEMA_signal_11224 ;
    wire new_AGEMA_signal_11225 ;
    wire new_AGEMA_signal_11226 ;
    wire new_AGEMA_signal_11227 ;
    wire new_AGEMA_signal_11228 ;
    wire new_AGEMA_signal_11229 ;
    wire new_AGEMA_signal_11230 ;
    wire new_AGEMA_signal_11231 ;
    wire new_AGEMA_signal_11232 ;
    wire new_AGEMA_signal_11233 ;
    wire new_AGEMA_signal_11234 ;
    wire new_AGEMA_signal_11235 ;
    wire new_AGEMA_signal_11236 ;
    wire new_AGEMA_signal_11237 ;
    wire new_AGEMA_signal_11238 ;
    wire new_AGEMA_signal_11239 ;
    wire new_AGEMA_signal_11240 ;
    wire new_AGEMA_signal_11241 ;
    wire new_AGEMA_signal_11242 ;
    wire new_AGEMA_signal_11243 ;
    wire new_AGEMA_signal_11244 ;
    wire new_AGEMA_signal_11245 ;
    wire new_AGEMA_signal_11246 ;
    wire new_AGEMA_signal_11247 ;
    wire new_AGEMA_signal_11248 ;
    wire new_AGEMA_signal_11249 ;
    wire new_AGEMA_signal_11250 ;
    wire new_AGEMA_signal_11251 ;
    wire new_AGEMA_signal_11252 ;
    wire new_AGEMA_signal_11253 ;
    wire new_AGEMA_signal_11254 ;
    wire new_AGEMA_signal_11255 ;
    wire new_AGEMA_signal_11256 ;
    wire new_AGEMA_signal_11257 ;
    wire new_AGEMA_signal_11258 ;
    wire new_AGEMA_signal_11259 ;
    wire new_AGEMA_signal_11260 ;
    wire new_AGEMA_signal_11261 ;
    wire new_AGEMA_signal_11262 ;
    wire new_AGEMA_signal_11263 ;
    wire new_AGEMA_signal_11264 ;
    wire new_AGEMA_signal_11265 ;
    wire new_AGEMA_signal_11266 ;
    wire new_AGEMA_signal_11267 ;
    wire new_AGEMA_signal_11268 ;
    wire new_AGEMA_signal_11269 ;
    wire new_AGEMA_signal_11270 ;
    wire new_AGEMA_signal_11271 ;
    wire new_AGEMA_signal_11272 ;
    wire new_AGEMA_signal_11273 ;
    wire new_AGEMA_signal_11274 ;
    wire new_AGEMA_signal_11275 ;
    wire new_AGEMA_signal_11276 ;
    wire new_AGEMA_signal_11277 ;
    wire new_AGEMA_signal_11278 ;
    wire new_AGEMA_signal_11279 ;
    wire new_AGEMA_signal_11280 ;
    wire new_AGEMA_signal_11281 ;
    wire new_AGEMA_signal_11282 ;
    wire new_AGEMA_signal_11283 ;
    wire new_AGEMA_signal_11284 ;
    wire new_AGEMA_signal_11285 ;
    wire new_AGEMA_signal_11286 ;
    wire new_AGEMA_signal_11287 ;
    wire new_AGEMA_signal_11288 ;
    wire new_AGEMA_signal_11289 ;
    wire new_AGEMA_signal_11290 ;
    wire new_AGEMA_signal_11291 ;
    wire new_AGEMA_signal_11292 ;
    wire new_AGEMA_signal_11293 ;
    wire new_AGEMA_signal_11294 ;
    wire new_AGEMA_signal_11295 ;
    wire new_AGEMA_signal_11296 ;
    wire new_AGEMA_signal_11297 ;
    wire new_AGEMA_signal_11298 ;
    wire new_AGEMA_signal_11299 ;
    wire new_AGEMA_signal_11300 ;
    wire new_AGEMA_signal_11301 ;
    wire new_AGEMA_signal_11302 ;
    wire new_AGEMA_signal_11303 ;
    wire new_AGEMA_signal_11304 ;
    wire new_AGEMA_signal_11305 ;
    wire new_AGEMA_signal_11306 ;
    wire new_AGEMA_signal_11307 ;
    wire new_AGEMA_signal_11308 ;
    wire new_AGEMA_signal_11309 ;
    wire new_AGEMA_signal_11310 ;
    wire new_AGEMA_signal_11311 ;
    wire new_AGEMA_signal_11312 ;
    wire new_AGEMA_signal_11313 ;
    wire new_AGEMA_signal_11314 ;
    wire new_AGEMA_signal_11315 ;
    wire new_AGEMA_signal_11316 ;
    wire new_AGEMA_signal_11317 ;
    wire new_AGEMA_signal_11318 ;
    wire new_AGEMA_signal_11319 ;
    wire new_AGEMA_signal_11320 ;
    wire new_AGEMA_signal_11321 ;
    wire new_AGEMA_signal_11322 ;
    wire new_AGEMA_signal_11323 ;
    wire new_AGEMA_signal_11324 ;
    wire new_AGEMA_signal_11325 ;
    wire new_AGEMA_signal_11326 ;
    wire new_AGEMA_signal_11327 ;
    wire new_AGEMA_signal_11328 ;
    wire new_AGEMA_signal_11329 ;
    wire new_AGEMA_signal_11330 ;
    wire new_AGEMA_signal_11331 ;
    wire new_AGEMA_signal_11332 ;
    wire new_AGEMA_signal_11333 ;
    wire new_AGEMA_signal_11334 ;
    wire new_AGEMA_signal_11335 ;
    wire new_AGEMA_signal_11336 ;
    wire new_AGEMA_signal_11337 ;
    wire new_AGEMA_signal_11338 ;
    wire new_AGEMA_signal_11339 ;
    wire new_AGEMA_signal_11340 ;
    wire new_AGEMA_signal_11341 ;
    wire new_AGEMA_signal_11342 ;
    wire new_AGEMA_signal_11343 ;
    wire new_AGEMA_signal_11344 ;
    wire new_AGEMA_signal_11345 ;
    wire new_AGEMA_signal_11346 ;
    wire new_AGEMA_signal_11347 ;
    wire new_AGEMA_signal_11348 ;
    wire new_AGEMA_signal_11349 ;
    wire new_AGEMA_signal_11350 ;
    wire new_AGEMA_signal_11351 ;
    wire new_AGEMA_signal_11352 ;
    wire new_AGEMA_signal_11353 ;
    wire new_AGEMA_signal_11354 ;
    wire new_AGEMA_signal_11355 ;
    wire new_AGEMA_signal_11356 ;
    wire new_AGEMA_signal_11357 ;
    wire new_AGEMA_signal_11358 ;
    wire new_AGEMA_signal_11359 ;
    wire new_AGEMA_signal_11360 ;
    wire new_AGEMA_signal_11361 ;
    wire new_AGEMA_signal_11362 ;
    wire new_AGEMA_signal_11363 ;
    wire new_AGEMA_signal_11364 ;
    wire new_AGEMA_signal_11365 ;
    wire new_AGEMA_signal_11366 ;
    wire new_AGEMA_signal_11367 ;
    wire new_AGEMA_signal_11368 ;
    wire new_AGEMA_signal_11369 ;
    wire new_AGEMA_signal_11370 ;
    wire new_AGEMA_signal_11371 ;
    wire new_AGEMA_signal_11372 ;
    wire new_AGEMA_signal_11373 ;
    wire new_AGEMA_signal_11374 ;
    wire new_AGEMA_signal_11375 ;
    wire new_AGEMA_signal_11376 ;
    wire new_AGEMA_signal_11377 ;
    wire new_AGEMA_signal_11378 ;
    wire new_AGEMA_signal_11379 ;
    wire new_AGEMA_signal_11380 ;
    wire new_AGEMA_signal_11381 ;
    wire new_AGEMA_signal_11382 ;
    wire new_AGEMA_signal_11383 ;
    wire new_AGEMA_signal_11384 ;
    wire new_AGEMA_signal_11385 ;
    wire new_AGEMA_signal_11386 ;
    wire new_AGEMA_signal_11387 ;
    wire new_AGEMA_signal_11388 ;
    wire new_AGEMA_signal_11389 ;
    wire new_AGEMA_signal_11390 ;
    wire new_AGEMA_signal_11391 ;
    wire new_AGEMA_signal_11392 ;
    wire new_AGEMA_signal_11393 ;
    wire new_AGEMA_signal_11394 ;
    wire new_AGEMA_signal_11395 ;
    wire new_AGEMA_signal_11396 ;
    wire new_AGEMA_signal_11397 ;
    wire new_AGEMA_signal_11398 ;
    wire new_AGEMA_signal_11399 ;
    wire new_AGEMA_signal_11400 ;
    wire new_AGEMA_signal_11401 ;
    wire new_AGEMA_signal_11402 ;
    wire new_AGEMA_signal_11403 ;
    wire new_AGEMA_signal_11404 ;
    wire new_AGEMA_signal_11405 ;
    wire new_AGEMA_signal_11406 ;
    wire new_AGEMA_signal_11407 ;
    wire new_AGEMA_signal_11408 ;
    wire new_AGEMA_signal_11409 ;
    wire new_AGEMA_signal_11410 ;
    wire new_AGEMA_signal_11411 ;
    wire new_AGEMA_signal_11412 ;
    wire new_AGEMA_signal_11413 ;
    wire new_AGEMA_signal_11414 ;
    wire new_AGEMA_signal_11415 ;
    wire new_AGEMA_signal_11416 ;
    wire new_AGEMA_signal_11417 ;
    wire new_AGEMA_signal_11418 ;
    wire new_AGEMA_signal_11419 ;
    wire new_AGEMA_signal_11420 ;
    wire new_AGEMA_signal_11421 ;
    wire new_AGEMA_signal_11422 ;
    wire new_AGEMA_signal_11423 ;
    wire new_AGEMA_signal_11424 ;
    wire new_AGEMA_signal_11425 ;
    wire new_AGEMA_signal_11426 ;
    wire new_AGEMA_signal_11427 ;
    wire new_AGEMA_signal_11428 ;
    wire new_AGEMA_signal_11429 ;
    wire new_AGEMA_signal_11430 ;
    wire new_AGEMA_signal_11431 ;
    wire new_AGEMA_signal_11432 ;
    wire new_AGEMA_signal_11433 ;
    wire new_AGEMA_signal_11434 ;
    wire new_AGEMA_signal_11435 ;
    wire new_AGEMA_signal_11436 ;
    wire new_AGEMA_signal_11437 ;
    wire new_AGEMA_signal_11438 ;
    wire new_AGEMA_signal_11439 ;
    wire new_AGEMA_signal_11440 ;
    wire new_AGEMA_signal_11441 ;
    wire new_AGEMA_signal_11442 ;
    wire new_AGEMA_signal_11443 ;
    wire new_AGEMA_signal_11444 ;
    wire new_AGEMA_signal_11445 ;
    wire new_AGEMA_signal_11446 ;
    wire new_AGEMA_signal_11447 ;
    wire new_AGEMA_signal_11448 ;
    wire new_AGEMA_signal_11449 ;
    wire new_AGEMA_signal_11450 ;
    wire new_AGEMA_signal_11451 ;
    wire new_AGEMA_signal_11452 ;
    wire new_AGEMA_signal_11453 ;
    wire new_AGEMA_signal_11454 ;
    wire new_AGEMA_signal_11455 ;
    wire new_AGEMA_signal_11456 ;
    wire new_AGEMA_signal_11457 ;
    wire new_AGEMA_signal_11458 ;
    wire new_AGEMA_signal_11459 ;
    wire new_AGEMA_signal_11460 ;
    wire new_AGEMA_signal_11461 ;
    wire new_AGEMA_signal_11462 ;
    wire new_AGEMA_signal_11463 ;
    wire new_AGEMA_signal_11464 ;
    wire new_AGEMA_signal_11465 ;
    wire new_AGEMA_signal_11466 ;
    wire new_AGEMA_signal_11467 ;
    wire new_AGEMA_signal_11468 ;
    wire new_AGEMA_signal_11469 ;
    wire new_AGEMA_signal_11470 ;
    wire new_AGEMA_signal_11471 ;
    wire new_AGEMA_signal_11472 ;
    wire new_AGEMA_signal_11473 ;
    wire new_AGEMA_signal_11474 ;
    wire new_AGEMA_signal_11475 ;
    wire new_AGEMA_signal_11476 ;
    wire new_AGEMA_signal_11477 ;
    wire new_AGEMA_signal_11478 ;
    wire new_AGEMA_signal_11479 ;
    wire new_AGEMA_signal_11480 ;
    wire new_AGEMA_signal_11481 ;
    wire new_AGEMA_signal_11482 ;
    wire new_AGEMA_signal_11483 ;
    wire new_AGEMA_signal_11484 ;
    wire new_AGEMA_signal_11485 ;
    wire new_AGEMA_signal_11486 ;
    wire new_AGEMA_signal_11487 ;
    wire new_AGEMA_signal_11488 ;
    wire new_AGEMA_signal_11489 ;
    wire new_AGEMA_signal_11490 ;
    wire new_AGEMA_signal_11491 ;
    wire new_AGEMA_signal_11492 ;
    wire new_AGEMA_signal_11493 ;
    wire new_AGEMA_signal_11494 ;
    wire new_AGEMA_signal_11495 ;
    wire new_AGEMA_signal_11496 ;
    wire new_AGEMA_signal_11497 ;
    wire new_AGEMA_signal_11498 ;
    wire new_AGEMA_signal_11499 ;
    wire new_AGEMA_signal_11500 ;
    wire new_AGEMA_signal_11501 ;
    wire new_AGEMA_signal_11502 ;
    wire new_AGEMA_signal_11503 ;
    wire new_AGEMA_signal_11504 ;
    wire new_AGEMA_signal_11505 ;
    wire new_AGEMA_signal_11506 ;
    wire new_AGEMA_signal_11507 ;
    wire new_AGEMA_signal_11508 ;
    wire new_AGEMA_signal_11509 ;
    wire new_AGEMA_signal_11510 ;
    wire new_AGEMA_signal_11511 ;
    wire new_AGEMA_signal_11512 ;
    wire new_AGEMA_signal_11513 ;
    wire new_AGEMA_signal_11514 ;
    wire new_AGEMA_signal_11515 ;
    wire new_AGEMA_signal_11516 ;
    wire new_AGEMA_signal_11517 ;
    wire new_AGEMA_signal_11518 ;
    wire new_AGEMA_signal_11519 ;
    wire new_AGEMA_signal_11520 ;
    wire new_AGEMA_signal_11521 ;
    wire new_AGEMA_signal_11522 ;
    wire new_AGEMA_signal_11523 ;
    wire new_AGEMA_signal_11524 ;
    wire new_AGEMA_signal_11525 ;
    wire new_AGEMA_signal_11526 ;
    wire new_AGEMA_signal_11527 ;
    wire new_AGEMA_signal_11528 ;
    wire new_AGEMA_signal_11529 ;
    wire new_AGEMA_signal_11530 ;
    wire new_AGEMA_signal_11531 ;
    wire new_AGEMA_signal_11532 ;
    wire new_AGEMA_signal_11533 ;
    wire new_AGEMA_signal_11534 ;
    wire new_AGEMA_signal_11535 ;
    wire new_AGEMA_signal_11536 ;
    wire new_AGEMA_signal_11537 ;
    wire new_AGEMA_signal_11538 ;
    wire new_AGEMA_signal_11539 ;
    wire new_AGEMA_signal_11540 ;
    wire new_AGEMA_signal_11541 ;
    wire new_AGEMA_signal_11542 ;
    wire new_AGEMA_signal_11543 ;
    wire new_AGEMA_signal_11544 ;
    wire new_AGEMA_signal_11545 ;
    wire new_AGEMA_signal_11546 ;
    wire new_AGEMA_signal_11547 ;
    wire new_AGEMA_signal_11548 ;
    wire new_AGEMA_signal_11549 ;
    wire new_AGEMA_signal_11550 ;
    wire new_AGEMA_signal_11551 ;
    wire new_AGEMA_signal_11552 ;
    wire new_AGEMA_signal_11553 ;
    wire new_AGEMA_signal_11554 ;
    wire new_AGEMA_signal_11555 ;
    wire new_AGEMA_signal_11556 ;
    wire new_AGEMA_signal_11557 ;
    wire new_AGEMA_signal_11558 ;
    wire new_AGEMA_signal_11559 ;
    wire new_AGEMA_signal_11560 ;
    wire new_AGEMA_signal_11561 ;
    wire new_AGEMA_signal_11562 ;
    wire new_AGEMA_signal_11563 ;
    wire new_AGEMA_signal_11564 ;
    wire new_AGEMA_signal_11565 ;
    wire new_AGEMA_signal_11566 ;
    wire new_AGEMA_signal_11567 ;
    wire new_AGEMA_signal_11568 ;
    wire new_AGEMA_signal_11569 ;
    wire new_AGEMA_signal_11570 ;
    wire new_AGEMA_signal_11571 ;
    wire new_AGEMA_signal_11572 ;
    wire new_AGEMA_signal_11573 ;
    wire new_AGEMA_signal_11574 ;
    wire new_AGEMA_signal_11575 ;
    wire new_AGEMA_signal_11576 ;
    wire new_AGEMA_signal_11577 ;
    wire new_AGEMA_signal_11578 ;
    wire new_AGEMA_signal_11579 ;
    wire new_AGEMA_signal_11580 ;
    wire new_AGEMA_signal_11581 ;
    wire new_AGEMA_signal_11582 ;
    wire new_AGEMA_signal_11583 ;
    wire new_AGEMA_signal_11584 ;
    wire new_AGEMA_signal_11585 ;
    wire new_AGEMA_signal_11586 ;
    wire new_AGEMA_signal_11587 ;
    wire new_AGEMA_signal_11588 ;
    wire new_AGEMA_signal_11589 ;
    wire new_AGEMA_signal_11590 ;
    wire new_AGEMA_signal_11591 ;
    wire new_AGEMA_signal_11592 ;
    wire new_AGEMA_signal_11593 ;
    wire new_AGEMA_signal_11594 ;
    wire new_AGEMA_signal_11595 ;
    wire new_AGEMA_signal_11596 ;
    wire new_AGEMA_signal_11597 ;
    wire new_AGEMA_signal_11598 ;
    wire new_AGEMA_signal_11599 ;
    wire new_AGEMA_signal_11600 ;
    wire new_AGEMA_signal_11601 ;
    wire new_AGEMA_signal_11602 ;
    wire new_AGEMA_signal_11603 ;
    wire new_AGEMA_signal_11604 ;
    wire new_AGEMA_signal_11605 ;
    wire new_AGEMA_signal_11606 ;
    wire new_AGEMA_signal_11607 ;
    wire new_AGEMA_signal_11608 ;
    wire new_AGEMA_signal_11609 ;
    wire new_AGEMA_signal_11610 ;
    wire new_AGEMA_signal_11611 ;
    wire new_AGEMA_signal_11615 ;
    wire new_AGEMA_signal_11616 ;
    wire new_AGEMA_signal_11617 ;
    wire new_AGEMA_signal_11618 ;
    wire new_AGEMA_signal_11619 ;
    wire new_AGEMA_signal_11620 ;
    wire new_AGEMA_signal_11621 ;
    wire new_AGEMA_signal_11622 ;
    wire new_AGEMA_signal_11623 ;
    wire new_AGEMA_signal_11624 ;
    wire new_AGEMA_signal_11625 ;
    wire new_AGEMA_signal_11626 ;
    wire new_AGEMA_signal_11627 ;
    wire new_AGEMA_signal_11628 ;
    wire new_AGEMA_signal_11629 ;
    wire new_AGEMA_signal_11630 ;
    wire new_AGEMA_signal_11631 ;
    wire new_AGEMA_signal_11632 ;
    wire new_AGEMA_signal_11633 ;
    wire new_AGEMA_signal_11634 ;
    wire new_AGEMA_signal_11635 ;
    wire new_AGEMA_signal_11636 ;
    wire new_AGEMA_signal_11637 ;
    wire new_AGEMA_signal_11638 ;
    wire new_AGEMA_signal_11639 ;
    wire new_AGEMA_signal_11640 ;
    wire new_AGEMA_signal_11641 ;
    wire new_AGEMA_signal_11645 ;
    wire new_AGEMA_signal_11646 ;
    wire new_AGEMA_signal_11647 ;
    wire new_AGEMA_signal_11651 ;
    wire new_AGEMA_signal_11652 ;
    wire new_AGEMA_signal_11653 ;
    wire new_AGEMA_signal_11657 ;
    wire new_AGEMA_signal_11658 ;
    wire new_AGEMA_signal_11659 ;
    wire new_AGEMA_signal_11663 ;
    wire new_AGEMA_signal_11664 ;
    wire new_AGEMA_signal_11665 ;
    wire new_AGEMA_signal_11669 ;
    wire new_AGEMA_signal_11670 ;
    wire new_AGEMA_signal_11671 ;
    wire new_AGEMA_signal_11675 ;
    wire new_AGEMA_signal_11676 ;
    wire new_AGEMA_signal_11677 ;
    wire new_AGEMA_signal_11681 ;
    wire new_AGEMA_signal_11682 ;
    wire new_AGEMA_signal_11683 ;
    wire new_AGEMA_signal_11684 ;
    wire new_AGEMA_signal_11685 ;
    wire new_AGEMA_signal_11686 ;
    wire new_AGEMA_signal_11687 ;
    wire new_AGEMA_signal_11688 ;
    wire new_AGEMA_signal_11689 ;
    wire new_AGEMA_signal_11690 ;
    wire new_AGEMA_signal_11691 ;
    wire new_AGEMA_signal_11692 ;
    wire new_AGEMA_signal_11693 ;
    wire new_AGEMA_signal_11694 ;
    wire new_AGEMA_signal_11695 ;
    wire new_AGEMA_signal_11696 ;
    wire new_AGEMA_signal_11697 ;
    wire new_AGEMA_signal_11698 ;
    wire new_AGEMA_signal_11699 ;
    wire new_AGEMA_signal_11700 ;
    wire new_AGEMA_signal_11701 ;
    wire new_AGEMA_signal_11702 ;
    wire new_AGEMA_signal_11703 ;
    wire new_AGEMA_signal_11704 ;
    wire new_AGEMA_signal_11705 ;
    wire new_AGEMA_signal_11706 ;
    wire new_AGEMA_signal_11707 ;
    wire new_AGEMA_signal_11708 ;
    wire new_AGEMA_signal_11709 ;
    wire new_AGEMA_signal_11710 ;
    wire new_AGEMA_signal_11711 ;
    wire new_AGEMA_signal_11712 ;
    wire new_AGEMA_signal_11713 ;
    wire new_AGEMA_signal_11714 ;
    wire new_AGEMA_signal_11715 ;
    wire new_AGEMA_signal_11716 ;
    wire new_AGEMA_signal_11717 ;
    wire new_AGEMA_signal_11718 ;
    wire new_AGEMA_signal_11719 ;
    wire new_AGEMA_signal_11720 ;
    wire new_AGEMA_signal_11721 ;
    wire new_AGEMA_signal_11722 ;
    wire new_AGEMA_signal_11723 ;
    wire new_AGEMA_signal_11724 ;
    wire new_AGEMA_signal_11725 ;
    wire new_AGEMA_signal_11726 ;
    wire new_AGEMA_signal_11727 ;
    wire new_AGEMA_signal_11728 ;
    wire new_AGEMA_signal_11729 ;
    wire new_AGEMA_signal_11730 ;
    wire new_AGEMA_signal_11731 ;
    wire new_AGEMA_signal_11732 ;
    wire new_AGEMA_signal_11733 ;
    wire new_AGEMA_signal_11734 ;
    wire new_AGEMA_signal_11735 ;
    wire new_AGEMA_signal_11736 ;
    wire new_AGEMA_signal_11737 ;
    wire new_AGEMA_signal_11738 ;
    wire new_AGEMA_signal_11739 ;
    wire new_AGEMA_signal_11740 ;
    wire new_AGEMA_signal_11741 ;
    wire new_AGEMA_signal_11742 ;
    wire new_AGEMA_signal_11743 ;
    wire new_AGEMA_signal_11744 ;
    wire new_AGEMA_signal_11745 ;
    wire new_AGEMA_signal_11746 ;
    wire new_AGEMA_signal_11747 ;
    wire new_AGEMA_signal_11748 ;
    wire new_AGEMA_signal_11749 ;
    wire new_AGEMA_signal_11750 ;
    wire new_AGEMA_signal_11751 ;
    wire new_AGEMA_signal_11752 ;
    wire new_AGEMA_signal_11753 ;
    wire new_AGEMA_signal_11754 ;
    wire new_AGEMA_signal_11755 ;
    wire new_AGEMA_signal_11756 ;
    wire new_AGEMA_signal_11757 ;
    wire new_AGEMA_signal_11758 ;
    wire new_AGEMA_signal_11759 ;
    wire new_AGEMA_signal_11760 ;
    wire new_AGEMA_signal_11761 ;
    wire new_AGEMA_signal_11762 ;
    wire new_AGEMA_signal_11763 ;
    wire new_AGEMA_signal_11764 ;
    wire new_AGEMA_signal_11765 ;
    wire new_AGEMA_signal_11766 ;
    wire new_AGEMA_signal_11767 ;
    wire new_AGEMA_signal_11768 ;
    wire new_AGEMA_signal_11769 ;
    wire new_AGEMA_signal_11770 ;
    wire new_AGEMA_signal_11771 ;
    wire new_AGEMA_signal_11772 ;
    wire new_AGEMA_signal_11773 ;
    wire new_AGEMA_signal_11774 ;
    wire new_AGEMA_signal_11775 ;
    wire new_AGEMA_signal_11776 ;

    /* cells in depth 0 */
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U31 ( .A0_t (ciphertext_s0_t[120]), .A0_f (ciphertext_s0_f[120]), .A1_t (ciphertext_s1_t[120]), .A1_f (ciphertext_s1_f[120]), .B0_t (keyStateIn[0]), .B0_f (new_AGEMA_signal_3432), .B1_t (new_AGEMA_signal_3433), .B1_f (new_AGEMA_signal_3434), .Z0_t (StateOutXORroundKey[0]), .Z0_f (new_AGEMA_signal_3435), .Z1_t (new_AGEMA_signal_3436), .Z1_f (new_AGEMA_signal_3437) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U32 ( .A0_t (ciphertext_s0_t[121]), .A0_f (ciphertext_s0_f[121]), .A1_t (ciphertext_s1_t[121]), .A1_f (ciphertext_s1_f[121]), .B0_t (keyStateIn[1]), .B0_f (new_AGEMA_signal_3441), .B1_t (new_AGEMA_signal_3442), .B1_f (new_AGEMA_signal_3443), .Z0_t (StateOutXORroundKey[1]), .Z0_f (new_AGEMA_signal_3444), .Z1_t (new_AGEMA_signal_3445), .Z1_f (new_AGEMA_signal_3446) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U33 ( .A0_t (ciphertext_s0_t[122]), .A0_f (ciphertext_s0_f[122]), .A1_t (ciphertext_s1_t[122]), .A1_f (ciphertext_s1_f[122]), .B0_t (keyStateIn[2]), .B0_f (new_AGEMA_signal_3450), .B1_t (new_AGEMA_signal_3451), .B1_f (new_AGEMA_signal_3452), .Z0_t (StateOutXORroundKey[2]), .Z0_f (new_AGEMA_signal_3453), .Z1_t (new_AGEMA_signal_3454), .Z1_f (new_AGEMA_signal_3455) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U34 ( .A0_t (ciphertext_s0_t[123]), .A0_f (ciphertext_s0_f[123]), .A1_t (ciphertext_s1_t[123]), .A1_f (ciphertext_s1_f[123]), .B0_t (keyStateIn[3]), .B0_f (new_AGEMA_signal_3459), .B1_t (new_AGEMA_signal_3460), .B1_f (new_AGEMA_signal_3461), .Z0_t (StateOutXORroundKey[3]), .Z0_f (new_AGEMA_signal_3462), .Z1_t (new_AGEMA_signal_3463), .Z1_f (new_AGEMA_signal_3464) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U35 ( .A0_t (ciphertext_s0_t[124]), .A0_f (ciphertext_s0_f[124]), .A1_t (ciphertext_s1_t[124]), .A1_f (ciphertext_s1_f[124]), .B0_t (keyStateIn[4]), .B0_f (new_AGEMA_signal_3468), .B1_t (new_AGEMA_signal_3469), .B1_f (new_AGEMA_signal_3470), .Z0_t (StateOutXORroundKey[4]), .Z0_f (new_AGEMA_signal_3471), .Z1_t (new_AGEMA_signal_3472), .Z1_f (new_AGEMA_signal_3473) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U36 ( .A0_t (ciphertext_s0_t[125]), .A0_f (ciphertext_s0_f[125]), .A1_t (ciphertext_s1_t[125]), .A1_f (ciphertext_s1_f[125]), .B0_t (keyStateIn[5]), .B0_f (new_AGEMA_signal_3477), .B1_t (new_AGEMA_signal_3478), .B1_f (new_AGEMA_signal_3479), .Z0_t (StateOutXORroundKey[5]), .Z0_f (new_AGEMA_signal_3480), .Z1_t (new_AGEMA_signal_3481), .Z1_f (new_AGEMA_signal_3482) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U37 ( .A0_t (ciphertext_s0_t[126]), .A0_f (ciphertext_s0_f[126]), .A1_t (ciphertext_s1_t[126]), .A1_f (ciphertext_s1_f[126]), .B0_t (keyStateIn[6]), .B0_f (new_AGEMA_signal_3486), .B1_t (new_AGEMA_signal_3487), .B1_f (new_AGEMA_signal_3488), .Z0_t (StateOutXORroundKey[6]), .Z0_f (new_AGEMA_signal_3489), .Z1_t (new_AGEMA_signal_3490), .Z1_f (new_AGEMA_signal_3491) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U38 ( .A0_t (ciphertext_s0_t[127]), .A0_f (ciphertext_s0_f[127]), .A1_t (ciphertext_s1_t[127]), .A1_f (ciphertext_s1_f[127]), .B0_t (keyStateIn[7]), .B0_f (new_AGEMA_signal_3495), .B1_t (new_AGEMA_signal_3496), .B1_f (new_AGEMA_signal_3497), .Z0_t (StateOutXORroundKey[7]), .Z0_f (new_AGEMA_signal_3498), .Z1_t (new_AGEMA_signal_3499), .Z1_f (new_AGEMA_signal_3500) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) U39 ( .A0_t (intFinal), .A0_f (new_AGEMA_signal_6594), .B0_t (finalStep), .B0_f (new_AGEMA_signal_7393), .Z0_t (n13), .Z0_f (new_AGEMA_signal_8139) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) U40 ( .A0_t (nReset), .A0_f (new_AGEMA_signal_3502), .B0_t (n13), .B0_f (new_AGEMA_signal_8139), .Z0_t (done_t), .Z0_f (done_f) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) U41 ( .A0_t (notFirst), .A0_f (new_AGEMA_signal_7366), .B0_t (selXOR), .B0_f (new_AGEMA_signal_5818), .Z0_t (intselXOR), .Z0_f (new_AGEMA_signal_7391) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) ctrl_U20 ( .A0_t (ctrl_n2), .A0_f (new_AGEMA_signal_3501), .B0_t (nReset), .B0_f (new_AGEMA_signal_3502), .Z0_t (selMC), .Z0_f (new_AGEMA_signal_3503) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) ctrl_U19 ( .A0_t (ctrl_n15), .A0_f (new_AGEMA_signal_6620), .B0_t (nReset), .B0_f (new_AGEMA_signal_3502), .Z0_t (ctrl_nRstSeq4), .Z0_f (new_AGEMA_signal_7392) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b0)) ctrl_U18 ( .A0_t (ctrl_seq6Out_4_), .A0_f (new_AGEMA_signal_3504), .B0_t (ctrl_seq6In_1_), .B0_f (new_AGEMA_signal_3505), .Z0_t (ctrl_n13), .Z0_f (new_AGEMA_signal_3506) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) ctrl_U17 ( .A0_t (ctrl_n15), .A0_f (new_AGEMA_signal_6620), .B0_t (ctrl_n11), .B0_f (new_AGEMA_signal_3509), .Z0_t (finalStep), .Z0_f (new_AGEMA_signal_7393) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) ctrl_U16 ( .A0_t (ctrl_seq4In_1_), .A0_f (new_AGEMA_signal_3507), .B0_t (ctrl_seq4Out_1_), .B0_f (new_AGEMA_signal_3508), .Z0_t (ctrl_n11), .Z0_f (new_AGEMA_signal_3509) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1), .NL(1'b1)) ctrl_U13 ( .A0_t (ctrl_n10), .A0_f (new_AGEMA_signal_6619), .B0_t (ctrl_n9), .B0_f (new_AGEMA_signal_7394), .Z0_t (ctrl_n2), .Z0_f (new_AGEMA_signal_3501) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) ctrl_U12 ( .A0_t (selXOR), .A0_f (new_AGEMA_signal_5818), .B0_t (ctrl_n2), .B0_f (new_AGEMA_signal_3501), .Z0_t (ctrl_n10), .Z0_f (new_AGEMA_signal_6619) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) ctrl_U11 ( .A0_t (ctrl_n7), .A0_f (new_AGEMA_signal_3513), .B0_t (ctrl_n6), .B0_f (new_AGEMA_signal_3511), .Z0_t (ctrl_n8), .Z0_f (new_AGEMA_signal_5817) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) ctrl_U10 ( .A0_t (ctrl_seq6In_3_), .A0_f (new_AGEMA_signal_3510), .B0_t (ctrl_seq6Out_4_), .B0_f (new_AGEMA_signal_3504), .Z0_t (ctrl_n6), .Z0_f (new_AGEMA_signal_3511) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) ctrl_U9 ( .A0_t (ctrl_seq6In_1_), .A0_f (new_AGEMA_signal_3505), .B0_t (ctrl_seq6In_4_), .B0_f (new_AGEMA_signal_3512), .Z0_t (ctrl_n7), .Z0_f (new_AGEMA_signal_3513) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) ctrl_U8 ( .A0_t (nReset), .A0_f (new_AGEMA_signal_3502), .B0_t (ctrl_n5), .B0_f (new_AGEMA_signal_3514), .Z0_t (selXOR), .Z0_f (new_AGEMA_signal_5818) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) ctrl_U7 ( .A0_t (ctrl_seq4Out_1_), .A0_f (new_AGEMA_signal_3508), .B0_t (ctrl_seq4In_1_), .B0_f (new_AGEMA_signal_3507), .Z0_t (ctrl_n5), .Z0_f (new_AGEMA_signal_3514) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) ctrl_U5 ( .A0_t (ctrl_seq6In_2_), .A0_f (new_AGEMA_signal_3516), .B0_t (ctrl_n8), .B0_f (new_AGEMA_signal_5817), .Z0_t (ctrl_n15), .Z0_f (new_AGEMA_signal_6620) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) ctrl_U4 ( .A0_t (nReset), .A0_f (new_AGEMA_signal_3502), .B0_t (ctrl_n15), .B0_f (new_AGEMA_signal_6620), .Z0_t (ctrl_n9), .Z0_f (new_AGEMA_signal_7394) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) ctrl_seq6_SFF_0_MUXInst_XOR1_U1 ( .A0_t (1'b1), .A0_f (1'b1), .B0_t (ctrl_n13), .B0_f (new_AGEMA_signal_3506), .Z0_t (ctrl_seq6_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_5819) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) ctrl_seq6_SFF_0_MUXInst_AND1_U1 ( .A0_t (nReset), .A0_f (new_AGEMA_signal_3502), .B0_t (ctrl_seq6_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_5819), .Z0_t (ctrl_seq6_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_6621) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1), .NL(1'b0)) ctrl_seq6_SFF_0_MUXInst_XOR2_U1 ( .A0_t (ctrl_seq6_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_6621), .B0_t (1'b1), .B0_f (1'b1), .Z0_t (ctrl_seq6In_1_), .Z0_f (new_AGEMA_signal_3505) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) ctrl_seq6_SFF_1_MUXInst_XOR1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .B0_t (ctrl_seq6In_1_), .B0_f (new_AGEMA_signal_3505), .Z0_t (ctrl_seq6_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_3515) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) ctrl_seq6_SFF_1_MUXInst_AND1_U1 ( .A0_t (nReset), .A0_f (new_AGEMA_signal_3502), .B0_t (ctrl_seq6_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_3515), .Z0_t (ctrl_seq6_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_5820) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1), .NL(1'b0)) ctrl_seq6_SFF_1_MUXInst_XOR2_U1 ( .A0_t (ctrl_seq6_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_5820), .B0_t (1'b0), .B0_f (1'b1), .Z0_t (ctrl_seq6In_2_), .Z0_f (new_AGEMA_signal_3516) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) ctrl_seq6_SFF_2_MUXInst_XOR1_U1 ( .A0_t (1'b1), .A0_f (1'b1), .B0_t (ctrl_seq6In_2_), .B0_f (new_AGEMA_signal_3516), .Z0_t (ctrl_seq6_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_3517) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) ctrl_seq6_SFF_2_MUXInst_AND1_U1 ( .A0_t (nReset), .A0_f (new_AGEMA_signal_3502), .B0_t (ctrl_seq6_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_3517), .Z0_t (ctrl_seq6_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_5821) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1), .NL(1'b0)) ctrl_seq6_SFF_2_MUXInst_XOR2_U1 ( .A0_t (ctrl_seq6_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_5821), .B0_t (1'b1), .B0_f (1'b1), .Z0_t (ctrl_seq6In_3_), .Z0_f (new_AGEMA_signal_3510) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) ctrl_seq6_SFF_3_MUXInst_XOR1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .B0_t (ctrl_seq6In_3_), .B0_f (new_AGEMA_signal_3510), .Z0_t (ctrl_seq6_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_3518) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) ctrl_seq6_SFF_3_MUXInst_AND1_U1 ( .A0_t (nReset), .A0_f (new_AGEMA_signal_3502), .B0_t (ctrl_seq6_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_3518), .Z0_t (ctrl_seq6_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_5822) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1), .NL(1'b0)) ctrl_seq6_SFF_3_MUXInst_XOR2_U1 ( .A0_t (ctrl_seq6_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_5822), .B0_t (1'b0), .B0_f (1'b1), .Z0_t (ctrl_seq6In_4_), .Z0_f (new_AGEMA_signal_3512) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) ctrl_seq6_SFF_4_MUXInst_XOR1_U1 ( .A0_t (1'b1), .A0_f (1'b1), .B0_t (ctrl_seq6In_4_), .B0_f (new_AGEMA_signal_3512), .Z0_t (ctrl_seq6_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_3519) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) ctrl_seq6_SFF_4_MUXInst_AND1_U1 ( .A0_t (nReset), .A0_f (new_AGEMA_signal_3502), .B0_t (ctrl_seq6_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_3519), .Z0_t (ctrl_seq6_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_5823) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1), .NL(1'b0)) ctrl_seq6_SFF_4_MUXInst_XOR2_U1 ( .A0_t (ctrl_seq6_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_5823), .B0_t (1'b1), .B0_f (1'b1), .Z0_t (ctrl_seq6Out_4_), .Z0_f (new_AGEMA_signal_3504) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) ctrl_seq4_SFF_0_MUXInst_XOR1_U1 ( .A0_t (1'b1), .A0_f (1'b1), .B0_t (ctrl_seq4Out_1_), .B0_f (new_AGEMA_signal_3508), .Z0_t (ctrl_seq4_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_3520) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) ctrl_seq4_SFF_0_MUXInst_AND1_U1 ( .A0_t (ctrl_nRstSeq4), .A0_f (new_AGEMA_signal_7392), .B0_t (ctrl_seq4_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_3520), .Z0_t (ctrl_seq4_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_8140) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1), .NL(1'b0)) ctrl_seq4_SFF_0_MUXInst_XOR2_U1 ( .A0_t (ctrl_seq4_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_8140), .B0_t (1'b1), .B0_f (1'b1), .Z0_t (ctrl_seq4In_1_), .Z0_f (new_AGEMA_signal_3507) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) ctrl_seq4_SFF_1_MUXInst_XOR1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .B0_t (ctrl_seq4In_1_), .B0_f (new_AGEMA_signal_3507), .Z0_t (ctrl_seq4_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_3521) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) ctrl_seq4_SFF_1_MUXInst_AND1_U1 ( .A0_t (ctrl_nRstSeq4), .A0_f (new_AGEMA_signal_7392), .B0_t (ctrl_seq4_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_3521), .Z0_t (ctrl_seq4_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_8141) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1), .NL(1'b0)) ctrl_seq4_SFF_1_MUXInst_XOR2_U1 ( .A0_t (ctrl_seq4_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_8141), .B0_t (1'b0), .B0_f (1'b1), .Z0_t (ctrl_seq4Out_1_), .Z0_f (new_AGEMA_signal_3508) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_0_XOR1_U1 ( .A0_t (SboxOut[0]), .A0_f (new_AGEMA_signal_11321), .A1_t (new_AGEMA_signal_11322), .A1_f (new_AGEMA_signal_11323), .B0_t (StateOutXORroundKey[0]), .B0_f (new_AGEMA_signal_3435), .B1_t (new_AGEMA_signal_3436), .B1_f (new_AGEMA_signal_3437), .Z0_t (MUX_StateIn_mux_inst_0_X), .Z0_f (new_AGEMA_signal_11324), .Z1_t (new_AGEMA_signal_11325), .Z1_f (new_AGEMA_signal_11326) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_0_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_6594), .B0_t (MUX_StateIn_mux_inst_0_X), .B0_f (new_AGEMA_signal_11324), .B1_t (new_AGEMA_signal_11325), .B1_f (new_AGEMA_signal_11326), .Z0_t (MUX_StateIn_mux_inst_0_Y), .Z0_f (new_AGEMA_signal_11351), .Z1_t (new_AGEMA_signal_11352), .Z1_f (new_AGEMA_signal_11353) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_0_XOR2_U1 ( .A0_t (MUX_StateIn_mux_inst_0_Y), .A0_f (new_AGEMA_signal_11351), .A1_t (new_AGEMA_signal_11352), .A1_f (new_AGEMA_signal_11353), .B0_t (SboxOut[0]), .B0_f (new_AGEMA_signal_11321), .B1_t (new_AGEMA_signal_11322), .B1_f (new_AGEMA_signal_11323), .Z0_t (StateIn[0]), .Z0_f (new_AGEMA_signal_11399), .Z1_t (new_AGEMA_signal_11400), .Z1_f (new_AGEMA_signal_11401) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_1_XOR1_U1 ( .A0_t (SboxOut[1]), .A0_f (new_AGEMA_signal_11348), .A1_t (new_AGEMA_signal_11349), .A1_f (new_AGEMA_signal_11350), .B0_t (StateOutXORroundKey[1]), .B0_f (new_AGEMA_signal_3444), .B1_t (new_AGEMA_signal_3445), .B1_f (new_AGEMA_signal_3446), .Z0_t (MUX_StateIn_mux_inst_1_X), .Z0_f (new_AGEMA_signal_11354), .Z1_t (new_AGEMA_signal_11355), .Z1_f (new_AGEMA_signal_11356) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_6594), .B0_t (MUX_StateIn_mux_inst_1_X), .B0_f (new_AGEMA_signal_11354), .B1_t (new_AGEMA_signal_11355), .B1_f (new_AGEMA_signal_11356), .Z0_t (MUX_StateIn_mux_inst_1_Y), .Z0_f (new_AGEMA_signal_11402), .Z1_t (new_AGEMA_signal_11403), .Z1_f (new_AGEMA_signal_11404) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_1_XOR2_U1 ( .A0_t (MUX_StateIn_mux_inst_1_Y), .A0_f (new_AGEMA_signal_11402), .A1_t (new_AGEMA_signal_11403), .A1_f (new_AGEMA_signal_11404), .B0_t (SboxOut[1]), .B0_f (new_AGEMA_signal_11348), .B1_t (new_AGEMA_signal_11349), .B1_f (new_AGEMA_signal_11350), .Z0_t (StateIn[1]), .Z0_f (new_AGEMA_signal_11447), .Z1_t (new_AGEMA_signal_11448), .Z1_f (new_AGEMA_signal_11449) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_2_XOR1_U1 ( .A0_t (SboxOut[2]), .A0_f (new_AGEMA_signal_11345), .A1_t (new_AGEMA_signal_11346), .A1_f (new_AGEMA_signal_11347), .B0_t (StateOutXORroundKey[2]), .B0_f (new_AGEMA_signal_3453), .B1_t (new_AGEMA_signal_3454), .B1_f (new_AGEMA_signal_3455), .Z0_t (MUX_StateIn_mux_inst_2_X), .Z0_f (new_AGEMA_signal_11357), .Z1_t (new_AGEMA_signal_11358), .Z1_f (new_AGEMA_signal_11359) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_2_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_6594), .B0_t (MUX_StateIn_mux_inst_2_X), .B0_f (new_AGEMA_signal_11357), .B1_t (new_AGEMA_signal_11358), .B1_f (new_AGEMA_signal_11359), .Z0_t (MUX_StateIn_mux_inst_2_Y), .Z0_f (new_AGEMA_signal_11405), .Z1_t (new_AGEMA_signal_11406), .Z1_f (new_AGEMA_signal_11407) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_2_XOR2_U1 ( .A0_t (MUX_StateIn_mux_inst_2_Y), .A0_f (new_AGEMA_signal_11405), .A1_t (new_AGEMA_signal_11406), .A1_f (new_AGEMA_signal_11407), .B0_t (SboxOut[2]), .B0_f (new_AGEMA_signal_11345), .B1_t (new_AGEMA_signal_11346), .B1_f (new_AGEMA_signal_11347), .Z0_t (StateIn[2]), .Z0_f (new_AGEMA_signal_11450), .Z1_t (new_AGEMA_signal_11451), .Z1_f (new_AGEMA_signal_11452) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_3_XOR1_U1 ( .A0_t (SboxOut[3]), .A0_f (new_AGEMA_signal_11342), .A1_t (new_AGEMA_signal_11343), .A1_f (new_AGEMA_signal_11344), .B0_t (StateOutXORroundKey[3]), .B0_f (new_AGEMA_signal_3462), .B1_t (new_AGEMA_signal_3463), .B1_f (new_AGEMA_signal_3464), .Z0_t (MUX_StateIn_mux_inst_3_X), .Z0_f (new_AGEMA_signal_11360), .Z1_t (new_AGEMA_signal_11361), .Z1_f (new_AGEMA_signal_11362) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_3_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_6594), .B0_t (MUX_StateIn_mux_inst_3_X), .B0_f (new_AGEMA_signal_11360), .B1_t (new_AGEMA_signal_11361), .B1_f (new_AGEMA_signal_11362), .Z0_t (MUX_StateIn_mux_inst_3_Y), .Z0_f (new_AGEMA_signal_11408), .Z1_t (new_AGEMA_signal_11409), .Z1_f (new_AGEMA_signal_11410) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_3_XOR2_U1 ( .A0_t (MUX_StateIn_mux_inst_3_Y), .A0_f (new_AGEMA_signal_11408), .A1_t (new_AGEMA_signal_11409), .A1_f (new_AGEMA_signal_11410), .B0_t (SboxOut[3]), .B0_f (new_AGEMA_signal_11342), .B1_t (new_AGEMA_signal_11343), .B1_f (new_AGEMA_signal_11344), .Z0_t (StateIn[3]), .Z0_f (new_AGEMA_signal_11453), .Z1_t (new_AGEMA_signal_11454), .Z1_f (new_AGEMA_signal_11455) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_4_XOR1_U1 ( .A0_t (SboxOut[4]), .A0_f (new_AGEMA_signal_11339), .A1_t (new_AGEMA_signal_11340), .A1_f (new_AGEMA_signal_11341), .B0_t (StateOutXORroundKey[4]), .B0_f (new_AGEMA_signal_3471), .B1_t (new_AGEMA_signal_3472), .B1_f (new_AGEMA_signal_3473), .Z0_t (MUX_StateIn_mux_inst_4_X), .Z0_f (new_AGEMA_signal_11363), .Z1_t (new_AGEMA_signal_11364), .Z1_f (new_AGEMA_signal_11365) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_4_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_6594), .B0_t (MUX_StateIn_mux_inst_4_X), .B0_f (new_AGEMA_signal_11363), .B1_t (new_AGEMA_signal_11364), .B1_f (new_AGEMA_signal_11365), .Z0_t (MUX_StateIn_mux_inst_4_Y), .Z0_f (new_AGEMA_signal_11411), .Z1_t (new_AGEMA_signal_11412), .Z1_f (new_AGEMA_signal_11413) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_4_XOR2_U1 ( .A0_t (MUX_StateIn_mux_inst_4_Y), .A0_f (new_AGEMA_signal_11411), .A1_t (new_AGEMA_signal_11412), .A1_f (new_AGEMA_signal_11413), .B0_t (SboxOut[4]), .B0_f (new_AGEMA_signal_11339), .B1_t (new_AGEMA_signal_11340), .B1_f (new_AGEMA_signal_11341), .Z0_t (StateIn[4]), .Z0_f (new_AGEMA_signal_11456), .Z1_t (new_AGEMA_signal_11457), .Z1_f (new_AGEMA_signal_11458) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_5_XOR1_U1 ( .A0_t (SboxOut[5]), .A0_f (new_AGEMA_signal_11336), .A1_t (new_AGEMA_signal_11337), .A1_f (new_AGEMA_signal_11338), .B0_t (StateOutXORroundKey[5]), .B0_f (new_AGEMA_signal_3480), .B1_t (new_AGEMA_signal_3481), .B1_f (new_AGEMA_signal_3482), .Z0_t (MUX_StateIn_mux_inst_5_X), .Z0_f (new_AGEMA_signal_11366), .Z1_t (new_AGEMA_signal_11367), .Z1_f (new_AGEMA_signal_11368) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_5_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_6594), .B0_t (MUX_StateIn_mux_inst_5_X), .B0_f (new_AGEMA_signal_11366), .B1_t (new_AGEMA_signal_11367), .B1_f (new_AGEMA_signal_11368), .Z0_t (MUX_StateIn_mux_inst_5_Y), .Z0_f (new_AGEMA_signal_11414), .Z1_t (new_AGEMA_signal_11415), .Z1_f (new_AGEMA_signal_11416) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_5_XOR2_U1 ( .A0_t (MUX_StateIn_mux_inst_5_Y), .A0_f (new_AGEMA_signal_11414), .A1_t (new_AGEMA_signal_11415), .A1_f (new_AGEMA_signal_11416), .B0_t (SboxOut[5]), .B0_f (new_AGEMA_signal_11336), .B1_t (new_AGEMA_signal_11337), .B1_f (new_AGEMA_signal_11338), .Z0_t (StateIn[5]), .Z0_f (new_AGEMA_signal_11459), .Z1_t (new_AGEMA_signal_11460), .Z1_f (new_AGEMA_signal_11461) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_6_XOR1_U1 ( .A0_t (SboxOut[6]), .A0_f (new_AGEMA_signal_11333), .A1_t (new_AGEMA_signal_11334), .A1_f (new_AGEMA_signal_11335), .B0_t (StateOutXORroundKey[6]), .B0_f (new_AGEMA_signal_3489), .B1_t (new_AGEMA_signal_3490), .B1_f (new_AGEMA_signal_3491), .Z0_t (MUX_StateIn_mux_inst_6_X), .Z0_f (new_AGEMA_signal_11369), .Z1_t (new_AGEMA_signal_11370), .Z1_f (new_AGEMA_signal_11371) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_6_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_6594), .B0_t (MUX_StateIn_mux_inst_6_X), .B0_f (new_AGEMA_signal_11369), .B1_t (new_AGEMA_signal_11370), .B1_f (new_AGEMA_signal_11371), .Z0_t (MUX_StateIn_mux_inst_6_Y), .Z0_f (new_AGEMA_signal_11417), .Z1_t (new_AGEMA_signal_11418), .Z1_f (new_AGEMA_signal_11419) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_6_XOR2_U1 ( .A0_t (MUX_StateIn_mux_inst_6_Y), .A0_f (new_AGEMA_signal_11417), .A1_t (new_AGEMA_signal_11418), .A1_f (new_AGEMA_signal_11419), .B0_t (SboxOut[6]), .B0_f (new_AGEMA_signal_11333), .B1_t (new_AGEMA_signal_11334), .B1_f (new_AGEMA_signal_11335), .Z0_t (StateIn[6]), .Z0_f (new_AGEMA_signal_11462), .Z1_t (new_AGEMA_signal_11463), .Z1_f (new_AGEMA_signal_11464) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_7_XOR1_U1 ( .A0_t (SboxOut[7]), .A0_f (new_AGEMA_signal_11330), .A1_t (new_AGEMA_signal_11331), .A1_f (new_AGEMA_signal_11332), .B0_t (StateOutXORroundKey[7]), .B0_f (new_AGEMA_signal_3498), .B1_t (new_AGEMA_signal_3499), .B1_f (new_AGEMA_signal_3500), .Z0_t (MUX_StateIn_mux_inst_7_X), .Z0_f (new_AGEMA_signal_11372), .Z1_t (new_AGEMA_signal_11373), .Z1_f (new_AGEMA_signal_11374) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_7_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_6594), .B0_t (MUX_StateIn_mux_inst_7_X), .B0_f (new_AGEMA_signal_11372), .B1_t (new_AGEMA_signal_11373), .B1_f (new_AGEMA_signal_11374), .Z0_t (MUX_StateIn_mux_inst_7_Y), .Z0_f (new_AGEMA_signal_11420), .Z1_t (new_AGEMA_signal_11421), .Z1_f (new_AGEMA_signal_11422) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_7_XOR2_U1 ( .A0_t (MUX_StateIn_mux_inst_7_Y), .A0_f (new_AGEMA_signal_11420), .A1_t (new_AGEMA_signal_11421), .A1_f (new_AGEMA_signal_11422), .B0_t (SboxOut[7]), .B0_f (new_AGEMA_signal_11330), .B1_t (new_AGEMA_signal_11331), .B1_f (new_AGEMA_signal_11332), .Z0_t (StateIn[7]), .Z0_f (new_AGEMA_signal_11465), .Z1_t (new_AGEMA_signal_11466), .Z1_f (new_AGEMA_signal_11467) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S00reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS00ser[0]), .A0_f (new_AGEMA_signal_6622), .A1_t (new_AGEMA_signal_6623), .A1_f (new_AGEMA_signal_6624), .B0_t (ciphertext_s0_t[120]), .B0_f (ciphertext_s0_f[120]), .B1_t (ciphertext_s1_t[120]), .B1_f (ciphertext_s1_f[120]), .Z0_t (stateArray_S00reg_gff_1_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_7395), .Z1_t (new_AGEMA_signal_7396), .Z1_f (new_AGEMA_signal_7397) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S00reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S00reg_gff_1_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_7395), .B1_t (new_AGEMA_signal_7396), .B1_f (new_AGEMA_signal_7397), .Z0_t (stateArray_S00reg_gff_1_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_8142), .Z1_t (new_AGEMA_signal_8143), .Z1_f (new_AGEMA_signal_8144) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S00reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (stateArray_S00reg_gff_1_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_8142), .A1_t (new_AGEMA_signal_8143), .A1_f (new_AGEMA_signal_8144), .B0_t (stateArray_inS00ser[0]), .B0_f (new_AGEMA_signal_6622), .B1_t (new_AGEMA_signal_6623), .B1_f (new_AGEMA_signal_6624), .Z0_t (ciphertext_s0_t[120]), .Z0_f (ciphertext_s0_f[120]), .Z1_t (ciphertext_s1_t[120]), .Z1_f (ciphertext_s1_f[120]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S00reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS00ser[1]), .A0_f (new_AGEMA_signal_6625), .A1_t (new_AGEMA_signal_6626), .A1_f (new_AGEMA_signal_6627), .B0_t (ciphertext_s0_t[121]), .B0_f (ciphertext_s0_f[121]), .B1_t (ciphertext_s1_t[121]), .B1_f (ciphertext_s1_f[121]), .Z0_t (stateArray_S00reg_gff_1_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_7398), .Z1_t (new_AGEMA_signal_7399), .Z1_f (new_AGEMA_signal_7400) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S00reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S00reg_gff_1_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_7398), .B1_t (new_AGEMA_signal_7399), .B1_f (new_AGEMA_signal_7400), .Z0_t (stateArray_S00reg_gff_1_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_8145), .Z1_t (new_AGEMA_signal_8146), .Z1_f (new_AGEMA_signal_8147) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S00reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (stateArray_S00reg_gff_1_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_8145), .A1_t (new_AGEMA_signal_8146), .A1_f (new_AGEMA_signal_8147), .B0_t (stateArray_inS00ser[1]), .B0_f (new_AGEMA_signal_6625), .B1_t (new_AGEMA_signal_6626), .B1_f (new_AGEMA_signal_6627), .Z0_t (ciphertext_s0_t[121]), .Z0_f (ciphertext_s0_f[121]), .Z1_t (ciphertext_s1_t[121]), .Z1_f (ciphertext_s1_f[121]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S00reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS00ser[2]), .A0_f (new_AGEMA_signal_6628), .A1_t (new_AGEMA_signal_6629), .A1_f (new_AGEMA_signal_6630), .B0_t (ciphertext_s0_t[122]), .B0_f (ciphertext_s0_f[122]), .B1_t (ciphertext_s1_t[122]), .B1_f (ciphertext_s1_f[122]), .Z0_t (stateArray_S00reg_gff_1_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_7401), .Z1_t (new_AGEMA_signal_7402), .Z1_f (new_AGEMA_signal_7403) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S00reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S00reg_gff_1_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_7401), .B1_t (new_AGEMA_signal_7402), .B1_f (new_AGEMA_signal_7403), .Z0_t (stateArray_S00reg_gff_1_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_8148), .Z1_t (new_AGEMA_signal_8149), .Z1_f (new_AGEMA_signal_8150) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S00reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (stateArray_S00reg_gff_1_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_8148), .A1_t (new_AGEMA_signal_8149), .A1_f (new_AGEMA_signal_8150), .B0_t (stateArray_inS00ser[2]), .B0_f (new_AGEMA_signal_6628), .B1_t (new_AGEMA_signal_6629), .B1_f (new_AGEMA_signal_6630), .Z0_t (ciphertext_s0_t[122]), .Z0_f (ciphertext_s0_f[122]), .Z1_t (ciphertext_s1_t[122]), .Z1_f (ciphertext_s1_f[122]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S00reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS00ser[3]), .A0_f (new_AGEMA_signal_6631), .A1_t (new_AGEMA_signal_6632), .A1_f (new_AGEMA_signal_6633), .B0_t (ciphertext_s0_t[123]), .B0_f (ciphertext_s0_f[123]), .B1_t (ciphertext_s1_t[123]), .B1_f (ciphertext_s1_f[123]), .Z0_t (stateArray_S00reg_gff_1_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_7404), .Z1_t (new_AGEMA_signal_7405), .Z1_f (new_AGEMA_signal_7406) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S00reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S00reg_gff_1_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_7404), .B1_t (new_AGEMA_signal_7405), .B1_f (new_AGEMA_signal_7406), .Z0_t (stateArray_S00reg_gff_1_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_8151), .Z1_t (new_AGEMA_signal_8152), .Z1_f (new_AGEMA_signal_8153) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S00reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (stateArray_S00reg_gff_1_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_8151), .A1_t (new_AGEMA_signal_8152), .A1_f (new_AGEMA_signal_8153), .B0_t (stateArray_inS00ser[3]), .B0_f (new_AGEMA_signal_6631), .B1_t (new_AGEMA_signal_6632), .B1_f (new_AGEMA_signal_6633), .Z0_t (ciphertext_s0_t[123]), .Z0_f (ciphertext_s0_f[123]), .Z1_t (ciphertext_s1_t[123]), .Z1_f (ciphertext_s1_f[123]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S00reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS00ser[4]), .A0_f (new_AGEMA_signal_6634), .A1_t (new_AGEMA_signal_6635), .A1_f (new_AGEMA_signal_6636), .B0_t (ciphertext_s0_t[124]), .B0_f (ciphertext_s0_f[124]), .B1_t (ciphertext_s1_t[124]), .B1_f (ciphertext_s1_f[124]), .Z0_t (stateArray_S00reg_gff_1_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_7407), .Z1_t (new_AGEMA_signal_7408), .Z1_f (new_AGEMA_signal_7409) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S00reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S00reg_gff_1_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_7407), .B1_t (new_AGEMA_signal_7408), .B1_f (new_AGEMA_signal_7409), .Z0_t (stateArray_S00reg_gff_1_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_8154), .Z1_t (new_AGEMA_signal_8155), .Z1_f (new_AGEMA_signal_8156) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S00reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (stateArray_S00reg_gff_1_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_8154), .A1_t (new_AGEMA_signal_8155), .A1_f (new_AGEMA_signal_8156), .B0_t (stateArray_inS00ser[4]), .B0_f (new_AGEMA_signal_6634), .B1_t (new_AGEMA_signal_6635), .B1_f (new_AGEMA_signal_6636), .Z0_t (ciphertext_s0_t[124]), .Z0_f (ciphertext_s0_f[124]), .Z1_t (ciphertext_s1_t[124]), .Z1_f (ciphertext_s1_f[124]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S00reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS00ser[5]), .A0_f (new_AGEMA_signal_6637), .A1_t (new_AGEMA_signal_6638), .A1_f (new_AGEMA_signal_6639), .B0_t (ciphertext_s0_t[125]), .B0_f (ciphertext_s0_f[125]), .B1_t (ciphertext_s1_t[125]), .B1_f (ciphertext_s1_f[125]), .Z0_t (stateArray_S00reg_gff_1_SFF_5_MUXInst_X), .Z0_f (new_AGEMA_signal_7410), .Z1_t (new_AGEMA_signal_7411), .Z1_f (new_AGEMA_signal_7412) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S00reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S00reg_gff_1_SFF_5_MUXInst_X), .B0_f (new_AGEMA_signal_7410), .B1_t (new_AGEMA_signal_7411), .B1_f (new_AGEMA_signal_7412), .Z0_t (stateArray_S00reg_gff_1_SFF_5_MUXInst_Y), .Z0_f (new_AGEMA_signal_8157), .Z1_t (new_AGEMA_signal_8158), .Z1_f (new_AGEMA_signal_8159) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S00reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (stateArray_S00reg_gff_1_SFF_5_MUXInst_Y), .A0_f (new_AGEMA_signal_8157), .A1_t (new_AGEMA_signal_8158), .A1_f (new_AGEMA_signal_8159), .B0_t (stateArray_inS00ser[5]), .B0_f (new_AGEMA_signal_6637), .B1_t (new_AGEMA_signal_6638), .B1_f (new_AGEMA_signal_6639), .Z0_t (ciphertext_s0_t[125]), .Z0_f (ciphertext_s0_f[125]), .Z1_t (ciphertext_s1_t[125]), .Z1_f (ciphertext_s1_f[125]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S00reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS00ser[6]), .A0_f (new_AGEMA_signal_6640), .A1_t (new_AGEMA_signal_6641), .A1_f (new_AGEMA_signal_6642), .B0_t (ciphertext_s0_t[126]), .B0_f (ciphertext_s0_f[126]), .B1_t (ciphertext_s1_t[126]), .B1_f (ciphertext_s1_f[126]), .Z0_t (stateArray_S00reg_gff_1_SFF_6_MUXInst_X), .Z0_f (new_AGEMA_signal_7413), .Z1_t (new_AGEMA_signal_7414), .Z1_f (new_AGEMA_signal_7415) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S00reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S00reg_gff_1_SFF_6_MUXInst_X), .B0_f (new_AGEMA_signal_7413), .B1_t (new_AGEMA_signal_7414), .B1_f (new_AGEMA_signal_7415), .Z0_t (stateArray_S00reg_gff_1_SFF_6_MUXInst_Y), .Z0_f (new_AGEMA_signal_8160), .Z1_t (new_AGEMA_signal_8161), .Z1_f (new_AGEMA_signal_8162) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S00reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (stateArray_S00reg_gff_1_SFF_6_MUXInst_Y), .A0_f (new_AGEMA_signal_8160), .A1_t (new_AGEMA_signal_8161), .A1_f (new_AGEMA_signal_8162), .B0_t (stateArray_inS00ser[6]), .B0_f (new_AGEMA_signal_6640), .B1_t (new_AGEMA_signal_6641), .B1_f (new_AGEMA_signal_6642), .Z0_t (ciphertext_s0_t[126]), .Z0_f (ciphertext_s0_f[126]), .Z1_t (ciphertext_s1_t[126]), .Z1_f (ciphertext_s1_f[126]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S00reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS00ser[7]), .A0_f (new_AGEMA_signal_6643), .A1_t (new_AGEMA_signal_6644), .A1_f (new_AGEMA_signal_6645), .B0_t (ciphertext_s0_t[127]), .B0_f (ciphertext_s0_f[127]), .B1_t (ciphertext_s1_t[127]), .B1_f (ciphertext_s1_f[127]), .Z0_t (stateArray_S00reg_gff_1_SFF_7_MUXInst_X), .Z0_f (new_AGEMA_signal_7416), .Z1_t (new_AGEMA_signal_7417), .Z1_f (new_AGEMA_signal_7418) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S00reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S00reg_gff_1_SFF_7_MUXInst_X), .B0_f (new_AGEMA_signal_7416), .B1_t (new_AGEMA_signal_7417), .B1_f (new_AGEMA_signal_7418), .Z0_t (stateArray_S00reg_gff_1_SFF_7_MUXInst_Y), .Z0_f (new_AGEMA_signal_8163), .Z1_t (new_AGEMA_signal_8164), .Z1_f (new_AGEMA_signal_8165) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S00reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (stateArray_S00reg_gff_1_SFF_7_MUXInst_Y), .A0_f (new_AGEMA_signal_8163), .A1_t (new_AGEMA_signal_8164), .A1_f (new_AGEMA_signal_8165), .B0_t (stateArray_inS00ser[7]), .B0_f (new_AGEMA_signal_6643), .B1_t (new_AGEMA_signal_6644), .B1_f (new_AGEMA_signal_6645), .Z0_t (ciphertext_s0_t[127]), .Z0_f (ciphertext_s0_f[127]), .Z1_t (ciphertext_s1_t[127]), .Z1_f (ciphertext_s1_f[127]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S01reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS01ser[0]), .A0_f (new_AGEMA_signal_6646), .A1_t (new_AGEMA_signal_6647), .A1_f (new_AGEMA_signal_6648), .B0_t (ciphertext_s0_t[88]), .B0_f (ciphertext_s0_f[88]), .B1_t (ciphertext_s1_t[88]), .B1_f (ciphertext_s1_f[88]), .Z0_t (stateArray_S01reg_gff_1_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_7419), .Z1_t (new_AGEMA_signal_7420), .Z1_f (new_AGEMA_signal_7421) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S01reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S01reg_gff_1_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_7419), .B1_t (new_AGEMA_signal_7420), .B1_f (new_AGEMA_signal_7421), .Z0_t (stateArray_S01reg_gff_1_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_8166), .Z1_t (new_AGEMA_signal_8167), .Z1_f (new_AGEMA_signal_8168) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S01reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (stateArray_S01reg_gff_1_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_8166), .A1_t (new_AGEMA_signal_8167), .A1_f (new_AGEMA_signal_8168), .B0_t (stateArray_inS01ser[0]), .B0_f (new_AGEMA_signal_6646), .B1_t (new_AGEMA_signal_6647), .B1_f (new_AGEMA_signal_6648), .Z0_t (ciphertext_s0_t[88]), .Z0_f (ciphertext_s0_f[88]), .Z1_t (ciphertext_s1_t[88]), .Z1_f (ciphertext_s1_f[88]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S01reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS01ser[1]), .A0_f (new_AGEMA_signal_6649), .A1_t (new_AGEMA_signal_6650), .A1_f (new_AGEMA_signal_6651), .B0_t (ciphertext_s0_t[89]), .B0_f (ciphertext_s0_f[89]), .B1_t (ciphertext_s1_t[89]), .B1_f (ciphertext_s1_f[89]), .Z0_t (stateArray_S01reg_gff_1_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_7422), .Z1_t (new_AGEMA_signal_7423), .Z1_f (new_AGEMA_signal_7424) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S01reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S01reg_gff_1_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_7422), .B1_t (new_AGEMA_signal_7423), .B1_f (new_AGEMA_signal_7424), .Z0_t (stateArray_S01reg_gff_1_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_8169), .Z1_t (new_AGEMA_signal_8170), .Z1_f (new_AGEMA_signal_8171) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S01reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (stateArray_S01reg_gff_1_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_8169), .A1_t (new_AGEMA_signal_8170), .A1_f (new_AGEMA_signal_8171), .B0_t (stateArray_inS01ser[1]), .B0_f (new_AGEMA_signal_6649), .B1_t (new_AGEMA_signal_6650), .B1_f (new_AGEMA_signal_6651), .Z0_t (ciphertext_s0_t[89]), .Z0_f (ciphertext_s0_f[89]), .Z1_t (ciphertext_s1_t[89]), .Z1_f (ciphertext_s1_f[89]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S01reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS01ser[2]), .A0_f (new_AGEMA_signal_6652), .A1_t (new_AGEMA_signal_6653), .A1_f (new_AGEMA_signal_6654), .B0_t (ciphertext_s0_t[90]), .B0_f (ciphertext_s0_f[90]), .B1_t (ciphertext_s1_t[90]), .B1_f (ciphertext_s1_f[90]), .Z0_t (stateArray_S01reg_gff_1_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_7425), .Z1_t (new_AGEMA_signal_7426), .Z1_f (new_AGEMA_signal_7427) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S01reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S01reg_gff_1_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_7425), .B1_t (new_AGEMA_signal_7426), .B1_f (new_AGEMA_signal_7427), .Z0_t (stateArray_S01reg_gff_1_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_8172), .Z1_t (new_AGEMA_signal_8173), .Z1_f (new_AGEMA_signal_8174) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S01reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (stateArray_S01reg_gff_1_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_8172), .A1_t (new_AGEMA_signal_8173), .A1_f (new_AGEMA_signal_8174), .B0_t (stateArray_inS01ser[2]), .B0_f (new_AGEMA_signal_6652), .B1_t (new_AGEMA_signal_6653), .B1_f (new_AGEMA_signal_6654), .Z0_t (ciphertext_s0_t[90]), .Z0_f (ciphertext_s0_f[90]), .Z1_t (ciphertext_s1_t[90]), .Z1_f (ciphertext_s1_f[90]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S01reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS01ser[3]), .A0_f (new_AGEMA_signal_6655), .A1_t (new_AGEMA_signal_6656), .A1_f (new_AGEMA_signal_6657), .B0_t (ciphertext_s0_t[91]), .B0_f (ciphertext_s0_f[91]), .B1_t (ciphertext_s1_t[91]), .B1_f (ciphertext_s1_f[91]), .Z0_t (stateArray_S01reg_gff_1_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_7428), .Z1_t (new_AGEMA_signal_7429), .Z1_f (new_AGEMA_signal_7430) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S01reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S01reg_gff_1_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_7428), .B1_t (new_AGEMA_signal_7429), .B1_f (new_AGEMA_signal_7430), .Z0_t (stateArray_S01reg_gff_1_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_8175), .Z1_t (new_AGEMA_signal_8176), .Z1_f (new_AGEMA_signal_8177) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S01reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (stateArray_S01reg_gff_1_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_8175), .A1_t (new_AGEMA_signal_8176), .A1_f (new_AGEMA_signal_8177), .B0_t (stateArray_inS01ser[3]), .B0_f (new_AGEMA_signal_6655), .B1_t (new_AGEMA_signal_6656), .B1_f (new_AGEMA_signal_6657), .Z0_t (ciphertext_s0_t[91]), .Z0_f (ciphertext_s0_f[91]), .Z1_t (ciphertext_s1_t[91]), .Z1_f (ciphertext_s1_f[91]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S01reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS01ser[4]), .A0_f (new_AGEMA_signal_6658), .A1_t (new_AGEMA_signal_6659), .A1_f (new_AGEMA_signal_6660), .B0_t (ciphertext_s0_t[92]), .B0_f (ciphertext_s0_f[92]), .B1_t (ciphertext_s1_t[92]), .B1_f (ciphertext_s1_f[92]), .Z0_t (stateArray_S01reg_gff_1_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_7431), .Z1_t (new_AGEMA_signal_7432), .Z1_f (new_AGEMA_signal_7433) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S01reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S01reg_gff_1_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_7431), .B1_t (new_AGEMA_signal_7432), .B1_f (new_AGEMA_signal_7433), .Z0_t (stateArray_S01reg_gff_1_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_8178), .Z1_t (new_AGEMA_signal_8179), .Z1_f (new_AGEMA_signal_8180) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S01reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (stateArray_S01reg_gff_1_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_8178), .A1_t (new_AGEMA_signal_8179), .A1_f (new_AGEMA_signal_8180), .B0_t (stateArray_inS01ser[4]), .B0_f (new_AGEMA_signal_6658), .B1_t (new_AGEMA_signal_6659), .B1_f (new_AGEMA_signal_6660), .Z0_t (ciphertext_s0_t[92]), .Z0_f (ciphertext_s0_f[92]), .Z1_t (ciphertext_s1_t[92]), .Z1_f (ciphertext_s1_f[92]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S01reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS01ser[5]), .A0_f (new_AGEMA_signal_6661), .A1_t (new_AGEMA_signal_6662), .A1_f (new_AGEMA_signal_6663), .B0_t (ciphertext_s0_t[93]), .B0_f (ciphertext_s0_f[93]), .B1_t (ciphertext_s1_t[93]), .B1_f (ciphertext_s1_f[93]), .Z0_t (stateArray_S01reg_gff_1_SFF_5_MUXInst_X), .Z0_f (new_AGEMA_signal_7434), .Z1_t (new_AGEMA_signal_7435), .Z1_f (new_AGEMA_signal_7436) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S01reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S01reg_gff_1_SFF_5_MUXInst_X), .B0_f (new_AGEMA_signal_7434), .B1_t (new_AGEMA_signal_7435), .B1_f (new_AGEMA_signal_7436), .Z0_t (stateArray_S01reg_gff_1_SFF_5_MUXInst_Y), .Z0_f (new_AGEMA_signal_8181), .Z1_t (new_AGEMA_signal_8182), .Z1_f (new_AGEMA_signal_8183) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S01reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (stateArray_S01reg_gff_1_SFF_5_MUXInst_Y), .A0_f (new_AGEMA_signal_8181), .A1_t (new_AGEMA_signal_8182), .A1_f (new_AGEMA_signal_8183), .B0_t (stateArray_inS01ser[5]), .B0_f (new_AGEMA_signal_6661), .B1_t (new_AGEMA_signal_6662), .B1_f (new_AGEMA_signal_6663), .Z0_t (ciphertext_s0_t[93]), .Z0_f (ciphertext_s0_f[93]), .Z1_t (ciphertext_s1_t[93]), .Z1_f (ciphertext_s1_f[93]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S01reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS01ser[6]), .A0_f (new_AGEMA_signal_6664), .A1_t (new_AGEMA_signal_6665), .A1_f (new_AGEMA_signal_6666), .B0_t (ciphertext_s0_t[94]), .B0_f (ciphertext_s0_f[94]), .B1_t (ciphertext_s1_t[94]), .B1_f (ciphertext_s1_f[94]), .Z0_t (stateArray_S01reg_gff_1_SFF_6_MUXInst_X), .Z0_f (new_AGEMA_signal_7437), .Z1_t (new_AGEMA_signal_7438), .Z1_f (new_AGEMA_signal_7439) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S01reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S01reg_gff_1_SFF_6_MUXInst_X), .B0_f (new_AGEMA_signal_7437), .B1_t (new_AGEMA_signal_7438), .B1_f (new_AGEMA_signal_7439), .Z0_t (stateArray_S01reg_gff_1_SFF_6_MUXInst_Y), .Z0_f (new_AGEMA_signal_8184), .Z1_t (new_AGEMA_signal_8185), .Z1_f (new_AGEMA_signal_8186) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S01reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (stateArray_S01reg_gff_1_SFF_6_MUXInst_Y), .A0_f (new_AGEMA_signal_8184), .A1_t (new_AGEMA_signal_8185), .A1_f (new_AGEMA_signal_8186), .B0_t (stateArray_inS01ser[6]), .B0_f (new_AGEMA_signal_6664), .B1_t (new_AGEMA_signal_6665), .B1_f (new_AGEMA_signal_6666), .Z0_t (ciphertext_s0_t[94]), .Z0_f (ciphertext_s0_f[94]), .Z1_t (ciphertext_s1_t[94]), .Z1_f (ciphertext_s1_f[94]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S01reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS01ser[7]), .A0_f (new_AGEMA_signal_6667), .A1_t (new_AGEMA_signal_6668), .A1_f (new_AGEMA_signal_6669), .B0_t (ciphertext_s0_t[95]), .B0_f (ciphertext_s0_f[95]), .B1_t (ciphertext_s1_t[95]), .B1_f (ciphertext_s1_f[95]), .Z0_t (stateArray_S01reg_gff_1_SFF_7_MUXInst_X), .Z0_f (new_AGEMA_signal_7440), .Z1_t (new_AGEMA_signal_7441), .Z1_f (new_AGEMA_signal_7442) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S01reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S01reg_gff_1_SFF_7_MUXInst_X), .B0_f (new_AGEMA_signal_7440), .B1_t (new_AGEMA_signal_7441), .B1_f (new_AGEMA_signal_7442), .Z0_t (stateArray_S01reg_gff_1_SFF_7_MUXInst_Y), .Z0_f (new_AGEMA_signal_8187), .Z1_t (new_AGEMA_signal_8188), .Z1_f (new_AGEMA_signal_8189) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S01reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (stateArray_S01reg_gff_1_SFF_7_MUXInst_Y), .A0_f (new_AGEMA_signal_8187), .A1_t (new_AGEMA_signal_8188), .A1_f (new_AGEMA_signal_8189), .B0_t (stateArray_inS01ser[7]), .B0_f (new_AGEMA_signal_6667), .B1_t (new_AGEMA_signal_6668), .B1_f (new_AGEMA_signal_6669), .Z0_t (ciphertext_s0_t[95]), .Z0_f (ciphertext_s0_f[95]), .Z1_t (ciphertext_s1_t[95]), .Z1_f (ciphertext_s1_f[95]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S02reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS02ser[0]), .A0_f (new_AGEMA_signal_6670), .A1_t (new_AGEMA_signal_6671), .A1_f (new_AGEMA_signal_6672), .B0_t (ciphertext_s0_t[56]), .B0_f (ciphertext_s0_f[56]), .B1_t (ciphertext_s1_t[56]), .B1_f (ciphertext_s1_f[56]), .Z0_t (stateArray_S02reg_gff_1_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_7443), .Z1_t (new_AGEMA_signal_7444), .Z1_f (new_AGEMA_signal_7445) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S02reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S02reg_gff_1_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_7443), .B1_t (new_AGEMA_signal_7444), .B1_f (new_AGEMA_signal_7445), .Z0_t (stateArray_S02reg_gff_1_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_8190), .Z1_t (new_AGEMA_signal_8191), .Z1_f (new_AGEMA_signal_8192) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S02reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (stateArray_S02reg_gff_1_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_8190), .A1_t (new_AGEMA_signal_8191), .A1_f (new_AGEMA_signal_8192), .B0_t (stateArray_inS02ser[0]), .B0_f (new_AGEMA_signal_6670), .B1_t (new_AGEMA_signal_6671), .B1_f (new_AGEMA_signal_6672), .Z0_t (ciphertext_s0_t[56]), .Z0_f (ciphertext_s0_f[56]), .Z1_t (ciphertext_s1_t[56]), .Z1_f (ciphertext_s1_f[56]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S02reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS02ser[1]), .A0_f (new_AGEMA_signal_6673), .A1_t (new_AGEMA_signal_6674), .A1_f (new_AGEMA_signal_6675), .B0_t (ciphertext_s0_t[57]), .B0_f (ciphertext_s0_f[57]), .B1_t (ciphertext_s1_t[57]), .B1_f (ciphertext_s1_f[57]), .Z0_t (stateArray_S02reg_gff_1_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_7446), .Z1_t (new_AGEMA_signal_7447), .Z1_f (new_AGEMA_signal_7448) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S02reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S02reg_gff_1_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_7446), .B1_t (new_AGEMA_signal_7447), .B1_f (new_AGEMA_signal_7448), .Z0_t (stateArray_S02reg_gff_1_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_8193), .Z1_t (new_AGEMA_signal_8194), .Z1_f (new_AGEMA_signal_8195) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S02reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (stateArray_S02reg_gff_1_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_8193), .A1_t (new_AGEMA_signal_8194), .A1_f (new_AGEMA_signal_8195), .B0_t (stateArray_inS02ser[1]), .B0_f (new_AGEMA_signal_6673), .B1_t (new_AGEMA_signal_6674), .B1_f (new_AGEMA_signal_6675), .Z0_t (ciphertext_s0_t[57]), .Z0_f (ciphertext_s0_f[57]), .Z1_t (ciphertext_s1_t[57]), .Z1_f (ciphertext_s1_f[57]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S02reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS02ser[2]), .A0_f (new_AGEMA_signal_6676), .A1_t (new_AGEMA_signal_6677), .A1_f (new_AGEMA_signal_6678), .B0_t (ciphertext_s0_t[58]), .B0_f (ciphertext_s0_f[58]), .B1_t (ciphertext_s1_t[58]), .B1_f (ciphertext_s1_f[58]), .Z0_t (stateArray_S02reg_gff_1_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_7449), .Z1_t (new_AGEMA_signal_7450), .Z1_f (new_AGEMA_signal_7451) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S02reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S02reg_gff_1_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_7449), .B1_t (new_AGEMA_signal_7450), .B1_f (new_AGEMA_signal_7451), .Z0_t (stateArray_S02reg_gff_1_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_8196), .Z1_t (new_AGEMA_signal_8197), .Z1_f (new_AGEMA_signal_8198) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S02reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (stateArray_S02reg_gff_1_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_8196), .A1_t (new_AGEMA_signal_8197), .A1_f (new_AGEMA_signal_8198), .B0_t (stateArray_inS02ser[2]), .B0_f (new_AGEMA_signal_6676), .B1_t (new_AGEMA_signal_6677), .B1_f (new_AGEMA_signal_6678), .Z0_t (ciphertext_s0_t[58]), .Z0_f (ciphertext_s0_f[58]), .Z1_t (ciphertext_s1_t[58]), .Z1_f (ciphertext_s1_f[58]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S02reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS02ser[3]), .A0_f (new_AGEMA_signal_6679), .A1_t (new_AGEMA_signal_6680), .A1_f (new_AGEMA_signal_6681), .B0_t (ciphertext_s0_t[59]), .B0_f (ciphertext_s0_f[59]), .B1_t (ciphertext_s1_t[59]), .B1_f (ciphertext_s1_f[59]), .Z0_t (stateArray_S02reg_gff_1_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_7452), .Z1_t (new_AGEMA_signal_7453), .Z1_f (new_AGEMA_signal_7454) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S02reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S02reg_gff_1_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_7452), .B1_t (new_AGEMA_signal_7453), .B1_f (new_AGEMA_signal_7454), .Z0_t (stateArray_S02reg_gff_1_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_8199), .Z1_t (new_AGEMA_signal_8200), .Z1_f (new_AGEMA_signal_8201) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S02reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (stateArray_S02reg_gff_1_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_8199), .A1_t (new_AGEMA_signal_8200), .A1_f (new_AGEMA_signal_8201), .B0_t (stateArray_inS02ser[3]), .B0_f (new_AGEMA_signal_6679), .B1_t (new_AGEMA_signal_6680), .B1_f (new_AGEMA_signal_6681), .Z0_t (ciphertext_s0_t[59]), .Z0_f (ciphertext_s0_f[59]), .Z1_t (ciphertext_s1_t[59]), .Z1_f (ciphertext_s1_f[59]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S02reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS02ser[4]), .A0_f (new_AGEMA_signal_6682), .A1_t (new_AGEMA_signal_6683), .A1_f (new_AGEMA_signal_6684), .B0_t (ciphertext_s0_t[60]), .B0_f (ciphertext_s0_f[60]), .B1_t (ciphertext_s1_t[60]), .B1_f (ciphertext_s1_f[60]), .Z0_t (stateArray_S02reg_gff_1_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_7455), .Z1_t (new_AGEMA_signal_7456), .Z1_f (new_AGEMA_signal_7457) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S02reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S02reg_gff_1_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_7455), .B1_t (new_AGEMA_signal_7456), .B1_f (new_AGEMA_signal_7457), .Z0_t (stateArray_S02reg_gff_1_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_8202), .Z1_t (new_AGEMA_signal_8203), .Z1_f (new_AGEMA_signal_8204) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S02reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (stateArray_S02reg_gff_1_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_8202), .A1_t (new_AGEMA_signal_8203), .A1_f (new_AGEMA_signal_8204), .B0_t (stateArray_inS02ser[4]), .B0_f (new_AGEMA_signal_6682), .B1_t (new_AGEMA_signal_6683), .B1_f (new_AGEMA_signal_6684), .Z0_t (ciphertext_s0_t[60]), .Z0_f (ciphertext_s0_f[60]), .Z1_t (ciphertext_s1_t[60]), .Z1_f (ciphertext_s1_f[60]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S02reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS02ser[5]), .A0_f (new_AGEMA_signal_6685), .A1_t (new_AGEMA_signal_6686), .A1_f (new_AGEMA_signal_6687), .B0_t (ciphertext_s0_t[61]), .B0_f (ciphertext_s0_f[61]), .B1_t (ciphertext_s1_t[61]), .B1_f (ciphertext_s1_f[61]), .Z0_t (stateArray_S02reg_gff_1_SFF_5_MUXInst_X), .Z0_f (new_AGEMA_signal_7458), .Z1_t (new_AGEMA_signal_7459), .Z1_f (new_AGEMA_signal_7460) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S02reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S02reg_gff_1_SFF_5_MUXInst_X), .B0_f (new_AGEMA_signal_7458), .B1_t (new_AGEMA_signal_7459), .B1_f (new_AGEMA_signal_7460), .Z0_t (stateArray_S02reg_gff_1_SFF_5_MUXInst_Y), .Z0_f (new_AGEMA_signal_8205), .Z1_t (new_AGEMA_signal_8206), .Z1_f (new_AGEMA_signal_8207) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S02reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (stateArray_S02reg_gff_1_SFF_5_MUXInst_Y), .A0_f (new_AGEMA_signal_8205), .A1_t (new_AGEMA_signal_8206), .A1_f (new_AGEMA_signal_8207), .B0_t (stateArray_inS02ser[5]), .B0_f (new_AGEMA_signal_6685), .B1_t (new_AGEMA_signal_6686), .B1_f (new_AGEMA_signal_6687), .Z0_t (ciphertext_s0_t[61]), .Z0_f (ciphertext_s0_f[61]), .Z1_t (ciphertext_s1_t[61]), .Z1_f (ciphertext_s1_f[61]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S02reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS02ser[6]), .A0_f (new_AGEMA_signal_6688), .A1_t (new_AGEMA_signal_6689), .A1_f (new_AGEMA_signal_6690), .B0_t (ciphertext_s0_t[62]), .B0_f (ciphertext_s0_f[62]), .B1_t (ciphertext_s1_t[62]), .B1_f (ciphertext_s1_f[62]), .Z0_t (stateArray_S02reg_gff_1_SFF_6_MUXInst_X), .Z0_f (new_AGEMA_signal_7461), .Z1_t (new_AGEMA_signal_7462), .Z1_f (new_AGEMA_signal_7463) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S02reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S02reg_gff_1_SFF_6_MUXInst_X), .B0_f (new_AGEMA_signal_7461), .B1_t (new_AGEMA_signal_7462), .B1_f (new_AGEMA_signal_7463), .Z0_t (stateArray_S02reg_gff_1_SFF_6_MUXInst_Y), .Z0_f (new_AGEMA_signal_8208), .Z1_t (new_AGEMA_signal_8209), .Z1_f (new_AGEMA_signal_8210) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S02reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (stateArray_S02reg_gff_1_SFF_6_MUXInst_Y), .A0_f (new_AGEMA_signal_8208), .A1_t (new_AGEMA_signal_8209), .A1_f (new_AGEMA_signal_8210), .B0_t (stateArray_inS02ser[6]), .B0_f (new_AGEMA_signal_6688), .B1_t (new_AGEMA_signal_6689), .B1_f (new_AGEMA_signal_6690), .Z0_t (ciphertext_s0_t[62]), .Z0_f (ciphertext_s0_f[62]), .Z1_t (ciphertext_s1_t[62]), .Z1_f (ciphertext_s1_f[62]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S02reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS02ser[7]), .A0_f (new_AGEMA_signal_6691), .A1_t (new_AGEMA_signal_6692), .A1_f (new_AGEMA_signal_6693), .B0_t (ciphertext_s0_t[63]), .B0_f (ciphertext_s0_f[63]), .B1_t (ciphertext_s1_t[63]), .B1_f (ciphertext_s1_f[63]), .Z0_t (stateArray_S02reg_gff_1_SFF_7_MUXInst_X), .Z0_f (new_AGEMA_signal_7464), .Z1_t (new_AGEMA_signal_7465), .Z1_f (new_AGEMA_signal_7466) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S02reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S02reg_gff_1_SFF_7_MUXInst_X), .B0_f (new_AGEMA_signal_7464), .B1_t (new_AGEMA_signal_7465), .B1_f (new_AGEMA_signal_7466), .Z0_t (stateArray_S02reg_gff_1_SFF_7_MUXInst_Y), .Z0_f (new_AGEMA_signal_8211), .Z1_t (new_AGEMA_signal_8212), .Z1_f (new_AGEMA_signal_8213) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S02reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (stateArray_S02reg_gff_1_SFF_7_MUXInst_Y), .A0_f (new_AGEMA_signal_8211), .A1_t (new_AGEMA_signal_8212), .A1_f (new_AGEMA_signal_8213), .B0_t (stateArray_inS02ser[7]), .B0_f (new_AGEMA_signal_6691), .B1_t (new_AGEMA_signal_6692), .B1_f (new_AGEMA_signal_6693), .Z0_t (ciphertext_s0_t[63]), .Z0_f (ciphertext_s0_f[63]), .Z1_t (ciphertext_s1_t[63]), .Z1_f (ciphertext_s1_f[63]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S03reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS03ser[0]), .A0_f (new_AGEMA_signal_10829), .A1_t (new_AGEMA_signal_10830), .A1_f (new_AGEMA_signal_10831), .B0_t (ciphertext_s0_t[24]), .B0_f (ciphertext_s0_f[24]), .B1_t (ciphertext_s1_t[24]), .B1_f (ciphertext_s1_f[24]), .Z0_t (stateArray_S03reg_gff_1_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_10940), .Z1_t (new_AGEMA_signal_10941), .Z1_f (new_AGEMA_signal_10942) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S03reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S03reg_gff_1_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_10940), .B1_t (new_AGEMA_signal_10941), .B1_f (new_AGEMA_signal_10942), .Z0_t (stateArray_S03reg_gff_1_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_11051), .Z1_t (new_AGEMA_signal_11052), .Z1_f (new_AGEMA_signal_11053) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S03reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (stateArray_S03reg_gff_1_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_11051), .A1_t (new_AGEMA_signal_11052), .A1_f (new_AGEMA_signal_11053), .B0_t (stateArray_inS03ser[0]), .B0_f (new_AGEMA_signal_10829), .B1_t (new_AGEMA_signal_10830), .B1_f (new_AGEMA_signal_10831), .Z0_t (ciphertext_s0_t[24]), .Z0_f (ciphertext_s0_f[24]), .Z1_t (ciphertext_s1_t[24]), .Z1_f (ciphertext_s1_f[24]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S03reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS03ser[1]), .A0_f (new_AGEMA_signal_10985), .A1_t (new_AGEMA_signal_10986), .A1_f (new_AGEMA_signal_10987), .B0_t (ciphertext_s0_t[25]), .B0_f (ciphertext_s0_f[25]), .B1_t (ciphertext_s1_t[25]), .B1_f (ciphertext_s1_f[25]), .Z0_t (stateArray_S03reg_gff_1_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_11054), .Z1_t (new_AGEMA_signal_11055), .Z1_f (new_AGEMA_signal_11056) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S03reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S03reg_gff_1_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_11054), .B1_t (new_AGEMA_signal_11055), .B1_f (new_AGEMA_signal_11056), .Z0_t (stateArray_S03reg_gff_1_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_11135), .Z1_t (new_AGEMA_signal_11136), .Z1_f (new_AGEMA_signal_11137) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S03reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (stateArray_S03reg_gff_1_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_11135), .A1_t (new_AGEMA_signal_11136), .A1_f (new_AGEMA_signal_11137), .B0_t (stateArray_inS03ser[1]), .B0_f (new_AGEMA_signal_10985), .B1_t (new_AGEMA_signal_10986), .B1_f (new_AGEMA_signal_10987), .Z0_t (ciphertext_s0_t[25]), .Z0_f (ciphertext_s0_f[25]), .Z1_t (ciphertext_s1_t[25]), .Z1_f (ciphertext_s1_f[25]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S03reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS03ser[2]), .A0_f (new_AGEMA_signal_10835), .A1_t (new_AGEMA_signal_10836), .A1_f (new_AGEMA_signal_10837), .B0_t (ciphertext_s0_t[26]), .B0_f (ciphertext_s0_f[26]), .B1_t (ciphertext_s1_t[26]), .B1_f (ciphertext_s1_f[26]), .Z0_t (stateArray_S03reg_gff_1_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_10943), .Z1_t (new_AGEMA_signal_10944), .Z1_f (new_AGEMA_signal_10945) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S03reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S03reg_gff_1_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_10943), .B1_t (new_AGEMA_signal_10944), .B1_f (new_AGEMA_signal_10945), .Z0_t (stateArray_S03reg_gff_1_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_11057), .Z1_t (new_AGEMA_signal_11058), .Z1_f (new_AGEMA_signal_11059) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S03reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (stateArray_S03reg_gff_1_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_11057), .A1_t (new_AGEMA_signal_11058), .A1_f (new_AGEMA_signal_11059), .B0_t (stateArray_inS03ser[2]), .B0_f (new_AGEMA_signal_10835), .B1_t (new_AGEMA_signal_10836), .B1_f (new_AGEMA_signal_10837), .Z0_t (ciphertext_s0_t[26]), .Z0_f (ciphertext_s0_f[26]), .Z1_t (ciphertext_s1_t[26]), .Z1_f (ciphertext_s1_f[26]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S03reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS03ser[3]), .A0_f (new_AGEMA_signal_10988), .A1_t (new_AGEMA_signal_10989), .A1_f (new_AGEMA_signal_10990), .B0_t (ciphertext_s0_t[27]), .B0_f (ciphertext_s0_f[27]), .B1_t (ciphertext_s1_t[27]), .B1_f (ciphertext_s1_f[27]), .Z0_t (stateArray_S03reg_gff_1_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_11060), .Z1_t (new_AGEMA_signal_11061), .Z1_f (new_AGEMA_signal_11062) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S03reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S03reg_gff_1_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_11060), .B1_t (new_AGEMA_signal_11061), .B1_f (new_AGEMA_signal_11062), .Z0_t (stateArray_S03reg_gff_1_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_11138), .Z1_t (new_AGEMA_signal_11139), .Z1_f (new_AGEMA_signal_11140) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S03reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (stateArray_S03reg_gff_1_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_11138), .A1_t (new_AGEMA_signal_11139), .A1_f (new_AGEMA_signal_11140), .B0_t (stateArray_inS03ser[3]), .B0_f (new_AGEMA_signal_10988), .B1_t (new_AGEMA_signal_10989), .B1_f (new_AGEMA_signal_10990), .Z0_t (ciphertext_s0_t[27]), .Z0_f (ciphertext_s0_f[27]), .Z1_t (ciphertext_s1_t[27]), .Z1_f (ciphertext_s1_f[27]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S03reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS03ser[4]), .A0_f (new_AGEMA_signal_10991), .A1_t (new_AGEMA_signal_10992), .A1_f (new_AGEMA_signal_10993), .B0_t (ciphertext_s0_t[28]), .B0_f (ciphertext_s0_f[28]), .B1_t (ciphertext_s1_t[28]), .B1_f (ciphertext_s1_f[28]), .Z0_t (stateArray_S03reg_gff_1_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_11063), .Z1_t (new_AGEMA_signal_11064), .Z1_f (new_AGEMA_signal_11065) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S03reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S03reg_gff_1_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_11063), .B1_t (new_AGEMA_signal_11064), .B1_f (new_AGEMA_signal_11065), .Z0_t (stateArray_S03reg_gff_1_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_11141), .Z1_t (new_AGEMA_signal_11142), .Z1_f (new_AGEMA_signal_11143) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S03reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (stateArray_S03reg_gff_1_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_11141), .A1_t (new_AGEMA_signal_11142), .A1_f (new_AGEMA_signal_11143), .B0_t (stateArray_inS03ser[4]), .B0_f (new_AGEMA_signal_10991), .B1_t (new_AGEMA_signal_10992), .B1_f (new_AGEMA_signal_10993), .Z0_t (ciphertext_s0_t[28]), .Z0_f (ciphertext_s0_f[28]), .Z1_t (ciphertext_s1_t[28]), .Z1_f (ciphertext_s1_f[28]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S03reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS03ser[5]), .A0_f (new_AGEMA_signal_10844), .A1_t (new_AGEMA_signal_10845), .A1_f (new_AGEMA_signal_10846), .B0_t (ciphertext_s0_t[29]), .B0_f (ciphertext_s0_f[29]), .B1_t (ciphertext_s1_t[29]), .B1_f (ciphertext_s1_f[29]), .Z0_t (stateArray_S03reg_gff_1_SFF_5_MUXInst_X), .Z0_f (new_AGEMA_signal_10946), .Z1_t (new_AGEMA_signal_10947), .Z1_f (new_AGEMA_signal_10948) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S03reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S03reg_gff_1_SFF_5_MUXInst_X), .B0_f (new_AGEMA_signal_10946), .B1_t (new_AGEMA_signal_10947), .B1_f (new_AGEMA_signal_10948), .Z0_t (stateArray_S03reg_gff_1_SFF_5_MUXInst_Y), .Z0_f (new_AGEMA_signal_11066), .Z1_t (new_AGEMA_signal_11067), .Z1_f (new_AGEMA_signal_11068) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S03reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (stateArray_S03reg_gff_1_SFF_5_MUXInst_Y), .A0_f (new_AGEMA_signal_11066), .A1_t (new_AGEMA_signal_11067), .A1_f (new_AGEMA_signal_11068), .B0_t (stateArray_inS03ser[5]), .B0_f (new_AGEMA_signal_10844), .B1_t (new_AGEMA_signal_10845), .B1_f (new_AGEMA_signal_10846), .Z0_t (ciphertext_s0_t[29]), .Z0_f (ciphertext_s0_f[29]), .Z1_t (ciphertext_s1_t[29]), .Z1_f (ciphertext_s1_f[29]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S03reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS03ser[6]), .A0_f (new_AGEMA_signal_10847), .A1_t (new_AGEMA_signal_10848), .A1_f (new_AGEMA_signal_10849), .B0_t (ciphertext_s0_t[30]), .B0_f (ciphertext_s0_f[30]), .B1_t (ciphertext_s1_t[30]), .B1_f (ciphertext_s1_f[30]), .Z0_t (stateArray_S03reg_gff_1_SFF_6_MUXInst_X), .Z0_f (new_AGEMA_signal_10949), .Z1_t (new_AGEMA_signal_10950), .Z1_f (new_AGEMA_signal_10951) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S03reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S03reg_gff_1_SFF_6_MUXInst_X), .B0_f (new_AGEMA_signal_10949), .B1_t (new_AGEMA_signal_10950), .B1_f (new_AGEMA_signal_10951), .Z0_t (stateArray_S03reg_gff_1_SFF_6_MUXInst_Y), .Z0_f (new_AGEMA_signal_11069), .Z1_t (new_AGEMA_signal_11070), .Z1_f (new_AGEMA_signal_11071) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S03reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (stateArray_S03reg_gff_1_SFF_6_MUXInst_Y), .A0_f (new_AGEMA_signal_11069), .A1_t (new_AGEMA_signal_11070), .A1_f (new_AGEMA_signal_11071), .B0_t (stateArray_inS03ser[6]), .B0_f (new_AGEMA_signal_10847), .B1_t (new_AGEMA_signal_10848), .B1_f (new_AGEMA_signal_10849), .Z0_t (ciphertext_s0_t[30]), .Z0_f (ciphertext_s0_f[30]), .Z1_t (ciphertext_s1_t[30]), .Z1_f (ciphertext_s1_f[30]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S03reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS03ser[7]), .A0_f (new_AGEMA_signal_10850), .A1_t (new_AGEMA_signal_10851), .A1_f (new_AGEMA_signal_10852), .B0_t (ciphertext_s0_t[31]), .B0_f (ciphertext_s0_f[31]), .B1_t (ciphertext_s1_t[31]), .B1_f (ciphertext_s1_f[31]), .Z0_t (stateArray_S03reg_gff_1_SFF_7_MUXInst_X), .Z0_f (new_AGEMA_signal_10952), .Z1_t (new_AGEMA_signal_10953), .Z1_f (new_AGEMA_signal_10954) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S03reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S03reg_gff_1_SFF_7_MUXInst_X), .B0_f (new_AGEMA_signal_10952), .B1_t (new_AGEMA_signal_10953), .B1_f (new_AGEMA_signal_10954), .Z0_t (stateArray_S03reg_gff_1_SFF_7_MUXInst_Y), .Z0_f (new_AGEMA_signal_11072), .Z1_t (new_AGEMA_signal_11073), .Z1_f (new_AGEMA_signal_11074) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S03reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (stateArray_S03reg_gff_1_SFF_7_MUXInst_Y), .A0_f (new_AGEMA_signal_11072), .A1_t (new_AGEMA_signal_11073), .A1_f (new_AGEMA_signal_11074), .B0_t (stateArray_inS03ser[7]), .B0_f (new_AGEMA_signal_10850), .B1_t (new_AGEMA_signal_10851), .B1_f (new_AGEMA_signal_10852), .Z0_t (ciphertext_s0_t[31]), .Z0_f (ciphertext_s0_f[31]), .Z1_t (ciphertext_s1_t[31]), .Z1_f (ciphertext_s1_f[31]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S10reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS10ser[0]), .A0_f (new_AGEMA_signal_6694), .A1_t (new_AGEMA_signal_6695), .A1_f (new_AGEMA_signal_6696), .B0_t (ciphertext_s0_t[80]), .B0_f (ciphertext_s0_f[80]), .B1_t (ciphertext_s1_t[80]), .B1_f (ciphertext_s1_f[80]), .Z0_t (stateArray_S10reg_gff_1_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_7467), .Z1_t (new_AGEMA_signal_7468), .Z1_f (new_AGEMA_signal_7469) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S10reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S10reg_gff_1_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_7467), .B1_t (new_AGEMA_signal_7468), .B1_f (new_AGEMA_signal_7469), .Z0_t (stateArray_S10reg_gff_1_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_8214), .Z1_t (new_AGEMA_signal_8215), .Z1_f (new_AGEMA_signal_8216) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S10reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (stateArray_S10reg_gff_1_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_8214), .A1_t (new_AGEMA_signal_8215), .A1_f (new_AGEMA_signal_8216), .B0_t (stateArray_inS10ser[0]), .B0_f (new_AGEMA_signal_6694), .B1_t (new_AGEMA_signal_6695), .B1_f (new_AGEMA_signal_6696), .Z0_t (ciphertext_s0_t[112]), .Z0_f (ciphertext_s0_f[112]), .Z1_t (ciphertext_s1_t[112]), .Z1_f (ciphertext_s1_f[112]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S10reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS10ser[1]), .A0_f (new_AGEMA_signal_6697), .A1_t (new_AGEMA_signal_6698), .A1_f (new_AGEMA_signal_6699), .B0_t (ciphertext_s0_t[81]), .B0_f (ciphertext_s0_f[81]), .B1_t (ciphertext_s1_t[81]), .B1_f (ciphertext_s1_f[81]), .Z0_t (stateArray_S10reg_gff_1_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_7470), .Z1_t (new_AGEMA_signal_7471), .Z1_f (new_AGEMA_signal_7472) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S10reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S10reg_gff_1_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_7470), .B1_t (new_AGEMA_signal_7471), .B1_f (new_AGEMA_signal_7472), .Z0_t (stateArray_S10reg_gff_1_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_8217), .Z1_t (new_AGEMA_signal_8218), .Z1_f (new_AGEMA_signal_8219) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S10reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (stateArray_S10reg_gff_1_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_8217), .A1_t (new_AGEMA_signal_8218), .A1_f (new_AGEMA_signal_8219), .B0_t (stateArray_inS10ser[1]), .B0_f (new_AGEMA_signal_6697), .B1_t (new_AGEMA_signal_6698), .B1_f (new_AGEMA_signal_6699), .Z0_t (ciphertext_s0_t[113]), .Z0_f (ciphertext_s0_f[113]), .Z1_t (ciphertext_s1_t[113]), .Z1_f (ciphertext_s1_f[113]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S10reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS10ser[2]), .A0_f (new_AGEMA_signal_6700), .A1_t (new_AGEMA_signal_6701), .A1_f (new_AGEMA_signal_6702), .B0_t (ciphertext_s0_t[82]), .B0_f (ciphertext_s0_f[82]), .B1_t (ciphertext_s1_t[82]), .B1_f (ciphertext_s1_f[82]), .Z0_t (stateArray_S10reg_gff_1_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_7473), .Z1_t (new_AGEMA_signal_7474), .Z1_f (new_AGEMA_signal_7475) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S10reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S10reg_gff_1_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_7473), .B1_t (new_AGEMA_signal_7474), .B1_f (new_AGEMA_signal_7475), .Z0_t (stateArray_S10reg_gff_1_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_8220), .Z1_t (new_AGEMA_signal_8221), .Z1_f (new_AGEMA_signal_8222) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S10reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (stateArray_S10reg_gff_1_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_8220), .A1_t (new_AGEMA_signal_8221), .A1_f (new_AGEMA_signal_8222), .B0_t (stateArray_inS10ser[2]), .B0_f (new_AGEMA_signal_6700), .B1_t (new_AGEMA_signal_6701), .B1_f (new_AGEMA_signal_6702), .Z0_t (ciphertext_s0_t[114]), .Z0_f (ciphertext_s0_f[114]), .Z1_t (ciphertext_s1_t[114]), .Z1_f (ciphertext_s1_f[114]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S10reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS10ser[3]), .A0_f (new_AGEMA_signal_6703), .A1_t (new_AGEMA_signal_6704), .A1_f (new_AGEMA_signal_6705), .B0_t (ciphertext_s0_t[83]), .B0_f (ciphertext_s0_f[83]), .B1_t (ciphertext_s1_t[83]), .B1_f (ciphertext_s1_f[83]), .Z0_t (stateArray_S10reg_gff_1_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_7476), .Z1_t (new_AGEMA_signal_7477), .Z1_f (new_AGEMA_signal_7478) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S10reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S10reg_gff_1_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_7476), .B1_t (new_AGEMA_signal_7477), .B1_f (new_AGEMA_signal_7478), .Z0_t (stateArray_S10reg_gff_1_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_8223), .Z1_t (new_AGEMA_signal_8224), .Z1_f (new_AGEMA_signal_8225) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S10reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (stateArray_S10reg_gff_1_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_8223), .A1_t (new_AGEMA_signal_8224), .A1_f (new_AGEMA_signal_8225), .B0_t (stateArray_inS10ser[3]), .B0_f (new_AGEMA_signal_6703), .B1_t (new_AGEMA_signal_6704), .B1_f (new_AGEMA_signal_6705), .Z0_t (ciphertext_s0_t[115]), .Z0_f (ciphertext_s0_f[115]), .Z1_t (ciphertext_s1_t[115]), .Z1_f (ciphertext_s1_f[115]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S10reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS10ser[4]), .A0_f (new_AGEMA_signal_6706), .A1_t (new_AGEMA_signal_6707), .A1_f (new_AGEMA_signal_6708), .B0_t (ciphertext_s0_t[84]), .B0_f (ciphertext_s0_f[84]), .B1_t (ciphertext_s1_t[84]), .B1_f (ciphertext_s1_f[84]), .Z0_t (stateArray_S10reg_gff_1_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_7479), .Z1_t (new_AGEMA_signal_7480), .Z1_f (new_AGEMA_signal_7481) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S10reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S10reg_gff_1_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_7479), .B1_t (new_AGEMA_signal_7480), .B1_f (new_AGEMA_signal_7481), .Z0_t (stateArray_S10reg_gff_1_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_8226), .Z1_t (new_AGEMA_signal_8227), .Z1_f (new_AGEMA_signal_8228) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S10reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (stateArray_S10reg_gff_1_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_8226), .A1_t (new_AGEMA_signal_8227), .A1_f (new_AGEMA_signal_8228), .B0_t (stateArray_inS10ser[4]), .B0_f (new_AGEMA_signal_6706), .B1_t (new_AGEMA_signal_6707), .B1_f (new_AGEMA_signal_6708), .Z0_t (ciphertext_s0_t[116]), .Z0_f (ciphertext_s0_f[116]), .Z1_t (ciphertext_s1_t[116]), .Z1_f (ciphertext_s1_f[116]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S10reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS10ser[5]), .A0_f (new_AGEMA_signal_6709), .A1_t (new_AGEMA_signal_6710), .A1_f (new_AGEMA_signal_6711), .B0_t (ciphertext_s0_t[85]), .B0_f (ciphertext_s0_f[85]), .B1_t (ciphertext_s1_t[85]), .B1_f (ciphertext_s1_f[85]), .Z0_t (stateArray_S10reg_gff_1_SFF_5_MUXInst_X), .Z0_f (new_AGEMA_signal_7482), .Z1_t (new_AGEMA_signal_7483), .Z1_f (new_AGEMA_signal_7484) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S10reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S10reg_gff_1_SFF_5_MUXInst_X), .B0_f (new_AGEMA_signal_7482), .B1_t (new_AGEMA_signal_7483), .B1_f (new_AGEMA_signal_7484), .Z0_t (stateArray_S10reg_gff_1_SFF_5_MUXInst_Y), .Z0_f (new_AGEMA_signal_8229), .Z1_t (new_AGEMA_signal_8230), .Z1_f (new_AGEMA_signal_8231) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S10reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (stateArray_S10reg_gff_1_SFF_5_MUXInst_Y), .A0_f (new_AGEMA_signal_8229), .A1_t (new_AGEMA_signal_8230), .A1_f (new_AGEMA_signal_8231), .B0_t (stateArray_inS10ser[5]), .B0_f (new_AGEMA_signal_6709), .B1_t (new_AGEMA_signal_6710), .B1_f (new_AGEMA_signal_6711), .Z0_t (ciphertext_s0_t[117]), .Z0_f (ciphertext_s0_f[117]), .Z1_t (ciphertext_s1_t[117]), .Z1_f (ciphertext_s1_f[117]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S10reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS10ser[6]), .A0_f (new_AGEMA_signal_6712), .A1_t (new_AGEMA_signal_6713), .A1_f (new_AGEMA_signal_6714), .B0_t (ciphertext_s0_t[86]), .B0_f (ciphertext_s0_f[86]), .B1_t (ciphertext_s1_t[86]), .B1_f (ciphertext_s1_f[86]), .Z0_t (stateArray_S10reg_gff_1_SFF_6_MUXInst_X), .Z0_f (new_AGEMA_signal_7485), .Z1_t (new_AGEMA_signal_7486), .Z1_f (new_AGEMA_signal_7487) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S10reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S10reg_gff_1_SFF_6_MUXInst_X), .B0_f (new_AGEMA_signal_7485), .B1_t (new_AGEMA_signal_7486), .B1_f (new_AGEMA_signal_7487), .Z0_t (stateArray_S10reg_gff_1_SFF_6_MUXInst_Y), .Z0_f (new_AGEMA_signal_8232), .Z1_t (new_AGEMA_signal_8233), .Z1_f (new_AGEMA_signal_8234) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S10reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (stateArray_S10reg_gff_1_SFF_6_MUXInst_Y), .A0_f (new_AGEMA_signal_8232), .A1_t (new_AGEMA_signal_8233), .A1_f (new_AGEMA_signal_8234), .B0_t (stateArray_inS10ser[6]), .B0_f (new_AGEMA_signal_6712), .B1_t (new_AGEMA_signal_6713), .B1_f (new_AGEMA_signal_6714), .Z0_t (ciphertext_s0_t[118]), .Z0_f (ciphertext_s0_f[118]), .Z1_t (ciphertext_s1_t[118]), .Z1_f (ciphertext_s1_f[118]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S10reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS10ser[7]), .A0_f (new_AGEMA_signal_6715), .A1_t (new_AGEMA_signal_6716), .A1_f (new_AGEMA_signal_6717), .B0_t (ciphertext_s0_t[87]), .B0_f (ciphertext_s0_f[87]), .B1_t (ciphertext_s1_t[87]), .B1_f (ciphertext_s1_f[87]), .Z0_t (stateArray_S10reg_gff_1_SFF_7_MUXInst_X), .Z0_f (new_AGEMA_signal_7488), .Z1_t (new_AGEMA_signal_7489), .Z1_f (new_AGEMA_signal_7490) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S10reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S10reg_gff_1_SFF_7_MUXInst_X), .B0_f (new_AGEMA_signal_7488), .B1_t (new_AGEMA_signal_7489), .B1_f (new_AGEMA_signal_7490), .Z0_t (stateArray_S10reg_gff_1_SFF_7_MUXInst_Y), .Z0_f (new_AGEMA_signal_8235), .Z1_t (new_AGEMA_signal_8236), .Z1_f (new_AGEMA_signal_8237) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S10reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (stateArray_S10reg_gff_1_SFF_7_MUXInst_Y), .A0_f (new_AGEMA_signal_8235), .A1_t (new_AGEMA_signal_8236), .A1_f (new_AGEMA_signal_8237), .B0_t (stateArray_inS10ser[7]), .B0_f (new_AGEMA_signal_6715), .B1_t (new_AGEMA_signal_6716), .B1_f (new_AGEMA_signal_6717), .Z0_t (ciphertext_s0_t[119]), .Z0_f (ciphertext_s0_f[119]), .Z1_t (ciphertext_s1_t[119]), .Z1_f (ciphertext_s1_f[119]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S11reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS11ser[0]), .A0_f (new_AGEMA_signal_6718), .A1_t (new_AGEMA_signal_6719), .A1_f (new_AGEMA_signal_6720), .B0_t (ciphertext_s0_t[48]), .B0_f (ciphertext_s0_f[48]), .B1_t (ciphertext_s1_t[48]), .B1_f (ciphertext_s1_f[48]), .Z0_t (stateArray_S11reg_gff_1_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_7491), .Z1_t (new_AGEMA_signal_7492), .Z1_f (new_AGEMA_signal_7493) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S11reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S11reg_gff_1_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_7491), .B1_t (new_AGEMA_signal_7492), .B1_f (new_AGEMA_signal_7493), .Z0_t (stateArray_S11reg_gff_1_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_8238), .Z1_t (new_AGEMA_signal_8239), .Z1_f (new_AGEMA_signal_8240) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S11reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (stateArray_S11reg_gff_1_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_8238), .A1_t (new_AGEMA_signal_8239), .A1_f (new_AGEMA_signal_8240), .B0_t (stateArray_inS11ser[0]), .B0_f (new_AGEMA_signal_6718), .B1_t (new_AGEMA_signal_6719), .B1_f (new_AGEMA_signal_6720), .Z0_t (ciphertext_s0_t[80]), .Z0_f (ciphertext_s0_f[80]), .Z1_t (ciphertext_s1_t[80]), .Z1_f (ciphertext_s1_f[80]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S11reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS11ser[1]), .A0_f (new_AGEMA_signal_6721), .A1_t (new_AGEMA_signal_6722), .A1_f (new_AGEMA_signal_6723), .B0_t (ciphertext_s0_t[49]), .B0_f (ciphertext_s0_f[49]), .B1_t (ciphertext_s1_t[49]), .B1_f (ciphertext_s1_f[49]), .Z0_t (stateArray_S11reg_gff_1_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_7494), .Z1_t (new_AGEMA_signal_7495), .Z1_f (new_AGEMA_signal_7496) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S11reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S11reg_gff_1_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_7494), .B1_t (new_AGEMA_signal_7495), .B1_f (new_AGEMA_signal_7496), .Z0_t (stateArray_S11reg_gff_1_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_8241), .Z1_t (new_AGEMA_signal_8242), .Z1_f (new_AGEMA_signal_8243) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S11reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (stateArray_S11reg_gff_1_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_8241), .A1_t (new_AGEMA_signal_8242), .A1_f (new_AGEMA_signal_8243), .B0_t (stateArray_inS11ser[1]), .B0_f (new_AGEMA_signal_6721), .B1_t (new_AGEMA_signal_6722), .B1_f (new_AGEMA_signal_6723), .Z0_t (ciphertext_s0_t[81]), .Z0_f (ciphertext_s0_f[81]), .Z1_t (ciphertext_s1_t[81]), .Z1_f (ciphertext_s1_f[81]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S11reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS11ser[2]), .A0_f (new_AGEMA_signal_6724), .A1_t (new_AGEMA_signal_6725), .A1_f (new_AGEMA_signal_6726), .B0_t (ciphertext_s0_t[50]), .B0_f (ciphertext_s0_f[50]), .B1_t (ciphertext_s1_t[50]), .B1_f (ciphertext_s1_f[50]), .Z0_t (stateArray_S11reg_gff_1_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_7497), .Z1_t (new_AGEMA_signal_7498), .Z1_f (new_AGEMA_signal_7499) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S11reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S11reg_gff_1_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_7497), .B1_t (new_AGEMA_signal_7498), .B1_f (new_AGEMA_signal_7499), .Z0_t (stateArray_S11reg_gff_1_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_8244), .Z1_t (new_AGEMA_signal_8245), .Z1_f (new_AGEMA_signal_8246) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S11reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (stateArray_S11reg_gff_1_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_8244), .A1_t (new_AGEMA_signal_8245), .A1_f (new_AGEMA_signal_8246), .B0_t (stateArray_inS11ser[2]), .B0_f (new_AGEMA_signal_6724), .B1_t (new_AGEMA_signal_6725), .B1_f (new_AGEMA_signal_6726), .Z0_t (ciphertext_s0_t[82]), .Z0_f (ciphertext_s0_f[82]), .Z1_t (ciphertext_s1_t[82]), .Z1_f (ciphertext_s1_f[82]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S11reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS11ser[3]), .A0_f (new_AGEMA_signal_6727), .A1_t (new_AGEMA_signal_6728), .A1_f (new_AGEMA_signal_6729), .B0_t (ciphertext_s0_t[51]), .B0_f (ciphertext_s0_f[51]), .B1_t (ciphertext_s1_t[51]), .B1_f (ciphertext_s1_f[51]), .Z0_t (stateArray_S11reg_gff_1_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_7500), .Z1_t (new_AGEMA_signal_7501), .Z1_f (new_AGEMA_signal_7502) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S11reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S11reg_gff_1_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_7500), .B1_t (new_AGEMA_signal_7501), .B1_f (new_AGEMA_signal_7502), .Z0_t (stateArray_S11reg_gff_1_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_8247), .Z1_t (new_AGEMA_signal_8248), .Z1_f (new_AGEMA_signal_8249) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S11reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (stateArray_S11reg_gff_1_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_8247), .A1_t (new_AGEMA_signal_8248), .A1_f (new_AGEMA_signal_8249), .B0_t (stateArray_inS11ser[3]), .B0_f (new_AGEMA_signal_6727), .B1_t (new_AGEMA_signal_6728), .B1_f (new_AGEMA_signal_6729), .Z0_t (ciphertext_s0_t[83]), .Z0_f (ciphertext_s0_f[83]), .Z1_t (ciphertext_s1_t[83]), .Z1_f (ciphertext_s1_f[83]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S11reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS11ser[4]), .A0_f (new_AGEMA_signal_6730), .A1_t (new_AGEMA_signal_6731), .A1_f (new_AGEMA_signal_6732), .B0_t (ciphertext_s0_t[52]), .B0_f (ciphertext_s0_f[52]), .B1_t (ciphertext_s1_t[52]), .B1_f (ciphertext_s1_f[52]), .Z0_t (stateArray_S11reg_gff_1_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_7503), .Z1_t (new_AGEMA_signal_7504), .Z1_f (new_AGEMA_signal_7505) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S11reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S11reg_gff_1_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_7503), .B1_t (new_AGEMA_signal_7504), .B1_f (new_AGEMA_signal_7505), .Z0_t (stateArray_S11reg_gff_1_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_8250), .Z1_t (new_AGEMA_signal_8251), .Z1_f (new_AGEMA_signal_8252) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S11reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (stateArray_S11reg_gff_1_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_8250), .A1_t (new_AGEMA_signal_8251), .A1_f (new_AGEMA_signal_8252), .B0_t (stateArray_inS11ser[4]), .B0_f (new_AGEMA_signal_6730), .B1_t (new_AGEMA_signal_6731), .B1_f (new_AGEMA_signal_6732), .Z0_t (ciphertext_s0_t[84]), .Z0_f (ciphertext_s0_f[84]), .Z1_t (ciphertext_s1_t[84]), .Z1_f (ciphertext_s1_f[84]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S11reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS11ser[5]), .A0_f (new_AGEMA_signal_6733), .A1_t (new_AGEMA_signal_6734), .A1_f (new_AGEMA_signal_6735), .B0_t (ciphertext_s0_t[53]), .B0_f (ciphertext_s0_f[53]), .B1_t (ciphertext_s1_t[53]), .B1_f (ciphertext_s1_f[53]), .Z0_t (stateArray_S11reg_gff_1_SFF_5_MUXInst_X), .Z0_f (new_AGEMA_signal_7506), .Z1_t (new_AGEMA_signal_7507), .Z1_f (new_AGEMA_signal_7508) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S11reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S11reg_gff_1_SFF_5_MUXInst_X), .B0_f (new_AGEMA_signal_7506), .B1_t (new_AGEMA_signal_7507), .B1_f (new_AGEMA_signal_7508), .Z0_t (stateArray_S11reg_gff_1_SFF_5_MUXInst_Y), .Z0_f (new_AGEMA_signal_8253), .Z1_t (new_AGEMA_signal_8254), .Z1_f (new_AGEMA_signal_8255) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S11reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (stateArray_S11reg_gff_1_SFF_5_MUXInst_Y), .A0_f (new_AGEMA_signal_8253), .A1_t (new_AGEMA_signal_8254), .A1_f (new_AGEMA_signal_8255), .B0_t (stateArray_inS11ser[5]), .B0_f (new_AGEMA_signal_6733), .B1_t (new_AGEMA_signal_6734), .B1_f (new_AGEMA_signal_6735), .Z0_t (ciphertext_s0_t[85]), .Z0_f (ciphertext_s0_f[85]), .Z1_t (ciphertext_s1_t[85]), .Z1_f (ciphertext_s1_f[85]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S11reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS11ser[6]), .A0_f (new_AGEMA_signal_6736), .A1_t (new_AGEMA_signal_6737), .A1_f (new_AGEMA_signal_6738), .B0_t (ciphertext_s0_t[54]), .B0_f (ciphertext_s0_f[54]), .B1_t (ciphertext_s1_t[54]), .B1_f (ciphertext_s1_f[54]), .Z0_t (stateArray_S11reg_gff_1_SFF_6_MUXInst_X), .Z0_f (new_AGEMA_signal_7509), .Z1_t (new_AGEMA_signal_7510), .Z1_f (new_AGEMA_signal_7511) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S11reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S11reg_gff_1_SFF_6_MUXInst_X), .B0_f (new_AGEMA_signal_7509), .B1_t (new_AGEMA_signal_7510), .B1_f (new_AGEMA_signal_7511), .Z0_t (stateArray_S11reg_gff_1_SFF_6_MUXInst_Y), .Z0_f (new_AGEMA_signal_8256), .Z1_t (new_AGEMA_signal_8257), .Z1_f (new_AGEMA_signal_8258) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S11reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (stateArray_S11reg_gff_1_SFF_6_MUXInst_Y), .A0_f (new_AGEMA_signal_8256), .A1_t (new_AGEMA_signal_8257), .A1_f (new_AGEMA_signal_8258), .B0_t (stateArray_inS11ser[6]), .B0_f (new_AGEMA_signal_6736), .B1_t (new_AGEMA_signal_6737), .B1_f (new_AGEMA_signal_6738), .Z0_t (ciphertext_s0_t[86]), .Z0_f (ciphertext_s0_f[86]), .Z1_t (ciphertext_s1_t[86]), .Z1_f (ciphertext_s1_f[86]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S11reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS11ser[7]), .A0_f (new_AGEMA_signal_6739), .A1_t (new_AGEMA_signal_6740), .A1_f (new_AGEMA_signal_6741), .B0_t (ciphertext_s0_t[55]), .B0_f (ciphertext_s0_f[55]), .B1_t (ciphertext_s1_t[55]), .B1_f (ciphertext_s1_f[55]), .Z0_t (stateArray_S11reg_gff_1_SFF_7_MUXInst_X), .Z0_f (new_AGEMA_signal_7512), .Z1_t (new_AGEMA_signal_7513), .Z1_f (new_AGEMA_signal_7514) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S11reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S11reg_gff_1_SFF_7_MUXInst_X), .B0_f (new_AGEMA_signal_7512), .B1_t (new_AGEMA_signal_7513), .B1_f (new_AGEMA_signal_7514), .Z0_t (stateArray_S11reg_gff_1_SFF_7_MUXInst_Y), .Z0_f (new_AGEMA_signal_8259), .Z1_t (new_AGEMA_signal_8260), .Z1_f (new_AGEMA_signal_8261) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S11reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (stateArray_S11reg_gff_1_SFF_7_MUXInst_Y), .A0_f (new_AGEMA_signal_8259), .A1_t (new_AGEMA_signal_8260), .A1_f (new_AGEMA_signal_8261), .B0_t (stateArray_inS11ser[7]), .B0_f (new_AGEMA_signal_6739), .B1_t (new_AGEMA_signal_6740), .B1_f (new_AGEMA_signal_6741), .Z0_t (ciphertext_s0_t[87]), .Z0_f (ciphertext_s0_f[87]), .Z1_t (ciphertext_s1_t[87]), .Z1_f (ciphertext_s1_f[87]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S12reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS12ser[0]), .A0_f (new_AGEMA_signal_6742), .A1_t (new_AGEMA_signal_6743), .A1_f (new_AGEMA_signal_6744), .B0_t (ciphertext_s0_t[16]), .B0_f (ciphertext_s0_f[16]), .B1_t (ciphertext_s1_t[16]), .B1_f (ciphertext_s1_f[16]), .Z0_t (stateArray_S12reg_gff_1_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_7515), .Z1_t (new_AGEMA_signal_7516), .Z1_f (new_AGEMA_signal_7517) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S12reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S12reg_gff_1_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_7515), .B1_t (new_AGEMA_signal_7516), .B1_f (new_AGEMA_signal_7517), .Z0_t (stateArray_S12reg_gff_1_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_8262), .Z1_t (new_AGEMA_signal_8263), .Z1_f (new_AGEMA_signal_8264) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S12reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (stateArray_S12reg_gff_1_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_8262), .A1_t (new_AGEMA_signal_8263), .A1_f (new_AGEMA_signal_8264), .B0_t (stateArray_inS12ser[0]), .B0_f (new_AGEMA_signal_6742), .B1_t (new_AGEMA_signal_6743), .B1_f (new_AGEMA_signal_6744), .Z0_t (ciphertext_s0_t[48]), .Z0_f (ciphertext_s0_f[48]), .Z1_t (ciphertext_s1_t[48]), .Z1_f (ciphertext_s1_f[48]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S12reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS12ser[1]), .A0_f (new_AGEMA_signal_6745), .A1_t (new_AGEMA_signal_6746), .A1_f (new_AGEMA_signal_6747), .B0_t (ciphertext_s0_t[17]), .B0_f (ciphertext_s0_f[17]), .B1_t (ciphertext_s1_t[17]), .B1_f (ciphertext_s1_f[17]), .Z0_t (stateArray_S12reg_gff_1_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_7518), .Z1_t (new_AGEMA_signal_7519), .Z1_f (new_AGEMA_signal_7520) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S12reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S12reg_gff_1_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_7518), .B1_t (new_AGEMA_signal_7519), .B1_f (new_AGEMA_signal_7520), .Z0_t (stateArray_S12reg_gff_1_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_8265), .Z1_t (new_AGEMA_signal_8266), .Z1_f (new_AGEMA_signal_8267) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S12reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (stateArray_S12reg_gff_1_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_8265), .A1_t (new_AGEMA_signal_8266), .A1_f (new_AGEMA_signal_8267), .B0_t (stateArray_inS12ser[1]), .B0_f (new_AGEMA_signal_6745), .B1_t (new_AGEMA_signal_6746), .B1_f (new_AGEMA_signal_6747), .Z0_t (ciphertext_s0_t[49]), .Z0_f (ciphertext_s0_f[49]), .Z1_t (ciphertext_s1_t[49]), .Z1_f (ciphertext_s1_f[49]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S12reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS12ser[2]), .A0_f (new_AGEMA_signal_6748), .A1_t (new_AGEMA_signal_6749), .A1_f (new_AGEMA_signal_6750), .B0_t (ciphertext_s0_t[18]), .B0_f (ciphertext_s0_f[18]), .B1_t (ciphertext_s1_t[18]), .B1_f (ciphertext_s1_f[18]), .Z0_t (stateArray_S12reg_gff_1_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_7521), .Z1_t (new_AGEMA_signal_7522), .Z1_f (new_AGEMA_signal_7523) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S12reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S12reg_gff_1_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_7521), .B1_t (new_AGEMA_signal_7522), .B1_f (new_AGEMA_signal_7523), .Z0_t (stateArray_S12reg_gff_1_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_8268), .Z1_t (new_AGEMA_signal_8269), .Z1_f (new_AGEMA_signal_8270) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S12reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (stateArray_S12reg_gff_1_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_8268), .A1_t (new_AGEMA_signal_8269), .A1_f (new_AGEMA_signal_8270), .B0_t (stateArray_inS12ser[2]), .B0_f (new_AGEMA_signal_6748), .B1_t (new_AGEMA_signal_6749), .B1_f (new_AGEMA_signal_6750), .Z0_t (ciphertext_s0_t[50]), .Z0_f (ciphertext_s0_f[50]), .Z1_t (ciphertext_s1_t[50]), .Z1_f (ciphertext_s1_f[50]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S12reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS12ser[3]), .A0_f (new_AGEMA_signal_6751), .A1_t (new_AGEMA_signal_6752), .A1_f (new_AGEMA_signal_6753), .B0_t (ciphertext_s0_t[19]), .B0_f (ciphertext_s0_f[19]), .B1_t (ciphertext_s1_t[19]), .B1_f (ciphertext_s1_f[19]), .Z0_t (stateArray_S12reg_gff_1_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_7524), .Z1_t (new_AGEMA_signal_7525), .Z1_f (new_AGEMA_signal_7526) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S12reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S12reg_gff_1_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_7524), .B1_t (new_AGEMA_signal_7525), .B1_f (new_AGEMA_signal_7526), .Z0_t (stateArray_S12reg_gff_1_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_8271), .Z1_t (new_AGEMA_signal_8272), .Z1_f (new_AGEMA_signal_8273) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S12reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (stateArray_S12reg_gff_1_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_8271), .A1_t (new_AGEMA_signal_8272), .A1_f (new_AGEMA_signal_8273), .B0_t (stateArray_inS12ser[3]), .B0_f (new_AGEMA_signal_6751), .B1_t (new_AGEMA_signal_6752), .B1_f (new_AGEMA_signal_6753), .Z0_t (ciphertext_s0_t[51]), .Z0_f (ciphertext_s0_f[51]), .Z1_t (ciphertext_s1_t[51]), .Z1_f (ciphertext_s1_f[51]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S12reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS12ser[4]), .A0_f (new_AGEMA_signal_6754), .A1_t (new_AGEMA_signal_6755), .A1_f (new_AGEMA_signal_6756), .B0_t (ciphertext_s0_t[20]), .B0_f (ciphertext_s0_f[20]), .B1_t (ciphertext_s1_t[20]), .B1_f (ciphertext_s1_f[20]), .Z0_t (stateArray_S12reg_gff_1_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_7527), .Z1_t (new_AGEMA_signal_7528), .Z1_f (new_AGEMA_signal_7529) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S12reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S12reg_gff_1_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_7527), .B1_t (new_AGEMA_signal_7528), .B1_f (new_AGEMA_signal_7529), .Z0_t (stateArray_S12reg_gff_1_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_8274), .Z1_t (new_AGEMA_signal_8275), .Z1_f (new_AGEMA_signal_8276) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S12reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (stateArray_S12reg_gff_1_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_8274), .A1_t (new_AGEMA_signal_8275), .A1_f (new_AGEMA_signal_8276), .B0_t (stateArray_inS12ser[4]), .B0_f (new_AGEMA_signal_6754), .B1_t (new_AGEMA_signal_6755), .B1_f (new_AGEMA_signal_6756), .Z0_t (ciphertext_s0_t[52]), .Z0_f (ciphertext_s0_f[52]), .Z1_t (ciphertext_s1_t[52]), .Z1_f (ciphertext_s1_f[52]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S12reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS12ser[5]), .A0_f (new_AGEMA_signal_6757), .A1_t (new_AGEMA_signal_6758), .A1_f (new_AGEMA_signal_6759), .B0_t (ciphertext_s0_t[21]), .B0_f (ciphertext_s0_f[21]), .B1_t (ciphertext_s1_t[21]), .B1_f (ciphertext_s1_f[21]), .Z0_t (stateArray_S12reg_gff_1_SFF_5_MUXInst_X), .Z0_f (new_AGEMA_signal_7530), .Z1_t (new_AGEMA_signal_7531), .Z1_f (new_AGEMA_signal_7532) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S12reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S12reg_gff_1_SFF_5_MUXInst_X), .B0_f (new_AGEMA_signal_7530), .B1_t (new_AGEMA_signal_7531), .B1_f (new_AGEMA_signal_7532), .Z0_t (stateArray_S12reg_gff_1_SFF_5_MUXInst_Y), .Z0_f (new_AGEMA_signal_8277), .Z1_t (new_AGEMA_signal_8278), .Z1_f (new_AGEMA_signal_8279) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S12reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (stateArray_S12reg_gff_1_SFF_5_MUXInst_Y), .A0_f (new_AGEMA_signal_8277), .A1_t (new_AGEMA_signal_8278), .A1_f (new_AGEMA_signal_8279), .B0_t (stateArray_inS12ser[5]), .B0_f (new_AGEMA_signal_6757), .B1_t (new_AGEMA_signal_6758), .B1_f (new_AGEMA_signal_6759), .Z0_t (ciphertext_s0_t[53]), .Z0_f (ciphertext_s0_f[53]), .Z1_t (ciphertext_s1_t[53]), .Z1_f (ciphertext_s1_f[53]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S12reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS12ser[6]), .A0_f (new_AGEMA_signal_6760), .A1_t (new_AGEMA_signal_6761), .A1_f (new_AGEMA_signal_6762), .B0_t (ciphertext_s0_t[22]), .B0_f (ciphertext_s0_f[22]), .B1_t (ciphertext_s1_t[22]), .B1_f (ciphertext_s1_f[22]), .Z0_t (stateArray_S12reg_gff_1_SFF_6_MUXInst_X), .Z0_f (new_AGEMA_signal_7533), .Z1_t (new_AGEMA_signal_7534), .Z1_f (new_AGEMA_signal_7535) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S12reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S12reg_gff_1_SFF_6_MUXInst_X), .B0_f (new_AGEMA_signal_7533), .B1_t (new_AGEMA_signal_7534), .B1_f (new_AGEMA_signal_7535), .Z0_t (stateArray_S12reg_gff_1_SFF_6_MUXInst_Y), .Z0_f (new_AGEMA_signal_8280), .Z1_t (new_AGEMA_signal_8281), .Z1_f (new_AGEMA_signal_8282) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S12reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (stateArray_S12reg_gff_1_SFF_6_MUXInst_Y), .A0_f (new_AGEMA_signal_8280), .A1_t (new_AGEMA_signal_8281), .A1_f (new_AGEMA_signal_8282), .B0_t (stateArray_inS12ser[6]), .B0_f (new_AGEMA_signal_6760), .B1_t (new_AGEMA_signal_6761), .B1_f (new_AGEMA_signal_6762), .Z0_t (ciphertext_s0_t[54]), .Z0_f (ciphertext_s0_f[54]), .Z1_t (ciphertext_s1_t[54]), .Z1_f (ciphertext_s1_f[54]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S12reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS12ser[7]), .A0_f (new_AGEMA_signal_6763), .A1_t (new_AGEMA_signal_6764), .A1_f (new_AGEMA_signal_6765), .B0_t (ciphertext_s0_t[23]), .B0_f (ciphertext_s0_f[23]), .B1_t (ciphertext_s1_t[23]), .B1_f (ciphertext_s1_f[23]), .Z0_t (stateArray_S12reg_gff_1_SFF_7_MUXInst_X), .Z0_f (new_AGEMA_signal_7536), .Z1_t (new_AGEMA_signal_7537), .Z1_f (new_AGEMA_signal_7538) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S12reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S12reg_gff_1_SFF_7_MUXInst_X), .B0_f (new_AGEMA_signal_7536), .B1_t (new_AGEMA_signal_7537), .B1_f (new_AGEMA_signal_7538), .Z0_t (stateArray_S12reg_gff_1_SFF_7_MUXInst_Y), .Z0_f (new_AGEMA_signal_8283), .Z1_t (new_AGEMA_signal_8284), .Z1_f (new_AGEMA_signal_8285) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S12reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (stateArray_S12reg_gff_1_SFF_7_MUXInst_Y), .A0_f (new_AGEMA_signal_8283), .A1_t (new_AGEMA_signal_8284), .A1_f (new_AGEMA_signal_8285), .B0_t (stateArray_inS12ser[7]), .B0_f (new_AGEMA_signal_6763), .B1_t (new_AGEMA_signal_6764), .B1_f (new_AGEMA_signal_6765), .Z0_t (ciphertext_s0_t[55]), .Z0_f (ciphertext_s0_f[55]), .Z1_t (ciphertext_s1_t[55]), .Z1_f (ciphertext_s1_f[55]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S13reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS13ser[0]), .A0_f (new_AGEMA_signal_10853), .A1_t (new_AGEMA_signal_10854), .A1_f (new_AGEMA_signal_10855), .B0_t (ciphertext_s0_t[112]), .B0_f (ciphertext_s0_f[112]), .B1_t (ciphertext_s1_t[112]), .B1_f (ciphertext_s1_f[112]), .Z0_t (stateArray_S13reg_gff_1_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_10955), .Z1_t (new_AGEMA_signal_10956), .Z1_f (new_AGEMA_signal_10957) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S13reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S13reg_gff_1_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_10955), .B1_t (new_AGEMA_signal_10956), .B1_f (new_AGEMA_signal_10957), .Z0_t (stateArray_S13reg_gff_1_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_11075), .Z1_t (new_AGEMA_signal_11076), .Z1_f (new_AGEMA_signal_11077) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S13reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (stateArray_S13reg_gff_1_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_11075), .A1_t (new_AGEMA_signal_11076), .A1_f (new_AGEMA_signal_11077), .B0_t (stateArray_inS13ser[0]), .B0_f (new_AGEMA_signal_10853), .B1_t (new_AGEMA_signal_10854), .B1_f (new_AGEMA_signal_10855), .Z0_t (ciphertext_s0_t[16]), .Z0_f (ciphertext_s0_f[16]), .Z1_t (ciphertext_s1_t[16]), .Z1_f (ciphertext_s1_f[16]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S13reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS13ser[1]), .A0_f (new_AGEMA_signal_10994), .A1_t (new_AGEMA_signal_10995), .A1_f (new_AGEMA_signal_10996), .B0_t (ciphertext_s0_t[113]), .B0_f (ciphertext_s0_f[113]), .B1_t (ciphertext_s1_t[113]), .B1_f (ciphertext_s1_f[113]), .Z0_t (stateArray_S13reg_gff_1_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_11078), .Z1_t (new_AGEMA_signal_11079), .Z1_f (new_AGEMA_signal_11080) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S13reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S13reg_gff_1_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_11078), .B1_t (new_AGEMA_signal_11079), .B1_f (new_AGEMA_signal_11080), .Z0_t (stateArray_S13reg_gff_1_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_11144), .Z1_t (new_AGEMA_signal_11145), .Z1_f (new_AGEMA_signal_11146) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S13reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (stateArray_S13reg_gff_1_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_11144), .A1_t (new_AGEMA_signal_11145), .A1_f (new_AGEMA_signal_11146), .B0_t (stateArray_inS13ser[1]), .B0_f (new_AGEMA_signal_10994), .B1_t (new_AGEMA_signal_10995), .B1_f (new_AGEMA_signal_10996), .Z0_t (ciphertext_s0_t[17]), .Z0_f (ciphertext_s0_f[17]), .Z1_t (ciphertext_s1_t[17]), .Z1_f (ciphertext_s1_f[17]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S13reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS13ser[2]), .A0_f (new_AGEMA_signal_10859), .A1_t (new_AGEMA_signal_10860), .A1_f (new_AGEMA_signal_10861), .B0_t (ciphertext_s0_t[114]), .B0_f (ciphertext_s0_f[114]), .B1_t (ciphertext_s1_t[114]), .B1_f (ciphertext_s1_f[114]), .Z0_t (stateArray_S13reg_gff_1_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_10958), .Z1_t (new_AGEMA_signal_10959), .Z1_f (new_AGEMA_signal_10960) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S13reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S13reg_gff_1_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_10958), .B1_t (new_AGEMA_signal_10959), .B1_f (new_AGEMA_signal_10960), .Z0_t (stateArray_S13reg_gff_1_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_11081), .Z1_t (new_AGEMA_signal_11082), .Z1_f (new_AGEMA_signal_11083) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S13reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (stateArray_S13reg_gff_1_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_11081), .A1_t (new_AGEMA_signal_11082), .A1_f (new_AGEMA_signal_11083), .B0_t (stateArray_inS13ser[2]), .B0_f (new_AGEMA_signal_10859), .B1_t (new_AGEMA_signal_10860), .B1_f (new_AGEMA_signal_10861), .Z0_t (ciphertext_s0_t[18]), .Z0_f (ciphertext_s0_f[18]), .Z1_t (ciphertext_s1_t[18]), .Z1_f (ciphertext_s1_f[18]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S13reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS13ser[3]), .A0_f (new_AGEMA_signal_10997), .A1_t (new_AGEMA_signal_10998), .A1_f (new_AGEMA_signal_10999), .B0_t (ciphertext_s0_t[115]), .B0_f (ciphertext_s0_f[115]), .B1_t (ciphertext_s1_t[115]), .B1_f (ciphertext_s1_f[115]), .Z0_t (stateArray_S13reg_gff_1_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_11084), .Z1_t (new_AGEMA_signal_11085), .Z1_f (new_AGEMA_signal_11086) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S13reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S13reg_gff_1_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_11084), .B1_t (new_AGEMA_signal_11085), .B1_f (new_AGEMA_signal_11086), .Z0_t (stateArray_S13reg_gff_1_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_11147), .Z1_t (new_AGEMA_signal_11148), .Z1_f (new_AGEMA_signal_11149) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S13reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (stateArray_S13reg_gff_1_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_11147), .A1_t (new_AGEMA_signal_11148), .A1_f (new_AGEMA_signal_11149), .B0_t (stateArray_inS13ser[3]), .B0_f (new_AGEMA_signal_10997), .B1_t (new_AGEMA_signal_10998), .B1_f (new_AGEMA_signal_10999), .Z0_t (ciphertext_s0_t[19]), .Z0_f (ciphertext_s0_f[19]), .Z1_t (ciphertext_s1_t[19]), .Z1_f (ciphertext_s1_f[19]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S13reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS13ser[4]), .A0_f (new_AGEMA_signal_11000), .A1_t (new_AGEMA_signal_11001), .A1_f (new_AGEMA_signal_11002), .B0_t (ciphertext_s0_t[116]), .B0_f (ciphertext_s0_f[116]), .B1_t (ciphertext_s1_t[116]), .B1_f (ciphertext_s1_f[116]), .Z0_t (stateArray_S13reg_gff_1_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_11087), .Z1_t (new_AGEMA_signal_11088), .Z1_f (new_AGEMA_signal_11089) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S13reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S13reg_gff_1_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_11087), .B1_t (new_AGEMA_signal_11088), .B1_f (new_AGEMA_signal_11089), .Z0_t (stateArray_S13reg_gff_1_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_11150), .Z1_t (new_AGEMA_signal_11151), .Z1_f (new_AGEMA_signal_11152) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S13reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (stateArray_S13reg_gff_1_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_11150), .A1_t (new_AGEMA_signal_11151), .A1_f (new_AGEMA_signal_11152), .B0_t (stateArray_inS13ser[4]), .B0_f (new_AGEMA_signal_11000), .B1_t (new_AGEMA_signal_11001), .B1_f (new_AGEMA_signal_11002), .Z0_t (ciphertext_s0_t[20]), .Z0_f (ciphertext_s0_f[20]), .Z1_t (ciphertext_s1_t[20]), .Z1_f (ciphertext_s1_f[20]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S13reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS13ser[5]), .A0_f (new_AGEMA_signal_10868), .A1_t (new_AGEMA_signal_10869), .A1_f (new_AGEMA_signal_10870), .B0_t (ciphertext_s0_t[117]), .B0_f (ciphertext_s0_f[117]), .B1_t (ciphertext_s1_t[117]), .B1_f (ciphertext_s1_f[117]), .Z0_t (stateArray_S13reg_gff_1_SFF_5_MUXInst_X), .Z0_f (new_AGEMA_signal_10961), .Z1_t (new_AGEMA_signal_10962), .Z1_f (new_AGEMA_signal_10963) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S13reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S13reg_gff_1_SFF_5_MUXInst_X), .B0_f (new_AGEMA_signal_10961), .B1_t (new_AGEMA_signal_10962), .B1_f (new_AGEMA_signal_10963), .Z0_t (stateArray_S13reg_gff_1_SFF_5_MUXInst_Y), .Z0_f (new_AGEMA_signal_11090), .Z1_t (new_AGEMA_signal_11091), .Z1_f (new_AGEMA_signal_11092) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S13reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (stateArray_S13reg_gff_1_SFF_5_MUXInst_Y), .A0_f (new_AGEMA_signal_11090), .A1_t (new_AGEMA_signal_11091), .A1_f (new_AGEMA_signal_11092), .B0_t (stateArray_inS13ser[5]), .B0_f (new_AGEMA_signal_10868), .B1_t (new_AGEMA_signal_10869), .B1_f (new_AGEMA_signal_10870), .Z0_t (ciphertext_s0_t[21]), .Z0_f (ciphertext_s0_f[21]), .Z1_t (ciphertext_s1_t[21]), .Z1_f (ciphertext_s1_f[21]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S13reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS13ser[6]), .A0_f (new_AGEMA_signal_10871), .A1_t (new_AGEMA_signal_10872), .A1_f (new_AGEMA_signal_10873), .B0_t (ciphertext_s0_t[118]), .B0_f (ciphertext_s0_f[118]), .B1_t (ciphertext_s1_t[118]), .B1_f (ciphertext_s1_f[118]), .Z0_t (stateArray_S13reg_gff_1_SFF_6_MUXInst_X), .Z0_f (new_AGEMA_signal_10964), .Z1_t (new_AGEMA_signal_10965), .Z1_f (new_AGEMA_signal_10966) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S13reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S13reg_gff_1_SFF_6_MUXInst_X), .B0_f (new_AGEMA_signal_10964), .B1_t (new_AGEMA_signal_10965), .B1_f (new_AGEMA_signal_10966), .Z0_t (stateArray_S13reg_gff_1_SFF_6_MUXInst_Y), .Z0_f (new_AGEMA_signal_11093), .Z1_t (new_AGEMA_signal_11094), .Z1_f (new_AGEMA_signal_11095) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S13reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (stateArray_S13reg_gff_1_SFF_6_MUXInst_Y), .A0_f (new_AGEMA_signal_11093), .A1_t (new_AGEMA_signal_11094), .A1_f (new_AGEMA_signal_11095), .B0_t (stateArray_inS13ser[6]), .B0_f (new_AGEMA_signal_10871), .B1_t (new_AGEMA_signal_10872), .B1_f (new_AGEMA_signal_10873), .Z0_t (ciphertext_s0_t[22]), .Z0_f (ciphertext_s0_f[22]), .Z1_t (ciphertext_s1_t[22]), .Z1_f (ciphertext_s1_f[22]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S13reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS13ser[7]), .A0_f (new_AGEMA_signal_10874), .A1_t (new_AGEMA_signal_10875), .A1_f (new_AGEMA_signal_10876), .B0_t (ciphertext_s0_t[119]), .B0_f (ciphertext_s0_f[119]), .B1_t (ciphertext_s1_t[119]), .B1_f (ciphertext_s1_f[119]), .Z0_t (stateArray_S13reg_gff_1_SFF_7_MUXInst_X), .Z0_f (new_AGEMA_signal_10967), .Z1_t (new_AGEMA_signal_10968), .Z1_f (new_AGEMA_signal_10969) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S13reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S13reg_gff_1_SFF_7_MUXInst_X), .B0_f (new_AGEMA_signal_10967), .B1_t (new_AGEMA_signal_10968), .B1_f (new_AGEMA_signal_10969), .Z0_t (stateArray_S13reg_gff_1_SFF_7_MUXInst_Y), .Z0_f (new_AGEMA_signal_11096), .Z1_t (new_AGEMA_signal_11097), .Z1_f (new_AGEMA_signal_11098) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S13reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (stateArray_S13reg_gff_1_SFF_7_MUXInst_Y), .A0_f (new_AGEMA_signal_11096), .A1_t (new_AGEMA_signal_11097), .A1_f (new_AGEMA_signal_11098), .B0_t (stateArray_inS13ser[7]), .B0_f (new_AGEMA_signal_10874), .B1_t (new_AGEMA_signal_10875), .B1_f (new_AGEMA_signal_10876), .Z0_t (ciphertext_s0_t[23]), .Z0_f (ciphertext_s0_f[23]), .Z1_t (ciphertext_s1_t[23]), .Z1_f (ciphertext_s1_f[23]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S20reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS20ser[0]), .A0_f (new_AGEMA_signal_6766), .A1_t (new_AGEMA_signal_6767), .A1_f (new_AGEMA_signal_6768), .B0_t (ciphertext_s0_t[40]), .B0_f (ciphertext_s0_f[40]), .B1_t (ciphertext_s1_t[40]), .B1_f (ciphertext_s1_f[40]), .Z0_t (stateArray_S20reg_gff_1_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_7539), .Z1_t (new_AGEMA_signal_7540), .Z1_f (new_AGEMA_signal_7541) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S20reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S20reg_gff_1_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_7539), .B1_t (new_AGEMA_signal_7540), .B1_f (new_AGEMA_signal_7541), .Z0_t (stateArray_S20reg_gff_1_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_8286), .Z1_t (new_AGEMA_signal_8287), .Z1_f (new_AGEMA_signal_8288) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S20reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (stateArray_S20reg_gff_1_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_8286), .A1_t (new_AGEMA_signal_8287), .A1_f (new_AGEMA_signal_8288), .B0_t (stateArray_inS20ser[0]), .B0_f (new_AGEMA_signal_6766), .B1_t (new_AGEMA_signal_6767), .B1_f (new_AGEMA_signal_6768), .Z0_t (ciphertext_s0_t[104]), .Z0_f (ciphertext_s0_f[104]), .Z1_t (ciphertext_s1_t[104]), .Z1_f (ciphertext_s1_f[104]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S20reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS20ser[1]), .A0_f (new_AGEMA_signal_6769), .A1_t (new_AGEMA_signal_6770), .A1_f (new_AGEMA_signal_6771), .B0_t (ciphertext_s0_t[41]), .B0_f (ciphertext_s0_f[41]), .B1_t (ciphertext_s1_t[41]), .B1_f (ciphertext_s1_f[41]), .Z0_t (stateArray_S20reg_gff_1_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_7542), .Z1_t (new_AGEMA_signal_7543), .Z1_f (new_AGEMA_signal_7544) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S20reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S20reg_gff_1_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_7542), .B1_t (new_AGEMA_signal_7543), .B1_f (new_AGEMA_signal_7544), .Z0_t (stateArray_S20reg_gff_1_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_8289), .Z1_t (new_AGEMA_signal_8290), .Z1_f (new_AGEMA_signal_8291) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S20reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (stateArray_S20reg_gff_1_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_8289), .A1_t (new_AGEMA_signal_8290), .A1_f (new_AGEMA_signal_8291), .B0_t (stateArray_inS20ser[1]), .B0_f (new_AGEMA_signal_6769), .B1_t (new_AGEMA_signal_6770), .B1_f (new_AGEMA_signal_6771), .Z0_t (ciphertext_s0_t[105]), .Z0_f (ciphertext_s0_f[105]), .Z1_t (ciphertext_s1_t[105]), .Z1_f (ciphertext_s1_f[105]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S20reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS20ser[2]), .A0_f (new_AGEMA_signal_6772), .A1_t (new_AGEMA_signal_6773), .A1_f (new_AGEMA_signal_6774), .B0_t (ciphertext_s0_t[42]), .B0_f (ciphertext_s0_f[42]), .B1_t (ciphertext_s1_t[42]), .B1_f (ciphertext_s1_f[42]), .Z0_t (stateArray_S20reg_gff_1_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_7545), .Z1_t (new_AGEMA_signal_7546), .Z1_f (new_AGEMA_signal_7547) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S20reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S20reg_gff_1_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_7545), .B1_t (new_AGEMA_signal_7546), .B1_f (new_AGEMA_signal_7547), .Z0_t (stateArray_S20reg_gff_1_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_8292), .Z1_t (new_AGEMA_signal_8293), .Z1_f (new_AGEMA_signal_8294) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S20reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (stateArray_S20reg_gff_1_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_8292), .A1_t (new_AGEMA_signal_8293), .A1_f (new_AGEMA_signal_8294), .B0_t (stateArray_inS20ser[2]), .B0_f (new_AGEMA_signal_6772), .B1_t (new_AGEMA_signal_6773), .B1_f (new_AGEMA_signal_6774), .Z0_t (ciphertext_s0_t[106]), .Z0_f (ciphertext_s0_f[106]), .Z1_t (ciphertext_s1_t[106]), .Z1_f (ciphertext_s1_f[106]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S20reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS20ser[3]), .A0_f (new_AGEMA_signal_6775), .A1_t (new_AGEMA_signal_6776), .A1_f (new_AGEMA_signal_6777), .B0_t (ciphertext_s0_t[43]), .B0_f (ciphertext_s0_f[43]), .B1_t (ciphertext_s1_t[43]), .B1_f (ciphertext_s1_f[43]), .Z0_t (stateArray_S20reg_gff_1_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_7548), .Z1_t (new_AGEMA_signal_7549), .Z1_f (new_AGEMA_signal_7550) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S20reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S20reg_gff_1_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_7548), .B1_t (new_AGEMA_signal_7549), .B1_f (new_AGEMA_signal_7550), .Z0_t (stateArray_S20reg_gff_1_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_8295), .Z1_t (new_AGEMA_signal_8296), .Z1_f (new_AGEMA_signal_8297) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S20reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (stateArray_S20reg_gff_1_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_8295), .A1_t (new_AGEMA_signal_8296), .A1_f (new_AGEMA_signal_8297), .B0_t (stateArray_inS20ser[3]), .B0_f (new_AGEMA_signal_6775), .B1_t (new_AGEMA_signal_6776), .B1_f (new_AGEMA_signal_6777), .Z0_t (ciphertext_s0_t[107]), .Z0_f (ciphertext_s0_f[107]), .Z1_t (ciphertext_s1_t[107]), .Z1_f (ciphertext_s1_f[107]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S20reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS20ser[4]), .A0_f (new_AGEMA_signal_6778), .A1_t (new_AGEMA_signal_6779), .A1_f (new_AGEMA_signal_6780), .B0_t (ciphertext_s0_t[44]), .B0_f (ciphertext_s0_f[44]), .B1_t (ciphertext_s1_t[44]), .B1_f (ciphertext_s1_f[44]), .Z0_t (stateArray_S20reg_gff_1_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_7551), .Z1_t (new_AGEMA_signal_7552), .Z1_f (new_AGEMA_signal_7553) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S20reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S20reg_gff_1_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_7551), .B1_t (new_AGEMA_signal_7552), .B1_f (new_AGEMA_signal_7553), .Z0_t (stateArray_S20reg_gff_1_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_8298), .Z1_t (new_AGEMA_signal_8299), .Z1_f (new_AGEMA_signal_8300) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S20reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (stateArray_S20reg_gff_1_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_8298), .A1_t (new_AGEMA_signal_8299), .A1_f (new_AGEMA_signal_8300), .B0_t (stateArray_inS20ser[4]), .B0_f (new_AGEMA_signal_6778), .B1_t (new_AGEMA_signal_6779), .B1_f (new_AGEMA_signal_6780), .Z0_t (ciphertext_s0_t[108]), .Z0_f (ciphertext_s0_f[108]), .Z1_t (ciphertext_s1_t[108]), .Z1_f (ciphertext_s1_f[108]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S20reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS20ser[5]), .A0_f (new_AGEMA_signal_6781), .A1_t (new_AGEMA_signal_6782), .A1_f (new_AGEMA_signal_6783), .B0_t (ciphertext_s0_t[45]), .B0_f (ciphertext_s0_f[45]), .B1_t (ciphertext_s1_t[45]), .B1_f (ciphertext_s1_f[45]), .Z0_t (stateArray_S20reg_gff_1_SFF_5_MUXInst_X), .Z0_f (new_AGEMA_signal_7554), .Z1_t (new_AGEMA_signal_7555), .Z1_f (new_AGEMA_signal_7556) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S20reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S20reg_gff_1_SFF_5_MUXInst_X), .B0_f (new_AGEMA_signal_7554), .B1_t (new_AGEMA_signal_7555), .B1_f (new_AGEMA_signal_7556), .Z0_t (stateArray_S20reg_gff_1_SFF_5_MUXInst_Y), .Z0_f (new_AGEMA_signal_8301), .Z1_t (new_AGEMA_signal_8302), .Z1_f (new_AGEMA_signal_8303) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S20reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (stateArray_S20reg_gff_1_SFF_5_MUXInst_Y), .A0_f (new_AGEMA_signal_8301), .A1_t (new_AGEMA_signal_8302), .A1_f (new_AGEMA_signal_8303), .B0_t (stateArray_inS20ser[5]), .B0_f (new_AGEMA_signal_6781), .B1_t (new_AGEMA_signal_6782), .B1_f (new_AGEMA_signal_6783), .Z0_t (ciphertext_s0_t[109]), .Z0_f (ciphertext_s0_f[109]), .Z1_t (ciphertext_s1_t[109]), .Z1_f (ciphertext_s1_f[109]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S20reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS20ser[6]), .A0_f (new_AGEMA_signal_6784), .A1_t (new_AGEMA_signal_6785), .A1_f (new_AGEMA_signal_6786), .B0_t (ciphertext_s0_t[46]), .B0_f (ciphertext_s0_f[46]), .B1_t (ciphertext_s1_t[46]), .B1_f (ciphertext_s1_f[46]), .Z0_t (stateArray_S20reg_gff_1_SFF_6_MUXInst_X), .Z0_f (new_AGEMA_signal_7557), .Z1_t (new_AGEMA_signal_7558), .Z1_f (new_AGEMA_signal_7559) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S20reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S20reg_gff_1_SFF_6_MUXInst_X), .B0_f (new_AGEMA_signal_7557), .B1_t (new_AGEMA_signal_7558), .B1_f (new_AGEMA_signal_7559), .Z0_t (stateArray_S20reg_gff_1_SFF_6_MUXInst_Y), .Z0_f (new_AGEMA_signal_8304), .Z1_t (new_AGEMA_signal_8305), .Z1_f (new_AGEMA_signal_8306) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S20reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (stateArray_S20reg_gff_1_SFF_6_MUXInst_Y), .A0_f (new_AGEMA_signal_8304), .A1_t (new_AGEMA_signal_8305), .A1_f (new_AGEMA_signal_8306), .B0_t (stateArray_inS20ser[6]), .B0_f (new_AGEMA_signal_6784), .B1_t (new_AGEMA_signal_6785), .B1_f (new_AGEMA_signal_6786), .Z0_t (ciphertext_s0_t[110]), .Z0_f (ciphertext_s0_f[110]), .Z1_t (ciphertext_s1_t[110]), .Z1_f (ciphertext_s1_f[110]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S20reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS20ser[7]), .A0_f (new_AGEMA_signal_6787), .A1_t (new_AGEMA_signal_6788), .A1_f (new_AGEMA_signal_6789), .B0_t (ciphertext_s0_t[47]), .B0_f (ciphertext_s0_f[47]), .B1_t (ciphertext_s1_t[47]), .B1_f (ciphertext_s1_f[47]), .Z0_t (stateArray_S20reg_gff_1_SFF_7_MUXInst_X), .Z0_f (new_AGEMA_signal_7560), .Z1_t (new_AGEMA_signal_7561), .Z1_f (new_AGEMA_signal_7562) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S20reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S20reg_gff_1_SFF_7_MUXInst_X), .B0_f (new_AGEMA_signal_7560), .B1_t (new_AGEMA_signal_7561), .B1_f (new_AGEMA_signal_7562), .Z0_t (stateArray_S20reg_gff_1_SFF_7_MUXInst_Y), .Z0_f (new_AGEMA_signal_8307), .Z1_t (new_AGEMA_signal_8308), .Z1_f (new_AGEMA_signal_8309) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S20reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (stateArray_S20reg_gff_1_SFF_7_MUXInst_Y), .A0_f (new_AGEMA_signal_8307), .A1_t (new_AGEMA_signal_8308), .A1_f (new_AGEMA_signal_8309), .B0_t (stateArray_inS20ser[7]), .B0_f (new_AGEMA_signal_6787), .B1_t (new_AGEMA_signal_6788), .B1_f (new_AGEMA_signal_6789), .Z0_t (ciphertext_s0_t[111]), .Z0_f (ciphertext_s0_f[111]), .Z1_t (ciphertext_s1_t[111]), .Z1_f (ciphertext_s1_f[111]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S21reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS21ser[0]), .A0_f (new_AGEMA_signal_6790), .A1_t (new_AGEMA_signal_6791), .A1_f (new_AGEMA_signal_6792), .B0_t (ciphertext_s0_t[8]), .B0_f (ciphertext_s0_f[8]), .B1_t (ciphertext_s1_t[8]), .B1_f (ciphertext_s1_f[8]), .Z0_t (stateArray_S21reg_gff_1_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_7563), .Z1_t (new_AGEMA_signal_7564), .Z1_f (new_AGEMA_signal_7565) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S21reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S21reg_gff_1_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_7563), .B1_t (new_AGEMA_signal_7564), .B1_f (new_AGEMA_signal_7565), .Z0_t (stateArray_S21reg_gff_1_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_8310), .Z1_t (new_AGEMA_signal_8311), .Z1_f (new_AGEMA_signal_8312) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S21reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (stateArray_S21reg_gff_1_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_8310), .A1_t (new_AGEMA_signal_8311), .A1_f (new_AGEMA_signal_8312), .B0_t (stateArray_inS21ser[0]), .B0_f (new_AGEMA_signal_6790), .B1_t (new_AGEMA_signal_6791), .B1_f (new_AGEMA_signal_6792), .Z0_t (ciphertext_s0_t[72]), .Z0_f (ciphertext_s0_f[72]), .Z1_t (ciphertext_s1_t[72]), .Z1_f (ciphertext_s1_f[72]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S21reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS21ser[1]), .A0_f (new_AGEMA_signal_6793), .A1_t (new_AGEMA_signal_6794), .A1_f (new_AGEMA_signal_6795), .B0_t (ciphertext_s0_t[9]), .B0_f (ciphertext_s0_f[9]), .B1_t (ciphertext_s1_t[9]), .B1_f (ciphertext_s1_f[9]), .Z0_t (stateArray_S21reg_gff_1_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_7566), .Z1_t (new_AGEMA_signal_7567), .Z1_f (new_AGEMA_signal_7568) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S21reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S21reg_gff_1_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_7566), .B1_t (new_AGEMA_signal_7567), .B1_f (new_AGEMA_signal_7568), .Z0_t (stateArray_S21reg_gff_1_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_8313), .Z1_t (new_AGEMA_signal_8314), .Z1_f (new_AGEMA_signal_8315) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S21reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (stateArray_S21reg_gff_1_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_8313), .A1_t (new_AGEMA_signal_8314), .A1_f (new_AGEMA_signal_8315), .B0_t (stateArray_inS21ser[1]), .B0_f (new_AGEMA_signal_6793), .B1_t (new_AGEMA_signal_6794), .B1_f (new_AGEMA_signal_6795), .Z0_t (ciphertext_s0_t[73]), .Z0_f (ciphertext_s0_f[73]), .Z1_t (ciphertext_s1_t[73]), .Z1_f (ciphertext_s1_f[73]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S21reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS21ser[2]), .A0_f (new_AGEMA_signal_6796), .A1_t (new_AGEMA_signal_6797), .A1_f (new_AGEMA_signal_6798), .B0_t (ciphertext_s0_t[10]), .B0_f (ciphertext_s0_f[10]), .B1_t (ciphertext_s1_t[10]), .B1_f (ciphertext_s1_f[10]), .Z0_t (stateArray_S21reg_gff_1_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_7569), .Z1_t (new_AGEMA_signal_7570), .Z1_f (new_AGEMA_signal_7571) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S21reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S21reg_gff_1_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_7569), .B1_t (new_AGEMA_signal_7570), .B1_f (new_AGEMA_signal_7571), .Z0_t (stateArray_S21reg_gff_1_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_8316), .Z1_t (new_AGEMA_signal_8317), .Z1_f (new_AGEMA_signal_8318) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S21reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (stateArray_S21reg_gff_1_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_8316), .A1_t (new_AGEMA_signal_8317), .A1_f (new_AGEMA_signal_8318), .B0_t (stateArray_inS21ser[2]), .B0_f (new_AGEMA_signal_6796), .B1_t (new_AGEMA_signal_6797), .B1_f (new_AGEMA_signal_6798), .Z0_t (ciphertext_s0_t[74]), .Z0_f (ciphertext_s0_f[74]), .Z1_t (ciphertext_s1_t[74]), .Z1_f (ciphertext_s1_f[74]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S21reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS21ser[3]), .A0_f (new_AGEMA_signal_6799), .A1_t (new_AGEMA_signal_6800), .A1_f (new_AGEMA_signal_6801), .B0_t (ciphertext_s0_t[11]), .B0_f (ciphertext_s0_f[11]), .B1_t (ciphertext_s1_t[11]), .B1_f (ciphertext_s1_f[11]), .Z0_t (stateArray_S21reg_gff_1_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_7572), .Z1_t (new_AGEMA_signal_7573), .Z1_f (new_AGEMA_signal_7574) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S21reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S21reg_gff_1_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_7572), .B1_t (new_AGEMA_signal_7573), .B1_f (new_AGEMA_signal_7574), .Z0_t (stateArray_S21reg_gff_1_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_8319), .Z1_t (new_AGEMA_signal_8320), .Z1_f (new_AGEMA_signal_8321) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S21reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (stateArray_S21reg_gff_1_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_8319), .A1_t (new_AGEMA_signal_8320), .A1_f (new_AGEMA_signal_8321), .B0_t (stateArray_inS21ser[3]), .B0_f (new_AGEMA_signal_6799), .B1_t (new_AGEMA_signal_6800), .B1_f (new_AGEMA_signal_6801), .Z0_t (ciphertext_s0_t[75]), .Z0_f (ciphertext_s0_f[75]), .Z1_t (ciphertext_s1_t[75]), .Z1_f (ciphertext_s1_f[75]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S21reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS21ser[4]), .A0_f (new_AGEMA_signal_6802), .A1_t (new_AGEMA_signal_6803), .A1_f (new_AGEMA_signal_6804), .B0_t (ciphertext_s0_t[12]), .B0_f (ciphertext_s0_f[12]), .B1_t (ciphertext_s1_t[12]), .B1_f (ciphertext_s1_f[12]), .Z0_t (stateArray_S21reg_gff_1_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_7575), .Z1_t (new_AGEMA_signal_7576), .Z1_f (new_AGEMA_signal_7577) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S21reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S21reg_gff_1_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_7575), .B1_t (new_AGEMA_signal_7576), .B1_f (new_AGEMA_signal_7577), .Z0_t (stateArray_S21reg_gff_1_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_8322), .Z1_t (new_AGEMA_signal_8323), .Z1_f (new_AGEMA_signal_8324) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S21reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (stateArray_S21reg_gff_1_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_8322), .A1_t (new_AGEMA_signal_8323), .A1_f (new_AGEMA_signal_8324), .B0_t (stateArray_inS21ser[4]), .B0_f (new_AGEMA_signal_6802), .B1_t (new_AGEMA_signal_6803), .B1_f (new_AGEMA_signal_6804), .Z0_t (ciphertext_s0_t[76]), .Z0_f (ciphertext_s0_f[76]), .Z1_t (ciphertext_s1_t[76]), .Z1_f (ciphertext_s1_f[76]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S21reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS21ser[5]), .A0_f (new_AGEMA_signal_6805), .A1_t (new_AGEMA_signal_6806), .A1_f (new_AGEMA_signal_6807), .B0_t (ciphertext_s0_t[13]), .B0_f (ciphertext_s0_f[13]), .B1_t (ciphertext_s1_t[13]), .B1_f (ciphertext_s1_f[13]), .Z0_t (stateArray_S21reg_gff_1_SFF_5_MUXInst_X), .Z0_f (new_AGEMA_signal_7578), .Z1_t (new_AGEMA_signal_7579), .Z1_f (new_AGEMA_signal_7580) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S21reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S21reg_gff_1_SFF_5_MUXInst_X), .B0_f (new_AGEMA_signal_7578), .B1_t (new_AGEMA_signal_7579), .B1_f (new_AGEMA_signal_7580), .Z0_t (stateArray_S21reg_gff_1_SFF_5_MUXInst_Y), .Z0_f (new_AGEMA_signal_8325), .Z1_t (new_AGEMA_signal_8326), .Z1_f (new_AGEMA_signal_8327) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S21reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (stateArray_S21reg_gff_1_SFF_5_MUXInst_Y), .A0_f (new_AGEMA_signal_8325), .A1_t (new_AGEMA_signal_8326), .A1_f (new_AGEMA_signal_8327), .B0_t (stateArray_inS21ser[5]), .B0_f (new_AGEMA_signal_6805), .B1_t (new_AGEMA_signal_6806), .B1_f (new_AGEMA_signal_6807), .Z0_t (ciphertext_s0_t[77]), .Z0_f (ciphertext_s0_f[77]), .Z1_t (ciphertext_s1_t[77]), .Z1_f (ciphertext_s1_f[77]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S21reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS21ser[6]), .A0_f (new_AGEMA_signal_6808), .A1_t (new_AGEMA_signal_6809), .A1_f (new_AGEMA_signal_6810), .B0_t (ciphertext_s0_t[14]), .B0_f (ciphertext_s0_f[14]), .B1_t (ciphertext_s1_t[14]), .B1_f (ciphertext_s1_f[14]), .Z0_t (stateArray_S21reg_gff_1_SFF_6_MUXInst_X), .Z0_f (new_AGEMA_signal_7581), .Z1_t (new_AGEMA_signal_7582), .Z1_f (new_AGEMA_signal_7583) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S21reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S21reg_gff_1_SFF_6_MUXInst_X), .B0_f (new_AGEMA_signal_7581), .B1_t (new_AGEMA_signal_7582), .B1_f (new_AGEMA_signal_7583), .Z0_t (stateArray_S21reg_gff_1_SFF_6_MUXInst_Y), .Z0_f (new_AGEMA_signal_8328), .Z1_t (new_AGEMA_signal_8329), .Z1_f (new_AGEMA_signal_8330) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S21reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (stateArray_S21reg_gff_1_SFF_6_MUXInst_Y), .A0_f (new_AGEMA_signal_8328), .A1_t (new_AGEMA_signal_8329), .A1_f (new_AGEMA_signal_8330), .B0_t (stateArray_inS21ser[6]), .B0_f (new_AGEMA_signal_6808), .B1_t (new_AGEMA_signal_6809), .B1_f (new_AGEMA_signal_6810), .Z0_t (ciphertext_s0_t[78]), .Z0_f (ciphertext_s0_f[78]), .Z1_t (ciphertext_s1_t[78]), .Z1_f (ciphertext_s1_f[78]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S21reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS21ser[7]), .A0_f (new_AGEMA_signal_6811), .A1_t (new_AGEMA_signal_6812), .A1_f (new_AGEMA_signal_6813), .B0_t (ciphertext_s0_t[15]), .B0_f (ciphertext_s0_f[15]), .B1_t (ciphertext_s1_t[15]), .B1_f (ciphertext_s1_f[15]), .Z0_t (stateArray_S21reg_gff_1_SFF_7_MUXInst_X), .Z0_f (new_AGEMA_signal_7584), .Z1_t (new_AGEMA_signal_7585), .Z1_f (new_AGEMA_signal_7586) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S21reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S21reg_gff_1_SFF_7_MUXInst_X), .B0_f (new_AGEMA_signal_7584), .B1_t (new_AGEMA_signal_7585), .B1_f (new_AGEMA_signal_7586), .Z0_t (stateArray_S21reg_gff_1_SFF_7_MUXInst_Y), .Z0_f (new_AGEMA_signal_8331), .Z1_t (new_AGEMA_signal_8332), .Z1_f (new_AGEMA_signal_8333) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S21reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (stateArray_S21reg_gff_1_SFF_7_MUXInst_Y), .A0_f (new_AGEMA_signal_8331), .A1_t (new_AGEMA_signal_8332), .A1_f (new_AGEMA_signal_8333), .B0_t (stateArray_inS21ser[7]), .B0_f (new_AGEMA_signal_6811), .B1_t (new_AGEMA_signal_6812), .B1_f (new_AGEMA_signal_6813), .Z0_t (ciphertext_s0_t[79]), .Z0_f (ciphertext_s0_f[79]), .Z1_t (ciphertext_s1_t[79]), .Z1_f (ciphertext_s1_f[79]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S22reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS22ser[0]), .A0_f (new_AGEMA_signal_6814), .A1_t (new_AGEMA_signal_6815), .A1_f (new_AGEMA_signal_6816), .B0_t (ciphertext_s0_t[104]), .B0_f (ciphertext_s0_f[104]), .B1_t (ciphertext_s1_t[104]), .B1_f (ciphertext_s1_f[104]), .Z0_t (stateArray_S22reg_gff_1_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_7587), .Z1_t (new_AGEMA_signal_7588), .Z1_f (new_AGEMA_signal_7589) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S22reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S22reg_gff_1_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_7587), .B1_t (new_AGEMA_signal_7588), .B1_f (new_AGEMA_signal_7589), .Z0_t (stateArray_S22reg_gff_1_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_8334), .Z1_t (new_AGEMA_signal_8335), .Z1_f (new_AGEMA_signal_8336) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S22reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (stateArray_S22reg_gff_1_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_8334), .A1_t (new_AGEMA_signal_8335), .A1_f (new_AGEMA_signal_8336), .B0_t (stateArray_inS22ser[0]), .B0_f (new_AGEMA_signal_6814), .B1_t (new_AGEMA_signal_6815), .B1_f (new_AGEMA_signal_6816), .Z0_t (ciphertext_s0_t[40]), .Z0_f (ciphertext_s0_f[40]), .Z1_t (ciphertext_s1_t[40]), .Z1_f (ciphertext_s1_f[40]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S22reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS22ser[1]), .A0_f (new_AGEMA_signal_6817), .A1_t (new_AGEMA_signal_6818), .A1_f (new_AGEMA_signal_6819), .B0_t (ciphertext_s0_t[105]), .B0_f (ciphertext_s0_f[105]), .B1_t (ciphertext_s1_t[105]), .B1_f (ciphertext_s1_f[105]), .Z0_t (stateArray_S22reg_gff_1_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_7590), .Z1_t (new_AGEMA_signal_7591), .Z1_f (new_AGEMA_signal_7592) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S22reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S22reg_gff_1_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_7590), .B1_t (new_AGEMA_signal_7591), .B1_f (new_AGEMA_signal_7592), .Z0_t (stateArray_S22reg_gff_1_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_8337), .Z1_t (new_AGEMA_signal_8338), .Z1_f (new_AGEMA_signal_8339) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S22reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (stateArray_S22reg_gff_1_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_8337), .A1_t (new_AGEMA_signal_8338), .A1_f (new_AGEMA_signal_8339), .B0_t (stateArray_inS22ser[1]), .B0_f (new_AGEMA_signal_6817), .B1_t (new_AGEMA_signal_6818), .B1_f (new_AGEMA_signal_6819), .Z0_t (ciphertext_s0_t[41]), .Z0_f (ciphertext_s0_f[41]), .Z1_t (ciphertext_s1_t[41]), .Z1_f (ciphertext_s1_f[41]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S22reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS22ser[2]), .A0_f (new_AGEMA_signal_6820), .A1_t (new_AGEMA_signal_6821), .A1_f (new_AGEMA_signal_6822), .B0_t (ciphertext_s0_t[106]), .B0_f (ciphertext_s0_f[106]), .B1_t (ciphertext_s1_t[106]), .B1_f (ciphertext_s1_f[106]), .Z0_t (stateArray_S22reg_gff_1_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_7593), .Z1_t (new_AGEMA_signal_7594), .Z1_f (new_AGEMA_signal_7595) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S22reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S22reg_gff_1_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_7593), .B1_t (new_AGEMA_signal_7594), .B1_f (new_AGEMA_signal_7595), .Z0_t (stateArray_S22reg_gff_1_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_8340), .Z1_t (new_AGEMA_signal_8341), .Z1_f (new_AGEMA_signal_8342) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S22reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (stateArray_S22reg_gff_1_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_8340), .A1_t (new_AGEMA_signal_8341), .A1_f (new_AGEMA_signal_8342), .B0_t (stateArray_inS22ser[2]), .B0_f (new_AGEMA_signal_6820), .B1_t (new_AGEMA_signal_6821), .B1_f (new_AGEMA_signal_6822), .Z0_t (ciphertext_s0_t[42]), .Z0_f (ciphertext_s0_f[42]), .Z1_t (ciphertext_s1_t[42]), .Z1_f (ciphertext_s1_f[42]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S22reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS22ser[3]), .A0_f (new_AGEMA_signal_6823), .A1_t (new_AGEMA_signal_6824), .A1_f (new_AGEMA_signal_6825), .B0_t (ciphertext_s0_t[107]), .B0_f (ciphertext_s0_f[107]), .B1_t (ciphertext_s1_t[107]), .B1_f (ciphertext_s1_f[107]), .Z0_t (stateArray_S22reg_gff_1_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_7596), .Z1_t (new_AGEMA_signal_7597), .Z1_f (new_AGEMA_signal_7598) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S22reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S22reg_gff_1_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_7596), .B1_t (new_AGEMA_signal_7597), .B1_f (new_AGEMA_signal_7598), .Z0_t (stateArray_S22reg_gff_1_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_8343), .Z1_t (new_AGEMA_signal_8344), .Z1_f (new_AGEMA_signal_8345) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S22reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (stateArray_S22reg_gff_1_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_8343), .A1_t (new_AGEMA_signal_8344), .A1_f (new_AGEMA_signal_8345), .B0_t (stateArray_inS22ser[3]), .B0_f (new_AGEMA_signal_6823), .B1_t (new_AGEMA_signal_6824), .B1_f (new_AGEMA_signal_6825), .Z0_t (ciphertext_s0_t[43]), .Z0_f (ciphertext_s0_f[43]), .Z1_t (ciphertext_s1_t[43]), .Z1_f (ciphertext_s1_f[43]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S22reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS22ser[4]), .A0_f (new_AGEMA_signal_6826), .A1_t (new_AGEMA_signal_6827), .A1_f (new_AGEMA_signal_6828), .B0_t (ciphertext_s0_t[108]), .B0_f (ciphertext_s0_f[108]), .B1_t (ciphertext_s1_t[108]), .B1_f (ciphertext_s1_f[108]), .Z0_t (stateArray_S22reg_gff_1_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_7599), .Z1_t (new_AGEMA_signal_7600), .Z1_f (new_AGEMA_signal_7601) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S22reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S22reg_gff_1_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_7599), .B1_t (new_AGEMA_signal_7600), .B1_f (new_AGEMA_signal_7601), .Z0_t (stateArray_S22reg_gff_1_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_8346), .Z1_t (new_AGEMA_signal_8347), .Z1_f (new_AGEMA_signal_8348) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S22reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (stateArray_S22reg_gff_1_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_8346), .A1_t (new_AGEMA_signal_8347), .A1_f (new_AGEMA_signal_8348), .B0_t (stateArray_inS22ser[4]), .B0_f (new_AGEMA_signal_6826), .B1_t (new_AGEMA_signal_6827), .B1_f (new_AGEMA_signal_6828), .Z0_t (ciphertext_s0_t[44]), .Z0_f (ciphertext_s0_f[44]), .Z1_t (ciphertext_s1_t[44]), .Z1_f (ciphertext_s1_f[44]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S22reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS22ser[5]), .A0_f (new_AGEMA_signal_6829), .A1_t (new_AGEMA_signal_6830), .A1_f (new_AGEMA_signal_6831), .B0_t (ciphertext_s0_t[109]), .B0_f (ciphertext_s0_f[109]), .B1_t (ciphertext_s1_t[109]), .B1_f (ciphertext_s1_f[109]), .Z0_t (stateArray_S22reg_gff_1_SFF_5_MUXInst_X), .Z0_f (new_AGEMA_signal_7602), .Z1_t (new_AGEMA_signal_7603), .Z1_f (new_AGEMA_signal_7604) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S22reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S22reg_gff_1_SFF_5_MUXInst_X), .B0_f (new_AGEMA_signal_7602), .B1_t (new_AGEMA_signal_7603), .B1_f (new_AGEMA_signal_7604), .Z0_t (stateArray_S22reg_gff_1_SFF_5_MUXInst_Y), .Z0_f (new_AGEMA_signal_8349), .Z1_t (new_AGEMA_signal_8350), .Z1_f (new_AGEMA_signal_8351) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S22reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (stateArray_S22reg_gff_1_SFF_5_MUXInst_Y), .A0_f (new_AGEMA_signal_8349), .A1_t (new_AGEMA_signal_8350), .A1_f (new_AGEMA_signal_8351), .B0_t (stateArray_inS22ser[5]), .B0_f (new_AGEMA_signal_6829), .B1_t (new_AGEMA_signal_6830), .B1_f (new_AGEMA_signal_6831), .Z0_t (ciphertext_s0_t[45]), .Z0_f (ciphertext_s0_f[45]), .Z1_t (ciphertext_s1_t[45]), .Z1_f (ciphertext_s1_f[45]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S22reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS22ser[6]), .A0_f (new_AGEMA_signal_6832), .A1_t (new_AGEMA_signal_6833), .A1_f (new_AGEMA_signal_6834), .B0_t (ciphertext_s0_t[110]), .B0_f (ciphertext_s0_f[110]), .B1_t (ciphertext_s1_t[110]), .B1_f (ciphertext_s1_f[110]), .Z0_t (stateArray_S22reg_gff_1_SFF_6_MUXInst_X), .Z0_f (new_AGEMA_signal_7605), .Z1_t (new_AGEMA_signal_7606), .Z1_f (new_AGEMA_signal_7607) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S22reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S22reg_gff_1_SFF_6_MUXInst_X), .B0_f (new_AGEMA_signal_7605), .B1_t (new_AGEMA_signal_7606), .B1_f (new_AGEMA_signal_7607), .Z0_t (stateArray_S22reg_gff_1_SFF_6_MUXInst_Y), .Z0_f (new_AGEMA_signal_8352), .Z1_t (new_AGEMA_signal_8353), .Z1_f (new_AGEMA_signal_8354) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S22reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (stateArray_S22reg_gff_1_SFF_6_MUXInst_Y), .A0_f (new_AGEMA_signal_8352), .A1_t (new_AGEMA_signal_8353), .A1_f (new_AGEMA_signal_8354), .B0_t (stateArray_inS22ser[6]), .B0_f (new_AGEMA_signal_6832), .B1_t (new_AGEMA_signal_6833), .B1_f (new_AGEMA_signal_6834), .Z0_t (ciphertext_s0_t[46]), .Z0_f (ciphertext_s0_f[46]), .Z1_t (ciphertext_s1_t[46]), .Z1_f (ciphertext_s1_f[46]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S22reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS22ser[7]), .A0_f (new_AGEMA_signal_6835), .A1_t (new_AGEMA_signal_6836), .A1_f (new_AGEMA_signal_6837), .B0_t (ciphertext_s0_t[111]), .B0_f (ciphertext_s0_f[111]), .B1_t (ciphertext_s1_t[111]), .B1_f (ciphertext_s1_f[111]), .Z0_t (stateArray_S22reg_gff_1_SFF_7_MUXInst_X), .Z0_f (new_AGEMA_signal_7608), .Z1_t (new_AGEMA_signal_7609), .Z1_f (new_AGEMA_signal_7610) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S22reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S22reg_gff_1_SFF_7_MUXInst_X), .B0_f (new_AGEMA_signal_7608), .B1_t (new_AGEMA_signal_7609), .B1_f (new_AGEMA_signal_7610), .Z0_t (stateArray_S22reg_gff_1_SFF_7_MUXInst_Y), .Z0_f (new_AGEMA_signal_8355), .Z1_t (new_AGEMA_signal_8356), .Z1_f (new_AGEMA_signal_8357) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S22reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (stateArray_S22reg_gff_1_SFF_7_MUXInst_Y), .A0_f (new_AGEMA_signal_8355), .A1_t (new_AGEMA_signal_8356), .A1_f (new_AGEMA_signal_8357), .B0_t (stateArray_inS22ser[7]), .B0_f (new_AGEMA_signal_6835), .B1_t (new_AGEMA_signal_6836), .B1_f (new_AGEMA_signal_6837), .Z0_t (ciphertext_s0_t[47]), .Z0_f (ciphertext_s0_f[47]), .Z1_t (ciphertext_s1_t[47]), .Z1_f (ciphertext_s1_f[47]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S23reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS23ser[0]), .A0_f (new_AGEMA_signal_10877), .A1_t (new_AGEMA_signal_10878), .A1_f (new_AGEMA_signal_10879), .B0_t (ciphertext_s0_t[72]), .B0_f (ciphertext_s0_f[72]), .B1_t (ciphertext_s1_t[72]), .B1_f (ciphertext_s1_f[72]), .Z0_t (stateArray_S23reg_gff_1_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_10970), .Z1_t (new_AGEMA_signal_10971), .Z1_f (new_AGEMA_signal_10972) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S23reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S23reg_gff_1_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_10970), .B1_t (new_AGEMA_signal_10971), .B1_f (new_AGEMA_signal_10972), .Z0_t (stateArray_S23reg_gff_1_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_11099), .Z1_t (new_AGEMA_signal_11100), .Z1_f (new_AGEMA_signal_11101) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S23reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (stateArray_S23reg_gff_1_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_11099), .A1_t (new_AGEMA_signal_11100), .A1_f (new_AGEMA_signal_11101), .B0_t (stateArray_inS23ser[0]), .B0_f (new_AGEMA_signal_10877), .B1_t (new_AGEMA_signal_10878), .B1_f (new_AGEMA_signal_10879), .Z0_t (ciphertext_s0_t[8]), .Z0_f (ciphertext_s0_f[8]), .Z1_t (ciphertext_s1_t[8]), .Z1_f (ciphertext_s1_f[8]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S23reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS23ser[1]), .A0_f (new_AGEMA_signal_11003), .A1_t (new_AGEMA_signal_11004), .A1_f (new_AGEMA_signal_11005), .B0_t (ciphertext_s0_t[73]), .B0_f (ciphertext_s0_f[73]), .B1_t (ciphertext_s1_t[73]), .B1_f (ciphertext_s1_f[73]), .Z0_t (stateArray_S23reg_gff_1_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_11102), .Z1_t (new_AGEMA_signal_11103), .Z1_f (new_AGEMA_signal_11104) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S23reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S23reg_gff_1_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_11102), .B1_t (new_AGEMA_signal_11103), .B1_f (new_AGEMA_signal_11104), .Z0_t (stateArray_S23reg_gff_1_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_11153), .Z1_t (new_AGEMA_signal_11154), .Z1_f (new_AGEMA_signal_11155) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S23reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (stateArray_S23reg_gff_1_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_11153), .A1_t (new_AGEMA_signal_11154), .A1_f (new_AGEMA_signal_11155), .B0_t (stateArray_inS23ser[1]), .B0_f (new_AGEMA_signal_11003), .B1_t (new_AGEMA_signal_11004), .B1_f (new_AGEMA_signal_11005), .Z0_t (ciphertext_s0_t[9]), .Z0_f (ciphertext_s0_f[9]), .Z1_t (ciphertext_s1_t[9]), .Z1_f (ciphertext_s1_f[9]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S23reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS23ser[2]), .A0_f (new_AGEMA_signal_10883), .A1_t (new_AGEMA_signal_10884), .A1_f (new_AGEMA_signal_10885), .B0_t (ciphertext_s0_t[74]), .B0_f (ciphertext_s0_f[74]), .B1_t (ciphertext_s1_t[74]), .B1_f (ciphertext_s1_f[74]), .Z0_t (stateArray_S23reg_gff_1_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_10973), .Z1_t (new_AGEMA_signal_10974), .Z1_f (new_AGEMA_signal_10975) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S23reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S23reg_gff_1_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_10973), .B1_t (new_AGEMA_signal_10974), .B1_f (new_AGEMA_signal_10975), .Z0_t (stateArray_S23reg_gff_1_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_11105), .Z1_t (new_AGEMA_signal_11106), .Z1_f (new_AGEMA_signal_11107) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S23reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (stateArray_S23reg_gff_1_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_11105), .A1_t (new_AGEMA_signal_11106), .A1_f (new_AGEMA_signal_11107), .B0_t (stateArray_inS23ser[2]), .B0_f (new_AGEMA_signal_10883), .B1_t (new_AGEMA_signal_10884), .B1_f (new_AGEMA_signal_10885), .Z0_t (ciphertext_s0_t[10]), .Z0_f (ciphertext_s0_f[10]), .Z1_t (ciphertext_s1_t[10]), .Z1_f (ciphertext_s1_f[10]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S23reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS23ser[3]), .A0_f (new_AGEMA_signal_11006), .A1_t (new_AGEMA_signal_11007), .A1_f (new_AGEMA_signal_11008), .B0_t (ciphertext_s0_t[75]), .B0_f (ciphertext_s0_f[75]), .B1_t (ciphertext_s1_t[75]), .B1_f (ciphertext_s1_f[75]), .Z0_t (stateArray_S23reg_gff_1_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_11108), .Z1_t (new_AGEMA_signal_11109), .Z1_f (new_AGEMA_signal_11110) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S23reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S23reg_gff_1_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_11108), .B1_t (new_AGEMA_signal_11109), .B1_f (new_AGEMA_signal_11110), .Z0_t (stateArray_S23reg_gff_1_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_11156), .Z1_t (new_AGEMA_signal_11157), .Z1_f (new_AGEMA_signal_11158) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S23reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (stateArray_S23reg_gff_1_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_11156), .A1_t (new_AGEMA_signal_11157), .A1_f (new_AGEMA_signal_11158), .B0_t (stateArray_inS23ser[3]), .B0_f (new_AGEMA_signal_11006), .B1_t (new_AGEMA_signal_11007), .B1_f (new_AGEMA_signal_11008), .Z0_t (ciphertext_s0_t[11]), .Z0_f (ciphertext_s0_f[11]), .Z1_t (ciphertext_s1_t[11]), .Z1_f (ciphertext_s1_f[11]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S23reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS23ser[4]), .A0_f (new_AGEMA_signal_11009), .A1_t (new_AGEMA_signal_11010), .A1_f (new_AGEMA_signal_11011), .B0_t (ciphertext_s0_t[76]), .B0_f (ciphertext_s0_f[76]), .B1_t (ciphertext_s1_t[76]), .B1_f (ciphertext_s1_f[76]), .Z0_t (stateArray_S23reg_gff_1_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_11111), .Z1_t (new_AGEMA_signal_11112), .Z1_f (new_AGEMA_signal_11113) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S23reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S23reg_gff_1_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_11111), .B1_t (new_AGEMA_signal_11112), .B1_f (new_AGEMA_signal_11113), .Z0_t (stateArray_S23reg_gff_1_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_11159), .Z1_t (new_AGEMA_signal_11160), .Z1_f (new_AGEMA_signal_11161) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S23reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (stateArray_S23reg_gff_1_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_11159), .A1_t (new_AGEMA_signal_11160), .A1_f (new_AGEMA_signal_11161), .B0_t (stateArray_inS23ser[4]), .B0_f (new_AGEMA_signal_11009), .B1_t (new_AGEMA_signal_11010), .B1_f (new_AGEMA_signal_11011), .Z0_t (ciphertext_s0_t[12]), .Z0_f (ciphertext_s0_f[12]), .Z1_t (ciphertext_s1_t[12]), .Z1_f (ciphertext_s1_f[12]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S23reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS23ser[5]), .A0_f (new_AGEMA_signal_10892), .A1_t (new_AGEMA_signal_10893), .A1_f (new_AGEMA_signal_10894), .B0_t (ciphertext_s0_t[77]), .B0_f (ciphertext_s0_f[77]), .B1_t (ciphertext_s1_t[77]), .B1_f (ciphertext_s1_f[77]), .Z0_t (stateArray_S23reg_gff_1_SFF_5_MUXInst_X), .Z0_f (new_AGEMA_signal_10976), .Z1_t (new_AGEMA_signal_10977), .Z1_f (new_AGEMA_signal_10978) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S23reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S23reg_gff_1_SFF_5_MUXInst_X), .B0_f (new_AGEMA_signal_10976), .B1_t (new_AGEMA_signal_10977), .B1_f (new_AGEMA_signal_10978), .Z0_t (stateArray_S23reg_gff_1_SFF_5_MUXInst_Y), .Z0_f (new_AGEMA_signal_11114), .Z1_t (new_AGEMA_signal_11115), .Z1_f (new_AGEMA_signal_11116) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S23reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (stateArray_S23reg_gff_1_SFF_5_MUXInst_Y), .A0_f (new_AGEMA_signal_11114), .A1_t (new_AGEMA_signal_11115), .A1_f (new_AGEMA_signal_11116), .B0_t (stateArray_inS23ser[5]), .B0_f (new_AGEMA_signal_10892), .B1_t (new_AGEMA_signal_10893), .B1_f (new_AGEMA_signal_10894), .Z0_t (ciphertext_s0_t[13]), .Z0_f (ciphertext_s0_f[13]), .Z1_t (ciphertext_s1_t[13]), .Z1_f (ciphertext_s1_f[13]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S23reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS23ser[6]), .A0_f (new_AGEMA_signal_10895), .A1_t (new_AGEMA_signal_10896), .A1_f (new_AGEMA_signal_10897), .B0_t (ciphertext_s0_t[78]), .B0_f (ciphertext_s0_f[78]), .B1_t (ciphertext_s1_t[78]), .B1_f (ciphertext_s1_f[78]), .Z0_t (stateArray_S23reg_gff_1_SFF_6_MUXInst_X), .Z0_f (new_AGEMA_signal_10979), .Z1_t (new_AGEMA_signal_10980), .Z1_f (new_AGEMA_signal_10981) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S23reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S23reg_gff_1_SFF_6_MUXInst_X), .B0_f (new_AGEMA_signal_10979), .B1_t (new_AGEMA_signal_10980), .B1_f (new_AGEMA_signal_10981), .Z0_t (stateArray_S23reg_gff_1_SFF_6_MUXInst_Y), .Z0_f (new_AGEMA_signal_11117), .Z1_t (new_AGEMA_signal_11118), .Z1_f (new_AGEMA_signal_11119) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S23reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (stateArray_S23reg_gff_1_SFF_6_MUXInst_Y), .A0_f (new_AGEMA_signal_11117), .A1_t (new_AGEMA_signal_11118), .A1_f (new_AGEMA_signal_11119), .B0_t (stateArray_inS23ser[6]), .B0_f (new_AGEMA_signal_10895), .B1_t (new_AGEMA_signal_10896), .B1_f (new_AGEMA_signal_10897), .Z0_t (ciphertext_s0_t[14]), .Z0_f (ciphertext_s0_f[14]), .Z1_t (ciphertext_s1_t[14]), .Z1_f (ciphertext_s1_f[14]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S23reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS23ser[7]), .A0_f (new_AGEMA_signal_10898), .A1_t (new_AGEMA_signal_10899), .A1_f (new_AGEMA_signal_10900), .B0_t (ciphertext_s0_t[79]), .B0_f (ciphertext_s0_f[79]), .B1_t (ciphertext_s1_t[79]), .B1_f (ciphertext_s1_f[79]), .Z0_t (stateArray_S23reg_gff_1_SFF_7_MUXInst_X), .Z0_f (new_AGEMA_signal_10982), .Z1_t (new_AGEMA_signal_10983), .Z1_f (new_AGEMA_signal_10984) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S23reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S23reg_gff_1_SFF_7_MUXInst_X), .B0_f (new_AGEMA_signal_10982), .B1_t (new_AGEMA_signal_10983), .B1_f (new_AGEMA_signal_10984), .Z0_t (stateArray_S23reg_gff_1_SFF_7_MUXInst_Y), .Z0_f (new_AGEMA_signal_11120), .Z1_t (new_AGEMA_signal_11121), .Z1_f (new_AGEMA_signal_11122) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S23reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (stateArray_S23reg_gff_1_SFF_7_MUXInst_Y), .A0_f (new_AGEMA_signal_11120), .A1_t (new_AGEMA_signal_11121), .A1_f (new_AGEMA_signal_11122), .B0_t (stateArray_inS23ser[7]), .B0_f (new_AGEMA_signal_10898), .B1_t (new_AGEMA_signal_10899), .B1_f (new_AGEMA_signal_10900), .Z0_t (ciphertext_s0_t[15]), .Z0_f (ciphertext_s0_f[15]), .Z1_t (ciphertext_s1_t[15]), .Z1_f (ciphertext_s1_f[15]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S30reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS30ser[0]), .A0_f (new_AGEMA_signal_6838), .A1_t (new_AGEMA_signal_6839), .A1_f (new_AGEMA_signal_6840), .B0_t (ciphertext_s0_t[0]), .B0_f (ciphertext_s0_f[0]), .B1_t (ciphertext_s1_t[0]), .B1_f (ciphertext_s1_f[0]), .Z0_t (stateArray_S30reg_gff_1_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_7611), .Z1_t (new_AGEMA_signal_7612), .Z1_f (new_AGEMA_signal_7613) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S30reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S30reg_gff_1_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_7611), .B1_t (new_AGEMA_signal_7612), .B1_f (new_AGEMA_signal_7613), .Z0_t (stateArray_S30reg_gff_1_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_8358), .Z1_t (new_AGEMA_signal_8359), .Z1_f (new_AGEMA_signal_8360) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S30reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (stateArray_S30reg_gff_1_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_8358), .A1_t (new_AGEMA_signal_8359), .A1_f (new_AGEMA_signal_8360), .B0_t (stateArray_inS30ser[0]), .B0_f (new_AGEMA_signal_6838), .B1_t (new_AGEMA_signal_6839), .B1_f (new_AGEMA_signal_6840), .Z0_t (ciphertext_s0_t[96]), .Z0_f (ciphertext_s0_f[96]), .Z1_t (ciphertext_s1_t[96]), .Z1_f (ciphertext_s1_f[96]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S30reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS30ser[1]), .A0_f (new_AGEMA_signal_6841), .A1_t (new_AGEMA_signal_6842), .A1_f (new_AGEMA_signal_6843), .B0_t (ciphertext_s0_t[1]), .B0_f (ciphertext_s0_f[1]), .B1_t (ciphertext_s1_t[1]), .B1_f (ciphertext_s1_f[1]), .Z0_t (stateArray_S30reg_gff_1_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_7614), .Z1_t (new_AGEMA_signal_7615), .Z1_f (new_AGEMA_signal_7616) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S30reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S30reg_gff_1_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_7614), .B1_t (new_AGEMA_signal_7615), .B1_f (new_AGEMA_signal_7616), .Z0_t (stateArray_S30reg_gff_1_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_8361), .Z1_t (new_AGEMA_signal_8362), .Z1_f (new_AGEMA_signal_8363) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S30reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (stateArray_S30reg_gff_1_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_8361), .A1_t (new_AGEMA_signal_8362), .A1_f (new_AGEMA_signal_8363), .B0_t (stateArray_inS30ser[1]), .B0_f (new_AGEMA_signal_6841), .B1_t (new_AGEMA_signal_6842), .B1_f (new_AGEMA_signal_6843), .Z0_t (ciphertext_s0_t[97]), .Z0_f (ciphertext_s0_f[97]), .Z1_t (ciphertext_s1_t[97]), .Z1_f (ciphertext_s1_f[97]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S30reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS30ser[2]), .A0_f (new_AGEMA_signal_6844), .A1_t (new_AGEMA_signal_6845), .A1_f (new_AGEMA_signal_6846), .B0_t (ciphertext_s0_t[2]), .B0_f (ciphertext_s0_f[2]), .B1_t (ciphertext_s1_t[2]), .B1_f (ciphertext_s1_f[2]), .Z0_t (stateArray_S30reg_gff_1_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_7617), .Z1_t (new_AGEMA_signal_7618), .Z1_f (new_AGEMA_signal_7619) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S30reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S30reg_gff_1_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_7617), .B1_t (new_AGEMA_signal_7618), .B1_f (new_AGEMA_signal_7619), .Z0_t (stateArray_S30reg_gff_1_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_8364), .Z1_t (new_AGEMA_signal_8365), .Z1_f (new_AGEMA_signal_8366) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S30reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (stateArray_S30reg_gff_1_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_8364), .A1_t (new_AGEMA_signal_8365), .A1_f (new_AGEMA_signal_8366), .B0_t (stateArray_inS30ser[2]), .B0_f (new_AGEMA_signal_6844), .B1_t (new_AGEMA_signal_6845), .B1_f (new_AGEMA_signal_6846), .Z0_t (ciphertext_s0_t[98]), .Z0_f (ciphertext_s0_f[98]), .Z1_t (ciphertext_s1_t[98]), .Z1_f (ciphertext_s1_f[98]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S30reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS30ser[3]), .A0_f (new_AGEMA_signal_6847), .A1_t (new_AGEMA_signal_6848), .A1_f (new_AGEMA_signal_6849), .B0_t (ciphertext_s0_t[3]), .B0_f (ciphertext_s0_f[3]), .B1_t (ciphertext_s1_t[3]), .B1_f (ciphertext_s1_f[3]), .Z0_t (stateArray_S30reg_gff_1_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_7620), .Z1_t (new_AGEMA_signal_7621), .Z1_f (new_AGEMA_signal_7622) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S30reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S30reg_gff_1_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_7620), .B1_t (new_AGEMA_signal_7621), .B1_f (new_AGEMA_signal_7622), .Z0_t (stateArray_S30reg_gff_1_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_8367), .Z1_t (new_AGEMA_signal_8368), .Z1_f (new_AGEMA_signal_8369) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S30reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (stateArray_S30reg_gff_1_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_8367), .A1_t (new_AGEMA_signal_8368), .A1_f (new_AGEMA_signal_8369), .B0_t (stateArray_inS30ser[3]), .B0_f (new_AGEMA_signal_6847), .B1_t (new_AGEMA_signal_6848), .B1_f (new_AGEMA_signal_6849), .Z0_t (ciphertext_s0_t[99]), .Z0_f (ciphertext_s0_f[99]), .Z1_t (ciphertext_s1_t[99]), .Z1_f (ciphertext_s1_f[99]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S30reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS30ser[4]), .A0_f (new_AGEMA_signal_6850), .A1_t (new_AGEMA_signal_6851), .A1_f (new_AGEMA_signal_6852), .B0_t (ciphertext_s0_t[4]), .B0_f (ciphertext_s0_f[4]), .B1_t (ciphertext_s1_t[4]), .B1_f (ciphertext_s1_f[4]), .Z0_t (stateArray_S30reg_gff_1_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_7623), .Z1_t (new_AGEMA_signal_7624), .Z1_f (new_AGEMA_signal_7625) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S30reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S30reg_gff_1_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_7623), .B1_t (new_AGEMA_signal_7624), .B1_f (new_AGEMA_signal_7625), .Z0_t (stateArray_S30reg_gff_1_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_8370), .Z1_t (new_AGEMA_signal_8371), .Z1_f (new_AGEMA_signal_8372) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S30reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (stateArray_S30reg_gff_1_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_8370), .A1_t (new_AGEMA_signal_8371), .A1_f (new_AGEMA_signal_8372), .B0_t (stateArray_inS30ser[4]), .B0_f (new_AGEMA_signal_6850), .B1_t (new_AGEMA_signal_6851), .B1_f (new_AGEMA_signal_6852), .Z0_t (ciphertext_s0_t[100]), .Z0_f (ciphertext_s0_f[100]), .Z1_t (ciphertext_s1_t[100]), .Z1_f (ciphertext_s1_f[100]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S30reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS30ser[5]), .A0_f (new_AGEMA_signal_6853), .A1_t (new_AGEMA_signal_6854), .A1_f (new_AGEMA_signal_6855), .B0_t (ciphertext_s0_t[5]), .B0_f (ciphertext_s0_f[5]), .B1_t (ciphertext_s1_t[5]), .B1_f (ciphertext_s1_f[5]), .Z0_t (stateArray_S30reg_gff_1_SFF_5_MUXInst_X), .Z0_f (new_AGEMA_signal_7626), .Z1_t (new_AGEMA_signal_7627), .Z1_f (new_AGEMA_signal_7628) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S30reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S30reg_gff_1_SFF_5_MUXInst_X), .B0_f (new_AGEMA_signal_7626), .B1_t (new_AGEMA_signal_7627), .B1_f (new_AGEMA_signal_7628), .Z0_t (stateArray_S30reg_gff_1_SFF_5_MUXInst_Y), .Z0_f (new_AGEMA_signal_8373), .Z1_t (new_AGEMA_signal_8374), .Z1_f (new_AGEMA_signal_8375) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S30reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (stateArray_S30reg_gff_1_SFF_5_MUXInst_Y), .A0_f (new_AGEMA_signal_8373), .A1_t (new_AGEMA_signal_8374), .A1_f (new_AGEMA_signal_8375), .B0_t (stateArray_inS30ser[5]), .B0_f (new_AGEMA_signal_6853), .B1_t (new_AGEMA_signal_6854), .B1_f (new_AGEMA_signal_6855), .Z0_t (ciphertext_s0_t[101]), .Z0_f (ciphertext_s0_f[101]), .Z1_t (ciphertext_s1_t[101]), .Z1_f (ciphertext_s1_f[101]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S30reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS30ser[6]), .A0_f (new_AGEMA_signal_6856), .A1_t (new_AGEMA_signal_6857), .A1_f (new_AGEMA_signal_6858), .B0_t (ciphertext_s0_t[6]), .B0_f (ciphertext_s0_f[6]), .B1_t (ciphertext_s1_t[6]), .B1_f (ciphertext_s1_f[6]), .Z0_t (stateArray_S30reg_gff_1_SFF_6_MUXInst_X), .Z0_f (new_AGEMA_signal_7629), .Z1_t (new_AGEMA_signal_7630), .Z1_f (new_AGEMA_signal_7631) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S30reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S30reg_gff_1_SFF_6_MUXInst_X), .B0_f (new_AGEMA_signal_7629), .B1_t (new_AGEMA_signal_7630), .B1_f (new_AGEMA_signal_7631), .Z0_t (stateArray_S30reg_gff_1_SFF_6_MUXInst_Y), .Z0_f (new_AGEMA_signal_8376), .Z1_t (new_AGEMA_signal_8377), .Z1_f (new_AGEMA_signal_8378) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S30reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (stateArray_S30reg_gff_1_SFF_6_MUXInst_Y), .A0_f (new_AGEMA_signal_8376), .A1_t (new_AGEMA_signal_8377), .A1_f (new_AGEMA_signal_8378), .B0_t (stateArray_inS30ser[6]), .B0_f (new_AGEMA_signal_6856), .B1_t (new_AGEMA_signal_6857), .B1_f (new_AGEMA_signal_6858), .Z0_t (ciphertext_s0_t[102]), .Z0_f (ciphertext_s0_f[102]), .Z1_t (ciphertext_s1_t[102]), .Z1_f (ciphertext_s1_f[102]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S30reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS30ser[7]), .A0_f (new_AGEMA_signal_6859), .A1_t (new_AGEMA_signal_6860), .A1_f (new_AGEMA_signal_6861), .B0_t (ciphertext_s0_t[7]), .B0_f (ciphertext_s0_f[7]), .B1_t (ciphertext_s1_t[7]), .B1_f (ciphertext_s1_f[7]), .Z0_t (stateArray_S30reg_gff_1_SFF_7_MUXInst_X), .Z0_f (new_AGEMA_signal_7632), .Z1_t (new_AGEMA_signal_7633), .Z1_f (new_AGEMA_signal_7634) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S30reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S30reg_gff_1_SFF_7_MUXInst_X), .B0_f (new_AGEMA_signal_7632), .B1_t (new_AGEMA_signal_7633), .B1_f (new_AGEMA_signal_7634), .Z0_t (stateArray_S30reg_gff_1_SFF_7_MUXInst_Y), .Z0_f (new_AGEMA_signal_8379), .Z1_t (new_AGEMA_signal_8380), .Z1_f (new_AGEMA_signal_8381) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S30reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (stateArray_S30reg_gff_1_SFF_7_MUXInst_Y), .A0_f (new_AGEMA_signal_8379), .A1_t (new_AGEMA_signal_8380), .A1_f (new_AGEMA_signal_8381), .B0_t (stateArray_inS30ser[7]), .B0_f (new_AGEMA_signal_6859), .B1_t (new_AGEMA_signal_6860), .B1_f (new_AGEMA_signal_6861), .Z0_t (ciphertext_s0_t[103]), .Z0_f (ciphertext_s0_f[103]), .Z1_t (ciphertext_s1_t[103]), .Z1_f (ciphertext_s1_f[103]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S31reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS31ser[0]), .A0_f (new_AGEMA_signal_6862), .A1_t (new_AGEMA_signal_6863), .A1_f (new_AGEMA_signal_6864), .B0_t (ciphertext_s0_t[96]), .B0_f (ciphertext_s0_f[96]), .B1_t (ciphertext_s1_t[96]), .B1_f (ciphertext_s1_f[96]), .Z0_t (stateArray_S31reg_gff_1_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_7635), .Z1_t (new_AGEMA_signal_7636), .Z1_f (new_AGEMA_signal_7637) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S31reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S31reg_gff_1_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_7635), .B1_t (new_AGEMA_signal_7636), .B1_f (new_AGEMA_signal_7637), .Z0_t (stateArray_S31reg_gff_1_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_8382), .Z1_t (new_AGEMA_signal_8383), .Z1_f (new_AGEMA_signal_8384) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S31reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (stateArray_S31reg_gff_1_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_8382), .A1_t (new_AGEMA_signal_8383), .A1_f (new_AGEMA_signal_8384), .B0_t (stateArray_inS31ser[0]), .B0_f (new_AGEMA_signal_6862), .B1_t (new_AGEMA_signal_6863), .B1_f (new_AGEMA_signal_6864), .Z0_t (ciphertext_s0_t[64]), .Z0_f (ciphertext_s0_f[64]), .Z1_t (ciphertext_s1_t[64]), .Z1_f (ciphertext_s1_f[64]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S31reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS31ser[1]), .A0_f (new_AGEMA_signal_6865), .A1_t (new_AGEMA_signal_6866), .A1_f (new_AGEMA_signal_6867), .B0_t (ciphertext_s0_t[97]), .B0_f (ciphertext_s0_f[97]), .B1_t (ciphertext_s1_t[97]), .B1_f (ciphertext_s1_f[97]), .Z0_t (stateArray_S31reg_gff_1_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_7638), .Z1_t (new_AGEMA_signal_7639), .Z1_f (new_AGEMA_signal_7640) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S31reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S31reg_gff_1_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_7638), .B1_t (new_AGEMA_signal_7639), .B1_f (new_AGEMA_signal_7640), .Z0_t (stateArray_S31reg_gff_1_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_8385), .Z1_t (new_AGEMA_signal_8386), .Z1_f (new_AGEMA_signal_8387) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S31reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (stateArray_S31reg_gff_1_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_8385), .A1_t (new_AGEMA_signal_8386), .A1_f (new_AGEMA_signal_8387), .B0_t (stateArray_inS31ser[1]), .B0_f (new_AGEMA_signal_6865), .B1_t (new_AGEMA_signal_6866), .B1_f (new_AGEMA_signal_6867), .Z0_t (ciphertext_s0_t[65]), .Z0_f (ciphertext_s0_f[65]), .Z1_t (ciphertext_s1_t[65]), .Z1_f (ciphertext_s1_f[65]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S31reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS31ser[2]), .A0_f (new_AGEMA_signal_6868), .A1_t (new_AGEMA_signal_6869), .A1_f (new_AGEMA_signal_6870), .B0_t (ciphertext_s0_t[98]), .B0_f (ciphertext_s0_f[98]), .B1_t (ciphertext_s1_t[98]), .B1_f (ciphertext_s1_f[98]), .Z0_t (stateArray_S31reg_gff_1_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_7641), .Z1_t (new_AGEMA_signal_7642), .Z1_f (new_AGEMA_signal_7643) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S31reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S31reg_gff_1_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_7641), .B1_t (new_AGEMA_signal_7642), .B1_f (new_AGEMA_signal_7643), .Z0_t (stateArray_S31reg_gff_1_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_8388), .Z1_t (new_AGEMA_signal_8389), .Z1_f (new_AGEMA_signal_8390) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S31reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (stateArray_S31reg_gff_1_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_8388), .A1_t (new_AGEMA_signal_8389), .A1_f (new_AGEMA_signal_8390), .B0_t (stateArray_inS31ser[2]), .B0_f (new_AGEMA_signal_6868), .B1_t (new_AGEMA_signal_6869), .B1_f (new_AGEMA_signal_6870), .Z0_t (ciphertext_s0_t[66]), .Z0_f (ciphertext_s0_f[66]), .Z1_t (ciphertext_s1_t[66]), .Z1_f (ciphertext_s1_f[66]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S31reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS31ser[3]), .A0_f (new_AGEMA_signal_6871), .A1_t (new_AGEMA_signal_6872), .A1_f (new_AGEMA_signal_6873), .B0_t (ciphertext_s0_t[99]), .B0_f (ciphertext_s0_f[99]), .B1_t (ciphertext_s1_t[99]), .B1_f (ciphertext_s1_f[99]), .Z0_t (stateArray_S31reg_gff_1_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_7644), .Z1_t (new_AGEMA_signal_7645), .Z1_f (new_AGEMA_signal_7646) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S31reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S31reg_gff_1_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_7644), .B1_t (new_AGEMA_signal_7645), .B1_f (new_AGEMA_signal_7646), .Z0_t (stateArray_S31reg_gff_1_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_8391), .Z1_t (new_AGEMA_signal_8392), .Z1_f (new_AGEMA_signal_8393) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S31reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (stateArray_S31reg_gff_1_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_8391), .A1_t (new_AGEMA_signal_8392), .A1_f (new_AGEMA_signal_8393), .B0_t (stateArray_inS31ser[3]), .B0_f (new_AGEMA_signal_6871), .B1_t (new_AGEMA_signal_6872), .B1_f (new_AGEMA_signal_6873), .Z0_t (ciphertext_s0_t[67]), .Z0_f (ciphertext_s0_f[67]), .Z1_t (ciphertext_s1_t[67]), .Z1_f (ciphertext_s1_f[67]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S31reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS31ser[4]), .A0_f (new_AGEMA_signal_6874), .A1_t (new_AGEMA_signal_6875), .A1_f (new_AGEMA_signal_6876), .B0_t (ciphertext_s0_t[100]), .B0_f (ciphertext_s0_f[100]), .B1_t (ciphertext_s1_t[100]), .B1_f (ciphertext_s1_f[100]), .Z0_t (stateArray_S31reg_gff_1_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_7647), .Z1_t (new_AGEMA_signal_7648), .Z1_f (new_AGEMA_signal_7649) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S31reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S31reg_gff_1_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_7647), .B1_t (new_AGEMA_signal_7648), .B1_f (new_AGEMA_signal_7649), .Z0_t (stateArray_S31reg_gff_1_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_8394), .Z1_t (new_AGEMA_signal_8395), .Z1_f (new_AGEMA_signal_8396) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S31reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (stateArray_S31reg_gff_1_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_8394), .A1_t (new_AGEMA_signal_8395), .A1_f (new_AGEMA_signal_8396), .B0_t (stateArray_inS31ser[4]), .B0_f (new_AGEMA_signal_6874), .B1_t (new_AGEMA_signal_6875), .B1_f (new_AGEMA_signal_6876), .Z0_t (ciphertext_s0_t[68]), .Z0_f (ciphertext_s0_f[68]), .Z1_t (ciphertext_s1_t[68]), .Z1_f (ciphertext_s1_f[68]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S31reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS31ser[5]), .A0_f (new_AGEMA_signal_6877), .A1_t (new_AGEMA_signal_6878), .A1_f (new_AGEMA_signal_6879), .B0_t (ciphertext_s0_t[101]), .B0_f (ciphertext_s0_f[101]), .B1_t (ciphertext_s1_t[101]), .B1_f (ciphertext_s1_f[101]), .Z0_t (stateArray_S31reg_gff_1_SFF_5_MUXInst_X), .Z0_f (new_AGEMA_signal_7650), .Z1_t (new_AGEMA_signal_7651), .Z1_f (new_AGEMA_signal_7652) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S31reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S31reg_gff_1_SFF_5_MUXInst_X), .B0_f (new_AGEMA_signal_7650), .B1_t (new_AGEMA_signal_7651), .B1_f (new_AGEMA_signal_7652), .Z0_t (stateArray_S31reg_gff_1_SFF_5_MUXInst_Y), .Z0_f (new_AGEMA_signal_8397), .Z1_t (new_AGEMA_signal_8398), .Z1_f (new_AGEMA_signal_8399) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S31reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (stateArray_S31reg_gff_1_SFF_5_MUXInst_Y), .A0_f (new_AGEMA_signal_8397), .A1_t (new_AGEMA_signal_8398), .A1_f (new_AGEMA_signal_8399), .B0_t (stateArray_inS31ser[5]), .B0_f (new_AGEMA_signal_6877), .B1_t (new_AGEMA_signal_6878), .B1_f (new_AGEMA_signal_6879), .Z0_t (ciphertext_s0_t[69]), .Z0_f (ciphertext_s0_f[69]), .Z1_t (ciphertext_s1_t[69]), .Z1_f (ciphertext_s1_f[69]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S31reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS31ser[6]), .A0_f (new_AGEMA_signal_6880), .A1_t (new_AGEMA_signal_6881), .A1_f (new_AGEMA_signal_6882), .B0_t (ciphertext_s0_t[102]), .B0_f (ciphertext_s0_f[102]), .B1_t (ciphertext_s1_t[102]), .B1_f (ciphertext_s1_f[102]), .Z0_t (stateArray_S31reg_gff_1_SFF_6_MUXInst_X), .Z0_f (new_AGEMA_signal_7653), .Z1_t (new_AGEMA_signal_7654), .Z1_f (new_AGEMA_signal_7655) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S31reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S31reg_gff_1_SFF_6_MUXInst_X), .B0_f (new_AGEMA_signal_7653), .B1_t (new_AGEMA_signal_7654), .B1_f (new_AGEMA_signal_7655), .Z0_t (stateArray_S31reg_gff_1_SFF_6_MUXInst_Y), .Z0_f (new_AGEMA_signal_8400), .Z1_t (new_AGEMA_signal_8401), .Z1_f (new_AGEMA_signal_8402) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S31reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (stateArray_S31reg_gff_1_SFF_6_MUXInst_Y), .A0_f (new_AGEMA_signal_8400), .A1_t (new_AGEMA_signal_8401), .A1_f (new_AGEMA_signal_8402), .B0_t (stateArray_inS31ser[6]), .B0_f (new_AGEMA_signal_6880), .B1_t (new_AGEMA_signal_6881), .B1_f (new_AGEMA_signal_6882), .Z0_t (ciphertext_s0_t[70]), .Z0_f (ciphertext_s0_f[70]), .Z1_t (ciphertext_s1_t[70]), .Z1_f (ciphertext_s1_f[70]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S31reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS31ser[7]), .A0_f (new_AGEMA_signal_6883), .A1_t (new_AGEMA_signal_6884), .A1_f (new_AGEMA_signal_6885), .B0_t (ciphertext_s0_t[103]), .B0_f (ciphertext_s0_f[103]), .B1_t (ciphertext_s1_t[103]), .B1_f (ciphertext_s1_f[103]), .Z0_t (stateArray_S31reg_gff_1_SFF_7_MUXInst_X), .Z0_f (new_AGEMA_signal_7656), .Z1_t (new_AGEMA_signal_7657), .Z1_f (new_AGEMA_signal_7658) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S31reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S31reg_gff_1_SFF_7_MUXInst_X), .B0_f (new_AGEMA_signal_7656), .B1_t (new_AGEMA_signal_7657), .B1_f (new_AGEMA_signal_7658), .Z0_t (stateArray_S31reg_gff_1_SFF_7_MUXInst_Y), .Z0_f (new_AGEMA_signal_8403), .Z1_t (new_AGEMA_signal_8404), .Z1_f (new_AGEMA_signal_8405) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S31reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (stateArray_S31reg_gff_1_SFF_7_MUXInst_Y), .A0_f (new_AGEMA_signal_8403), .A1_t (new_AGEMA_signal_8404), .A1_f (new_AGEMA_signal_8405), .B0_t (stateArray_inS31ser[7]), .B0_f (new_AGEMA_signal_6883), .B1_t (new_AGEMA_signal_6884), .B1_f (new_AGEMA_signal_6885), .Z0_t (ciphertext_s0_t[71]), .Z0_f (ciphertext_s0_f[71]), .Z1_t (ciphertext_s1_t[71]), .Z1_f (ciphertext_s1_f[71]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S32reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS32ser[0]), .A0_f (new_AGEMA_signal_6886), .A1_t (new_AGEMA_signal_6887), .A1_f (new_AGEMA_signal_6888), .B0_t (ciphertext_s0_t[64]), .B0_f (ciphertext_s0_f[64]), .B1_t (ciphertext_s1_t[64]), .B1_f (ciphertext_s1_f[64]), .Z0_t (stateArray_S32reg_gff_1_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_7659), .Z1_t (new_AGEMA_signal_7660), .Z1_f (new_AGEMA_signal_7661) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S32reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S32reg_gff_1_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_7659), .B1_t (new_AGEMA_signal_7660), .B1_f (new_AGEMA_signal_7661), .Z0_t (stateArray_S32reg_gff_1_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_8406), .Z1_t (new_AGEMA_signal_8407), .Z1_f (new_AGEMA_signal_8408) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S32reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (stateArray_S32reg_gff_1_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_8406), .A1_t (new_AGEMA_signal_8407), .A1_f (new_AGEMA_signal_8408), .B0_t (stateArray_inS32ser[0]), .B0_f (new_AGEMA_signal_6886), .B1_t (new_AGEMA_signal_6887), .B1_f (new_AGEMA_signal_6888), .Z0_t (ciphertext_s0_t[32]), .Z0_f (ciphertext_s0_f[32]), .Z1_t (ciphertext_s1_t[32]), .Z1_f (ciphertext_s1_f[32]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S32reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS32ser[1]), .A0_f (new_AGEMA_signal_6889), .A1_t (new_AGEMA_signal_6890), .A1_f (new_AGEMA_signal_6891), .B0_t (ciphertext_s0_t[65]), .B0_f (ciphertext_s0_f[65]), .B1_t (ciphertext_s1_t[65]), .B1_f (ciphertext_s1_f[65]), .Z0_t (stateArray_S32reg_gff_1_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_7662), .Z1_t (new_AGEMA_signal_7663), .Z1_f (new_AGEMA_signal_7664) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S32reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S32reg_gff_1_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_7662), .B1_t (new_AGEMA_signal_7663), .B1_f (new_AGEMA_signal_7664), .Z0_t (stateArray_S32reg_gff_1_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_8409), .Z1_t (new_AGEMA_signal_8410), .Z1_f (new_AGEMA_signal_8411) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S32reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (stateArray_S32reg_gff_1_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_8409), .A1_t (new_AGEMA_signal_8410), .A1_f (new_AGEMA_signal_8411), .B0_t (stateArray_inS32ser[1]), .B0_f (new_AGEMA_signal_6889), .B1_t (new_AGEMA_signal_6890), .B1_f (new_AGEMA_signal_6891), .Z0_t (ciphertext_s0_t[33]), .Z0_f (ciphertext_s0_f[33]), .Z1_t (ciphertext_s1_t[33]), .Z1_f (ciphertext_s1_f[33]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S32reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS32ser[2]), .A0_f (new_AGEMA_signal_6892), .A1_t (new_AGEMA_signal_6893), .A1_f (new_AGEMA_signal_6894), .B0_t (ciphertext_s0_t[66]), .B0_f (ciphertext_s0_f[66]), .B1_t (ciphertext_s1_t[66]), .B1_f (ciphertext_s1_f[66]), .Z0_t (stateArray_S32reg_gff_1_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_7665), .Z1_t (new_AGEMA_signal_7666), .Z1_f (new_AGEMA_signal_7667) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S32reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S32reg_gff_1_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_7665), .B1_t (new_AGEMA_signal_7666), .B1_f (new_AGEMA_signal_7667), .Z0_t (stateArray_S32reg_gff_1_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_8412), .Z1_t (new_AGEMA_signal_8413), .Z1_f (new_AGEMA_signal_8414) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S32reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (stateArray_S32reg_gff_1_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_8412), .A1_t (new_AGEMA_signal_8413), .A1_f (new_AGEMA_signal_8414), .B0_t (stateArray_inS32ser[2]), .B0_f (new_AGEMA_signal_6892), .B1_t (new_AGEMA_signal_6893), .B1_f (new_AGEMA_signal_6894), .Z0_t (ciphertext_s0_t[34]), .Z0_f (ciphertext_s0_f[34]), .Z1_t (ciphertext_s1_t[34]), .Z1_f (ciphertext_s1_f[34]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S32reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS32ser[3]), .A0_f (new_AGEMA_signal_6895), .A1_t (new_AGEMA_signal_6896), .A1_f (new_AGEMA_signal_6897), .B0_t (ciphertext_s0_t[67]), .B0_f (ciphertext_s0_f[67]), .B1_t (ciphertext_s1_t[67]), .B1_f (ciphertext_s1_f[67]), .Z0_t (stateArray_S32reg_gff_1_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_7668), .Z1_t (new_AGEMA_signal_7669), .Z1_f (new_AGEMA_signal_7670) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S32reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S32reg_gff_1_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_7668), .B1_t (new_AGEMA_signal_7669), .B1_f (new_AGEMA_signal_7670), .Z0_t (stateArray_S32reg_gff_1_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_8415), .Z1_t (new_AGEMA_signal_8416), .Z1_f (new_AGEMA_signal_8417) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S32reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (stateArray_S32reg_gff_1_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_8415), .A1_t (new_AGEMA_signal_8416), .A1_f (new_AGEMA_signal_8417), .B0_t (stateArray_inS32ser[3]), .B0_f (new_AGEMA_signal_6895), .B1_t (new_AGEMA_signal_6896), .B1_f (new_AGEMA_signal_6897), .Z0_t (ciphertext_s0_t[35]), .Z0_f (ciphertext_s0_f[35]), .Z1_t (ciphertext_s1_t[35]), .Z1_f (ciphertext_s1_f[35]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S32reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS32ser[4]), .A0_f (new_AGEMA_signal_6898), .A1_t (new_AGEMA_signal_6899), .A1_f (new_AGEMA_signal_6900), .B0_t (ciphertext_s0_t[68]), .B0_f (ciphertext_s0_f[68]), .B1_t (ciphertext_s1_t[68]), .B1_f (ciphertext_s1_f[68]), .Z0_t (stateArray_S32reg_gff_1_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_7671), .Z1_t (new_AGEMA_signal_7672), .Z1_f (new_AGEMA_signal_7673) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S32reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S32reg_gff_1_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_7671), .B1_t (new_AGEMA_signal_7672), .B1_f (new_AGEMA_signal_7673), .Z0_t (stateArray_S32reg_gff_1_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_8418), .Z1_t (new_AGEMA_signal_8419), .Z1_f (new_AGEMA_signal_8420) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S32reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (stateArray_S32reg_gff_1_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_8418), .A1_t (new_AGEMA_signal_8419), .A1_f (new_AGEMA_signal_8420), .B0_t (stateArray_inS32ser[4]), .B0_f (new_AGEMA_signal_6898), .B1_t (new_AGEMA_signal_6899), .B1_f (new_AGEMA_signal_6900), .Z0_t (ciphertext_s0_t[36]), .Z0_f (ciphertext_s0_f[36]), .Z1_t (ciphertext_s1_t[36]), .Z1_f (ciphertext_s1_f[36]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S32reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS32ser[5]), .A0_f (new_AGEMA_signal_6901), .A1_t (new_AGEMA_signal_6902), .A1_f (new_AGEMA_signal_6903), .B0_t (ciphertext_s0_t[69]), .B0_f (ciphertext_s0_f[69]), .B1_t (ciphertext_s1_t[69]), .B1_f (ciphertext_s1_f[69]), .Z0_t (stateArray_S32reg_gff_1_SFF_5_MUXInst_X), .Z0_f (new_AGEMA_signal_7674), .Z1_t (new_AGEMA_signal_7675), .Z1_f (new_AGEMA_signal_7676) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S32reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S32reg_gff_1_SFF_5_MUXInst_X), .B0_f (new_AGEMA_signal_7674), .B1_t (new_AGEMA_signal_7675), .B1_f (new_AGEMA_signal_7676), .Z0_t (stateArray_S32reg_gff_1_SFF_5_MUXInst_Y), .Z0_f (new_AGEMA_signal_8421), .Z1_t (new_AGEMA_signal_8422), .Z1_f (new_AGEMA_signal_8423) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S32reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (stateArray_S32reg_gff_1_SFF_5_MUXInst_Y), .A0_f (new_AGEMA_signal_8421), .A1_t (new_AGEMA_signal_8422), .A1_f (new_AGEMA_signal_8423), .B0_t (stateArray_inS32ser[5]), .B0_f (new_AGEMA_signal_6901), .B1_t (new_AGEMA_signal_6902), .B1_f (new_AGEMA_signal_6903), .Z0_t (ciphertext_s0_t[37]), .Z0_f (ciphertext_s0_f[37]), .Z1_t (ciphertext_s1_t[37]), .Z1_f (ciphertext_s1_f[37]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S32reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS32ser[6]), .A0_f (new_AGEMA_signal_6904), .A1_t (new_AGEMA_signal_6905), .A1_f (new_AGEMA_signal_6906), .B0_t (ciphertext_s0_t[70]), .B0_f (ciphertext_s0_f[70]), .B1_t (ciphertext_s1_t[70]), .B1_f (ciphertext_s1_f[70]), .Z0_t (stateArray_S32reg_gff_1_SFF_6_MUXInst_X), .Z0_f (new_AGEMA_signal_7677), .Z1_t (new_AGEMA_signal_7678), .Z1_f (new_AGEMA_signal_7679) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S32reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S32reg_gff_1_SFF_6_MUXInst_X), .B0_f (new_AGEMA_signal_7677), .B1_t (new_AGEMA_signal_7678), .B1_f (new_AGEMA_signal_7679), .Z0_t (stateArray_S32reg_gff_1_SFF_6_MUXInst_Y), .Z0_f (new_AGEMA_signal_8424), .Z1_t (new_AGEMA_signal_8425), .Z1_f (new_AGEMA_signal_8426) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S32reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (stateArray_S32reg_gff_1_SFF_6_MUXInst_Y), .A0_f (new_AGEMA_signal_8424), .A1_t (new_AGEMA_signal_8425), .A1_f (new_AGEMA_signal_8426), .B0_t (stateArray_inS32ser[6]), .B0_f (new_AGEMA_signal_6904), .B1_t (new_AGEMA_signal_6905), .B1_f (new_AGEMA_signal_6906), .Z0_t (ciphertext_s0_t[38]), .Z0_f (ciphertext_s0_f[38]), .Z1_t (ciphertext_s1_t[38]), .Z1_f (ciphertext_s1_f[38]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S32reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS32ser[7]), .A0_f (new_AGEMA_signal_6907), .A1_t (new_AGEMA_signal_6908), .A1_f (new_AGEMA_signal_6909), .B0_t (ciphertext_s0_t[71]), .B0_f (ciphertext_s0_f[71]), .B1_t (ciphertext_s1_t[71]), .B1_f (ciphertext_s1_f[71]), .Z0_t (stateArray_S32reg_gff_1_SFF_7_MUXInst_X), .Z0_f (new_AGEMA_signal_7680), .Z1_t (new_AGEMA_signal_7681), .Z1_f (new_AGEMA_signal_7682) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S32reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S32reg_gff_1_SFF_7_MUXInst_X), .B0_f (new_AGEMA_signal_7680), .B1_t (new_AGEMA_signal_7681), .B1_f (new_AGEMA_signal_7682), .Z0_t (stateArray_S32reg_gff_1_SFF_7_MUXInst_Y), .Z0_f (new_AGEMA_signal_8427), .Z1_t (new_AGEMA_signal_8428), .Z1_f (new_AGEMA_signal_8429) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S32reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (stateArray_S32reg_gff_1_SFF_7_MUXInst_Y), .A0_f (new_AGEMA_signal_8427), .A1_t (new_AGEMA_signal_8428), .A1_f (new_AGEMA_signal_8429), .B0_t (stateArray_inS32ser[7]), .B0_f (new_AGEMA_signal_6907), .B1_t (new_AGEMA_signal_6908), .B1_f (new_AGEMA_signal_6909), .Z0_t (ciphertext_s0_t[39]), .Z0_f (ciphertext_s0_f[39]), .Z1_t (ciphertext_s1_t[39]), .Z1_f (ciphertext_s1_f[39]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S33reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS33ser[0]), .A0_f (new_AGEMA_signal_11684), .A1_t (new_AGEMA_signal_11685), .A1_f (new_AGEMA_signal_11686), .B0_t (ciphertext_s0_t[32]), .B0_f (ciphertext_s0_f[32]), .B1_t (ciphertext_s1_t[32]), .B1_f (ciphertext_s1_f[32]), .Z0_t (stateArray_S33reg_gff_1_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_11708), .Z1_t (new_AGEMA_signal_11709), .Z1_f (new_AGEMA_signal_11710) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S33reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S33reg_gff_1_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_11708), .B1_t (new_AGEMA_signal_11709), .B1_f (new_AGEMA_signal_11710), .Z0_t (stateArray_S33reg_gff_1_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_11732), .Z1_t (new_AGEMA_signal_11733), .Z1_f (new_AGEMA_signal_11734) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S33reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (stateArray_S33reg_gff_1_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_11732), .A1_t (new_AGEMA_signal_11733), .A1_f (new_AGEMA_signal_11734), .B0_t (stateArray_inS33ser[0]), .B0_f (new_AGEMA_signal_11684), .B1_t (new_AGEMA_signal_11685), .B1_f (new_AGEMA_signal_11686), .Z0_t (ciphertext_s0_t[0]), .Z0_f (ciphertext_s0_f[0]), .Z1_t (ciphertext_s1_t[0]), .Z1_f (ciphertext_s1_f[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S33reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS33ser[1]), .A0_f (new_AGEMA_signal_11711), .A1_t (new_AGEMA_signal_11712), .A1_f (new_AGEMA_signal_11713), .B0_t (ciphertext_s0_t[33]), .B0_f (ciphertext_s0_f[33]), .B1_t (ciphertext_s1_t[33]), .B1_f (ciphertext_s1_f[33]), .Z0_t (stateArray_S33reg_gff_1_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_11735), .Z1_t (new_AGEMA_signal_11736), .Z1_f (new_AGEMA_signal_11737) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S33reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S33reg_gff_1_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_11735), .B1_t (new_AGEMA_signal_11736), .B1_f (new_AGEMA_signal_11737), .Z0_t (stateArray_S33reg_gff_1_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_11756), .Z1_t (new_AGEMA_signal_11757), .Z1_f (new_AGEMA_signal_11758) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S33reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (stateArray_S33reg_gff_1_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_11756), .A1_t (new_AGEMA_signal_11757), .A1_f (new_AGEMA_signal_11758), .B0_t (stateArray_inS33ser[1]), .B0_f (new_AGEMA_signal_11711), .B1_t (new_AGEMA_signal_11712), .B1_f (new_AGEMA_signal_11713), .Z0_t (ciphertext_s0_t[1]), .Z0_f (ciphertext_s0_f[1]), .Z1_t (ciphertext_s1_t[1]), .Z1_f (ciphertext_s1_f[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S33reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS33ser[2]), .A0_f (new_AGEMA_signal_11714), .A1_t (new_AGEMA_signal_11715), .A1_f (new_AGEMA_signal_11716), .B0_t (ciphertext_s0_t[34]), .B0_f (ciphertext_s0_f[34]), .B1_t (ciphertext_s1_t[34]), .B1_f (ciphertext_s1_f[34]), .Z0_t (stateArray_S33reg_gff_1_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_11738), .Z1_t (new_AGEMA_signal_11739), .Z1_f (new_AGEMA_signal_11740) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S33reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S33reg_gff_1_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_11738), .B1_t (new_AGEMA_signal_11739), .B1_f (new_AGEMA_signal_11740), .Z0_t (stateArray_S33reg_gff_1_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_11759), .Z1_t (new_AGEMA_signal_11760), .Z1_f (new_AGEMA_signal_11761) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S33reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (stateArray_S33reg_gff_1_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_11759), .A1_t (new_AGEMA_signal_11760), .A1_f (new_AGEMA_signal_11761), .B0_t (stateArray_inS33ser[2]), .B0_f (new_AGEMA_signal_11714), .B1_t (new_AGEMA_signal_11715), .B1_f (new_AGEMA_signal_11716), .Z0_t (ciphertext_s0_t[2]), .Z0_f (ciphertext_s0_f[2]), .Z1_t (ciphertext_s1_t[2]), .Z1_f (ciphertext_s1_f[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S33reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS33ser[3]), .A0_f (new_AGEMA_signal_11717), .A1_t (new_AGEMA_signal_11718), .A1_f (new_AGEMA_signal_11719), .B0_t (ciphertext_s0_t[35]), .B0_f (ciphertext_s0_f[35]), .B1_t (ciphertext_s1_t[35]), .B1_f (ciphertext_s1_f[35]), .Z0_t (stateArray_S33reg_gff_1_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_11741), .Z1_t (new_AGEMA_signal_11742), .Z1_f (new_AGEMA_signal_11743) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S33reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S33reg_gff_1_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_11741), .B1_t (new_AGEMA_signal_11742), .B1_f (new_AGEMA_signal_11743), .Z0_t (stateArray_S33reg_gff_1_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_11762), .Z1_t (new_AGEMA_signal_11763), .Z1_f (new_AGEMA_signal_11764) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S33reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (stateArray_S33reg_gff_1_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_11762), .A1_t (new_AGEMA_signal_11763), .A1_f (new_AGEMA_signal_11764), .B0_t (stateArray_inS33ser[3]), .B0_f (new_AGEMA_signal_11717), .B1_t (new_AGEMA_signal_11718), .B1_f (new_AGEMA_signal_11719), .Z0_t (ciphertext_s0_t[3]), .Z0_f (ciphertext_s0_f[3]), .Z1_t (ciphertext_s1_t[3]), .Z1_f (ciphertext_s1_f[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S33reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS33ser[4]), .A0_f (new_AGEMA_signal_11720), .A1_t (new_AGEMA_signal_11721), .A1_f (new_AGEMA_signal_11722), .B0_t (ciphertext_s0_t[36]), .B0_f (ciphertext_s0_f[36]), .B1_t (ciphertext_s1_t[36]), .B1_f (ciphertext_s1_f[36]), .Z0_t (stateArray_S33reg_gff_1_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_11744), .Z1_t (new_AGEMA_signal_11745), .Z1_f (new_AGEMA_signal_11746) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S33reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S33reg_gff_1_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_11744), .B1_t (new_AGEMA_signal_11745), .B1_f (new_AGEMA_signal_11746), .Z0_t (stateArray_S33reg_gff_1_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_11765), .Z1_t (new_AGEMA_signal_11766), .Z1_f (new_AGEMA_signal_11767) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S33reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (stateArray_S33reg_gff_1_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_11765), .A1_t (new_AGEMA_signal_11766), .A1_f (new_AGEMA_signal_11767), .B0_t (stateArray_inS33ser[4]), .B0_f (new_AGEMA_signal_11720), .B1_t (new_AGEMA_signal_11721), .B1_f (new_AGEMA_signal_11722), .Z0_t (ciphertext_s0_t[4]), .Z0_f (ciphertext_s0_f[4]), .Z1_t (ciphertext_s1_t[4]), .Z1_f (ciphertext_s1_f[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S33reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS33ser[5]), .A0_f (new_AGEMA_signal_11723), .A1_t (new_AGEMA_signal_11724), .A1_f (new_AGEMA_signal_11725), .B0_t (ciphertext_s0_t[37]), .B0_f (ciphertext_s0_f[37]), .B1_t (ciphertext_s1_t[37]), .B1_f (ciphertext_s1_f[37]), .Z0_t (stateArray_S33reg_gff_1_SFF_5_MUXInst_X), .Z0_f (new_AGEMA_signal_11747), .Z1_t (new_AGEMA_signal_11748), .Z1_f (new_AGEMA_signal_11749) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S33reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S33reg_gff_1_SFF_5_MUXInst_X), .B0_f (new_AGEMA_signal_11747), .B1_t (new_AGEMA_signal_11748), .B1_f (new_AGEMA_signal_11749), .Z0_t (stateArray_S33reg_gff_1_SFF_5_MUXInst_Y), .Z0_f (new_AGEMA_signal_11768), .Z1_t (new_AGEMA_signal_11769), .Z1_f (new_AGEMA_signal_11770) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S33reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (stateArray_S33reg_gff_1_SFF_5_MUXInst_Y), .A0_f (new_AGEMA_signal_11768), .A1_t (new_AGEMA_signal_11769), .A1_f (new_AGEMA_signal_11770), .B0_t (stateArray_inS33ser[5]), .B0_f (new_AGEMA_signal_11723), .B1_t (new_AGEMA_signal_11724), .B1_f (new_AGEMA_signal_11725), .Z0_t (ciphertext_s0_t[5]), .Z0_f (ciphertext_s0_f[5]), .Z1_t (ciphertext_s1_t[5]), .Z1_f (ciphertext_s1_f[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S33reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS33ser[6]), .A0_f (new_AGEMA_signal_11726), .A1_t (new_AGEMA_signal_11727), .A1_f (new_AGEMA_signal_11728), .B0_t (ciphertext_s0_t[38]), .B0_f (ciphertext_s0_f[38]), .B1_t (ciphertext_s1_t[38]), .B1_f (ciphertext_s1_f[38]), .Z0_t (stateArray_S33reg_gff_1_SFF_6_MUXInst_X), .Z0_f (new_AGEMA_signal_11750), .Z1_t (new_AGEMA_signal_11751), .Z1_f (new_AGEMA_signal_11752) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S33reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S33reg_gff_1_SFF_6_MUXInst_X), .B0_f (new_AGEMA_signal_11750), .B1_t (new_AGEMA_signal_11751), .B1_f (new_AGEMA_signal_11752), .Z0_t (stateArray_S33reg_gff_1_SFF_6_MUXInst_Y), .Z0_f (new_AGEMA_signal_11771), .Z1_t (new_AGEMA_signal_11772), .Z1_f (new_AGEMA_signal_11773) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S33reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (stateArray_S33reg_gff_1_SFF_6_MUXInst_Y), .A0_f (new_AGEMA_signal_11771), .A1_t (new_AGEMA_signal_11772), .A1_f (new_AGEMA_signal_11773), .B0_t (stateArray_inS33ser[6]), .B0_f (new_AGEMA_signal_11726), .B1_t (new_AGEMA_signal_11727), .B1_f (new_AGEMA_signal_11728), .Z0_t (ciphertext_s0_t[6]), .Z0_f (ciphertext_s0_f[6]), .Z1_t (ciphertext_s1_t[6]), .Z1_f (ciphertext_s1_f[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S33reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS33ser[7]), .A0_f (new_AGEMA_signal_11729), .A1_t (new_AGEMA_signal_11730), .A1_f (new_AGEMA_signal_11731), .B0_t (ciphertext_s0_t[39]), .B0_f (ciphertext_s0_f[39]), .B1_t (ciphertext_s1_t[39]), .B1_f (ciphertext_s1_f[39]), .Z0_t (stateArray_S33reg_gff_1_SFF_7_MUXInst_X), .Z0_f (new_AGEMA_signal_11753), .Z1_t (new_AGEMA_signal_11754), .Z1_f (new_AGEMA_signal_11755) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S33reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (stateArray_S33reg_gff_1_SFF_7_MUXInst_X), .B0_f (new_AGEMA_signal_11753), .B1_t (new_AGEMA_signal_11754), .B1_f (new_AGEMA_signal_11755), .Z0_t (stateArray_S33reg_gff_1_SFF_7_MUXInst_Y), .Z0_f (new_AGEMA_signal_11774), .Z1_t (new_AGEMA_signal_11775), .Z1_f (new_AGEMA_signal_11776) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S33reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (stateArray_S33reg_gff_1_SFF_7_MUXInst_Y), .A0_f (new_AGEMA_signal_11774), .A1_t (new_AGEMA_signal_11775), .A1_f (new_AGEMA_signal_11776), .B0_t (stateArray_inS33ser[7]), .B0_f (new_AGEMA_signal_11729), .B1_t (new_AGEMA_signal_11730), .B1_f (new_AGEMA_signal_11731), .Z0_t (ciphertext_s0_t[7]), .Z0_f (ciphertext_s0_f[7]), .Z1_t (ciphertext_s1_t[7]), .Z1_f (ciphertext_s1_f[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS00ser_mux_inst_0_XOR1_U1 ( .A0_t (plaintext_s0_t[120]), .A0_f (plaintext_s0_f[120]), .A1_t (plaintext_s1_t[120]), .A1_f (plaintext_s1_f[120]), .B0_t (ciphertext_s0_t[88]), .B0_f (ciphertext_s0_f[88]), .B1_t (ciphertext_s1_t[88]), .B1_f (ciphertext_s1_f[88]), .Z0_t (stateArray_MUX_inS00ser_mux_inst_0_X), .Z0_f (new_AGEMA_signal_3528), .Z1_t (new_AGEMA_signal_3529), .Z1_f (new_AGEMA_signal_3530) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS00ser_mux_inst_0_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS00ser_mux_inst_0_X), .B0_f (new_AGEMA_signal_3528), .B1_t (new_AGEMA_signal_3529), .B1_f (new_AGEMA_signal_3530), .Z0_t (stateArray_MUX_inS00ser_mux_inst_0_Y), .Z0_f (new_AGEMA_signal_5824), .Z1_t (new_AGEMA_signal_5825), .Z1_f (new_AGEMA_signal_5826) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS00ser_mux_inst_0_XOR2_U1 ( .A0_t (stateArray_MUX_inS00ser_mux_inst_0_Y), .A0_f (new_AGEMA_signal_5824), .A1_t (new_AGEMA_signal_5825), .A1_f (new_AGEMA_signal_5826), .B0_t (plaintext_s0_t[120]), .B0_f (plaintext_s0_f[120]), .B1_t (plaintext_s1_t[120]), .B1_f (plaintext_s1_f[120]), .Z0_t (stateArray_inS00ser[0]), .Z0_f (new_AGEMA_signal_6622), .Z1_t (new_AGEMA_signal_6623), .Z1_f (new_AGEMA_signal_6624) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS00ser_mux_inst_1_XOR1_U1 ( .A0_t (plaintext_s0_t[121]), .A0_f (plaintext_s0_f[121]), .A1_t (plaintext_s1_t[121]), .A1_f (plaintext_s1_f[121]), .B0_t (ciphertext_s0_t[89]), .B0_f (ciphertext_s0_f[89]), .B1_t (ciphertext_s1_t[89]), .B1_f (ciphertext_s1_f[89]), .Z0_t (stateArray_MUX_inS00ser_mux_inst_1_X), .Z0_f (new_AGEMA_signal_3537), .Z1_t (new_AGEMA_signal_3538), .Z1_f (new_AGEMA_signal_3539) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS00ser_mux_inst_1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS00ser_mux_inst_1_X), .B0_f (new_AGEMA_signal_3537), .B1_t (new_AGEMA_signal_3538), .B1_f (new_AGEMA_signal_3539), .Z0_t (stateArray_MUX_inS00ser_mux_inst_1_Y), .Z0_f (new_AGEMA_signal_5827), .Z1_t (new_AGEMA_signal_5828), .Z1_f (new_AGEMA_signal_5829) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS00ser_mux_inst_1_XOR2_U1 ( .A0_t (stateArray_MUX_inS00ser_mux_inst_1_Y), .A0_f (new_AGEMA_signal_5827), .A1_t (new_AGEMA_signal_5828), .A1_f (new_AGEMA_signal_5829), .B0_t (plaintext_s0_t[121]), .B0_f (plaintext_s0_f[121]), .B1_t (plaintext_s1_t[121]), .B1_f (plaintext_s1_f[121]), .Z0_t (stateArray_inS00ser[1]), .Z0_f (new_AGEMA_signal_6625), .Z1_t (new_AGEMA_signal_6626), .Z1_f (new_AGEMA_signal_6627) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS00ser_mux_inst_2_XOR1_U1 ( .A0_t (plaintext_s0_t[122]), .A0_f (plaintext_s0_f[122]), .A1_t (plaintext_s1_t[122]), .A1_f (plaintext_s1_f[122]), .B0_t (ciphertext_s0_t[90]), .B0_f (ciphertext_s0_f[90]), .B1_t (ciphertext_s1_t[90]), .B1_f (ciphertext_s1_f[90]), .Z0_t (stateArray_MUX_inS00ser_mux_inst_2_X), .Z0_f (new_AGEMA_signal_3546), .Z1_t (new_AGEMA_signal_3547), .Z1_f (new_AGEMA_signal_3548) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS00ser_mux_inst_2_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS00ser_mux_inst_2_X), .B0_f (new_AGEMA_signal_3546), .B1_t (new_AGEMA_signal_3547), .B1_f (new_AGEMA_signal_3548), .Z0_t (stateArray_MUX_inS00ser_mux_inst_2_Y), .Z0_f (new_AGEMA_signal_5830), .Z1_t (new_AGEMA_signal_5831), .Z1_f (new_AGEMA_signal_5832) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS00ser_mux_inst_2_XOR2_U1 ( .A0_t (stateArray_MUX_inS00ser_mux_inst_2_Y), .A0_f (new_AGEMA_signal_5830), .A1_t (new_AGEMA_signal_5831), .A1_f (new_AGEMA_signal_5832), .B0_t (plaintext_s0_t[122]), .B0_f (plaintext_s0_f[122]), .B1_t (plaintext_s1_t[122]), .B1_f (plaintext_s1_f[122]), .Z0_t (stateArray_inS00ser[2]), .Z0_f (new_AGEMA_signal_6628), .Z1_t (new_AGEMA_signal_6629), .Z1_f (new_AGEMA_signal_6630) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS00ser_mux_inst_3_XOR1_U1 ( .A0_t (plaintext_s0_t[123]), .A0_f (plaintext_s0_f[123]), .A1_t (plaintext_s1_t[123]), .A1_f (plaintext_s1_f[123]), .B0_t (ciphertext_s0_t[91]), .B0_f (ciphertext_s0_f[91]), .B1_t (ciphertext_s1_t[91]), .B1_f (ciphertext_s1_f[91]), .Z0_t (stateArray_MUX_inS00ser_mux_inst_3_X), .Z0_f (new_AGEMA_signal_3555), .Z1_t (new_AGEMA_signal_3556), .Z1_f (new_AGEMA_signal_3557) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS00ser_mux_inst_3_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS00ser_mux_inst_3_X), .B0_f (new_AGEMA_signal_3555), .B1_t (new_AGEMA_signal_3556), .B1_f (new_AGEMA_signal_3557), .Z0_t (stateArray_MUX_inS00ser_mux_inst_3_Y), .Z0_f (new_AGEMA_signal_5833), .Z1_t (new_AGEMA_signal_5834), .Z1_f (new_AGEMA_signal_5835) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS00ser_mux_inst_3_XOR2_U1 ( .A0_t (stateArray_MUX_inS00ser_mux_inst_3_Y), .A0_f (new_AGEMA_signal_5833), .A1_t (new_AGEMA_signal_5834), .A1_f (new_AGEMA_signal_5835), .B0_t (plaintext_s0_t[123]), .B0_f (plaintext_s0_f[123]), .B1_t (plaintext_s1_t[123]), .B1_f (plaintext_s1_f[123]), .Z0_t (stateArray_inS00ser[3]), .Z0_f (new_AGEMA_signal_6631), .Z1_t (new_AGEMA_signal_6632), .Z1_f (new_AGEMA_signal_6633) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS00ser_mux_inst_4_XOR1_U1 ( .A0_t (plaintext_s0_t[124]), .A0_f (plaintext_s0_f[124]), .A1_t (plaintext_s1_t[124]), .A1_f (plaintext_s1_f[124]), .B0_t (ciphertext_s0_t[92]), .B0_f (ciphertext_s0_f[92]), .B1_t (ciphertext_s1_t[92]), .B1_f (ciphertext_s1_f[92]), .Z0_t (stateArray_MUX_inS00ser_mux_inst_4_X), .Z0_f (new_AGEMA_signal_3564), .Z1_t (new_AGEMA_signal_3565), .Z1_f (new_AGEMA_signal_3566) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS00ser_mux_inst_4_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS00ser_mux_inst_4_X), .B0_f (new_AGEMA_signal_3564), .B1_t (new_AGEMA_signal_3565), .B1_f (new_AGEMA_signal_3566), .Z0_t (stateArray_MUX_inS00ser_mux_inst_4_Y), .Z0_f (new_AGEMA_signal_5836), .Z1_t (new_AGEMA_signal_5837), .Z1_f (new_AGEMA_signal_5838) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS00ser_mux_inst_4_XOR2_U1 ( .A0_t (stateArray_MUX_inS00ser_mux_inst_4_Y), .A0_f (new_AGEMA_signal_5836), .A1_t (new_AGEMA_signal_5837), .A1_f (new_AGEMA_signal_5838), .B0_t (plaintext_s0_t[124]), .B0_f (plaintext_s0_f[124]), .B1_t (plaintext_s1_t[124]), .B1_f (plaintext_s1_f[124]), .Z0_t (stateArray_inS00ser[4]), .Z0_f (new_AGEMA_signal_6634), .Z1_t (new_AGEMA_signal_6635), .Z1_f (new_AGEMA_signal_6636) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS00ser_mux_inst_5_XOR1_U1 ( .A0_t (plaintext_s0_t[125]), .A0_f (plaintext_s0_f[125]), .A1_t (plaintext_s1_t[125]), .A1_f (plaintext_s1_f[125]), .B0_t (ciphertext_s0_t[93]), .B0_f (ciphertext_s0_f[93]), .B1_t (ciphertext_s1_t[93]), .B1_f (ciphertext_s1_f[93]), .Z0_t (stateArray_MUX_inS00ser_mux_inst_5_X), .Z0_f (new_AGEMA_signal_3573), .Z1_t (new_AGEMA_signal_3574), .Z1_f (new_AGEMA_signal_3575) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS00ser_mux_inst_5_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS00ser_mux_inst_5_X), .B0_f (new_AGEMA_signal_3573), .B1_t (new_AGEMA_signal_3574), .B1_f (new_AGEMA_signal_3575), .Z0_t (stateArray_MUX_inS00ser_mux_inst_5_Y), .Z0_f (new_AGEMA_signal_5839), .Z1_t (new_AGEMA_signal_5840), .Z1_f (new_AGEMA_signal_5841) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS00ser_mux_inst_5_XOR2_U1 ( .A0_t (stateArray_MUX_inS00ser_mux_inst_5_Y), .A0_f (new_AGEMA_signal_5839), .A1_t (new_AGEMA_signal_5840), .A1_f (new_AGEMA_signal_5841), .B0_t (plaintext_s0_t[125]), .B0_f (plaintext_s0_f[125]), .B1_t (plaintext_s1_t[125]), .B1_f (plaintext_s1_f[125]), .Z0_t (stateArray_inS00ser[5]), .Z0_f (new_AGEMA_signal_6637), .Z1_t (new_AGEMA_signal_6638), .Z1_f (new_AGEMA_signal_6639) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS00ser_mux_inst_6_XOR1_U1 ( .A0_t (plaintext_s0_t[126]), .A0_f (plaintext_s0_f[126]), .A1_t (plaintext_s1_t[126]), .A1_f (plaintext_s1_f[126]), .B0_t (ciphertext_s0_t[94]), .B0_f (ciphertext_s0_f[94]), .B1_t (ciphertext_s1_t[94]), .B1_f (ciphertext_s1_f[94]), .Z0_t (stateArray_MUX_inS00ser_mux_inst_6_X), .Z0_f (new_AGEMA_signal_3582), .Z1_t (new_AGEMA_signal_3583), .Z1_f (new_AGEMA_signal_3584) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS00ser_mux_inst_6_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS00ser_mux_inst_6_X), .B0_f (new_AGEMA_signal_3582), .B1_t (new_AGEMA_signal_3583), .B1_f (new_AGEMA_signal_3584), .Z0_t (stateArray_MUX_inS00ser_mux_inst_6_Y), .Z0_f (new_AGEMA_signal_5842), .Z1_t (new_AGEMA_signal_5843), .Z1_f (new_AGEMA_signal_5844) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS00ser_mux_inst_6_XOR2_U1 ( .A0_t (stateArray_MUX_inS00ser_mux_inst_6_Y), .A0_f (new_AGEMA_signal_5842), .A1_t (new_AGEMA_signal_5843), .A1_f (new_AGEMA_signal_5844), .B0_t (plaintext_s0_t[126]), .B0_f (plaintext_s0_f[126]), .B1_t (plaintext_s1_t[126]), .B1_f (plaintext_s1_f[126]), .Z0_t (stateArray_inS00ser[6]), .Z0_f (new_AGEMA_signal_6640), .Z1_t (new_AGEMA_signal_6641), .Z1_f (new_AGEMA_signal_6642) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS00ser_mux_inst_7_XOR1_U1 ( .A0_t (plaintext_s0_t[127]), .A0_f (plaintext_s0_f[127]), .A1_t (plaintext_s1_t[127]), .A1_f (plaintext_s1_f[127]), .B0_t (ciphertext_s0_t[95]), .B0_f (ciphertext_s0_f[95]), .B1_t (ciphertext_s1_t[95]), .B1_f (ciphertext_s1_f[95]), .Z0_t (stateArray_MUX_inS00ser_mux_inst_7_X), .Z0_f (new_AGEMA_signal_3591), .Z1_t (new_AGEMA_signal_3592), .Z1_f (new_AGEMA_signal_3593) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS00ser_mux_inst_7_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS00ser_mux_inst_7_X), .B0_f (new_AGEMA_signal_3591), .B1_t (new_AGEMA_signal_3592), .B1_f (new_AGEMA_signal_3593), .Z0_t (stateArray_MUX_inS00ser_mux_inst_7_Y), .Z0_f (new_AGEMA_signal_5845), .Z1_t (new_AGEMA_signal_5846), .Z1_f (new_AGEMA_signal_5847) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS00ser_mux_inst_7_XOR2_U1 ( .A0_t (stateArray_MUX_inS00ser_mux_inst_7_Y), .A0_f (new_AGEMA_signal_5845), .A1_t (new_AGEMA_signal_5846), .A1_f (new_AGEMA_signal_5847), .B0_t (plaintext_s0_t[127]), .B0_f (plaintext_s0_f[127]), .B1_t (plaintext_s1_t[127]), .B1_f (plaintext_s1_f[127]), .Z0_t (stateArray_inS00ser[7]), .Z0_f (new_AGEMA_signal_6643), .Z1_t (new_AGEMA_signal_6644), .Z1_f (new_AGEMA_signal_6645) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS01ser_mux_inst_0_XOR1_U1 ( .A0_t (plaintext_s0_t[88]), .A0_f (plaintext_s0_f[88]), .A1_t (plaintext_s1_t[88]), .A1_f (plaintext_s1_f[88]), .B0_t (ciphertext_s0_t[56]), .B0_f (ciphertext_s0_f[56]), .B1_t (ciphertext_s1_t[56]), .B1_f (ciphertext_s1_f[56]), .Z0_t (stateArray_MUX_inS01ser_mux_inst_0_X), .Z0_f (new_AGEMA_signal_3600), .Z1_t (new_AGEMA_signal_3601), .Z1_f (new_AGEMA_signal_3602) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS01ser_mux_inst_0_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS01ser_mux_inst_0_X), .B0_f (new_AGEMA_signal_3600), .B1_t (new_AGEMA_signal_3601), .B1_f (new_AGEMA_signal_3602), .Z0_t (stateArray_MUX_inS01ser_mux_inst_0_Y), .Z0_f (new_AGEMA_signal_5848), .Z1_t (new_AGEMA_signal_5849), .Z1_f (new_AGEMA_signal_5850) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS01ser_mux_inst_0_XOR2_U1 ( .A0_t (stateArray_MUX_inS01ser_mux_inst_0_Y), .A0_f (new_AGEMA_signal_5848), .A1_t (new_AGEMA_signal_5849), .A1_f (new_AGEMA_signal_5850), .B0_t (plaintext_s0_t[88]), .B0_f (plaintext_s0_f[88]), .B1_t (plaintext_s1_t[88]), .B1_f (plaintext_s1_f[88]), .Z0_t (stateArray_inS01ser[0]), .Z0_f (new_AGEMA_signal_6646), .Z1_t (new_AGEMA_signal_6647), .Z1_f (new_AGEMA_signal_6648) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS01ser_mux_inst_1_XOR1_U1 ( .A0_t (plaintext_s0_t[89]), .A0_f (plaintext_s0_f[89]), .A1_t (plaintext_s1_t[89]), .A1_f (plaintext_s1_f[89]), .B0_t (ciphertext_s0_t[57]), .B0_f (ciphertext_s0_f[57]), .B1_t (ciphertext_s1_t[57]), .B1_f (ciphertext_s1_f[57]), .Z0_t (stateArray_MUX_inS01ser_mux_inst_1_X), .Z0_f (new_AGEMA_signal_3609), .Z1_t (new_AGEMA_signal_3610), .Z1_f (new_AGEMA_signal_3611) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS01ser_mux_inst_1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS01ser_mux_inst_1_X), .B0_f (new_AGEMA_signal_3609), .B1_t (new_AGEMA_signal_3610), .B1_f (new_AGEMA_signal_3611), .Z0_t (stateArray_MUX_inS01ser_mux_inst_1_Y), .Z0_f (new_AGEMA_signal_5851), .Z1_t (new_AGEMA_signal_5852), .Z1_f (new_AGEMA_signal_5853) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS01ser_mux_inst_1_XOR2_U1 ( .A0_t (stateArray_MUX_inS01ser_mux_inst_1_Y), .A0_f (new_AGEMA_signal_5851), .A1_t (new_AGEMA_signal_5852), .A1_f (new_AGEMA_signal_5853), .B0_t (plaintext_s0_t[89]), .B0_f (plaintext_s0_f[89]), .B1_t (plaintext_s1_t[89]), .B1_f (plaintext_s1_f[89]), .Z0_t (stateArray_inS01ser[1]), .Z0_f (new_AGEMA_signal_6649), .Z1_t (new_AGEMA_signal_6650), .Z1_f (new_AGEMA_signal_6651) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS01ser_mux_inst_2_XOR1_U1 ( .A0_t (plaintext_s0_t[90]), .A0_f (plaintext_s0_f[90]), .A1_t (plaintext_s1_t[90]), .A1_f (plaintext_s1_f[90]), .B0_t (ciphertext_s0_t[58]), .B0_f (ciphertext_s0_f[58]), .B1_t (ciphertext_s1_t[58]), .B1_f (ciphertext_s1_f[58]), .Z0_t (stateArray_MUX_inS01ser_mux_inst_2_X), .Z0_f (new_AGEMA_signal_3618), .Z1_t (new_AGEMA_signal_3619), .Z1_f (new_AGEMA_signal_3620) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS01ser_mux_inst_2_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS01ser_mux_inst_2_X), .B0_f (new_AGEMA_signal_3618), .B1_t (new_AGEMA_signal_3619), .B1_f (new_AGEMA_signal_3620), .Z0_t (stateArray_MUX_inS01ser_mux_inst_2_Y), .Z0_f (new_AGEMA_signal_5854), .Z1_t (new_AGEMA_signal_5855), .Z1_f (new_AGEMA_signal_5856) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS01ser_mux_inst_2_XOR2_U1 ( .A0_t (stateArray_MUX_inS01ser_mux_inst_2_Y), .A0_f (new_AGEMA_signal_5854), .A1_t (new_AGEMA_signal_5855), .A1_f (new_AGEMA_signal_5856), .B0_t (plaintext_s0_t[90]), .B0_f (plaintext_s0_f[90]), .B1_t (plaintext_s1_t[90]), .B1_f (plaintext_s1_f[90]), .Z0_t (stateArray_inS01ser[2]), .Z0_f (new_AGEMA_signal_6652), .Z1_t (new_AGEMA_signal_6653), .Z1_f (new_AGEMA_signal_6654) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS01ser_mux_inst_3_XOR1_U1 ( .A0_t (plaintext_s0_t[91]), .A0_f (plaintext_s0_f[91]), .A1_t (plaintext_s1_t[91]), .A1_f (plaintext_s1_f[91]), .B0_t (ciphertext_s0_t[59]), .B0_f (ciphertext_s0_f[59]), .B1_t (ciphertext_s1_t[59]), .B1_f (ciphertext_s1_f[59]), .Z0_t (stateArray_MUX_inS01ser_mux_inst_3_X), .Z0_f (new_AGEMA_signal_3627), .Z1_t (new_AGEMA_signal_3628), .Z1_f (new_AGEMA_signal_3629) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS01ser_mux_inst_3_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS01ser_mux_inst_3_X), .B0_f (new_AGEMA_signal_3627), .B1_t (new_AGEMA_signal_3628), .B1_f (new_AGEMA_signal_3629), .Z0_t (stateArray_MUX_inS01ser_mux_inst_3_Y), .Z0_f (new_AGEMA_signal_5857), .Z1_t (new_AGEMA_signal_5858), .Z1_f (new_AGEMA_signal_5859) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS01ser_mux_inst_3_XOR2_U1 ( .A0_t (stateArray_MUX_inS01ser_mux_inst_3_Y), .A0_f (new_AGEMA_signal_5857), .A1_t (new_AGEMA_signal_5858), .A1_f (new_AGEMA_signal_5859), .B0_t (plaintext_s0_t[91]), .B0_f (plaintext_s0_f[91]), .B1_t (plaintext_s1_t[91]), .B1_f (plaintext_s1_f[91]), .Z0_t (stateArray_inS01ser[3]), .Z0_f (new_AGEMA_signal_6655), .Z1_t (new_AGEMA_signal_6656), .Z1_f (new_AGEMA_signal_6657) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS01ser_mux_inst_4_XOR1_U1 ( .A0_t (plaintext_s0_t[92]), .A0_f (plaintext_s0_f[92]), .A1_t (plaintext_s1_t[92]), .A1_f (plaintext_s1_f[92]), .B0_t (ciphertext_s0_t[60]), .B0_f (ciphertext_s0_f[60]), .B1_t (ciphertext_s1_t[60]), .B1_f (ciphertext_s1_f[60]), .Z0_t (stateArray_MUX_inS01ser_mux_inst_4_X), .Z0_f (new_AGEMA_signal_3636), .Z1_t (new_AGEMA_signal_3637), .Z1_f (new_AGEMA_signal_3638) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS01ser_mux_inst_4_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS01ser_mux_inst_4_X), .B0_f (new_AGEMA_signal_3636), .B1_t (new_AGEMA_signal_3637), .B1_f (new_AGEMA_signal_3638), .Z0_t (stateArray_MUX_inS01ser_mux_inst_4_Y), .Z0_f (new_AGEMA_signal_5860), .Z1_t (new_AGEMA_signal_5861), .Z1_f (new_AGEMA_signal_5862) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS01ser_mux_inst_4_XOR2_U1 ( .A0_t (stateArray_MUX_inS01ser_mux_inst_4_Y), .A0_f (new_AGEMA_signal_5860), .A1_t (new_AGEMA_signal_5861), .A1_f (new_AGEMA_signal_5862), .B0_t (plaintext_s0_t[92]), .B0_f (plaintext_s0_f[92]), .B1_t (plaintext_s1_t[92]), .B1_f (plaintext_s1_f[92]), .Z0_t (stateArray_inS01ser[4]), .Z0_f (new_AGEMA_signal_6658), .Z1_t (new_AGEMA_signal_6659), .Z1_f (new_AGEMA_signal_6660) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS01ser_mux_inst_5_XOR1_U1 ( .A0_t (plaintext_s0_t[93]), .A0_f (plaintext_s0_f[93]), .A1_t (plaintext_s1_t[93]), .A1_f (plaintext_s1_f[93]), .B0_t (ciphertext_s0_t[61]), .B0_f (ciphertext_s0_f[61]), .B1_t (ciphertext_s1_t[61]), .B1_f (ciphertext_s1_f[61]), .Z0_t (stateArray_MUX_inS01ser_mux_inst_5_X), .Z0_f (new_AGEMA_signal_3645), .Z1_t (new_AGEMA_signal_3646), .Z1_f (new_AGEMA_signal_3647) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS01ser_mux_inst_5_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS01ser_mux_inst_5_X), .B0_f (new_AGEMA_signal_3645), .B1_t (new_AGEMA_signal_3646), .B1_f (new_AGEMA_signal_3647), .Z0_t (stateArray_MUX_inS01ser_mux_inst_5_Y), .Z0_f (new_AGEMA_signal_5863), .Z1_t (new_AGEMA_signal_5864), .Z1_f (new_AGEMA_signal_5865) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS01ser_mux_inst_5_XOR2_U1 ( .A0_t (stateArray_MUX_inS01ser_mux_inst_5_Y), .A0_f (new_AGEMA_signal_5863), .A1_t (new_AGEMA_signal_5864), .A1_f (new_AGEMA_signal_5865), .B0_t (plaintext_s0_t[93]), .B0_f (plaintext_s0_f[93]), .B1_t (plaintext_s1_t[93]), .B1_f (plaintext_s1_f[93]), .Z0_t (stateArray_inS01ser[5]), .Z0_f (new_AGEMA_signal_6661), .Z1_t (new_AGEMA_signal_6662), .Z1_f (new_AGEMA_signal_6663) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS01ser_mux_inst_6_XOR1_U1 ( .A0_t (plaintext_s0_t[94]), .A0_f (plaintext_s0_f[94]), .A1_t (plaintext_s1_t[94]), .A1_f (plaintext_s1_f[94]), .B0_t (ciphertext_s0_t[62]), .B0_f (ciphertext_s0_f[62]), .B1_t (ciphertext_s1_t[62]), .B1_f (ciphertext_s1_f[62]), .Z0_t (stateArray_MUX_inS01ser_mux_inst_6_X), .Z0_f (new_AGEMA_signal_3654), .Z1_t (new_AGEMA_signal_3655), .Z1_f (new_AGEMA_signal_3656) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS01ser_mux_inst_6_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS01ser_mux_inst_6_X), .B0_f (new_AGEMA_signal_3654), .B1_t (new_AGEMA_signal_3655), .B1_f (new_AGEMA_signal_3656), .Z0_t (stateArray_MUX_inS01ser_mux_inst_6_Y), .Z0_f (new_AGEMA_signal_5866), .Z1_t (new_AGEMA_signal_5867), .Z1_f (new_AGEMA_signal_5868) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS01ser_mux_inst_6_XOR2_U1 ( .A0_t (stateArray_MUX_inS01ser_mux_inst_6_Y), .A0_f (new_AGEMA_signal_5866), .A1_t (new_AGEMA_signal_5867), .A1_f (new_AGEMA_signal_5868), .B0_t (plaintext_s0_t[94]), .B0_f (plaintext_s0_f[94]), .B1_t (plaintext_s1_t[94]), .B1_f (plaintext_s1_f[94]), .Z0_t (stateArray_inS01ser[6]), .Z0_f (new_AGEMA_signal_6664), .Z1_t (new_AGEMA_signal_6665), .Z1_f (new_AGEMA_signal_6666) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS01ser_mux_inst_7_XOR1_U1 ( .A0_t (plaintext_s0_t[95]), .A0_f (plaintext_s0_f[95]), .A1_t (plaintext_s1_t[95]), .A1_f (plaintext_s1_f[95]), .B0_t (ciphertext_s0_t[63]), .B0_f (ciphertext_s0_f[63]), .B1_t (ciphertext_s1_t[63]), .B1_f (ciphertext_s1_f[63]), .Z0_t (stateArray_MUX_inS01ser_mux_inst_7_X), .Z0_f (new_AGEMA_signal_3663), .Z1_t (new_AGEMA_signal_3664), .Z1_f (new_AGEMA_signal_3665) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS01ser_mux_inst_7_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS01ser_mux_inst_7_X), .B0_f (new_AGEMA_signal_3663), .B1_t (new_AGEMA_signal_3664), .B1_f (new_AGEMA_signal_3665), .Z0_t (stateArray_MUX_inS01ser_mux_inst_7_Y), .Z0_f (new_AGEMA_signal_5869), .Z1_t (new_AGEMA_signal_5870), .Z1_f (new_AGEMA_signal_5871) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS01ser_mux_inst_7_XOR2_U1 ( .A0_t (stateArray_MUX_inS01ser_mux_inst_7_Y), .A0_f (new_AGEMA_signal_5869), .A1_t (new_AGEMA_signal_5870), .A1_f (new_AGEMA_signal_5871), .B0_t (plaintext_s0_t[95]), .B0_f (plaintext_s0_f[95]), .B1_t (plaintext_s1_t[95]), .B1_f (plaintext_s1_f[95]), .Z0_t (stateArray_inS01ser[7]), .Z0_f (new_AGEMA_signal_6667), .Z1_t (new_AGEMA_signal_6668), .Z1_f (new_AGEMA_signal_6669) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS02ser_mux_inst_0_XOR1_U1 ( .A0_t (plaintext_s0_t[56]), .A0_f (plaintext_s0_f[56]), .A1_t (plaintext_s1_t[56]), .A1_f (plaintext_s1_f[56]), .B0_t (ciphertext_s0_t[24]), .B0_f (ciphertext_s0_f[24]), .B1_t (ciphertext_s1_t[24]), .B1_f (ciphertext_s1_f[24]), .Z0_t (stateArray_MUX_inS02ser_mux_inst_0_X), .Z0_f (new_AGEMA_signal_3672), .Z1_t (new_AGEMA_signal_3673), .Z1_f (new_AGEMA_signal_3674) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS02ser_mux_inst_0_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS02ser_mux_inst_0_X), .B0_f (new_AGEMA_signal_3672), .B1_t (new_AGEMA_signal_3673), .B1_f (new_AGEMA_signal_3674), .Z0_t (stateArray_MUX_inS02ser_mux_inst_0_Y), .Z0_f (new_AGEMA_signal_5872), .Z1_t (new_AGEMA_signal_5873), .Z1_f (new_AGEMA_signal_5874) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS02ser_mux_inst_0_XOR2_U1 ( .A0_t (stateArray_MUX_inS02ser_mux_inst_0_Y), .A0_f (new_AGEMA_signal_5872), .A1_t (new_AGEMA_signal_5873), .A1_f (new_AGEMA_signal_5874), .B0_t (plaintext_s0_t[56]), .B0_f (plaintext_s0_f[56]), .B1_t (plaintext_s1_t[56]), .B1_f (plaintext_s1_f[56]), .Z0_t (stateArray_inS02ser[0]), .Z0_f (new_AGEMA_signal_6670), .Z1_t (new_AGEMA_signal_6671), .Z1_f (new_AGEMA_signal_6672) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS02ser_mux_inst_1_XOR1_U1 ( .A0_t (plaintext_s0_t[57]), .A0_f (plaintext_s0_f[57]), .A1_t (plaintext_s1_t[57]), .A1_f (plaintext_s1_f[57]), .B0_t (ciphertext_s0_t[25]), .B0_f (ciphertext_s0_f[25]), .B1_t (ciphertext_s1_t[25]), .B1_f (ciphertext_s1_f[25]), .Z0_t (stateArray_MUX_inS02ser_mux_inst_1_X), .Z0_f (new_AGEMA_signal_3681), .Z1_t (new_AGEMA_signal_3682), .Z1_f (new_AGEMA_signal_3683) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS02ser_mux_inst_1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS02ser_mux_inst_1_X), .B0_f (new_AGEMA_signal_3681), .B1_t (new_AGEMA_signal_3682), .B1_f (new_AGEMA_signal_3683), .Z0_t (stateArray_MUX_inS02ser_mux_inst_1_Y), .Z0_f (new_AGEMA_signal_5875), .Z1_t (new_AGEMA_signal_5876), .Z1_f (new_AGEMA_signal_5877) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS02ser_mux_inst_1_XOR2_U1 ( .A0_t (stateArray_MUX_inS02ser_mux_inst_1_Y), .A0_f (new_AGEMA_signal_5875), .A1_t (new_AGEMA_signal_5876), .A1_f (new_AGEMA_signal_5877), .B0_t (plaintext_s0_t[57]), .B0_f (plaintext_s0_f[57]), .B1_t (plaintext_s1_t[57]), .B1_f (plaintext_s1_f[57]), .Z0_t (stateArray_inS02ser[1]), .Z0_f (new_AGEMA_signal_6673), .Z1_t (new_AGEMA_signal_6674), .Z1_f (new_AGEMA_signal_6675) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS02ser_mux_inst_2_XOR1_U1 ( .A0_t (plaintext_s0_t[58]), .A0_f (plaintext_s0_f[58]), .A1_t (plaintext_s1_t[58]), .A1_f (plaintext_s1_f[58]), .B0_t (ciphertext_s0_t[26]), .B0_f (ciphertext_s0_f[26]), .B1_t (ciphertext_s1_t[26]), .B1_f (ciphertext_s1_f[26]), .Z0_t (stateArray_MUX_inS02ser_mux_inst_2_X), .Z0_f (new_AGEMA_signal_3690), .Z1_t (new_AGEMA_signal_3691), .Z1_f (new_AGEMA_signal_3692) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS02ser_mux_inst_2_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS02ser_mux_inst_2_X), .B0_f (new_AGEMA_signal_3690), .B1_t (new_AGEMA_signal_3691), .B1_f (new_AGEMA_signal_3692), .Z0_t (stateArray_MUX_inS02ser_mux_inst_2_Y), .Z0_f (new_AGEMA_signal_5878), .Z1_t (new_AGEMA_signal_5879), .Z1_f (new_AGEMA_signal_5880) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS02ser_mux_inst_2_XOR2_U1 ( .A0_t (stateArray_MUX_inS02ser_mux_inst_2_Y), .A0_f (new_AGEMA_signal_5878), .A1_t (new_AGEMA_signal_5879), .A1_f (new_AGEMA_signal_5880), .B0_t (plaintext_s0_t[58]), .B0_f (plaintext_s0_f[58]), .B1_t (plaintext_s1_t[58]), .B1_f (plaintext_s1_f[58]), .Z0_t (stateArray_inS02ser[2]), .Z0_f (new_AGEMA_signal_6676), .Z1_t (new_AGEMA_signal_6677), .Z1_f (new_AGEMA_signal_6678) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS02ser_mux_inst_3_XOR1_U1 ( .A0_t (plaintext_s0_t[59]), .A0_f (plaintext_s0_f[59]), .A1_t (plaintext_s1_t[59]), .A1_f (plaintext_s1_f[59]), .B0_t (ciphertext_s0_t[27]), .B0_f (ciphertext_s0_f[27]), .B1_t (ciphertext_s1_t[27]), .B1_f (ciphertext_s1_f[27]), .Z0_t (stateArray_MUX_inS02ser_mux_inst_3_X), .Z0_f (new_AGEMA_signal_3699), .Z1_t (new_AGEMA_signal_3700), .Z1_f (new_AGEMA_signal_3701) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS02ser_mux_inst_3_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS02ser_mux_inst_3_X), .B0_f (new_AGEMA_signal_3699), .B1_t (new_AGEMA_signal_3700), .B1_f (new_AGEMA_signal_3701), .Z0_t (stateArray_MUX_inS02ser_mux_inst_3_Y), .Z0_f (new_AGEMA_signal_5881), .Z1_t (new_AGEMA_signal_5882), .Z1_f (new_AGEMA_signal_5883) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS02ser_mux_inst_3_XOR2_U1 ( .A0_t (stateArray_MUX_inS02ser_mux_inst_3_Y), .A0_f (new_AGEMA_signal_5881), .A1_t (new_AGEMA_signal_5882), .A1_f (new_AGEMA_signal_5883), .B0_t (plaintext_s0_t[59]), .B0_f (plaintext_s0_f[59]), .B1_t (plaintext_s1_t[59]), .B1_f (plaintext_s1_f[59]), .Z0_t (stateArray_inS02ser[3]), .Z0_f (new_AGEMA_signal_6679), .Z1_t (new_AGEMA_signal_6680), .Z1_f (new_AGEMA_signal_6681) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS02ser_mux_inst_4_XOR1_U1 ( .A0_t (plaintext_s0_t[60]), .A0_f (plaintext_s0_f[60]), .A1_t (plaintext_s1_t[60]), .A1_f (plaintext_s1_f[60]), .B0_t (ciphertext_s0_t[28]), .B0_f (ciphertext_s0_f[28]), .B1_t (ciphertext_s1_t[28]), .B1_f (ciphertext_s1_f[28]), .Z0_t (stateArray_MUX_inS02ser_mux_inst_4_X), .Z0_f (new_AGEMA_signal_3708), .Z1_t (new_AGEMA_signal_3709), .Z1_f (new_AGEMA_signal_3710) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS02ser_mux_inst_4_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS02ser_mux_inst_4_X), .B0_f (new_AGEMA_signal_3708), .B1_t (new_AGEMA_signal_3709), .B1_f (new_AGEMA_signal_3710), .Z0_t (stateArray_MUX_inS02ser_mux_inst_4_Y), .Z0_f (new_AGEMA_signal_5884), .Z1_t (new_AGEMA_signal_5885), .Z1_f (new_AGEMA_signal_5886) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS02ser_mux_inst_4_XOR2_U1 ( .A0_t (stateArray_MUX_inS02ser_mux_inst_4_Y), .A0_f (new_AGEMA_signal_5884), .A1_t (new_AGEMA_signal_5885), .A1_f (new_AGEMA_signal_5886), .B0_t (plaintext_s0_t[60]), .B0_f (plaintext_s0_f[60]), .B1_t (plaintext_s1_t[60]), .B1_f (plaintext_s1_f[60]), .Z0_t (stateArray_inS02ser[4]), .Z0_f (new_AGEMA_signal_6682), .Z1_t (new_AGEMA_signal_6683), .Z1_f (new_AGEMA_signal_6684) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS02ser_mux_inst_5_XOR1_U1 ( .A0_t (plaintext_s0_t[61]), .A0_f (plaintext_s0_f[61]), .A1_t (plaintext_s1_t[61]), .A1_f (plaintext_s1_f[61]), .B0_t (ciphertext_s0_t[29]), .B0_f (ciphertext_s0_f[29]), .B1_t (ciphertext_s1_t[29]), .B1_f (ciphertext_s1_f[29]), .Z0_t (stateArray_MUX_inS02ser_mux_inst_5_X), .Z0_f (new_AGEMA_signal_3717), .Z1_t (new_AGEMA_signal_3718), .Z1_f (new_AGEMA_signal_3719) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS02ser_mux_inst_5_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS02ser_mux_inst_5_X), .B0_f (new_AGEMA_signal_3717), .B1_t (new_AGEMA_signal_3718), .B1_f (new_AGEMA_signal_3719), .Z0_t (stateArray_MUX_inS02ser_mux_inst_5_Y), .Z0_f (new_AGEMA_signal_5887), .Z1_t (new_AGEMA_signal_5888), .Z1_f (new_AGEMA_signal_5889) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS02ser_mux_inst_5_XOR2_U1 ( .A0_t (stateArray_MUX_inS02ser_mux_inst_5_Y), .A0_f (new_AGEMA_signal_5887), .A1_t (new_AGEMA_signal_5888), .A1_f (new_AGEMA_signal_5889), .B0_t (plaintext_s0_t[61]), .B0_f (plaintext_s0_f[61]), .B1_t (plaintext_s1_t[61]), .B1_f (plaintext_s1_f[61]), .Z0_t (stateArray_inS02ser[5]), .Z0_f (new_AGEMA_signal_6685), .Z1_t (new_AGEMA_signal_6686), .Z1_f (new_AGEMA_signal_6687) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS02ser_mux_inst_6_XOR1_U1 ( .A0_t (plaintext_s0_t[62]), .A0_f (plaintext_s0_f[62]), .A1_t (plaintext_s1_t[62]), .A1_f (plaintext_s1_f[62]), .B0_t (ciphertext_s0_t[30]), .B0_f (ciphertext_s0_f[30]), .B1_t (ciphertext_s1_t[30]), .B1_f (ciphertext_s1_f[30]), .Z0_t (stateArray_MUX_inS02ser_mux_inst_6_X), .Z0_f (new_AGEMA_signal_3726), .Z1_t (new_AGEMA_signal_3727), .Z1_f (new_AGEMA_signal_3728) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS02ser_mux_inst_6_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS02ser_mux_inst_6_X), .B0_f (new_AGEMA_signal_3726), .B1_t (new_AGEMA_signal_3727), .B1_f (new_AGEMA_signal_3728), .Z0_t (stateArray_MUX_inS02ser_mux_inst_6_Y), .Z0_f (new_AGEMA_signal_5890), .Z1_t (new_AGEMA_signal_5891), .Z1_f (new_AGEMA_signal_5892) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS02ser_mux_inst_6_XOR2_U1 ( .A0_t (stateArray_MUX_inS02ser_mux_inst_6_Y), .A0_f (new_AGEMA_signal_5890), .A1_t (new_AGEMA_signal_5891), .A1_f (new_AGEMA_signal_5892), .B0_t (plaintext_s0_t[62]), .B0_f (plaintext_s0_f[62]), .B1_t (plaintext_s1_t[62]), .B1_f (plaintext_s1_f[62]), .Z0_t (stateArray_inS02ser[6]), .Z0_f (new_AGEMA_signal_6688), .Z1_t (new_AGEMA_signal_6689), .Z1_f (new_AGEMA_signal_6690) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS02ser_mux_inst_7_XOR1_U1 ( .A0_t (plaintext_s0_t[63]), .A0_f (plaintext_s0_f[63]), .A1_t (plaintext_s1_t[63]), .A1_f (plaintext_s1_f[63]), .B0_t (ciphertext_s0_t[31]), .B0_f (ciphertext_s0_f[31]), .B1_t (ciphertext_s1_t[31]), .B1_f (ciphertext_s1_f[31]), .Z0_t (stateArray_MUX_inS02ser_mux_inst_7_X), .Z0_f (new_AGEMA_signal_3735), .Z1_t (new_AGEMA_signal_3736), .Z1_f (new_AGEMA_signal_3737) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS02ser_mux_inst_7_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS02ser_mux_inst_7_X), .B0_f (new_AGEMA_signal_3735), .B1_t (new_AGEMA_signal_3736), .B1_f (new_AGEMA_signal_3737), .Z0_t (stateArray_MUX_inS02ser_mux_inst_7_Y), .Z0_f (new_AGEMA_signal_5893), .Z1_t (new_AGEMA_signal_5894), .Z1_f (new_AGEMA_signal_5895) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS02ser_mux_inst_7_XOR2_U1 ( .A0_t (stateArray_MUX_inS02ser_mux_inst_7_Y), .A0_f (new_AGEMA_signal_5893), .A1_t (new_AGEMA_signal_5894), .A1_f (new_AGEMA_signal_5895), .B0_t (plaintext_s0_t[63]), .B0_f (plaintext_s0_f[63]), .B1_t (plaintext_s1_t[63]), .B1_f (plaintext_s1_f[63]), .Z0_t (stateArray_inS02ser[7]), .Z0_f (new_AGEMA_signal_6691), .Z1_t (new_AGEMA_signal_6692), .Z1_f (new_AGEMA_signal_6693) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS10_MC_mux_inst_0_XOR1_U1 ( .A0_t (ciphertext_s0_t[112]), .A0_f (ciphertext_s0_f[112]), .A1_t (ciphertext_s1_t[112]), .A1_f (ciphertext_s1_f[112]), .B0_t (StateInMC[24]), .B0_f (new_AGEMA_signal_9376), .B1_t (new_AGEMA_signal_9377), .B1_f (new_AGEMA_signal_9378), .Z0_t (stateArray_MUX_outS10_MC_mux_inst_0_X), .Z0_f (new_AGEMA_signal_9795), .Z1_t (new_AGEMA_signal_9796), .Z1_f (new_AGEMA_signal_9797) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS10_MC_mux_inst_0_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (stateArray_MUX_outS10_MC_mux_inst_0_X), .B0_f (new_AGEMA_signal_9795), .B1_t (new_AGEMA_signal_9796), .B1_f (new_AGEMA_signal_9797), .Z0_t (stateArray_MUX_outS10_MC_mux_inst_0_Y), .Z0_f (new_AGEMA_signal_10307), .Z1_t (new_AGEMA_signal_10308), .Z1_f (new_AGEMA_signal_10309) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS10_MC_mux_inst_0_XOR2_U1 ( .A0_t (stateArray_MUX_outS10_MC_mux_inst_0_Y), .A0_f (new_AGEMA_signal_10307), .A1_t (new_AGEMA_signal_10308), .A1_f (new_AGEMA_signal_10309), .B0_t (ciphertext_s0_t[112]), .B0_f (ciphertext_s0_f[112]), .B1_t (ciphertext_s1_t[112]), .B1_f (ciphertext_s1_f[112]), .Z0_t (stateArray_outS10ser_MC[0]), .Z0_f (new_AGEMA_signal_10430), .Z1_t (new_AGEMA_signal_10431), .Z1_f (new_AGEMA_signal_10432) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS10_MC_mux_inst_1_XOR1_U1 ( .A0_t (ciphertext_s0_t[113]), .A0_f (ciphertext_s0_f[113]), .A1_t (ciphertext_s1_t[113]), .A1_f (ciphertext_s1_f[113]), .B0_t (StateInMC[25]), .B0_f (new_AGEMA_signal_9867), .B1_t (new_AGEMA_signal_9868), .B1_f (new_AGEMA_signal_9869), .Z0_t (stateArray_MUX_outS10_MC_mux_inst_1_X), .Z0_f (new_AGEMA_signal_10310), .Z1_t (new_AGEMA_signal_10311), .Z1_f (new_AGEMA_signal_10312) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS10_MC_mux_inst_1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (stateArray_MUX_outS10_MC_mux_inst_1_X), .B0_f (new_AGEMA_signal_10310), .B1_t (new_AGEMA_signal_10311), .B1_f (new_AGEMA_signal_10312), .Z0_t (stateArray_MUX_outS10_MC_mux_inst_1_Y), .Z0_f (new_AGEMA_signal_10433), .Z1_t (new_AGEMA_signal_10434), .Z1_f (new_AGEMA_signal_10435) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS10_MC_mux_inst_1_XOR2_U1 ( .A0_t (stateArray_MUX_outS10_MC_mux_inst_1_Y), .A0_f (new_AGEMA_signal_10433), .A1_t (new_AGEMA_signal_10434), .A1_f (new_AGEMA_signal_10435), .B0_t (ciphertext_s0_t[113]), .B0_f (ciphertext_s0_f[113]), .B1_t (ciphertext_s1_t[113]), .B1_f (ciphertext_s1_f[113]), .Z0_t (stateArray_outS10ser_MC[1]), .Z0_f (new_AGEMA_signal_10541), .Z1_t (new_AGEMA_signal_10542), .Z1_f (new_AGEMA_signal_10543) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS10_MC_mux_inst_2_XOR1_U1 ( .A0_t (ciphertext_s0_t[114]), .A0_f (ciphertext_s0_f[114]), .A1_t (ciphertext_s1_t[114]), .A1_f (ciphertext_s1_f[114]), .B0_t (StateInMC[26]), .B0_f (new_AGEMA_signal_9382), .B1_t (new_AGEMA_signal_9383), .B1_f (new_AGEMA_signal_9384), .Z0_t (stateArray_MUX_outS10_MC_mux_inst_2_X), .Z0_f (new_AGEMA_signal_9798), .Z1_t (new_AGEMA_signal_9799), .Z1_f (new_AGEMA_signal_9800) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS10_MC_mux_inst_2_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (stateArray_MUX_outS10_MC_mux_inst_2_X), .B0_f (new_AGEMA_signal_9798), .B1_t (new_AGEMA_signal_9799), .B1_f (new_AGEMA_signal_9800), .Z0_t (stateArray_MUX_outS10_MC_mux_inst_2_Y), .Z0_f (new_AGEMA_signal_10313), .Z1_t (new_AGEMA_signal_10314), .Z1_f (new_AGEMA_signal_10315) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS10_MC_mux_inst_2_XOR2_U1 ( .A0_t (stateArray_MUX_outS10_MC_mux_inst_2_Y), .A0_f (new_AGEMA_signal_10313), .A1_t (new_AGEMA_signal_10314), .A1_f (new_AGEMA_signal_10315), .B0_t (ciphertext_s0_t[114]), .B0_f (ciphertext_s0_f[114]), .B1_t (ciphertext_s1_t[114]), .B1_f (ciphertext_s1_f[114]), .Z0_t (stateArray_outS10ser_MC[2]), .Z0_f (new_AGEMA_signal_10436), .Z1_t (new_AGEMA_signal_10437), .Z1_f (new_AGEMA_signal_10438) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS10_MC_mux_inst_3_XOR1_U1 ( .A0_t (ciphertext_s0_t[115]), .A0_f (ciphertext_s0_f[115]), .A1_t (ciphertext_s1_t[115]), .A1_f (ciphertext_s1_f[115]), .B0_t (StateInMC[27]), .B0_f (new_AGEMA_signal_9870), .B1_t (new_AGEMA_signal_9871), .B1_f (new_AGEMA_signal_9872), .Z0_t (stateArray_MUX_outS10_MC_mux_inst_3_X), .Z0_f (new_AGEMA_signal_10316), .Z1_t (new_AGEMA_signal_10317), .Z1_f (new_AGEMA_signal_10318) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS10_MC_mux_inst_3_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (stateArray_MUX_outS10_MC_mux_inst_3_X), .B0_f (new_AGEMA_signal_10316), .B1_t (new_AGEMA_signal_10317), .B1_f (new_AGEMA_signal_10318), .Z0_t (stateArray_MUX_outS10_MC_mux_inst_3_Y), .Z0_f (new_AGEMA_signal_10439), .Z1_t (new_AGEMA_signal_10440), .Z1_f (new_AGEMA_signal_10441) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS10_MC_mux_inst_3_XOR2_U1 ( .A0_t (stateArray_MUX_outS10_MC_mux_inst_3_Y), .A0_f (new_AGEMA_signal_10439), .A1_t (new_AGEMA_signal_10440), .A1_f (new_AGEMA_signal_10441), .B0_t (ciphertext_s0_t[115]), .B0_f (ciphertext_s0_f[115]), .B1_t (ciphertext_s1_t[115]), .B1_f (ciphertext_s1_f[115]), .Z0_t (stateArray_outS10ser_MC[3]), .Z0_f (new_AGEMA_signal_10544), .Z1_t (new_AGEMA_signal_10545), .Z1_f (new_AGEMA_signal_10546) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS10_MC_mux_inst_4_XOR1_U1 ( .A0_t (ciphertext_s0_t[116]), .A0_f (ciphertext_s0_f[116]), .A1_t (ciphertext_s1_t[116]), .A1_f (ciphertext_s1_f[116]), .B0_t (StateInMC[28]), .B0_f (new_AGEMA_signal_9873), .B1_t (new_AGEMA_signal_9874), .B1_f (new_AGEMA_signal_9875), .Z0_t (stateArray_MUX_outS10_MC_mux_inst_4_X), .Z0_f (new_AGEMA_signal_10319), .Z1_t (new_AGEMA_signal_10320), .Z1_f (new_AGEMA_signal_10321) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS10_MC_mux_inst_4_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (stateArray_MUX_outS10_MC_mux_inst_4_X), .B0_f (new_AGEMA_signal_10319), .B1_t (new_AGEMA_signal_10320), .B1_f (new_AGEMA_signal_10321), .Z0_t (stateArray_MUX_outS10_MC_mux_inst_4_Y), .Z0_f (new_AGEMA_signal_10442), .Z1_t (new_AGEMA_signal_10443), .Z1_f (new_AGEMA_signal_10444) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS10_MC_mux_inst_4_XOR2_U1 ( .A0_t (stateArray_MUX_outS10_MC_mux_inst_4_Y), .A0_f (new_AGEMA_signal_10442), .A1_t (new_AGEMA_signal_10443), .A1_f (new_AGEMA_signal_10444), .B0_t (ciphertext_s0_t[116]), .B0_f (ciphertext_s0_f[116]), .B1_t (ciphertext_s1_t[116]), .B1_f (ciphertext_s1_f[116]), .Z0_t (stateArray_outS10ser_MC[4]), .Z0_f (new_AGEMA_signal_10547), .Z1_t (new_AGEMA_signal_10548), .Z1_f (new_AGEMA_signal_10549) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS10_MC_mux_inst_5_XOR1_U1 ( .A0_t (ciphertext_s0_t[117]), .A0_f (ciphertext_s0_f[117]), .A1_t (ciphertext_s1_t[117]), .A1_f (ciphertext_s1_f[117]), .B0_t (StateInMC[29]), .B0_f (new_AGEMA_signal_9391), .B1_t (new_AGEMA_signal_9392), .B1_f (new_AGEMA_signal_9393), .Z0_t (stateArray_MUX_outS10_MC_mux_inst_5_X), .Z0_f (new_AGEMA_signal_9801), .Z1_t (new_AGEMA_signal_9802), .Z1_f (new_AGEMA_signal_9803) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS10_MC_mux_inst_5_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (stateArray_MUX_outS10_MC_mux_inst_5_X), .B0_f (new_AGEMA_signal_9801), .B1_t (new_AGEMA_signal_9802), .B1_f (new_AGEMA_signal_9803), .Z0_t (stateArray_MUX_outS10_MC_mux_inst_5_Y), .Z0_f (new_AGEMA_signal_10322), .Z1_t (new_AGEMA_signal_10323), .Z1_f (new_AGEMA_signal_10324) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS10_MC_mux_inst_5_XOR2_U1 ( .A0_t (stateArray_MUX_outS10_MC_mux_inst_5_Y), .A0_f (new_AGEMA_signal_10322), .A1_t (new_AGEMA_signal_10323), .A1_f (new_AGEMA_signal_10324), .B0_t (ciphertext_s0_t[117]), .B0_f (ciphertext_s0_f[117]), .B1_t (ciphertext_s1_t[117]), .B1_f (ciphertext_s1_f[117]), .Z0_t (stateArray_outS10ser_MC[5]), .Z0_f (new_AGEMA_signal_10445), .Z1_t (new_AGEMA_signal_10446), .Z1_f (new_AGEMA_signal_10447) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS10_MC_mux_inst_6_XOR1_U1 ( .A0_t (ciphertext_s0_t[118]), .A0_f (ciphertext_s0_f[118]), .A1_t (ciphertext_s1_t[118]), .A1_f (ciphertext_s1_f[118]), .B0_t (StateInMC[30]), .B0_f (new_AGEMA_signal_9394), .B1_t (new_AGEMA_signal_9395), .B1_f (new_AGEMA_signal_9396), .Z0_t (stateArray_MUX_outS10_MC_mux_inst_6_X), .Z0_f (new_AGEMA_signal_9804), .Z1_t (new_AGEMA_signal_9805), .Z1_f (new_AGEMA_signal_9806) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS10_MC_mux_inst_6_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (stateArray_MUX_outS10_MC_mux_inst_6_X), .B0_f (new_AGEMA_signal_9804), .B1_t (new_AGEMA_signal_9805), .B1_f (new_AGEMA_signal_9806), .Z0_t (stateArray_MUX_outS10_MC_mux_inst_6_Y), .Z0_f (new_AGEMA_signal_10325), .Z1_t (new_AGEMA_signal_10326), .Z1_f (new_AGEMA_signal_10327) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS10_MC_mux_inst_6_XOR2_U1 ( .A0_t (stateArray_MUX_outS10_MC_mux_inst_6_Y), .A0_f (new_AGEMA_signal_10325), .A1_t (new_AGEMA_signal_10326), .A1_f (new_AGEMA_signal_10327), .B0_t (ciphertext_s0_t[118]), .B0_f (ciphertext_s0_f[118]), .B1_t (ciphertext_s1_t[118]), .B1_f (ciphertext_s1_f[118]), .Z0_t (stateArray_outS10ser_MC[6]), .Z0_f (new_AGEMA_signal_10448), .Z1_t (new_AGEMA_signal_10449), .Z1_f (new_AGEMA_signal_10450) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS10_MC_mux_inst_7_XOR1_U1 ( .A0_t (ciphertext_s0_t[119]), .A0_f (ciphertext_s0_f[119]), .A1_t (ciphertext_s1_t[119]), .A1_f (ciphertext_s1_f[119]), .B0_t (StateInMC[31]), .B0_f (new_AGEMA_signal_9397), .B1_t (new_AGEMA_signal_9398), .B1_f (new_AGEMA_signal_9399), .Z0_t (stateArray_MUX_outS10_MC_mux_inst_7_X), .Z0_f (new_AGEMA_signal_9807), .Z1_t (new_AGEMA_signal_9808), .Z1_f (new_AGEMA_signal_9809) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS10_MC_mux_inst_7_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (stateArray_MUX_outS10_MC_mux_inst_7_X), .B0_f (new_AGEMA_signal_9807), .B1_t (new_AGEMA_signal_9808), .B1_f (new_AGEMA_signal_9809), .Z0_t (stateArray_MUX_outS10_MC_mux_inst_7_Y), .Z0_f (new_AGEMA_signal_10328), .Z1_t (new_AGEMA_signal_10329), .Z1_f (new_AGEMA_signal_10330) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS10_MC_mux_inst_7_XOR2_U1 ( .A0_t (stateArray_MUX_outS10_MC_mux_inst_7_Y), .A0_f (new_AGEMA_signal_10328), .A1_t (new_AGEMA_signal_10329), .A1_f (new_AGEMA_signal_10330), .B0_t (ciphertext_s0_t[119]), .B0_f (ciphertext_s0_f[119]), .B1_t (ciphertext_s1_t[119]), .B1_f (ciphertext_s1_f[119]), .Z0_t (stateArray_outS10ser_MC[7]), .Z0_f (new_AGEMA_signal_10451), .Z1_t (new_AGEMA_signal_10452), .Z1_f (new_AGEMA_signal_10453) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_0_XOR1_U1 ( .A0_t (plaintext_s0_t[24]), .A0_f (plaintext_s0_f[24]), .A1_t (plaintext_s1_t[24]), .A1_f (plaintext_s1_f[24]), .B0_t (stateArray_outS10ser_MC[0]), .B0_f (new_AGEMA_signal_10430), .B1_t (new_AGEMA_signal_10431), .B1_f (new_AGEMA_signal_10432), .Z0_t (stateArray_MUX_inS03ser_mux_inst_0_X), .Z0_f (new_AGEMA_signal_10553), .Z1_t (new_AGEMA_signal_10554), .Z1_f (new_AGEMA_signal_10555) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_0_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS03ser_mux_inst_0_X), .B0_f (new_AGEMA_signal_10553), .B1_t (new_AGEMA_signal_10554), .B1_f (new_AGEMA_signal_10555), .Z0_t (stateArray_MUX_inS03ser_mux_inst_0_Y), .Z0_f (new_AGEMA_signal_10694), .Z1_t (new_AGEMA_signal_10695), .Z1_f (new_AGEMA_signal_10696) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_0_XOR2_U1 ( .A0_t (stateArray_MUX_inS03ser_mux_inst_0_Y), .A0_f (new_AGEMA_signal_10694), .A1_t (new_AGEMA_signal_10695), .A1_f (new_AGEMA_signal_10696), .B0_t (plaintext_s0_t[24]), .B0_f (plaintext_s0_f[24]), .B1_t (plaintext_s1_t[24]), .B1_f (plaintext_s1_f[24]), .Z0_t (stateArray_inS03ser[0]), .Z0_f (new_AGEMA_signal_10829), .Z1_t (new_AGEMA_signal_10830), .Z1_f (new_AGEMA_signal_10831) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_1_XOR1_U1 ( .A0_t (plaintext_s0_t[25]), .A0_f (plaintext_s0_f[25]), .A1_t (plaintext_s1_t[25]), .A1_f (plaintext_s1_f[25]), .B0_t (stateArray_outS10ser_MC[1]), .B0_f (new_AGEMA_signal_10541), .B1_t (new_AGEMA_signal_10542), .B1_f (new_AGEMA_signal_10543), .Z0_t (stateArray_MUX_inS03ser_mux_inst_1_X), .Z0_f (new_AGEMA_signal_10700), .Z1_t (new_AGEMA_signal_10701), .Z1_f (new_AGEMA_signal_10702) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS03ser_mux_inst_1_X), .B0_f (new_AGEMA_signal_10700), .B1_t (new_AGEMA_signal_10701), .B1_f (new_AGEMA_signal_10702), .Z0_t (stateArray_MUX_inS03ser_mux_inst_1_Y), .Z0_f (new_AGEMA_signal_10832), .Z1_t (new_AGEMA_signal_10833), .Z1_f (new_AGEMA_signal_10834) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_1_XOR2_U1 ( .A0_t (stateArray_MUX_inS03ser_mux_inst_1_Y), .A0_f (new_AGEMA_signal_10832), .A1_t (new_AGEMA_signal_10833), .A1_f (new_AGEMA_signal_10834), .B0_t (plaintext_s0_t[25]), .B0_f (plaintext_s0_f[25]), .B1_t (plaintext_s1_t[25]), .B1_f (plaintext_s1_f[25]), .Z0_t (stateArray_inS03ser[1]), .Z0_f (new_AGEMA_signal_10985), .Z1_t (new_AGEMA_signal_10986), .Z1_f (new_AGEMA_signal_10987) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_2_XOR1_U1 ( .A0_t (plaintext_s0_t[26]), .A0_f (plaintext_s0_f[26]), .A1_t (plaintext_s1_t[26]), .A1_f (plaintext_s1_f[26]), .B0_t (stateArray_outS10ser_MC[2]), .B0_f (new_AGEMA_signal_10436), .B1_t (new_AGEMA_signal_10437), .B1_f (new_AGEMA_signal_10438), .Z0_t (stateArray_MUX_inS03ser_mux_inst_2_X), .Z0_f (new_AGEMA_signal_10559), .Z1_t (new_AGEMA_signal_10560), .Z1_f (new_AGEMA_signal_10561) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_2_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS03ser_mux_inst_2_X), .B0_f (new_AGEMA_signal_10559), .B1_t (new_AGEMA_signal_10560), .B1_f (new_AGEMA_signal_10561), .Z0_t (stateArray_MUX_inS03ser_mux_inst_2_Y), .Z0_f (new_AGEMA_signal_10703), .Z1_t (new_AGEMA_signal_10704), .Z1_f (new_AGEMA_signal_10705) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_2_XOR2_U1 ( .A0_t (stateArray_MUX_inS03ser_mux_inst_2_Y), .A0_f (new_AGEMA_signal_10703), .A1_t (new_AGEMA_signal_10704), .A1_f (new_AGEMA_signal_10705), .B0_t (plaintext_s0_t[26]), .B0_f (plaintext_s0_f[26]), .B1_t (plaintext_s1_t[26]), .B1_f (plaintext_s1_f[26]), .Z0_t (stateArray_inS03ser[2]), .Z0_f (new_AGEMA_signal_10835), .Z1_t (new_AGEMA_signal_10836), .Z1_f (new_AGEMA_signal_10837) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_3_XOR1_U1 ( .A0_t (plaintext_s0_t[27]), .A0_f (plaintext_s0_f[27]), .A1_t (plaintext_s1_t[27]), .A1_f (plaintext_s1_f[27]), .B0_t (stateArray_outS10ser_MC[3]), .B0_f (new_AGEMA_signal_10544), .B1_t (new_AGEMA_signal_10545), .B1_f (new_AGEMA_signal_10546), .Z0_t (stateArray_MUX_inS03ser_mux_inst_3_X), .Z0_f (new_AGEMA_signal_10709), .Z1_t (new_AGEMA_signal_10710), .Z1_f (new_AGEMA_signal_10711) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_3_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS03ser_mux_inst_3_X), .B0_f (new_AGEMA_signal_10709), .B1_t (new_AGEMA_signal_10710), .B1_f (new_AGEMA_signal_10711), .Z0_t (stateArray_MUX_inS03ser_mux_inst_3_Y), .Z0_f (new_AGEMA_signal_10838), .Z1_t (new_AGEMA_signal_10839), .Z1_f (new_AGEMA_signal_10840) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_3_XOR2_U1 ( .A0_t (stateArray_MUX_inS03ser_mux_inst_3_Y), .A0_f (new_AGEMA_signal_10838), .A1_t (new_AGEMA_signal_10839), .A1_f (new_AGEMA_signal_10840), .B0_t (plaintext_s0_t[27]), .B0_f (plaintext_s0_f[27]), .B1_t (plaintext_s1_t[27]), .B1_f (plaintext_s1_f[27]), .Z0_t (stateArray_inS03ser[3]), .Z0_f (new_AGEMA_signal_10988), .Z1_t (new_AGEMA_signal_10989), .Z1_f (new_AGEMA_signal_10990) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_4_XOR1_U1 ( .A0_t (plaintext_s0_t[28]), .A0_f (plaintext_s0_f[28]), .A1_t (plaintext_s1_t[28]), .A1_f (plaintext_s1_f[28]), .B0_t (stateArray_outS10ser_MC[4]), .B0_f (new_AGEMA_signal_10547), .B1_t (new_AGEMA_signal_10548), .B1_f (new_AGEMA_signal_10549), .Z0_t (stateArray_MUX_inS03ser_mux_inst_4_X), .Z0_f (new_AGEMA_signal_10715), .Z1_t (new_AGEMA_signal_10716), .Z1_f (new_AGEMA_signal_10717) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_4_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS03ser_mux_inst_4_X), .B0_f (new_AGEMA_signal_10715), .B1_t (new_AGEMA_signal_10716), .B1_f (new_AGEMA_signal_10717), .Z0_t (stateArray_MUX_inS03ser_mux_inst_4_Y), .Z0_f (new_AGEMA_signal_10841), .Z1_t (new_AGEMA_signal_10842), .Z1_f (new_AGEMA_signal_10843) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_4_XOR2_U1 ( .A0_t (stateArray_MUX_inS03ser_mux_inst_4_Y), .A0_f (new_AGEMA_signal_10841), .A1_t (new_AGEMA_signal_10842), .A1_f (new_AGEMA_signal_10843), .B0_t (plaintext_s0_t[28]), .B0_f (plaintext_s0_f[28]), .B1_t (plaintext_s1_t[28]), .B1_f (plaintext_s1_f[28]), .Z0_t (stateArray_inS03ser[4]), .Z0_f (new_AGEMA_signal_10991), .Z1_t (new_AGEMA_signal_10992), .Z1_f (new_AGEMA_signal_10993) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_5_XOR1_U1 ( .A0_t (plaintext_s0_t[29]), .A0_f (plaintext_s0_f[29]), .A1_t (plaintext_s1_t[29]), .A1_f (plaintext_s1_f[29]), .B0_t (stateArray_outS10ser_MC[5]), .B0_f (new_AGEMA_signal_10445), .B1_t (new_AGEMA_signal_10446), .B1_f (new_AGEMA_signal_10447), .Z0_t (stateArray_MUX_inS03ser_mux_inst_5_X), .Z0_f (new_AGEMA_signal_10565), .Z1_t (new_AGEMA_signal_10566), .Z1_f (new_AGEMA_signal_10567) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_5_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS03ser_mux_inst_5_X), .B0_f (new_AGEMA_signal_10565), .B1_t (new_AGEMA_signal_10566), .B1_f (new_AGEMA_signal_10567), .Z0_t (stateArray_MUX_inS03ser_mux_inst_5_Y), .Z0_f (new_AGEMA_signal_10718), .Z1_t (new_AGEMA_signal_10719), .Z1_f (new_AGEMA_signal_10720) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_5_XOR2_U1 ( .A0_t (stateArray_MUX_inS03ser_mux_inst_5_Y), .A0_f (new_AGEMA_signal_10718), .A1_t (new_AGEMA_signal_10719), .A1_f (new_AGEMA_signal_10720), .B0_t (plaintext_s0_t[29]), .B0_f (plaintext_s0_f[29]), .B1_t (plaintext_s1_t[29]), .B1_f (plaintext_s1_f[29]), .Z0_t (stateArray_inS03ser[5]), .Z0_f (new_AGEMA_signal_10844), .Z1_t (new_AGEMA_signal_10845), .Z1_f (new_AGEMA_signal_10846) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_6_XOR1_U1 ( .A0_t (plaintext_s0_t[30]), .A0_f (plaintext_s0_f[30]), .A1_t (plaintext_s1_t[30]), .A1_f (plaintext_s1_f[30]), .B0_t (stateArray_outS10ser_MC[6]), .B0_f (new_AGEMA_signal_10448), .B1_t (new_AGEMA_signal_10449), .B1_f (new_AGEMA_signal_10450), .Z0_t (stateArray_MUX_inS03ser_mux_inst_6_X), .Z0_f (new_AGEMA_signal_10571), .Z1_t (new_AGEMA_signal_10572), .Z1_f (new_AGEMA_signal_10573) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_6_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS03ser_mux_inst_6_X), .B0_f (new_AGEMA_signal_10571), .B1_t (new_AGEMA_signal_10572), .B1_f (new_AGEMA_signal_10573), .Z0_t (stateArray_MUX_inS03ser_mux_inst_6_Y), .Z0_f (new_AGEMA_signal_10721), .Z1_t (new_AGEMA_signal_10722), .Z1_f (new_AGEMA_signal_10723) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_6_XOR2_U1 ( .A0_t (stateArray_MUX_inS03ser_mux_inst_6_Y), .A0_f (new_AGEMA_signal_10721), .A1_t (new_AGEMA_signal_10722), .A1_f (new_AGEMA_signal_10723), .B0_t (plaintext_s0_t[30]), .B0_f (plaintext_s0_f[30]), .B1_t (plaintext_s1_t[30]), .B1_f (plaintext_s1_f[30]), .Z0_t (stateArray_inS03ser[6]), .Z0_f (new_AGEMA_signal_10847), .Z1_t (new_AGEMA_signal_10848), .Z1_f (new_AGEMA_signal_10849) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_7_XOR1_U1 ( .A0_t (plaintext_s0_t[31]), .A0_f (plaintext_s0_f[31]), .A1_t (plaintext_s1_t[31]), .A1_f (plaintext_s1_f[31]), .B0_t (stateArray_outS10ser_MC[7]), .B0_f (new_AGEMA_signal_10451), .B1_t (new_AGEMA_signal_10452), .B1_f (new_AGEMA_signal_10453), .Z0_t (stateArray_MUX_inS03ser_mux_inst_7_X), .Z0_f (new_AGEMA_signal_10577), .Z1_t (new_AGEMA_signal_10578), .Z1_f (new_AGEMA_signal_10579) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_7_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS03ser_mux_inst_7_X), .B0_f (new_AGEMA_signal_10577), .B1_t (new_AGEMA_signal_10578), .B1_f (new_AGEMA_signal_10579), .Z0_t (stateArray_MUX_inS03ser_mux_inst_7_Y), .Z0_f (new_AGEMA_signal_10724), .Z1_t (new_AGEMA_signal_10725), .Z1_f (new_AGEMA_signal_10726) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_7_XOR2_U1 ( .A0_t (stateArray_MUX_inS03ser_mux_inst_7_Y), .A0_f (new_AGEMA_signal_10724), .A1_t (new_AGEMA_signal_10725), .A1_f (new_AGEMA_signal_10726), .B0_t (plaintext_s0_t[31]), .B0_f (plaintext_s0_f[31]), .B1_t (plaintext_s1_t[31]), .B1_f (plaintext_s1_f[31]), .Z0_t (stateArray_inS03ser[7]), .Z0_f (new_AGEMA_signal_10850), .Z1_t (new_AGEMA_signal_10851), .Z1_f (new_AGEMA_signal_10852) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS10ser_mux_inst_0_XOR1_U1 ( .A0_t (plaintext_s0_t[112]), .A0_f (plaintext_s0_f[112]), .A1_t (plaintext_s1_t[112]), .A1_f (plaintext_s1_f[112]), .B0_t (ciphertext_s0_t[80]), .B0_f (ciphertext_s0_f[80]), .B1_t (ciphertext_s1_t[80]), .B1_f (ciphertext_s1_f[80]), .Z0_t (stateArray_MUX_inS10ser_mux_inst_0_X), .Z0_f (new_AGEMA_signal_3744), .Z1_t (new_AGEMA_signal_3745), .Z1_f (new_AGEMA_signal_3746) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS10ser_mux_inst_0_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS10ser_mux_inst_0_X), .B0_f (new_AGEMA_signal_3744), .B1_t (new_AGEMA_signal_3745), .B1_f (new_AGEMA_signal_3746), .Z0_t (stateArray_MUX_inS10ser_mux_inst_0_Y), .Z0_f (new_AGEMA_signal_5896), .Z1_t (new_AGEMA_signal_5897), .Z1_f (new_AGEMA_signal_5898) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS10ser_mux_inst_0_XOR2_U1 ( .A0_t (stateArray_MUX_inS10ser_mux_inst_0_Y), .A0_f (new_AGEMA_signal_5896), .A1_t (new_AGEMA_signal_5897), .A1_f (new_AGEMA_signal_5898), .B0_t (plaintext_s0_t[112]), .B0_f (plaintext_s0_f[112]), .B1_t (plaintext_s1_t[112]), .B1_f (plaintext_s1_f[112]), .Z0_t (stateArray_inS10ser[0]), .Z0_f (new_AGEMA_signal_6694), .Z1_t (new_AGEMA_signal_6695), .Z1_f (new_AGEMA_signal_6696) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS10ser_mux_inst_1_XOR1_U1 ( .A0_t (plaintext_s0_t[113]), .A0_f (plaintext_s0_f[113]), .A1_t (plaintext_s1_t[113]), .A1_f (plaintext_s1_f[113]), .B0_t (ciphertext_s0_t[81]), .B0_f (ciphertext_s0_f[81]), .B1_t (ciphertext_s1_t[81]), .B1_f (ciphertext_s1_f[81]), .Z0_t (stateArray_MUX_inS10ser_mux_inst_1_X), .Z0_f (new_AGEMA_signal_3753), .Z1_t (new_AGEMA_signal_3754), .Z1_f (new_AGEMA_signal_3755) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS10ser_mux_inst_1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS10ser_mux_inst_1_X), .B0_f (new_AGEMA_signal_3753), .B1_t (new_AGEMA_signal_3754), .B1_f (new_AGEMA_signal_3755), .Z0_t (stateArray_MUX_inS10ser_mux_inst_1_Y), .Z0_f (new_AGEMA_signal_5899), .Z1_t (new_AGEMA_signal_5900), .Z1_f (new_AGEMA_signal_5901) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS10ser_mux_inst_1_XOR2_U1 ( .A0_t (stateArray_MUX_inS10ser_mux_inst_1_Y), .A0_f (new_AGEMA_signal_5899), .A1_t (new_AGEMA_signal_5900), .A1_f (new_AGEMA_signal_5901), .B0_t (plaintext_s0_t[113]), .B0_f (plaintext_s0_f[113]), .B1_t (plaintext_s1_t[113]), .B1_f (plaintext_s1_f[113]), .Z0_t (stateArray_inS10ser[1]), .Z0_f (new_AGEMA_signal_6697), .Z1_t (new_AGEMA_signal_6698), .Z1_f (new_AGEMA_signal_6699) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS10ser_mux_inst_2_XOR1_U1 ( .A0_t (plaintext_s0_t[114]), .A0_f (plaintext_s0_f[114]), .A1_t (plaintext_s1_t[114]), .A1_f (plaintext_s1_f[114]), .B0_t (ciphertext_s0_t[82]), .B0_f (ciphertext_s0_f[82]), .B1_t (ciphertext_s1_t[82]), .B1_f (ciphertext_s1_f[82]), .Z0_t (stateArray_MUX_inS10ser_mux_inst_2_X), .Z0_f (new_AGEMA_signal_3762), .Z1_t (new_AGEMA_signal_3763), .Z1_f (new_AGEMA_signal_3764) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS10ser_mux_inst_2_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS10ser_mux_inst_2_X), .B0_f (new_AGEMA_signal_3762), .B1_t (new_AGEMA_signal_3763), .B1_f (new_AGEMA_signal_3764), .Z0_t (stateArray_MUX_inS10ser_mux_inst_2_Y), .Z0_f (new_AGEMA_signal_5902), .Z1_t (new_AGEMA_signal_5903), .Z1_f (new_AGEMA_signal_5904) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS10ser_mux_inst_2_XOR2_U1 ( .A0_t (stateArray_MUX_inS10ser_mux_inst_2_Y), .A0_f (new_AGEMA_signal_5902), .A1_t (new_AGEMA_signal_5903), .A1_f (new_AGEMA_signal_5904), .B0_t (plaintext_s0_t[114]), .B0_f (plaintext_s0_f[114]), .B1_t (plaintext_s1_t[114]), .B1_f (plaintext_s1_f[114]), .Z0_t (stateArray_inS10ser[2]), .Z0_f (new_AGEMA_signal_6700), .Z1_t (new_AGEMA_signal_6701), .Z1_f (new_AGEMA_signal_6702) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS10ser_mux_inst_3_XOR1_U1 ( .A0_t (plaintext_s0_t[115]), .A0_f (plaintext_s0_f[115]), .A1_t (plaintext_s1_t[115]), .A1_f (plaintext_s1_f[115]), .B0_t (ciphertext_s0_t[83]), .B0_f (ciphertext_s0_f[83]), .B1_t (ciphertext_s1_t[83]), .B1_f (ciphertext_s1_f[83]), .Z0_t (stateArray_MUX_inS10ser_mux_inst_3_X), .Z0_f (new_AGEMA_signal_3771), .Z1_t (new_AGEMA_signal_3772), .Z1_f (new_AGEMA_signal_3773) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS10ser_mux_inst_3_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS10ser_mux_inst_3_X), .B0_f (new_AGEMA_signal_3771), .B1_t (new_AGEMA_signal_3772), .B1_f (new_AGEMA_signal_3773), .Z0_t (stateArray_MUX_inS10ser_mux_inst_3_Y), .Z0_f (new_AGEMA_signal_5905), .Z1_t (new_AGEMA_signal_5906), .Z1_f (new_AGEMA_signal_5907) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS10ser_mux_inst_3_XOR2_U1 ( .A0_t (stateArray_MUX_inS10ser_mux_inst_3_Y), .A0_f (new_AGEMA_signal_5905), .A1_t (new_AGEMA_signal_5906), .A1_f (new_AGEMA_signal_5907), .B0_t (plaintext_s0_t[115]), .B0_f (plaintext_s0_f[115]), .B1_t (plaintext_s1_t[115]), .B1_f (plaintext_s1_f[115]), .Z0_t (stateArray_inS10ser[3]), .Z0_f (new_AGEMA_signal_6703), .Z1_t (new_AGEMA_signal_6704), .Z1_f (new_AGEMA_signal_6705) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS10ser_mux_inst_4_XOR1_U1 ( .A0_t (plaintext_s0_t[116]), .A0_f (plaintext_s0_f[116]), .A1_t (plaintext_s1_t[116]), .A1_f (plaintext_s1_f[116]), .B0_t (ciphertext_s0_t[84]), .B0_f (ciphertext_s0_f[84]), .B1_t (ciphertext_s1_t[84]), .B1_f (ciphertext_s1_f[84]), .Z0_t (stateArray_MUX_inS10ser_mux_inst_4_X), .Z0_f (new_AGEMA_signal_3780), .Z1_t (new_AGEMA_signal_3781), .Z1_f (new_AGEMA_signal_3782) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS10ser_mux_inst_4_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS10ser_mux_inst_4_X), .B0_f (new_AGEMA_signal_3780), .B1_t (new_AGEMA_signal_3781), .B1_f (new_AGEMA_signal_3782), .Z0_t (stateArray_MUX_inS10ser_mux_inst_4_Y), .Z0_f (new_AGEMA_signal_5908), .Z1_t (new_AGEMA_signal_5909), .Z1_f (new_AGEMA_signal_5910) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS10ser_mux_inst_4_XOR2_U1 ( .A0_t (stateArray_MUX_inS10ser_mux_inst_4_Y), .A0_f (new_AGEMA_signal_5908), .A1_t (new_AGEMA_signal_5909), .A1_f (new_AGEMA_signal_5910), .B0_t (plaintext_s0_t[116]), .B0_f (plaintext_s0_f[116]), .B1_t (plaintext_s1_t[116]), .B1_f (plaintext_s1_f[116]), .Z0_t (stateArray_inS10ser[4]), .Z0_f (new_AGEMA_signal_6706), .Z1_t (new_AGEMA_signal_6707), .Z1_f (new_AGEMA_signal_6708) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS10ser_mux_inst_5_XOR1_U1 ( .A0_t (plaintext_s0_t[117]), .A0_f (plaintext_s0_f[117]), .A1_t (plaintext_s1_t[117]), .A1_f (plaintext_s1_f[117]), .B0_t (ciphertext_s0_t[85]), .B0_f (ciphertext_s0_f[85]), .B1_t (ciphertext_s1_t[85]), .B1_f (ciphertext_s1_f[85]), .Z0_t (stateArray_MUX_inS10ser_mux_inst_5_X), .Z0_f (new_AGEMA_signal_3789), .Z1_t (new_AGEMA_signal_3790), .Z1_f (new_AGEMA_signal_3791) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS10ser_mux_inst_5_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS10ser_mux_inst_5_X), .B0_f (new_AGEMA_signal_3789), .B1_t (new_AGEMA_signal_3790), .B1_f (new_AGEMA_signal_3791), .Z0_t (stateArray_MUX_inS10ser_mux_inst_5_Y), .Z0_f (new_AGEMA_signal_5911), .Z1_t (new_AGEMA_signal_5912), .Z1_f (new_AGEMA_signal_5913) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS10ser_mux_inst_5_XOR2_U1 ( .A0_t (stateArray_MUX_inS10ser_mux_inst_5_Y), .A0_f (new_AGEMA_signal_5911), .A1_t (new_AGEMA_signal_5912), .A1_f (new_AGEMA_signal_5913), .B0_t (plaintext_s0_t[117]), .B0_f (plaintext_s0_f[117]), .B1_t (plaintext_s1_t[117]), .B1_f (plaintext_s1_f[117]), .Z0_t (stateArray_inS10ser[5]), .Z0_f (new_AGEMA_signal_6709), .Z1_t (new_AGEMA_signal_6710), .Z1_f (new_AGEMA_signal_6711) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS10ser_mux_inst_6_XOR1_U1 ( .A0_t (plaintext_s0_t[118]), .A0_f (plaintext_s0_f[118]), .A1_t (plaintext_s1_t[118]), .A1_f (plaintext_s1_f[118]), .B0_t (ciphertext_s0_t[86]), .B0_f (ciphertext_s0_f[86]), .B1_t (ciphertext_s1_t[86]), .B1_f (ciphertext_s1_f[86]), .Z0_t (stateArray_MUX_inS10ser_mux_inst_6_X), .Z0_f (new_AGEMA_signal_3798), .Z1_t (new_AGEMA_signal_3799), .Z1_f (new_AGEMA_signal_3800) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS10ser_mux_inst_6_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS10ser_mux_inst_6_X), .B0_f (new_AGEMA_signal_3798), .B1_t (new_AGEMA_signal_3799), .B1_f (new_AGEMA_signal_3800), .Z0_t (stateArray_MUX_inS10ser_mux_inst_6_Y), .Z0_f (new_AGEMA_signal_5914), .Z1_t (new_AGEMA_signal_5915), .Z1_f (new_AGEMA_signal_5916) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS10ser_mux_inst_6_XOR2_U1 ( .A0_t (stateArray_MUX_inS10ser_mux_inst_6_Y), .A0_f (new_AGEMA_signal_5914), .A1_t (new_AGEMA_signal_5915), .A1_f (new_AGEMA_signal_5916), .B0_t (plaintext_s0_t[118]), .B0_f (plaintext_s0_f[118]), .B1_t (plaintext_s1_t[118]), .B1_f (plaintext_s1_f[118]), .Z0_t (stateArray_inS10ser[6]), .Z0_f (new_AGEMA_signal_6712), .Z1_t (new_AGEMA_signal_6713), .Z1_f (new_AGEMA_signal_6714) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS10ser_mux_inst_7_XOR1_U1 ( .A0_t (plaintext_s0_t[119]), .A0_f (plaintext_s0_f[119]), .A1_t (plaintext_s1_t[119]), .A1_f (plaintext_s1_f[119]), .B0_t (ciphertext_s0_t[87]), .B0_f (ciphertext_s0_f[87]), .B1_t (ciphertext_s1_t[87]), .B1_f (ciphertext_s1_f[87]), .Z0_t (stateArray_MUX_inS10ser_mux_inst_7_X), .Z0_f (new_AGEMA_signal_3807), .Z1_t (new_AGEMA_signal_3808), .Z1_f (new_AGEMA_signal_3809) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS10ser_mux_inst_7_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS10ser_mux_inst_7_X), .B0_f (new_AGEMA_signal_3807), .B1_t (new_AGEMA_signal_3808), .B1_f (new_AGEMA_signal_3809), .Z0_t (stateArray_MUX_inS10ser_mux_inst_7_Y), .Z0_f (new_AGEMA_signal_5917), .Z1_t (new_AGEMA_signal_5918), .Z1_f (new_AGEMA_signal_5919) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS10ser_mux_inst_7_XOR2_U1 ( .A0_t (stateArray_MUX_inS10ser_mux_inst_7_Y), .A0_f (new_AGEMA_signal_5917), .A1_t (new_AGEMA_signal_5918), .A1_f (new_AGEMA_signal_5919), .B0_t (plaintext_s0_t[119]), .B0_f (plaintext_s0_f[119]), .B1_t (plaintext_s1_t[119]), .B1_f (plaintext_s1_f[119]), .Z0_t (stateArray_inS10ser[7]), .Z0_f (new_AGEMA_signal_6715), .Z1_t (new_AGEMA_signal_6716), .Z1_f (new_AGEMA_signal_6717) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS11ser_mux_inst_0_XOR1_U1 ( .A0_t (plaintext_s0_t[80]), .A0_f (plaintext_s0_f[80]), .A1_t (plaintext_s1_t[80]), .A1_f (plaintext_s1_f[80]), .B0_t (ciphertext_s0_t[48]), .B0_f (ciphertext_s0_f[48]), .B1_t (ciphertext_s1_t[48]), .B1_f (ciphertext_s1_f[48]), .Z0_t (stateArray_MUX_inS11ser_mux_inst_0_X), .Z0_f (new_AGEMA_signal_3816), .Z1_t (new_AGEMA_signal_3817), .Z1_f (new_AGEMA_signal_3818) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS11ser_mux_inst_0_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS11ser_mux_inst_0_X), .B0_f (new_AGEMA_signal_3816), .B1_t (new_AGEMA_signal_3817), .B1_f (new_AGEMA_signal_3818), .Z0_t (stateArray_MUX_inS11ser_mux_inst_0_Y), .Z0_f (new_AGEMA_signal_5920), .Z1_t (new_AGEMA_signal_5921), .Z1_f (new_AGEMA_signal_5922) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS11ser_mux_inst_0_XOR2_U1 ( .A0_t (stateArray_MUX_inS11ser_mux_inst_0_Y), .A0_f (new_AGEMA_signal_5920), .A1_t (new_AGEMA_signal_5921), .A1_f (new_AGEMA_signal_5922), .B0_t (plaintext_s0_t[80]), .B0_f (plaintext_s0_f[80]), .B1_t (plaintext_s1_t[80]), .B1_f (plaintext_s1_f[80]), .Z0_t (stateArray_inS11ser[0]), .Z0_f (new_AGEMA_signal_6718), .Z1_t (new_AGEMA_signal_6719), .Z1_f (new_AGEMA_signal_6720) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS11ser_mux_inst_1_XOR1_U1 ( .A0_t (plaintext_s0_t[81]), .A0_f (plaintext_s0_f[81]), .A1_t (plaintext_s1_t[81]), .A1_f (plaintext_s1_f[81]), .B0_t (ciphertext_s0_t[49]), .B0_f (ciphertext_s0_f[49]), .B1_t (ciphertext_s1_t[49]), .B1_f (ciphertext_s1_f[49]), .Z0_t (stateArray_MUX_inS11ser_mux_inst_1_X), .Z0_f (new_AGEMA_signal_3825), .Z1_t (new_AGEMA_signal_3826), .Z1_f (new_AGEMA_signal_3827) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS11ser_mux_inst_1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS11ser_mux_inst_1_X), .B0_f (new_AGEMA_signal_3825), .B1_t (new_AGEMA_signal_3826), .B1_f (new_AGEMA_signal_3827), .Z0_t (stateArray_MUX_inS11ser_mux_inst_1_Y), .Z0_f (new_AGEMA_signal_5923), .Z1_t (new_AGEMA_signal_5924), .Z1_f (new_AGEMA_signal_5925) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS11ser_mux_inst_1_XOR2_U1 ( .A0_t (stateArray_MUX_inS11ser_mux_inst_1_Y), .A0_f (new_AGEMA_signal_5923), .A1_t (new_AGEMA_signal_5924), .A1_f (new_AGEMA_signal_5925), .B0_t (plaintext_s0_t[81]), .B0_f (plaintext_s0_f[81]), .B1_t (plaintext_s1_t[81]), .B1_f (plaintext_s1_f[81]), .Z0_t (stateArray_inS11ser[1]), .Z0_f (new_AGEMA_signal_6721), .Z1_t (new_AGEMA_signal_6722), .Z1_f (new_AGEMA_signal_6723) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS11ser_mux_inst_2_XOR1_U1 ( .A0_t (plaintext_s0_t[82]), .A0_f (plaintext_s0_f[82]), .A1_t (plaintext_s1_t[82]), .A1_f (plaintext_s1_f[82]), .B0_t (ciphertext_s0_t[50]), .B0_f (ciphertext_s0_f[50]), .B1_t (ciphertext_s1_t[50]), .B1_f (ciphertext_s1_f[50]), .Z0_t (stateArray_MUX_inS11ser_mux_inst_2_X), .Z0_f (new_AGEMA_signal_3834), .Z1_t (new_AGEMA_signal_3835), .Z1_f (new_AGEMA_signal_3836) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS11ser_mux_inst_2_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS11ser_mux_inst_2_X), .B0_f (new_AGEMA_signal_3834), .B1_t (new_AGEMA_signal_3835), .B1_f (new_AGEMA_signal_3836), .Z0_t (stateArray_MUX_inS11ser_mux_inst_2_Y), .Z0_f (new_AGEMA_signal_5926), .Z1_t (new_AGEMA_signal_5927), .Z1_f (new_AGEMA_signal_5928) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS11ser_mux_inst_2_XOR2_U1 ( .A0_t (stateArray_MUX_inS11ser_mux_inst_2_Y), .A0_f (new_AGEMA_signal_5926), .A1_t (new_AGEMA_signal_5927), .A1_f (new_AGEMA_signal_5928), .B0_t (plaintext_s0_t[82]), .B0_f (plaintext_s0_f[82]), .B1_t (plaintext_s1_t[82]), .B1_f (plaintext_s1_f[82]), .Z0_t (stateArray_inS11ser[2]), .Z0_f (new_AGEMA_signal_6724), .Z1_t (new_AGEMA_signal_6725), .Z1_f (new_AGEMA_signal_6726) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS11ser_mux_inst_3_XOR1_U1 ( .A0_t (plaintext_s0_t[83]), .A0_f (plaintext_s0_f[83]), .A1_t (plaintext_s1_t[83]), .A1_f (plaintext_s1_f[83]), .B0_t (ciphertext_s0_t[51]), .B0_f (ciphertext_s0_f[51]), .B1_t (ciphertext_s1_t[51]), .B1_f (ciphertext_s1_f[51]), .Z0_t (stateArray_MUX_inS11ser_mux_inst_3_X), .Z0_f (new_AGEMA_signal_3843), .Z1_t (new_AGEMA_signal_3844), .Z1_f (new_AGEMA_signal_3845) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS11ser_mux_inst_3_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS11ser_mux_inst_3_X), .B0_f (new_AGEMA_signal_3843), .B1_t (new_AGEMA_signal_3844), .B1_f (new_AGEMA_signal_3845), .Z0_t (stateArray_MUX_inS11ser_mux_inst_3_Y), .Z0_f (new_AGEMA_signal_5929), .Z1_t (new_AGEMA_signal_5930), .Z1_f (new_AGEMA_signal_5931) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS11ser_mux_inst_3_XOR2_U1 ( .A0_t (stateArray_MUX_inS11ser_mux_inst_3_Y), .A0_f (new_AGEMA_signal_5929), .A1_t (new_AGEMA_signal_5930), .A1_f (new_AGEMA_signal_5931), .B0_t (plaintext_s0_t[83]), .B0_f (plaintext_s0_f[83]), .B1_t (plaintext_s1_t[83]), .B1_f (plaintext_s1_f[83]), .Z0_t (stateArray_inS11ser[3]), .Z0_f (new_AGEMA_signal_6727), .Z1_t (new_AGEMA_signal_6728), .Z1_f (new_AGEMA_signal_6729) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS11ser_mux_inst_4_XOR1_U1 ( .A0_t (plaintext_s0_t[84]), .A0_f (plaintext_s0_f[84]), .A1_t (plaintext_s1_t[84]), .A1_f (plaintext_s1_f[84]), .B0_t (ciphertext_s0_t[52]), .B0_f (ciphertext_s0_f[52]), .B1_t (ciphertext_s1_t[52]), .B1_f (ciphertext_s1_f[52]), .Z0_t (stateArray_MUX_inS11ser_mux_inst_4_X), .Z0_f (new_AGEMA_signal_3852), .Z1_t (new_AGEMA_signal_3853), .Z1_f (new_AGEMA_signal_3854) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS11ser_mux_inst_4_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS11ser_mux_inst_4_X), .B0_f (new_AGEMA_signal_3852), .B1_t (new_AGEMA_signal_3853), .B1_f (new_AGEMA_signal_3854), .Z0_t (stateArray_MUX_inS11ser_mux_inst_4_Y), .Z0_f (new_AGEMA_signal_5932), .Z1_t (new_AGEMA_signal_5933), .Z1_f (new_AGEMA_signal_5934) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS11ser_mux_inst_4_XOR2_U1 ( .A0_t (stateArray_MUX_inS11ser_mux_inst_4_Y), .A0_f (new_AGEMA_signal_5932), .A1_t (new_AGEMA_signal_5933), .A1_f (new_AGEMA_signal_5934), .B0_t (plaintext_s0_t[84]), .B0_f (plaintext_s0_f[84]), .B1_t (plaintext_s1_t[84]), .B1_f (plaintext_s1_f[84]), .Z0_t (stateArray_inS11ser[4]), .Z0_f (new_AGEMA_signal_6730), .Z1_t (new_AGEMA_signal_6731), .Z1_f (new_AGEMA_signal_6732) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS11ser_mux_inst_5_XOR1_U1 ( .A0_t (plaintext_s0_t[85]), .A0_f (plaintext_s0_f[85]), .A1_t (plaintext_s1_t[85]), .A1_f (plaintext_s1_f[85]), .B0_t (ciphertext_s0_t[53]), .B0_f (ciphertext_s0_f[53]), .B1_t (ciphertext_s1_t[53]), .B1_f (ciphertext_s1_f[53]), .Z0_t (stateArray_MUX_inS11ser_mux_inst_5_X), .Z0_f (new_AGEMA_signal_3861), .Z1_t (new_AGEMA_signal_3862), .Z1_f (new_AGEMA_signal_3863) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS11ser_mux_inst_5_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS11ser_mux_inst_5_X), .B0_f (new_AGEMA_signal_3861), .B1_t (new_AGEMA_signal_3862), .B1_f (new_AGEMA_signal_3863), .Z0_t (stateArray_MUX_inS11ser_mux_inst_5_Y), .Z0_f (new_AGEMA_signal_5935), .Z1_t (new_AGEMA_signal_5936), .Z1_f (new_AGEMA_signal_5937) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS11ser_mux_inst_5_XOR2_U1 ( .A0_t (stateArray_MUX_inS11ser_mux_inst_5_Y), .A0_f (new_AGEMA_signal_5935), .A1_t (new_AGEMA_signal_5936), .A1_f (new_AGEMA_signal_5937), .B0_t (plaintext_s0_t[85]), .B0_f (plaintext_s0_f[85]), .B1_t (plaintext_s1_t[85]), .B1_f (plaintext_s1_f[85]), .Z0_t (stateArray_inS11ser[5]), .Z0_f (new_AGEMA_signal_6733), .Z1_t (new_AGEMA_signal_6734), .Z1_f (new_AGEMA_signal_6735) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS11ser_mux_inst_6_XOR1_U1 ( .A0_t (plaintext_s0_t[86]), .A0_f (plaintext_s0_f[86]), .A1_t (plaintext_s1_t[86]), .A1_f (plaintext_s1_f[86]), .B0_t (ciphertext_s0_t[54]), .B0_f (ciphertext_s0_f[54]), .B1_t (ciphertext_s1_t[54]), .B1_f (ciphertext_s1_f[54]), .Z0_t (stateArray_MUX_inS11ser_mux_inst_6_X), .Z0_f (new_AGEMA_signal_3870), .Z1_t (new_AGEMA_signal_3871), .Z1_f (new_AGEMA_signal_3872) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS11ser_mux_inst_6_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS11ser_mux_inst_6_X), .B0_f (new_AGEMA_signal_3870), .B1_t (new_AGEMA_signal_3871), .B1_f (new_AGEMA_signal_3872), .Z0_t (stateArray_MUX_inS11ser_mux_inst_6_Y), .Z0_f (new_AGEMA_signal_5938), .Z1_t (new_AGEMA_signal_5939), .Z1_f (new_AGEMA_signal_5940) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS11ser_mux_inst_6_XOR2_U1 ( .A0_t (stateArray_MUX_inS11ser_mux_inst_6_Y), .A0_f (new_AGEMA_signal_5938), .A1_t (new_AGEMA_signal_5939), .A1_f (new_AGEMA_signal_5940), .B0_t (plaintext_s0_t[86]), .B0_f (plaintext_s0_f[86]), .B1_t (plaintext_s1_t[86]), .B1_f (plaintext_s1_f[86]), .Z0_t (stateArray_inS11ser[6]), .Z0_f (new_AGEMA_signal_6736), .Z1_t (new_AGEMA_signal_6737), .Z1_f (new_AGEMA_signal_6738) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS11ser_mux_inst_7_XOR1_U1 ( .A0_t (plaintext_s0_t[87]), .A0_f (plaintext_s0_f[87]), .A1_t (plaintext_s1_t[87]), .A1_f (plaintext_s1_f[87]), .B0_t (ciphertext_s0_t[55]), .B0_f (ciphertext_s0_f[55]), .B1_t (ciphertext_s1_t[55]), .B1_f (ciphertext_s1_f[55]), .Z0_t (stateArray_MUX_inS11ser_mux_inst_7_X), .Z0_f (new_AGEMA_signal_3879), .Z1_t (new_AGEMA_signal_3880), .Z1_f (new_AGEMA_signal_3881) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS11ser_mux_inst_7_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS11ser_mux_inst_7_X), .B0_f (new_AGEMA_signal_3879), .B1_t (new_AGEMA_signal_3880), .B1_f (new_AGEMA_signal_3881), .Z0_t (stateArray_MUX_inS11ser_mux_inst_7_Y), .Z0_f (new_AGEMA_signal_5941), .Z1_t (new_AGEMA_signal_5942), .Z1_f (new_AGEMA_signal_5943) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS11ser_mux_inst_7_XOR2_U1 ( .A0_t (stateArray_MUX_inS11ser_mux_inst_7_Y), .A0_f (new_AGEMA_signal_5941), .A1_t (new_AGEMA_signal_5942), .A1_f (new_AGEMA_signal_5943), .B0_t (plaintext_s0_t[87]), .B0_f (plaintext_s0_f[87]), .B1_t (plaintext_s1_t[87]), .B1_f (plaintext_s1_f[87]), .Z0_t (stateArray_inS11ser[7]), .Z0_f (new_AGEMA_signal_6739), .Z1_t (new_AGEMA_signal_6740), .Z1_f (new_AGEMA_signal_6741) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS12ser_mux_inst_0_XOR1_U1 ( .A0_t (plaintext_s0_t[48]), .A0_f (plaintext_s0_f[48]), .A1_t (plaintext_s1_t[48]), .A1_f (plaintext_s1_f[48]), .B0_t (ciphertext_s0_t[16]), .B0_f (ciphertext_s0_f[16]), .B1_t (ciphertext_s1_t[16]), .B1_f (ciphertext_s1_f[16]), .Z0_t (stateArray_MUX_inS12ser_mux_inst_0_X), .Z0_f (new_AGEMA_signal_3888), .Z1_t (new_AGEMA_signal_3889), .Z1_f (new_AGEMA_signal_3890) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS12ser_mux_inst_0_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS12ser_mux_inst_0_X), .B0_f (new_AGEMA_signal_3888), .B1_t (new_AGEMA_signal_3889), .B1_f (new_AGEMA_signal_3890), .Z0_t (stateArray_MUX_inS12ser_mux_inst_0_Y), .Z0_f (new_AGEMA_signal_5944), .Z1_t (new_AGEMA_signal_5945), .Z1_f (new_AGEMA_signal_5946) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS12ser_mux_inst_0_XOR2_U1 ( .A0_t (stateArray_MUX_inS12ser_mux_inst_0_Y), .A0_f (new_AGEMA_signal_5944), .A1_t (new_AGEMA_signal_5945), .A1_f (new_AGEMA_signal_5946), .B0_t (plaintext_s0_t[48]), .B0_f (plaintext_s0_f[48]), .B1_t (plaintext_s1_t[48]), .B1_f (plaintext_s1_f[48]), .Z0_t (stateArray_inS12ser[0]), .Z0_f (new_AGEMA_signal_6742), .Z1_t (new_AGEMA_signal_6743), .Z1_f (new_AGEMA_signal_6744) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS12ser_mux_inst_1_XOR1_U1 ( .A0_t (plaintext_s0_t[49]), .A0_f (plaintext_s0_f[49]), .A1_t (plaintext_s1_t[49]), .A1_f (plaintext_s1_f[49]), .B0_t (ciphertext_s0_t[17]), .B0_f (ciphertext_s0_f[17]), .B1_t (ciphertext_s1_t[17]), .B1_f (ciphertext_s1_f[17]), .Z0_t (stateArray_MUX_inS12ser_mux_inst_1_X), .Z0_f (new_AGEMA_signal_3897), .Z1_t (new_AGEMA_signal_3898), .Z1_f (new_AGEMA_signal_3899) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS12ser_mux_inst_1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS12ser_mux_inst_1_X), .B0_f (new_AGEMA_signal_3897), .B1_t (new_AGEMA_signal_3898), .B1_f (new_AGEMA_signal_3899), .Z0_t (stateArray_MUX_inS12ser_mux_inst_1_Y), .Z0_f (new_AGEMA_signal_5947), .Z1_t (new_AGEMA_signal_5948), .Z1_f (new_AGEMA_signal_5949) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS12ser_mux_inst_1_XOR2_U1 ( .A0_t (stateArray_MUX_inS12ser_mux_inst_1_Y), .A0_f (new_AGEMA_signal_5947), .A1_t (new_AGEMA_signal_5948), .A1_f (new_AGEMA_signal_5949), .B0_t (plaintext_s0_t[49]), .B0_f (plaintext_s0_f[49]), .B1_t (plaintext_s1_t[49]), .B1_f (plaintext_s1_f[49]), .Z0_t (stateArray_inS12ser[1]), .Z0_f (new_AGEMA_signal_6745), .Z1_t (new_AGEMA_signal_6746), .Z1_f (new_AGEMA_signal_6747) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS12ser_mux_inst_2_XOR1_U1 ( .A0_t (plaintext_s0_t[50]), .A0_f (plaintext_s0_f[50]), .A1_t (plaintext_s1_t[50]), .A1_f (plaintext_s1_f[50]), .B0_t (ciphertext_s0_t[18]), .B0_f (ciphertext_s0_f[18]), .B1_t (ciphertext_s1_t[18]), .B1_f (ciphertext_s1_f[18]), .Z0_t (stateArray_MUX_inS12ser_mux_inst_2_X), .Z0_f (new_AGEMA_signal_3906), .Z1_t (new_AGEMA_signal_3907), .Z1_f (new_AGEMA_signal_3908) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS12ser_mux_inst_2_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS12ser_mux_inst_2_X), .B0_f (new_AGEMA_signal_3906), .B1_t (new_AGEMA_signal_3907), .B1_f (new_AGEMA_signal_3908), .Z0_t (stateArray_MUX_inS12ser_mux_inst_2_Y), .Z0_f (new_AGEMA_signal_5950), .Z1_t (new_AGEMA_signal_5951), .Z1_f (new_AGEMA_signal_5952) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS12ser_mux_inst_2_XOR2_U1 ( .A0_t (stateArray_MUX_inS12ser_mux_inst_2_Y), .A0_f (new_AGEMA_signal_5950), .A1_t (new_AGEMA_signal_5951), .A1_f (new_AGEMA_signal_5952), .B0_t (plaintext_s0_t[50]), .B0_f (plaintext_s0_f[50]), .B1_t (plaintext_s1_t[50]), .B1_f (plaintext_s1_f[50]), .Z0_t (stateArray_inS12ser[2]), .Z0_f (new_AGEMA_signal_6748), .Z1_t (new_AGEMA_signal_6749), .Z1_f (new_AGEMA_signal_6750) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS12ser_mux_inst_3_XOR1_U1 ( .A0_t (plaintext_s0_t[51]), .A0_f (plaintext_s0_f[51]), .A1_t (plaintext_s1_t[51]), .A1_f (plaintext_s1_f[51]), .B0_t (ciphertext_s0_t[19]), .B0_f (ciphertext_s0_f[19]), .B1_t (ciphertext_s1_t[19]), .B1_f (ciphertext_s1_f[19]), .Z0_t (stateArray_MUX_inS12ser_mux_inst_3_X), .Z0_f (new_AGEMA_signal_3915), .Z1_t (new_AGEMA_signal_3916), .Z1_f (new_AGEMA_signal_3917) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS12ser_mux_inst_3_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS12ser_mux_inst_3_X), .B0_f (new_AGEMA_signal_3915), .B1_t (new_AGEMA_signal_3916), .B1_f (new_AGEMA_signal_3917), .Z0_t (stateArray_MUX_inS12ser_mux_inst_3_Y), .Z0_f (new_AGEMA_signal_5953), .Z1_t (new_AGEMA_signal_5954), .Z1_f (new_AGEMA_signal_5955) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS12ser_mux_inst_3_XOR2_U1 ( .A0_t (stateArray_MUX_inS12ser_mux_inst_3_Y), .A0_f (new_AGEMA_signal_5953), .A1_t (new_AGEMA_signal_5954), .A1_f (new_AGEMA_signal_5955), .B0_t (plaintext_s0_t[51]), .B0_f (plaintext_s0_f[51]), .B1_t (plaintext_s1_t[51]), .B1_f (plaintext_s1_f[51]), .Z0_t (stateArray_inS12ser[3]), .Z0_f (new_AGEMA_signal_6751), .Z1_t (new_AGEMA_signal_6752), .Z1_f (new_AGEMA_signal_6753) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS12ser_mux_inst_4_XOR1_U1 ( .A0_t (plaintext_s0_t[52]), .A0_f (plaintext_s0_f[52]), .A1_t (plaintext_s1_t[52]), .A1_f (plaintext_s1_f[52]), .B0_t (ciphertext_s0_t[20]), .B0_f (ciphertext_s0_f[20]), .B1_t (ciphertext_s1_t[20]), .B1_f (ciphertext_s1_f[20]), .Z0_t (stateArray_MUX_inS12ser_mux_inst_4_X), .Z0_f (new_AGEMA_signal_3924), .Z1_t (new_AGEMA_signal_3925), .Z1_f (new_AGEMA_signal_3926) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS12ser_mux_inst_4_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS12ser_mux_inst_4_X), .B0_f (new_AGEMA_signal_3924), .B1_t (new_AGEMA_signal_3925), .B1_f (new_AGEMA_signal_3926), .Z0_t (stateArray_MUX_inS12ser_mux_inst_4_Y), .Z0_f (new_AGEMA_signal_5956), .Z1_t (new_AGEMA_signal_5957), .Z1_f (new_AGEMA_signal_5958) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS12ser_mux_inst_4_XOR2_U1 ( .A0_t (stateArray_MUX_inS12ser_mux_inst_4_Y), .A0_f (new_AGEMA_signal_5956), .A1_t (new_AGEMA_signal_5957), .A1_f (new_AGEMA_signal_5958), .B0_t (plaintext_s0_t[52]), .B0_f (plaintext_s0_f[52]), .B1_t (plaintext_s1_t[52]), .B1_f (plaintext_s1_f[52]), .Z0_t (stateArray_inS12ser[4]), .Z0_f (new_AGEMA_signal_6754), .Z1_t (new_AGEMA_signal_6755), .Z1_f (new_AGEMA_signal_6756) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS12ser_mux_inst_5_XOR1_U1 ( .A0_t (plaintext_s0_t[53]), .A0_f (plaintext_s0_f[53]), .A1_t (plaintext_s1_t[53]), .A1_f (plaintext_s1_f[53]), .B0_t (ciphertext_s0_t[21]), .B0_f (ciphertext_s0_f[21]), .B1_t (ciphertext_s1_t[21]), .B1_f (ciphertext_s1_f[21]), .Z0_t (stateArray_MUX_inS12ser_mux_inst_5_X), .Z0_f (new_AGEMA_signal_3933), .Z1_t (new_AGEMA_signal_3934), .Z1_f (new_AGEMA_signal_3935) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS12ser_mux_inst_5_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS12ser_mux_inst_5_X), .B0_f (new_AGEMA_signal_3933), .B1_t (new_AGEMA_signal_3934), .B1_f (new_AGEMA_signal_3935), .Z0_t (stateArray_MUX_inS12ser_mux_inst_5_Y), .Z0_f (new_AGEMA_signal_5959), .Z1_t (new_AGEMA_signal_5960), .Z1_f (new_AGEMA_signal_5961) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS12ser_mux_inst_5_XOR2_U1 ( .A0_t (stateArray_MUX_inS12ser_mux_inst_5_Y), .A0_f (new_AGEMA_signal_5959), .A1_t (new_AGEMA_signal_5960), .A1_f (new_AGEMA_signal_5961), .B0_t (plaintext_s0_t[53]), .B0_f (plaintext_s0_f[53]), .B1_t (plaintext_s1_t[53]), .B1_f (plaintext_s1_f[53]), .Z0_t (stateArray_inS12ser[5]), .Z0_f (new_AGEMA_signal_6757), .Z1_t (new_AGEMA_signal_6758), .Z1_f (new_AGEMA_signal_6759) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS12ser_mux_inst_6_XOR1_U1 ( .A0_t (plaintext_s0_t[54]), .A0_f (plaintext_s0_f[54]), .A1_t (plaintext_s1_t[54]), .A1_f (plaintext_s1_f[54]), .B0_t (ciphertext_s0_t[22]), .B0_f (ciphertext_s0_f[22]), .B1_t (ciphertext_s1_t[22]), .B1_f (ciphertext_s1_f[22]), .Z0_t (stateArray_MUX_inS12ser_mux_inst_6_X), .Z0_f (new_AGEMA_signal_3942), .Z1_t (new_AGEMA_signal_3943), .Z1_f (new_AGEMA_signal_3944) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS12ser_mux_inst_6_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS12ser_mux_inst_6_X), .B0_f (new_AGEMA_signal_3942), .B1_t (new_AGEMA_signal_3943), .B1_f (new_AGEMA_signal_3944), .Z0_t (stateArray_MUX_inS12ser_mux_inst_6_Y), .Z0_f (new_AGEMA_signal_5962), .Z1_t (new_AGEMA_signal_5963), .Z1_f (new_AGEMA_signal_5964) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS12ser_mux_inst_6_XOR2_U1 ( .A0_t (stateArray_MUX_inS12ser_mux_inst_6_Y), .A0_f (new_AGEMA_signal_5962), .A1_t (new_AGEMA_signal_5963), .A1_f (new_AGEMA_signal_5964), .B0_t (plaintext_s0_t[54]), .B0_f (plaintext_s0_f[54]), .B1_t (plaintext_s1_t[54]), .B1_f (plaintext_s1_f[54]), .Z0_t (stateArray_inS12ser[6]), .Z0_f (new_AGEMA_signal_6760), .Z1_t (new_AGEMA_signal_6761), .Z1_f (new_AGEMA_signal_6762) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS12ser_mux_inst_7_XOR1_U1 ( .A0_t (plaintext_s0_t[55]), .A0_f (plaintext_s0_f[55]), .A1_t (plaintext_s1_t[55]), .A1_f (plaintext_s1_f[55]), .B0_t (ciphertext_s0_t[23]), .B0_f (ciphertext_s0_f[23]), .B1_t (ciphertext_s1_t[23]), .B1_f (ciphertext_s1_f[23]), .Z0_t (stateArray_MUX_inS12ser_mux_inst_7_X), .Z0_f (new_AGEMA_signal_3951), .Z1_t (new_AGEMA_signal_3952), .Z1_f (new_AGEMA_signal_3953) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS12ser_mux_inst_7_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS12ser_mux_inst_7_X), .B0_f (new_AGEMA_signal_3951), .B1_t (new_AGEMA_signal_3952), .B1_f (new_AGEMA_signal_3953), .Z0_t (stateArray_MUX_inS12ser_mux_inst_7_Y), .Z0_f (new_AGEMA_signal_5965), .Z1_t (new_AGEMA_signal_5966), .Z1_f (new_AGEMA_signal_5967) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS12ser_mux_inst_7_XOR2_U1 ( .A0_t (stateArray_MUX_inS12ser_mux_inst_7_Y), .A0_f (new_AGEMA_signal_5965), .A1_t (new_AGEMA_signal_5966), .A1_f (new_AGEMA_signal_5967), .B0_t (plaintext_s0_t[55]), .B0_f (plaintext_s0_f[55]), .B1_t (plaintext_s1_t[55]), .B1_f (plaintext_s1_f[55]), .Z0_t (stateArray_inS12ser[7]), .Z0_f (new_AGEMA_signal_6763), .Z1_t (new_AGEMA_signal_6764), .Z1_f (new_AGEMA_signal_6765) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS20_MC_mux_inst_0_XOR1_U1 ( .A0_t (ciphertext_s0_t[104]), .A0_f (ciphertext_s0_f[104]), .A1_t (ciphertext_s1_t[104]), .A1_f (ciphertext_s1_f[104]), .B0_t (StateInMC[16]), .B0_f (new_AGEMA_signal_9352), .B1_t (new_AGEMA_signal_9353), .B1_f (new_AGEMA_signal_9354), .Z0_t (stateArray_MUX_outS20_MC_mux_inst_0_X), .Z0_f (new_AGEMA_signal_9810), .Z1_t (new_AGEMA_signal_9811), .Z1_f (new_AGEMA_signal_9812) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS20_MC_mux_inst_0_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (stateArray_MUX_outS20_MC_mux_inst_0_X), .B0_f (new_AGEMA_signal_9810), .B1_t (new_AGEMA_signal_9811), .B1_f (new_AGEMA_signal_9812), .Z0_t (stateArray_MUX_outS20_MC_mux_inst_0_Y), .Z0_f (new_AGEMA_signal_10331), .Z1_t (new_AGEMA_signal_10332), .Z1_f (new_AGEMA_signal_10333) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS20_MC_mux_inst_0_XOR2_U1 ( .A0_t (stateArray_MUX_outS20_MC_mux_inst_0_Y), .A0_f (new_AGEMA_signal_10331), .A1_t (new_AGEMA_signal_10332), .A1_f (new_AGEMA_signal_10333), .B0_t (ciphertext_s0_t[104]), .B0_f (ciphertext_s0_f[104]), .B1_t (ciphertext_s1_t[104]), .B1_f (ciphertext_s1_f[104]), .Z0_t (stateArray_outS20ser_MC[0]), .Z0_f (new_AGEMA_signal_10454), .Z1_t (new_AGEMA_signal_10455), .Z1_f (new_AGEMA_signal_10456) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS20_MC_mux_inst_1_XOR1_U1 ( .A0_t (ciphertext_s0_t[105]), .A0_f (ciphertext_s0_f[105]), .A1_t (ciphertext_s1_t[105]), .A1_f (ciphertext_s1_f[105]), .B0_t (StateInMC[17]), .B0_f (new_AGEMA_signal_9858), .B1_t (new_AGEMA_signal_9859), .B1_f (new_AGEMA_signal_9860), .Z0_t (stateArray_MUX_outS20_MC_mux_inst_1_X), .Z0_f (new_AGEMA_signal_10334), .Z1_t (new_AGEMA_signal_10335), .Z1_f (new_AGEMA_signal_10336) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS20_MC_mux_inst_1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (stateArray_MUX_outS20_MC_mux_inst_1_X), .B0_f (new_AGEMA_signal_10334), .B1_t (new_AGEMA_signal_10335), .B1_f (new_AGEMA_signal_10336), .Z0_t (stateArray_MUX_outS20_MC_mux_inst_1_Y), .Z0_f (new_AGEMA_signal_10457), .Z1_t (new_AGEMA_signal_10458), .Z1_f (new_AGEMA_signal_10459) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS20_MC_mux_inst_1_XOR2_U1 ( .A0_t (stateArray_MUX_outS20_MC_mux_inst_1_Y), .A0_f (new_AGEMA_signal_10457), .A1_t (new_AGEMA_signal_10458), .A1_f (new_AGEMA_signal_10459), .B0_t (ciphertext_s0_t[105]), .B0_f (ciphertext_s0_f[105]), .B1_t (ciphertext_s1_t[105]), .B1_f (ciphertext_s1_f[105]), .Z0_t (stateArray_outS20ser_MC[1]), .Z0_f (new_AGEMA_signal_10580), .Z1_t (new_AGEMA_signal_10581), .Z1_f (new_AGEMA_signal_10582) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS20_MC_mux_inst_2_XOR1_U1 ( .A0_t (ciphertext_s0_t[106]), .A0_f (ciphertext_s0_f[106]), .A1_t (ciphertext_s1_t[106]), .A1_f (ciphertext_s1_f[106]), .B0_t (StateInMC[18]), .B0_f (new_AGEMA_signal_9358), .B1_t (new_AGEMA_signal_9359), .B1_f (new_AGEMA_signal_9360), .Z0_t (stateArray_MUX_outS20_MC_mux_inst_2_X), .Z0_f (new_AGEMA_signal_9813), .Z1_t (new_AGEMA_signal_9814), .Z1_f (new_AGEMA_signal_9815) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS20_MC_mux_inst_2_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (stateArray_MUX_outS20_MC_mux_inst_2_X), .B0_f (new_AGEMA_signal_9813), .B1_t (new_AGEMA_signal_9814), .B1_f (new_AGEMA_signal_9815), .Z0_t (stateArray_MUX_outS20_MC_mux_inst_2_Y), .Z0_f (new_AGEMA_signal_10337), .Z1_t (new_AGEMA_signal_10338), .Z1_f (new_AGEMA_signal_10339) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS20_MC_mux_inst_2_XOR2_U1 ( .A0_t (stateArray_MUX_outS20_MC_mux_inst_2_Y), .A0_f (new_AGEMA_signal_10337), .A1_t (new_AGEMA_signal_10338), .A1_f (new_AGEMA_signal_10339), .B0_t (ciphertext_s0_t[106]), .B0_f (ciphertext_s0_f[106]), .B1_t (ciphertext_s1_t[106]), .B1_f (ciphertext_s1_f[106]), .Z0_t (stateArray_outS20ser_MC[2]), .Z0_f (new_AGEMA_signal_10460), .Z1_t (new_AGEMA_signal_10461), .Z1_f (new_AGEMA_signal_10462) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS20_MC_mux_inst_3_XOR1_U1 ( .A0_t (ciphertext_s0_t[107]), .A0_f (ciphertext_s0_f[107]), .A1_t (ciphertext_s1_t[107]), .A1_f (ciphertext_s1_f[107]), .B0_t (StateInMC[19]), .B0_f (new_AGEMA_signal_9861), .B1_t (new_AGEMA_signal_9862), .B1_f (new_AGEMA_signal_9863), .Z0_t (stateArray_MUX_outS20_MC_mux_inst_3_X), .Z0_f (new_AGEMA_signal_10340), .Z1_t (new_AGEMA_signal_10341), .Z1_f (new_AGEMA_signal_10342) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS20_MC_mux_inst_3_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (stateArray_MUX_outS20_MC_mux_inst_3_X), .B0_f (new_AGEMA_signal_10340), .B1_t (new_AGEMA_signal_10341), .B1_f (new_AGEMA_signal_10342), .Z0_t (stateArray_MUX_outS20_MC_mux_inst_3_Y), .Z0_f (new_AGEMA_signal_10463), .Z1_t (new_AGEMA_signal_10464), .Z1_f (new_AGEMA_signal_10465) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS20_MC_mux_inst_3_XOR2_U1 ( .A0_t (stateArray_MUX_outS20_MC_mux_inst_3_Y), .A0_f (new_AGEMA_signal_10463), .A1_t (new_AGEMA_signal_10464), .A1_f (new_AGEMA_signal_10465), .B0_t (ciphertext_s0_t[107]), .B0_f (ciphertext_s0_f[107]), .B1_t (ciphertext_s1_t[107]), .B1_f (ciphertext_s1_f[107]), .Z0_t (stateArray_outS20ser_MC[3]), .Z0_f (new_AGEMA_signal_10583), .Z1_t (new_AGEMA_signal_10584), .Z1_f (new_AGEMA_signal_10585) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS20_MC_mux_inst_4_XOR1_U1 ( .A0_t (ciphertext_s0_t[108]), .A0_f (ciphertext_s0_f[108]), .A1_t (ciphertext_s1_t[108]), .A1_f (ciphertext_s1_f[108]), .B0_t (StateInMC[20]), .B0_f (new_AGEMA_signal_9864), .B1_t (new_AGEMA_signal_9865), .B1_f (new_AGEMA_signal_9866), .Z0_t (stateArray_MUX_outS20_MC_mux_inst_4_X), .Z0_f (new_AGEMA_signal_10343), .Z1_t (new_AGEMA_signal_10344), .Z1_f (new_AGEMA_signal_10345) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS20_MC_mux_inst_4_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (stateArray_MUX_outS20_MC_mux_inst_4_X), .B0_f (new_AGEMA_signal_10343), .B1_t (new_AGEMA_signal_10344), .B1_f (new_AGEMA_signal_10345), .Z0_t (stateArray_MUX_outS20_MC_mux_inst_4_Y), .Z0_f (new_AGEMA_signal_10466), .Z1_t (new_AGEMA_signal_10467), .Z1_f (new_AGEMA_signal_10468) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS20_MC_mux_inst_4_XOR2_U1 ( .A0_t (stateArray_MUX_outS20_MC_mux_inst_4_Y), .A0_f (new_AGEMA_signal_10466), .A1_t (new_AGEMA_signal_10467), .A1_f (new_AGEMA_signal_10468), .B0_t (ciphertext_s0_t[108]), .B0_f (ciphertext_s0_f[108]), .B1_t (ciphertext_s1_t[108]), .B1_f (ciphertext_s1_f[108]), .Z0_t (stateArray_outS20ser_MC[4]), .Z0_f (new_AGEMA_signal_10586), .Z1_t (new_AGEMA_signal_10587), .Z1_f (new_AGEMA_signal_10588) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS20_MC_mux_inst_5_XOR1_U1 ( .A0_t (ciphertext_s0_t[109]), .A0_f (ciphertext_s0_f[109]), .A1_t (ciphertext_s1_t[109]), .A1_f (ciphertext_s1_f[109]), .B0_t (StateInMC[21]), .B0_f (new_AGEMA_signal_9367), .B1_t (new_AGEMA_signal_9368), .B1_f (new_AGEMA_signal_9369), .Z0_t (stateArray_MUX_outS20_MC_mux_inst_5_X), .Z0_f (new_AGEMA_signal_9816), .Z1_t (new_AGEMA_signal_9817), .Z1_f (new_AGEMA_signal_9818) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS20_MC_mux_inst_5_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (stateArray_MUX_outS20_MC_mux_inst_5_X), .B0_f (new_AGEMA_signal_9816), .B1_t (new_AGEMA_signal_9817), .B1_f (new_AGEMA_signal_9818), .Z0_t (stateArray_MUX_outS20_MC_mux_inst_5_Y), .Z0_f (new_AGEMA_signal_10346), .Z1_t (new_AGEMA_signal_10347), .Z1_f (new_AGEMA_signal_10348) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS20_MC_mux_inst_5_XOR2_U1 ( .A0_t (stateArray_MUX_outS20_MC_mux_inst_5_Y), .A0_f (new_AGEMA_signal_10346), .A1_t (new_AGEMA_signal_10347), .A1_f (new_AGEMA_signal_10348), .B0_t (ciphertext_s0_t[109]), .B0_f (ciphertext_s0_f[109]), .B1_t (ciphertext_s1_t[109]), .B1_f (ciphertext_s1_f[109]), .Z0_t (stateArray_outS20ser_MC[5]), .Z0_f (new_AGEMA_signal_10469), .Z1_t (new_AGEMA_signal_10470), .Z1_f (new_AGEMA_signal_10471) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS20_MC_mux_inst_6_XOR1_U1 ( .A0_t (ciphertext_s0_t[110]), .A0_f (ciphertext_s0_f[110]), .A1_t (ciphertext_s1_t[110]), .A1_f (ciphertext_s1_f[110]), .B0_t (StateInMC[22]), .B0_f (new_AGEMA_signal_9370), .B1_t (new_AGEMA_signal_9371), .B1_f (new_AGEMA_signal_9372), .Z0_t (stateArray_MUX_outS20_MC_mux_inst_6_X), .Z0_f (new_AGEMA_signal_9819), .Z1_t (new_AGEMA_signal_9820), .Z1_f (new_AGEMA_signal_9821) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS20_MC_mux_inst_6_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (stateArray_MUX_outS20_MC_mux_inst_6_X), .B0_f (new_AGEMA_signal_9819), .B1_t (new_AGEMA_signal_9820), .B1_f (new_AGEMA_signal_9821), .Z0_t (stateArray_MUX_outS20_MC_mux_inst_6_Y), .Z0_f (new_AGEMA_signal_10349), .Z1_t (new_AGEMA_signal_10350), .Z1_f (new_AGEMA_signal_10351) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS20_MC_mux_inst_6_XOR2_U1 ( .A0_t (stateArray_MUX_outS20_MC_mux_inst_6_Y), .A0_f (new_AGEMA_signal_10349), .A1_t (new_AGEMA_signal_10350), .A1_f (new_AGEMA_signal_10351), .B0_t (ciphertext_s0_t[110]), .B0_f (ciphertext_s0_f[110]), .B1_t (ciphertext_s1_t[110]), .B1_f (ciphertext_s1_f[110]), .Z0_t (stateArray_outS20ser_MC[6]), .Z0_f (new_AGEMA_signal_10472), .Z1_t (new_AGEMA_signal_10473), .Z1_f (new_AGEMA_signal_10474) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS20_MC_mux_inst_7_XOR1_U1 ( .A0_t (ciphertext_s0_t[111]), .A0_f (ciphertext_s0_f[111]), .A1_t (ciphertext_s1_t[111]), .A1_f (ciphertext_s1_f[111]), .B0_t (StateInMC[23]), .B0_f (new_AGEMA_signal_9373), .B1_t (new_AGEMA_signal_9374), .B1_f (new_AGEMA_signal_9375), .Z0_t (stateArray_MUX_outS20_MC_mux_inst_7_X), .Z0_f (new_AGEMA_signal_9822), .Z1_t (new_AGEMA_signal_9823), .Z1_f (new_AGEMA_signal_9824) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS20_MC_mux_inst_7_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (stateArray_MUX_outS20_MC_mux_inst_7_X), .B0_f (new_AGEMA_signal_9822), .B1_t (new_AGEMA_signal_9823), .B1_f (new_AGEMA_signal_9824), .Z0_t (stateArray_MUX_outS20_MC_mux_inst_7_Y), .Z0_f (new_AGEMA_signal_10352), .Z1_t (new_AGEMA_signal_10353), .Z1_f (new_AGEMA_signal_10354) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS20_MC_mux_inst_7_XOR2_U1 ( .A0_t (stateArray_MUX_outS20_MC_mux_inst_7_Y), .A0_f (new_AGEMA_signal_10352), .A1_t (new_AGEMA_signal_10353), .A1_f (new_AGEMA_signal_10354), .B0_t (ciphertext_s0_t[111]), .B0_f (ciphertext_s0_f[111]), .B1_t (ciphertext_s1_t[111]), .B1_f (ciphertext_s1_f[111]), .Z0_t (stateArray_outS20ser_MC[7]), .Z0_f (new_AGEMA_signal_10475), .Z1_t (new_AGEMA_signal_10476), .Z1_f (new_AGEMA_signal_10477) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_0_XOR1_U1 ( .A0_t (plaintext_s0_t[16]), .A0_f (plaintext_s0_f[16]), .A1_t (plaintext_s1_t[16]), .A1_f (plaintext_s1_f[16]), .B0_t (stateArray_outS20ser_MC[0]), .B0_f (new_AGEMA_signal_10454), .B1_t (new_AGEMA_signal_10455), .B1_f (new_AGEMA_signal_10456), .Z0_t (stateArray_MUX_inS13ser_mux_inst_0_X), .Z0_f (new_AGEMA_signal_10592), .Z1_t (new_AGEMA_signal_10593), .Z1_f (new_AGEMA_signal_10594) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_0_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS13ser_mux_inst_0_X), .B0_f (new_AGEMA_signal_10592), .B1_t (new_AGEMA_signal_10593), .B1_f (new_AGEMA_signal_10594), .Z0_t (stateArray_MUX_inS13ser_mux_inst_0_Y), .Z0_f (new_AGEMA_signal_10727), .Z1_t (new_AGEMA_signal_10728), .Z1_f (new_AGEMA_signal_10729) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_0_XOR2_U1 ( .A0_t (stateArray_MUX_inS13ser_mux_inst_0_Y), .A0_f (new_AGEMA_signal_10727), .A1_t (new_AGEMA_signal_10728), .A1_f (new_AGEMA_signal_10729), .B0_t (plaintext_s0_t[16]), .B0_f (plaintext_s0_f[16]), .B1_t (plaintext_s1_t[16]), .B1_f (plaintext_s1_f[16]), .Z0_t (stateArray_inS13ser[0]), .Z0_f (new_AGEMA_signal_10853), .Z1_t (new_AGEMA_signal_10854), .Z1_f (new_AGEMA_signal_10855) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_1_XOR1_U1 ( .A0_t (plaintext_s0_t[17]), .A0_f (plaintext_s0_f[17]), .A1_t (plaintext_s1_t[17]), .A1_f (plaintext_s1_f[17]), .B0_t (stateArray_outS20ser_MC[1]), .B0_f (new_AGEMA_signal_10580), .B1_t (new_AGEMA_signal_10581), .B1_f (new_AGEMA_signal_10582), .Z0_t (stateArray_MUX_inS13ser_mux_inst_1_X), .Z0_f (new_AGEMA_signal_10733), .Z1_t (new_AGEMA_signal_10734), .Z1_f (new_AGEMA_signal_10735) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS13ser_mux_inst_1_X), .B0_f (new_AGEMA_signal_10733), .B1_t (new_AGEMA_signal_10734), .B1_f (new_AGEMA_signal_10735), .Z0_t (stateArray_MUX_inS13ser_mux_inst_1_Y), .Z0_f (new_AGEMA_signal_10856), .Z1_t (new_AGEMA_signal_10857), .Z1_f (new_AGEMA_signal_10858) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_1_XOR2_U1 ( .A0_t (stateArray_MUX_inS13ser_mux_inst_1_Y), .A0_f (new_AGEMA_signal_10856), .A1_t (new_AGEMA_signal_10857), .A1_f (new_AGEMA_signal_10858), .B0_t (plaintext_s0_t[17]), .B0_f (plaintext_s0_f[17]), .B1_t (plaintext_s1_t[17]), .B1_f (plaintext_s1_f[17]), .Z0_t (stateArray_inS13ser[1]), .Z0_f (new_AGEMA_signal_10994), .Z1_t (new_AGEMA_signal_10995), .Z1_f (new_AGEMA_signal_10996) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_2_XOR1_U1 ( .A0_t (plaintext_s0_t[18]), .A0_f (plaintext_s0_f[18]), .A1_t (plaintext_s1_t[18]), .A1_f (plaintext_s1_f[18]), .B0_t (stateArray_outS20ser_MC[2]), .B0_f (new_AGEMA_signal_10460), .B1_t (new_AGEMA_signal_10461), .B1_f (new_AGEMA_signal_10462), .Z0_t (stateArray_MUX_inS13ser_mux_inst_2_X), .Z0_f (new_AGEMA_signal_10598), .Z1_t (new_AGEMA_signal_10599), .Z1_f (new_AGEMA_signal_10600) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_2_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS13ser_mux_inst_2_X), .B0_f (new_AGEMA_signal_10598), .B1_t (new_AGEMA_signal_10599), .B1_f (new_AGEMA_signal_10600), .Z0_t (stateArray_MUX_inS13ser_mux_inst_2_Y), .Z0_f (new_AGEMA_signal_10736), .Z1_t (new_AGEMA_signal_10737), .Z1_f (new_AGEMA_signal_10738) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_2_XOR2_U1 ( .A0_t (stateArray_MUX_inS13ser_mux_inst_2_Y), .A0_f (new_AGEMA_signal_10736), .A1_t (new_AGEMA_signal_10737), .A1_f (new_AGEMA_signal_10738), .B0_t (plaintext_s0_t[18]), .B0_f (plaintext_s0_f[18]), .B1_t (plaintext_s1_t[18]), .B1_f (plaintext_s1_f[18]), .Z0_t (stateArray_inS13ser[2]), .Z0_f (new_AGEMA_signal_10859), .Z1_t (new_AGEMA_signal_10860), .Z1_f (new_AGEMA_signal_10861) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_3_XOR1_U1 ( .A0_t (plaintext_s0_t[19]), .A0_f (plaintext_s0_f[19]), .A1_t (plaintext_s1_t[19]), .A1_f (plaintext_s1_f[19]), .B0_t (stateArray_outS20ser_MC[3]), .B0_f (new_AGEMA_signal_10583), .B1_t (new_AGEMA_signal_10584), .B1_f (new_AGEMA_signal_10585), .Z0_t (stateArray_MUX_inS13ser_mux_inst_3_X), .Z0_f (new_AGEMA_signal_10742), .Z1_t (new_AGEMA_signal_10743), .Z1_f (new_AGEMA_signal_10744) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_3_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS13ser_mux_inst_3_X), .B0_f (new_AGEMA_signal_10742), .B1_t (new_AGEMA_signal_10743), .B1_f (new_AGEMA_signal_10744), .Z0_t (stateArray_MUX_inS13ser_mux_inst_3_Y), .Z0_f (new_AGEMA_signal_10862), .Z1_t (new_AGEMA_signal_10863), .Z1_f (new_AGEMA_signal_10864) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_3_XOR2_U1 ( .A0_t (stateArray_MUX_inS13ser_mux_inst_3_Y), .A0_f (new_AGEMA_signal_10862), .A1_t (new_AGEMA_signal_10863), .A1_f (new_AGEMA_signal_10864), .B0_t (plaintext_s0_t[19]), .B0_f (plaintext_s0_f[19]), .B1_t (plaintext_s1_t[19]), .B1_f (plaintext_s1_f[19]), .Z0_t (stateArray_inS13ser[3]), .Z0_f (new_AGEMA_signal_10997), .Z1_t (new_AGEMA_signal_10998), .Z1_f (new_AGEMA_signal_10999) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_4_XOR1_U1 ( .A0_t (plaintext_s0_t[20]), .A0_f (plaintext_s0_f[20]), .A1_t (plaintext_s1_t[20]), .A1_f (plaintext_s1_f[20]), .B0_t (stateArray_outS20ser_MC[4]), .B0_f (new_AGEMA_signal_10586), .B1_t (new_AGEMA_signal_10587), .B1_f (new_AGEMA_signal_10588), .Z0_t (stateArray_MUX_inS13ser_mux_inst_4_X), .Z0_f (new_AGEMA_signal_10748), .Z1_t (new_AGEMA_signal_10749), .Z1_f (new_AGEMA_signal_10750) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_4_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS13ser_mux_inst_4_X), .B0_f (new_AGEMA_signal_10748), .B1_t (new_AGEMA_signal_10749), .B1_f (new_AGEMA_signal_10750), .Z0_t (stateArray_MUX_inS13ser_mux_inst_4_Y), .Z0_f (new_AGEMA_signal_10865), .Z1_t (new_AGEMA_signal_10866), .Z1_f (new_AGEMA_signal_10867) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_4_XOR2_U1 ( .A0_t (stateArray_MUX_inS13ser_mux_inst_4_Y), .A0_f (new_AGEMA_signal_10865), .A1_t (new_AGEMA_signal_10866), .A1_f (new_AGEMA_signal_10867), .B0_t (plaintext_s0_t[20]), .B0_f (plaintext_s0_f[20]), .B1_t (plaintext_s1_t[20]), .B1_f (plaintext_s1_f[20]), .Z0_t (stateArray_inS13ser[4]), .Z0_f (new_AGEMA_signal_11000), .Z1_t (new_AGEMA_signal_11001), .Z1_f (new_AGEMA_signal_11002) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_5_XOR1_U1 ( .A0_t (plaintext_s0_t[21]), .A0_f (plaintext_s0_f[21]), .A1_t (plaintext_s1_t[21]), .A1_f (plaintext_s1_f[21]), .B0_t (stateArray_outS20ser_MC[5]), .B0_f (new_AGEMA_signal_10469), .B1_t (new_AGEMA_signal_10470), .B1_f (new_AGEMA_signal_10471), .Z0_t (stateArray_MUX_inS13ser_mux_inst_5_X), .Z0_f (new_AGEMA_signal_10604), .Z1_t (new_AGEMA_signal_10605), .Z1_f (new_AGEMA_signal_10606) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_5_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS13ser_mux_inst_5_X), .B0_f (new_AGEMA_signal_10604), .B1_t (new_AGEMA_signal_10605), .B1_f (new_AGEMA_signal_10606), .Z0_t (stateArray_MUX_inS13ser_mux_inst_5_Y), .Z0_f (new_AGEMA_signal_10751), .Z1_t (new_AGEMA_signal_10752), .Z1_f (new_AGEMA_signal_10753) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_5_XOR2_U1 ( .A0_t (stateArray_MUX_inS13ser_mux_inst_5_Y), .A0_f (new_AGEMA_signal_10751), .A1_t (new_AGEMA_signal_10752), .A1_f (new_AGEMA_signal_10753), .B0_t (plaintext_s0_t[21]), .B0_f (plaintext_s0_f[21]), .B1_t (plaintext_s1_t[21]), .B1_f (plaintext_s1_f[21]), .Z0_t (stateArray_inS13ser[5]), .Z0_f (new_AGEMA_signal_10868), .Z1_t (new_AGEMA_signal_10869), .Z1_f (new_AGEMA_signal_10870) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_6_XOR1_U1 ( .A0_t (plaintext_s0_t[22]), .A0_f (plaintext_s0_f[22]), .A1_t (plaintext_s1_t[22]), .A1_f (plaintext_s1_f[22]), .B0_t (stateArray_outS20ser_MC[6]), .B0_f (new_AGEMA_signal_10472), .B1_t (new_AGEMA_signal_10473), .B1_f (new_AGEMA_signal_10474), .Z0_t (stateArray_MUX_inS13ser_mux_inst_6_X), .Z0_f (new_AGEMA_signal_10610), .Z1_t (new_AGEMA_signal_10611), .Z1_f (new_AGEMA_signal_10612) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_6_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS13ser_mux_inst_6_X), .B0_f (new_AGEMA_signal_10610), .B1_t (new_AGEMA_signal_10611), .B1_f (new_AGEMA_signal_10612), .Z0_t (stateArray_MUX_inS13ser_mux_inst_6_Y), .Z0_f (new_AGEMA_signal_10754), .Z1_t (new_AGEMA_signal_10755), .Z1_f (new_AGEMA_signal_10756) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_6_XOR2_U1 ( .A0_t (stateArray_MUX_inS13ser_mux_inst_6_Y), .A0_f (new_AGEMA_signal_10754), .A1_t (new_AGEMA_signal_10755), .A1_f (new_AGEMA_signal_10756), .B0_t (plaintext_s0_t[22]), .B0_f (plaintext_s0_f[22]), .B1_t (plaintext_s1_t[22]), .B1_f (plaintext_s1_f[22]), .Z0_t (stateArray_inS13ser[6]), .Z0_f (new_AGEMA_signal_10871), .Z1_t (new_AGEMA_signal_10872), .Z1_f (new_AGEMA_signal_10873) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_7_XOR1_U1 ( .A0_t (plaintext_s0_t[23]), .A0_f (plaintext_s0_f[23]), .A1_t (plaintext_s1_t[23]), .A1_f (plaintext_s1_f[23]), .B0_t (stateArray_outS20ser_MC[7]), .B0_f (new_AGEMA_signal_10475), .B1_t (new_AGEMA_signal_10476), .B1_f (new_AGEMA_signal_10477), .Z0_t (stateArray_MUX_inS13ser_mux_inst_7_X), .Z0_f (new_AGEMA_signal_10616), .Z1_t (new_AGEMA_signal_10617), .Z1_f (new_AGEMA_signal_10618) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_7_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS13ser_mux_inst_7_X), .B0_f (new_AGEMA_signal_10616), .B1_t (new_AGEMA_signal_10617), .B1_f (new_AGEMA_signal_10618), .Z0_t (stateArray_MUX_inS13ser_mux_inst_7_Y), .Z0_f (new_AGEMA_signal_10757), .Z1_t (new_AGEMA_signal_10758), .Z1_f (new_AGEMA_signal_10759) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_7_XOR2_U1 ( .A0_t (stateArray_MUX_inS13ser_mux_inst_7_Y), .A0_f (new_AGEMA_signal_10757), .A1_t (new_AGEMA_signal_10758), .A1_f (new_AGEMA_signal_10759), .B0_t (plaintext_s0_t[23]), .B0_f (plaintext_s0_f[23]), .B1_t (plaintext_s1_t[23]), .B1_f (plaintext_s1_f[23]), .Z0_t (stateArray_inS13ser[7]), .Z0_f (new_AGEMA_signal_10874), .Z1_t (new_AGEMA_signal_10875), .Z1_f (new_AGEMA_signal_10876) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS20ser_mux_inst_0_XOR1_U1 ( .A0_t (plaintext_s0_t[104]), .A0_f (plaintext_s0_f[104]), .A1_t (plaintext_s1_t[104]), .A1_f (plaintext_s1_f[104]), .B0_t (ciphertext_s0_t[72]), .B0_f (ciphertext_s0_f[72]), .B1_t (ciphertext_s1_t[72]), .B1_f (ciphertext_s1_f[72]), .Z0_t (stateArray_MUX_inS20ser_mux_inst_0_X), .Z0_f (new_AGEMA_signal_3960), .Z1_t (new_AGEMA_signal_3961), .Z1_f (new_AGEMA_signal_3962) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS20ser_mux_inst_0_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS20ser_mux_inst_0_X), .B0_f (new_AGEMA_signal_3960), .B1_t (new_AGEMA_signal_3961), .B1_f (new_AGEMA_signal_3962), .Z0_t (stateArray_MUX_inS20ser_mux_inst_0_Y), .Z0_f (new_AGEMA_signal_5968), .Z1_t (new_AGEMA_signal_5969), .Z1_f (new_AGEMA_signal_5970) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS20ser_mux_inst_0_XOR2_U1 ( .A0_t (stateArray_MUX_inS20ser_mux_inst_0_Y), .A0_f (new_AGEMA_signal_5968), .A1_t (new_AGEMA_signal_5969), .A1_f (new_AGEMA_signal_5970), .B0_t (plaintext_s0_t[104]), .B0_f (plaintext_s0_f[104]), .B1_t (plaintext_s1_t[104]), .B1_f (plaintext_s1_f[104]), .Z0_t (stateArray_inS20ser[0]), .Z0_f (new_AGEMA_signal_6766), .Z1_t (new_AGEMA_signal_6767), .Z1_f (new_AGEMA_signal_6768) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS20ser_mux_inst_1_XOR1_U1 ( .A0_t (plaintext_s0_t[105]), .A0_f (plaintext_s0_f[105]), .A1_t (plaintext_s1_t[105]), .A1_f (plaintext_s1_f[105]), .B0_t (ciphertext_s0_t[73]), .B0_f (ciphertext_s0_f[73]), .B1_t (ciphertext_s1_t[73]), .B1_f (ciphertext_s1_f[73]), .Z0_t (stateArray_MUX_inS20ser_mux_inst_1_X), .Z0_f (new_AGEMA_signal_3969), .Z1_t (new_AGEMA_signal_3970), .Z1_f (new_AGEMA_signal_3971) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS20ser_mux_inst_1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS20ser_mux_inst_1_X), .B0_f (new_AGEMA_signal_3969), .B1_t (new_AGEMA_signal_3970), .B1_f (new_AGEMA_signal_3971), .Z0_t (stateArray_MUX_inS20ser_mux_inst_1_Y), .Z0_f (new_AGEMA_signal_5971), .Z1_t (new_AGEMA_signal_5972), .Z1_f (new_AGEMA_signal_5973) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS20ser_mux_inst_1_XOR2_U1 ( .A0_t (stateArray_MUX_inS20ser_mux_inst_1_Y), .A0_f (new_AGEMA_signal_5971), .A1_t (new_AGEMA_signal_5972), .A1_f (new_AGEMA_signal_5973), .B0_t (plaintext_s0_t[105]), .B0_f (plaintext_s0_f[105]), .B1_t (plaintext_s1_t[105]), .B1_f (plaintext_s1_f[105]), .Z0_t (stateArray_inS20ser[1]), .Z0_f (new_AGEMA_signal_6769), .Z1_t (new_AGEMA_signal_6770), .Z1_f (new_AGEMA_signal_6771) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS20ser_mux_inst_2_XOR1_U1 ( .A0_t (plaintext_s0_t[106]), .A0_f (plaintext_s0_f[106]), .A1_t (plaintext_s1_t[106]), .A1_f (plaintext_s1_f[106]), .B0_t (ciphertext_s0_t[74]), .B0_f (ciphertext_s0_f[74]), .B1_t (ciphertext_s1_t[74]), .B1_f (ciphertext_s1_f[74]), .Z0_t (stateArray_MUX_inS20ser_mux_inst_2_X), .Z0_f (new_AGEMA_signal_3978), .Z1_t (new_AGEMA_signal_3979), .Z1_f (new_AGEMA_signal_3980) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS20ser_mux_inst_2_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS20ser_mux_inst_2_X), .B0_f (new_AGEMA_signal_3978), .B1_t (new_AGEMA_signal_3979), .B1_f (new_AGEMA_signal_3980), .Z0_t (stateArray_MUX_inS20ser_mux_inst_2_Y), .Z0_f (new_AGEMA_signal_5974), .Z1_t (new_AGEMA_signal_5975), .Z1_f (new_AGEMA_signal_5976) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS20ser_mux_inst_2_XOR2_U1 ( .A0_t (stateArray_MUX_inS20ser_mux_inst_2_Y), .A0_f (new_AGEMA_signal_5974), .A1_t (new_AGEMA_signal_5975), .A1_f (new_AGEMA_signal_5976), .B0_t (plaintext_s0_t[106]), .B0_f (plaintext_s0_f[106]), .B1_t (plaintext_s1_t[106]), .B1_f (plaintext_s1_f[106]), .Z0_t (stateArray_inS20ser[2]), .Z0_f (new_AGEMA_signal_6772), .Z1_t (new_AGEMA_signal_6773), .Z1_f (new_AGEMA_signal_6774) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS20ser_mux_inst_3_XOR1_U1 ( .A0_t (plaintext_s0_t[107]), .A0_f (plaintext_s0_f[107]), .A1_t (plaintext_s1_t[107]), .A1_f (plaintext_s1_f[107]), .B0_t (ciphertext_s0_t[75]), .B0_f (ciphertext_s0_f[75]), .B1_t (ciphertext_s1_t[75]), .B1_f (ciphertext_s1_f[75]), .Z0_t (stateArray_MUX_inS20ser_mux_inst_3_X), .Z0_f (new_AGEMA_signal_3987), .Z1_t (new_AGEMA_signal_3988), .Z1_f (new_AGEMA_signal_3989) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS20ser_mux_inst_3_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS20ser_mux_inst_3_X), .B0_f (new_AGEMA_signal_3987), .B1_t (new_AGEMA_signal_3988), .B1_f (new_AGEMA_signal_3989), .Z0_t (stateArray_MUX_inS20ser_mux_inst_3_Y), .Z0_f (new_AGEMA_signal_5977), .Z1_t (new_AGEMA_signal_5978), .Z1_f (new_AGEMA_signal_5979) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS20ser_mux_inst_3_XOR2_U1 ( .A0_t (stateArray_MUX_inS20ser_mux_inst_3_Y), .A0_f (new_AGEMA_signal_5977), .A1_t (new_AGEMA_signal_5978), .A1_f (new_AGEMA_signal_5979), .B0_t (plaintext_s0_t[107]), .B0_f (plaintext_s0_f[107]), .B1_t (plaintext_s1_t[107]), .B1_f (plaintext_s1_f[107]), .Z0_t (stateArray_inS20ser[3]), .Z0_f (new_AGEMA_signal_6775), .Z1_t (new_AGEMA_signal_6776), .Z1_f (new_AGEMA_signal_6777) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS20ser_mux_inst_4_XOR1_U1 ( .A0_t (plaintext_s0_t[108]), .A0_f (plaintext_s0_f[108]), .A1_t (plaintext_s1_t[108]), .A1_f (plaintext_s1_f[108]), .B0_t (ciphertext_s0_t[76]), .B0_f (ciphertext_s0_f[76]), .B1_t (ciphertext_s1_t[76]), .B1_f (ciphertext_s1_f[76]), .Z0_t (stateArray_MUX_inS20ser_mux_inst_4_X), .Z0_f (new_AGEMA_signal_3996), .Z1_t (new_AGEMA_signal_3997), .Z1_f (new_AGEMA_signal_3998) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS20ser_mux_inst_4_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS20ser_mux_inst_4_X), .B0_f (new_AGEMA_signal_3996), .B1_t (new_AGEMA_signal_3997), .B1_f (new_AGEMA_signal_3998), .Z0_t (stateArray_MUX_inS20ser_mux_inst_4_Y), .Z0_f (new_AGEMA_signal_5980), .Z1_t (new_AGEMA_signal_5981), .Z1_f (new_AGEMA_signal_5982) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS20ser_mux_inst_4_XOR2_U1 ( .A0_t (stateArray_MUX_inS20ser_mux_inst_4_Y), .A0_f (new_AGEMA_signal_5980), .A1_t (new_AGEMA_signal_5981), .A1_f (new_AGEMA_signal_5982), .B0_t (plaintext_s0_t[108]), .B0_f (plaintext_s0_f[108]), .B1_t (plaintext_s1_t[108]), .B1_f (plaintext_s1_f[108]), .Z0_t (stateArray_inS20ser[4]), .Z0_f (new_AGEMA_signal_6778), .Z1_t (new_AGEMA_signal_6779), .Z1_f (new_AGEMA_signal_6780) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS20ser_mux_inst_5_XOR1_U1 ( .A0_t (plaintext_s0_t[109]), .A0_f (plaintext_s0_f[109]), .A1_t (plaintext_s1_t[109]), .A1_f (plaintext_s1_f[109]), .B0_t (ciphertext_s0_t[77]), .B0_f (ciphertext_s0_f[77]), .B1_t (ciphertext_s1_t[77]), .B1_f (ciphertext_s1_f[77]), .Z0_t (stateArray_MUX_inS20ser_mux_inst_5_X), .Z0_f (new_AGEMA_signal_4005), .Z1_t (new_AGEMA_signal_4006), .Z1_f (new_AGEMA_signal_4007) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS20ser_mux_inst_5_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS20ser_mux_inst_5_X), .B0_f (new_AGEMA_signal_4005), .B1_t (new_AGEMA_signal_4006), .B1_f (new_AGEMA_signal_4007), .Z0_t (stateArray_MUX_inS20ser_mux_inst_5_Y), .Z0_f (new_AGEMA_signal_5983), .Z1_t (new_AGEMA_signal_5984), .Z1_f (new_AGEMA_signal_5985) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS20ser_mux_inst_5_XOR2_U1 ( .A0_t (stateArray_MUX_inS20ser_mux_inst_5_Y), .A0_f (new_AGEMA_signal_5983), .A1_t (new_AGEMA_signal_5984), .A1_f (new_AGEMA_signal_5985), .B0_t (plaintext_s0_t[109]), .B0_f (plaintext_s0_f[109]), .B1_t (plaintext_s1_t[109]), .B1_f (plaintext_s1_f[109]), .Z0_t (stateArray_inS20ser[5]), .Z0_f (new_AGEMA_signal_6781), .Z1_t (new_AGEMA_signal_6782), .Z1_f (new_AGEMA_signal_6783) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS20ser_mux_inst_6_XOR1_U1 ( .A0_t (plaintext_s0_t[110]), .A0_f (plaintext_s0_f[110]), .A1_t (plaintext_s1_t[110]), .A1_f (plaintext_s1_f[110]), .B0_t (ciphertext_s0_t[78]), .B0_f (ciphertext_s0_f[78]), .B1_t (ciphertext_s1_t[78]), .B1_f (ciphertext_s1_f[78]), .Z0_t (stateArray_MUX_inS20ser_mux_inst_6_X), .Z0_f (new_AGEMA_signal_4014), .Z1_t (new_AGEMA_signal_4015), .Z1_f (new_AGEMA_signal_4016) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS20ser_mux_inst_6_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS20ser_mux_inst_6_X), .B0_f (new_AGEMA_signal_4014), .B1_t (new_AGEMA_signal_4015), .B1_f (new_AGEMA_signal_4016), .Z0_t (stateArray_MUX_inS20ser_mux_inst_6_Y), .Z0_f (new_AGEMA_signal_5986), .Z1_t (new_AGEMA_signal_5987), .Z1_f (new_AGEMA_signal_5988) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS20ser_mux_inst_6_XOR2_U1 ( .A0_t (stateArray_MUX_inS20ser_mux_inst_6_Y), .A0_f (new_AGEMA_signal_5986), .A1_t (new_AGEMA_signal_5987), .A1_f (new_AGEMA_signal_5988), .B0_t (plaintext_s0_t[110]), .B0_f (plaintext_s0_f[110]), .B1_t (plaintext_s1_t[110]), .B1_f (plaintext_s1_f[110]), .Z0_t (stateArray_inS20ser[6]), .Z0_f (new_AGEMA_signal_6784), .Z1_t (new_AGEMA_signal_6785), .Z1_f (new_AGEMA_signal_6786) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS20ser_mux_inst_7_XOR1_U1 ( .A0_t (plaintext_s0_t[111]), .A0_f (plaintext_s0_f[111]), .A1_t (plaintext_s1_t[111]), .A1_f (plaintext_s1_f[111]), .B0_t (ciphertext_s0_t[79]), .B0_f (ciphertext_s0_f[79]), .B1_t (ciphertext_s1_t[79]), .B1_f (ciphertext_s1_f[79]), .Z0_t (stateArray_MUX_inS20ser_mux_inst_7_X), .Z0_f (new_AGEMA_signal_4023), .Z1_t (new_AGEMA_signal_4024), .Z1_f (new_AGEMA_signal_4025) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS20ser_mux_inst_7_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS20ser_mux_inst_7_X), .B0_f (new_AGEMA_signal_4023), .B1_t (new_AGEMA_signal_4024), .B1_f (new_AGEMA_signal_4025), .Z0_t (stateArray_MUX_inS20ser_mux_inst_7_Y), .Z0_f (new_AGEMA_signal_5989), .Z1_t (new_AGEMA_signal_5990), .Z1_f (new_AGEMA_signal_5991) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS20ser_mux_inst_7_XOR2_U1 ( .A0_t (stateArray_MUX_inS20ser_mux_inst_7_Y), .A0_f (new_AGEMA_signal_5989), .A1_t (new_AGEMA_signal_5990), .A1_f (new_AGEMA_signal_5991), .B0_t (plaintext_s0_t[111]), .B0_f (plaintext_s0_f[111]), .B1_t (plaintext_s1_t[111]), .B1_f (plaintext_s1_f[111]), .Z0_t (stateArray_inS20ser[7]), .Z0_f (new_AGEMA_signal_6787), .Z1_t (new_AGEMA_signal_6788), .Z1_f (new_AGEMA_signal_6789) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS21ser_mux_inst_0_XOR1_U1 ( .A0_t (plaintext_s0_t[72]), .A0_f (plaintext_s0_f[72]), .A1_t (plaintext_s1_t[72]), .A1_f (plaintext_s1_f[72]), .B0_t (ciphertext_s0_t[40]), .B0_f (ciphertext_s0_f[40]), .B1_t (ciphertext_s1_t[40]), .B1_f (ciphertext_s1_f[40]), .Z0_t (stateArray_MUX_inS21ser_mux_inst_0_X), .Z0_f (new_AGEMA_signal_4032), .Z1_t (new_AGEMA_signal_4033), .Z1_f (new_AGEMA_signal_4034) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS21ser_mux_inst_0_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS21ser_mux_inst_0_X), .B0_f (new_AGEMA_signal_4032), .B1_t (new_AGEMA_signal_4033), .B1_f (new_AGEMA_signal_4034), .Z0_t (stateArray_MUX_inS21ser_mux_inst_0_Y), .Z0_f (new_AGEMA_signal_5992), .Z1_t (new_AGEMA_signal_5993), .Z1_f (new_AGEMA_signal_5994) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS21ser_mux_inst_0_XOR2_U1 ( .A0_t (stateArray_MUX_inS21ser_mux_inst_0_Y), .A0_f (new_AGEMA_signal_5992), .A1_t (new_AGEMA_signal_5993), .A1_f (new_AGEMA_signal_5994), .B0_t (plaintext_s0_t[72]), .B0_f (plaintext_s0_f[72]), .B1_t (plaintext_s1_t[72]), .B1_f (plaintext_s1_f[72]), .Z0_t (stateArray_inS21ser[0]), .Z0_f (new_AGEMA_signal_6790), .Z1_t (new_AGEMA_signal_6791), .Z1_f (new_AGEMA_signal_6792) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS21ser_mux_inst_1_XOR1_U1 ( .A0_t (plaintext_s0_t[73]), .A0_f (plaintext_s0_f[73]), .A1_t (plaintext_s1_t[73]), .A1_f (plaintext_s1_f[73]), .B0_t (ciphertext_s0_t[41]), .B0_f (ciphertext_s0_f[41]), .B1_t (ciphertext_s1_t[41]), .B1_f (ciphertext_s1_f[41]), .Z0_t (stateArray_MUX_inS21ser_mux_inst_1_X), .Z0_f (new_AGEMA_signal_4041), .Z1_t (new_AGEMA_signal_4042), .Z1_f (new_AGEMA_signal_4043) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS21ser_mux_inst_1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS21ser_mux_inst_1_X), .B0_f (new_AGEMA_signal_4041), .B1_t (new_AGEMA_signal_4042), .B1_f (new_AGEMA_signal_4043), .Z0_t (stateArray_MUX_inS21ser_mux_inst_1_Y), .Z0_f (new_AGEMA_signal_5995), .Z1_t (new_AGEMA_signal_5996), .Z1_f (new_AGEMA_signal_5997) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS21ser_mux_inst_1_XOR2_U1 ( .A0_t (stateArray_MUX_inS21ser_mux_inst_1_Y), .A0_f (new_AGEMA_signal_5995), .A1_t (new_AGEMA_signal_5996), .A1_f (new_AGEMA_signal_5997), .B0_t (plaintext_s0_t[73]), .B0_f (plaintext_s0_f[73]), .B1_t (plaintext_s1_t[73]), .B1_f (plaintext_s1_f[73]), .Z0_t (stateArray_inS21ser[1]), .Z0_f (new_AGEMA_signal_6793), .Z1_t (new_AGEMA_signal_6794), .Z1_f (new_AGEMA_signal_6795) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS21ser_mux_inst_2_XOR1_U1 ( .A0_t (plaintext_s0_t[74]), .A0_f (plaintext_s0_f[74]), .A1_t (plaintext_s1_t[74]), .A1_f (plaintext_s1_f[74]), .B0_t (ciphertext_s0_t[42]), .B0_f (ciphertext_s0_f[42]), .B1_t (ciphertext_s1_t[42]), .B1_f (ciphertext_s1_f[42]), .Z0_t (stateArray_MUX_inS21ser_mux_inst_2_X), .Z0_f (new_AGEMA_signal_4050), .Z1_t (new_AGEMA_signal_4051), .Z1_f (new_AGEMA_signal_4052) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS21ser_mux_inst_2_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS21ser_mux_inst_2_X), .B0_f (new_AGEMA_signal_4050), .B1_t (new_AGEMA_signal_4051), .B1_f (new_AGEMA_signal_4052), .Z0_t (stateArray_MUX_inS21ser_mux_inst_2_Y), .Z0_f (new_AGEMA_signal_5998), .Z1_t (new_AGEMA_signal_5999), .Z1_f (new_AGEMA_signal_6000) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS21ser_mux_inst_2_XOR2_U1 ( .A0_t (stateArray_MUX_inS21ser_mux_inst_2_Y), .A0_f (new_AGEMA_signal_5998), .A1_t (new_AGEMA_signal_5999), .A1_f (new_AGEMA_signal_6000), .B0_t (plaintext_s0_t[74]), .B0_f (plaintext_s0_f[74]), .B1_t (plaintext_s1_t[74]), .B1_f (plaintext_s1_f[74]), .Z0_t (stateArray_inS21ser[2]), .Z0_f (new_AGEMA_signal_6796), .Z1_t (new_AGEMA_signal_6797), .Z1_f (new_AGEMA_signal_6798) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS21ser_mux_inst_3_XOR1_U1 ( .A0_t (plaintext_s0_t[75]), .A0_f (plaintext_s0_f[75]), .A1_t (plaintext_s1_t[75]), .A1_f (plaintext_s1_f[75]), .B0_t (ciphertext_s0_t[43]), .B0_f (ciphertext_s0_f[43]), .B1_t (ciphertext_s1_t[43]), .B1_f (ciphertext_s1_f[43]), .Z0_t (stateArray_MUX_inS21ser_mux_inst_3_X), .Z0_f (new_AGEMA_signal_4059), .Z1_t (new_AGEMA_signal_4060), .Z1_f (new_AGEMA_signal_4061) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS21ser_mux_inst_3_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS21ser_mux_inst_3_X), .B0_f (new_AGEMA_signal_4059), .B1_t (new_AGEMA_signal_4060), .B1_f (new_AGEMA_signal_4061), .Z0_t (stateArray_MUX_inS21ser_mux_inst_3_Y), .Z0_f (new_AGEMA_signal_6001), .Z1_t (new_AGEMA_signal_6002), .Z1_f (new_AGEMA_signal_6003) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS21ser_mux_inst_3_XOR2_U1 ( .A0_t (stateArray_MUX_inS21ser_mux_inst_3_Y), .A0_f (new_AGEMA_signal_6001), .A1_t (new_AGEMA_signal_6002), .A1_f (new_AGEMA_signal_6003), .B0_t (plaintext_s0_t[75]), .B0_f (plaintext_s0_f[75]), .B1_t (plaintext_s1_t[75]), .B1_f (plaintext_s1_f[75]), .Z0_t (stateArray_inS21ser[3]), .Z0_f (new_AGEMA_signal_6799), .Z1_t (new_AGEMA_signal_6800), .Z1_f (new_AGEMA_signal_6801) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS21ser_mux_inst_4_XOR1_U1 ( .A0_t (plaintext_s0_t[76]), .A0_f (plaintext_s0_f[76]), .A1_t (plaintext_s1_t[76]), .A1_f (plaintext_s1_f[76]), .B0_t (ciphertext_s0_t[44]), .B0_f (ciphertext_s0_f[44]), .B1_t (ciphertext_s1_t[44]), .B1_f (ciphertext_s1_f[44]), .Z0_t (stateArray_MUX_inS21ser_mux_inst_4_X), .Z0_f (new_AGEMA_signal_4068), .Z1_t (new_AGEMA_signal_4069), .Z1_f (new_AGEMA_signal_4070) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS21ser_mux_inst_4_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS21ser_mux_inst_4_X), .B0_f (new_AGEMA_signal_4068), .B1_t (new_AGEMA_signal_4069), .B1_f (new_AGEMA_signal_4070), .Z0_t (stateArray_MUX_inS21ser_mux_inst_4_Y), .Z0_f (new_AGEMA_signal_6004), .Z1_t (new_AGEMA_signal_6005), .Z1_f (new_AGEMA_signal_6006) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS21ser_mux_inst_4_XOR2_U1 ( .A0_t (stateArray_MUX_inS21ser_mux_inst_4_Y), .A0_f (new_AGEMA_signal_6004), .A1_t (new_AGEMA_signal_6005), .A1_f (new_AGEMA_signal_6006), .B0_t (plaintext_s0_t[76]), .B0_f (plaintext_s0_f[76]), .B1_t (plaintext_s1_t[76]), .B1_f (plaintext_s1_f[76]), .Z0_t (stateArray_inS21ser[4]), .Z0_f (new_AGEMA_signal_6802), .Z1_t (new_AGEMA_signal_6803), .Z1_f (new_AGEMA_signal_6804) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS21ser_mux_inst_5_XOR1_U1 ( .A0_t (plaintext_s0_t[77]), .A0_f (plaintext_s0_f[77]), .A1_t (plaintext_s1_t[77]), .A1_f (plaintext_s1_f[77]), .B0_t (ciphertext_s0_t[45]), .B0_f (ciphertext_s0_f[45]), .B1_t (ciphertext_s1_t[45]), .B1_f (ciphertext_s1_f[45]), .Z0_t (stateArray_MUX_inS21ser_mux_inst_5_X), .Z0_f (new_AGEMA_signal_4077), .Z1_t (new_AGEMA_signal_4078), .Z1_f (new_AGEMA_signal_4079) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS21ser_mux_inst_5_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS21ser_mux_inst_5_X), .B0_f (new_AGEMA_signal_4077), .B1_t (new_AGEMA_signal_4078), .B1_f (new_AGEMA_signal_4079), .Z0_t (stateArray_MUX_inS21ser_mux_inst_5_Y), .Z0_f (new_AGEMA_signal_6007), .Z1_t (new_AGEMA_signal_6008), .Z1_f (new_AGEMA_signal_6009) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS21ser_mux_inst_5_XOR2_U1 ( .A0_t (stateArray_MUX_inS21ser_mux_inst_5_Y), .A0_f (new_AGEMA_signal_6007), .A1_t (new_AGEMA_signal_6008), .A1_f (new_AGEMA_signal_6009), .B0_t (plaintext_s0_t[77]), .B0_f (plaintext_s0_f[77]), .B1_t (plaintext_s1_t[77]), .B1_f (plaintext_s1_f[77]), .Z0_t (stateArray_inS21ser[5]), .Z0_f (new_AGEMA_signal_6805), .Z1_t (new_AGEMA_signal_6806), .Z1_f (new_AGEMA_signal_6807) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS21ser_mux_inst_6_XOR1_U1 ( .A0_t (plaintext_s0_t[78]), .A0_f (plaintext_s0_f[78]), .A1_t (plaintext_s1_t[78]), .A1_f (plaintext_s1_f[78]), .B0_t (ciphertext_s0_t[46]), .B0_f (ciphertext_s0_f[46]), .B1_t (ciphertext_s1_t[46]), .B1_f (ciphertext_s1_f[46]), .Z0_t (stateArray_MUX_inS21ser_mux_inst_6_X), .Z0_f (new_AGEMA_signal_4086), .Z1_t (new_AGEMA_signal_4087), .Z1_f (new_AGEMA_signal_4088) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS21ser_mux_inst_6_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS21ser_mux_inst_6_X), .B0_f (new_AGEMA_signal_4086), .B1_t (new_AGEMA_signal_4087), .B1_f (new_AGEMA_signal_4088), .Z0_t (stateArray_MUX_inS21ser_mux_inst_6_Y), .Z0_f (new_AGEMA_signal_6010), .Z1_t (new_AGEMA_signal_6011), .Z1_f (new_AGEMA_signal_6012) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS21ser_mux_inst_6_XOR2_U1 ( .A0_t (stateArray_MUX_inS21ser_mux_inst_6_Y), .A0_f (new_AGEMA_signal_6010), .A1_t (new_AGEMA_signal_6011), .A1_f (new_AGEMA_signal_6012), .B0_t (plaintext_s0_t[78]), .B0_f (plaintext_s0_f[78]), .B1_t (plaintext_s1_t[78]), .B1_f (plaintext_s1_f[78]), .Z0_t (stateArray_inS21ser[6]), .Z0_f (new_AGEMA_signal_6808), .Z1_t (new_AGEMA_signal_6809), .Z1_f (new_AGEMA_signal_6810) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS21ser_mux_inst_7_XOR1_U1 ( .A0_t (plaintext_s0_t[79]), .A0_f (plaintext_s0_f[79]), .A1_t (plaintext_s1_t[79]), .A1_f (plaintext_s1_f[79]), .B0_t (ciphertext_s0_t[47]), .B0_f (ciphertext_s0_f[47]), .B1_t (ciphertext_s1_t[47]), .B1_f (ciphertext_s1_f[47]), .Z0_t (stateArray_MUX_inS21ser_mux_inst_7_X), .Z0_f (new_AGEMA_signal_4095), .Z1_t (new_AGEMA_signal_4096), .Z1_f (new_AGEMA_signal_4097) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS21ser_mux_inst_7_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS21ser_mux_inst_7_X), .B0_f (new_AGEMA_signal_4095), .B1_t (new_AGEMA_signal_4096), .B1_f (new_AGEMA_signal_4097), .Z0_t (stateArray_MUX_inS21ser_mux_inst_7_Y), .Z0_f (new_AGEMA_signal_6013), .Z1_t (new_AGEMA_signal_6014), .Z1_f (new_AGEMA_signal_6015) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS21ser_mux_inst_7_XOR2_U1 ( .A0_t (stateArray_MUX_inS21ser_mux_inst_7_Y), .A0_f (new_AGEMA_signal_6013), .A1_t (new_AGEMA_signal_6014), .A1_f (new_AGEMA_signal_6015), .B0_t (plaintext_s0_t[79]), .B0_f (plaintext_s0_f[79]), .B1_t (plaintext_s1_t[79]), .B1_f (plaintext_s1_f[79]), .Z0_t (stateArray_inS21ser[7]), .Z0_f (new_AGEMA_signal_6811), .Z1_t (new_AGEMA_signal_6812), .Z1_f (new_AGEMA_signal_6813) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS22ser_mux_inst_0_XOR1_U1 ( .A0_t (plaintext_s0_t[40]), .A0_f (plaintext_s0_f[40]), .A1_t (plaintext_s1_t[40]), .A1_f (plaintext_s1_f[40]), .B0_t (ciphertext_s0_t[8]), .B0_f (ciphertext_s0_f[8]), .B1_t (ciphertext_s1_t[8]), .B1_f (ciphertext_s1_f[8]), .Z0_t (stateArray_MUX_inS22ser_mux_inst_0_X), .Z0_f (new_AGEMA_signal_4104), .Z1_t (new_AGEMA_signal_4105), .Z1_f (new_AGEMA_signal_4106) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS22ser_mux_inst_0_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS22ser_mux_inst_0_X), .B0_f (new_AGEMA_signal_4104), .B1_t (new_AGEMA_signal_4105), .B1_f (new_AGEMA_signal_4106), .Z0_t (stateArray_MUX_inS22ser_mux_inst_0_Y), .Z0_f (new_AGEMA_signal_6016), .Z1_t (new_AGEMA_signal_6017), .Z1_f (new_AGEMA_signal_6018) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS22ser_mux_inst_0_XOR2_U1 ( .A0_t (stateArray_MUX_inS22ser_mux_inst_0_Y), .A0_f (new_AGEMA_signal_6016), .A1_t (new_AGEMA_signal_6017), .A1_f (new_AGEMA_signal_6018), .B0_t (plaintext_s0_t[40]), .B0_f (plaintext_s0_f[40]), .B1_t (plaintext_s1_t[40]), .B1_f (plaintext_s1_f[40]), .Z0_t (stateArray_inS22ser[0]), .Z0_f (new_AGEMA_signal_6814), .Z1_t (new_AGEMA_signal_6815), .Z1_f (new_AGEMA_signal_6816) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS22ser_mux_inst_1_XOR1_U1 ( .A0_t (plaintext_s0_t[41]), .A0_f (plaintext_s0_f[41]), .A1_t (plaintext_s1_t[41]), .A1_f (plaintext_s1_f[41]), .B0_t (ciphertext_s0_t[9]), .B0_f (ciphertext_s0_f[9]), .B1_t (ciphertext_s1_t[9]), .B1_f (ciphertext_s1_f[9]), .Z0_t (stateArray_MUX_inS22ser_mux_inst_1_X), .Z0_f (new_AGEMA_signal_4113), .Z1_t (new_AGEMA_signal_4114), .Z1_f (new_AGEMA_signal_4115) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS22ser_mux_inst_1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS22ser_mux_inst_1_X), .B0_f (new_AGEMA_signal_4113), .B1_t (new_AGEMA_signal_4114), .B1_f (new_AGEMA_signal_4115), .Z0_t (stateArray_MUX_inS22ser_mux_inst_1_Y), .Z0_f (new_AGEMA_signal_6019), .Z1_t (new_AGEMA_signal_6020), .Z1_f (new_AGEMA_signal_6021) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS22ser_mux_inst_1_XOR2_U1 ( .A0_t (stateArray_MUX_inS22ser_mux_inst_1_Y), .A0_f (new_AGEMA_signal_6019), .A1_t (new_AGEMA_signal_6020), .A1_f (new_AGEMA_signal_6021), .B0_t (plaintext_s0_t[41]), .B0_f (plaintext_s0_f[41]), .B1_t (plaintext_s1_t[41]), .B1_f (plaintext_s1_f[41]), .Z0_t (stateArray_inS22ser[1]), .Z0_f (new_AGEMA_signal_6817), .Z1_t (new_AGEMA_signal_6818), .Z1_f (new_AGEMA_signal_6819) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS22ser_mux_inst_2_XOR1_U1 ( .A0_t (plaintext_s0_t[42]), .A0_f (plaintext_s0_f[42]), .A1_t (plaintext_s1_t[42]), .A1_f (plaintext_s1_f[42]), .B0_t (ciphertext_s0_t[10]), .B0_f (ciphertext_s0_f[10]), .B1_t (ciphertext_s1_t[10]), .B1_f (ciphertext_s1_f[10]), .Z0_t (stateArray_MUX_inS22ser_mux_inst_2_X), .Z0_f (new_AGEMA_signal_4122), .Z1_t (new_AGEMA_signal_4123), .Z1_f (new_AGEMA_signal_4124) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS22ser_mux_inst_2_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS22ser_mux_inst_2_X), .B0_f (new_AGEMA_signal_4122), .B1_t (new_AGEMA_signal_4123), .B1_f (new_AGEMA_signal_4124), .Z0_t (stateArray_MUX_inS22ser_mux_inst_2_Y), .Z0_f (new_AGEMA_signal_6022), .Z1_t (new_AGEMA_signal_6023), .Z1_f (new_AGEMA_signal_6024) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS22ser_mux_inst_2_XOR2_U1 ( .A0_t (stateArray_MUX_inS22ser_mux_inst_2_Y), .A0_f (new_AGEMA_signal_6022), .A1_t (new_AGEMA_signal_6023), .A1_f (new_AGEMA_signal_6024), .B0_t (plaintext_s0_t[42]), .B0_f (plaintext_s0_f[42]), .B1_t (plaintext_s1_t[42]), .B1_f (plaintext_s1_f[42]), .Z0_t (stateArray_inS22ser[2]), .Z0_f (new_AGEMA_signal_6820), .Z1_t (new_AGEMA_signal_6821), .Z1_f (new_AGEMA_signal_6822) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS22ser_mux_inst_3_XOR1_U1 ( .A0_t (plaintext_s0_t[43]), .A0_f (plaintext_s0_f[43]), .A1_t (plaintext_s1_t[43]), .A1_f (plaintext_s1_f[43]), .B0_t (ciphertext_s0_t[11]), .B0_f (ciphertext_s0_f[11]), .B1_t (ciphertext_s1_t[11]), .B1_f (ciphertext_s1_f[11]), .Z0_t (stateArray_MUX_inS22ser_mux_inst_3_X), .Z0_f (new_AGEMA_signal_4131), .Z1_t (new_AGEMA_signal_4132), .Z1_f (new_AGEMA_signal_4133) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS22ser_mux_inst_3_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS22ser_mux_inst_3_X), .B0_f (new_AGEMA_signal_4131), .B1_t (new_AGEMA_signal_4132), .B1_f (new_AGEMA_signal_4133), .Z0_t (stateArray_MUX_inS22ser_mux_inst_3_Y), .Z0_f (new_AGEMA_signal_6025), .Z1_t (new_AGEMA_signal_6026), .Z1_f (new_AGEMA_signal_6027) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS22ser_mux_inst_3_XOR2_U1 ( .A0_t (stateArray_MUX_inS22ser_mux_inst_3_Y), .A0_f (new_AGEMA_signal_6025), .A1_t (new_AGEMA_signal_6026), .A1_f (new_AGEMA_signal_6027), .B0_t (plaintext_s0_t[43]), .B0_f (plaintext_s0_f[43]), .B1_t (plaintext_s1_t[43]), .B1_f (plaintext_s1_f[43]), .Z0_t (stateArray_inS22ser[3]), .Z0_f (new_AGEMA_signal_6823), .Z1_t (new_AGEMA_signal_6824), .Z1_f (new_AGEMA_signal_6825) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS22ser_mux_inst_4_XOR1_U1 ( .A0_t (plaintext_s0_t[44]), .A0_f (plaintext_s0_f[44]), .A1_t (plaintext_s1_t[44]), .A1_f (plaintext_s1_f[44]), .B0_t (ciphertext_s0_t[12]), .B0_f (ciphertext_s0_f[12]), .B1_t (ciphertext_s1_t[12]), .B1_f (ciphertext_s1_f[12]), .Z0_t (stateArray_MUX_inS22ser_mux_inst_4_X), .Z0_f (new_AGEMA_signal_4140), .Z1_t (new_AGEMA_signal_4141), .Z1_f (new_AGEMA_signal_4142) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS22ser_mux_inst_4_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS22ser_mux_inst_4_X), .B0_f (new_AGEMA_signal_4140), .B1_t (new_AGEMA_signal_4141), .B1_f (new_AGEMA_signal_4142), .Z0_t (stateArray_MUX_inS22ser_mux_inst_4_Y), .Z0_f (new_AGEMA_signal_6028), .Z1_t (new_AGEMA_signal_6029), .Z1_f (new_AGEMA_signal_6030) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS22ser_mux_inst_4_XOR2_U1 ( .A0_t (stateArray_MUX_inS22ser_mux_inst_4_Y), .A0_f (new_AGEMA_signal_6028), .A1_t (new_AGEMA_signal_6029), .A1_f (new_AGEMA_signal_6030), .B0_t (plaintext_s0_t[44]), .B0_f (plaintext_s0_f[44]), .B1_t (plaintext_s1_t[44]), .B1_f (plaintext_s1_f[44]), .Z0_t (stateArray_inS22ser[4]), .Z0_f (new_AGEMA_signal_6826), .Z1_t (new_AGEMA_signal_6827), .Z1_f (new_AGEMA_signal_6828) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS22ser_mux_inst_5_XOR1_U1 ( .A0_t (plaintext_s0_t[45]), .A0_f (plaintext_s0_f[45]), .A1_t (plaintext_s1_t[45]), .A1_f (plaintext_s1_f[45]), .B0_t (ciphertext_s0_t[13]), .B0_f (ciphertext_s0_f[13]), .B1_t (ciphertext_s1_t[13]), .B1_f (ciphertext_s1_f[13]), .Z0_t (stateArray_MUX_inS22ser_mux_inst_5_X), .Z0_f (new_AGEMA_signal_4149), .Z1_t (new_AGEMA_signal_4150), .Z1_f (new_AGEMA_signal_4151) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS22ser_mux_inst_5_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS22ser_mux_inst_5_X), .B0_f (new_AGEMA_signal_4149), .B1_t (new_AGEMA_signal_4150), .B1_f (new_AGEMA_signal_4151), .Z0_t (stateArray_MUX_inS22ser_mux_inst_5_Y), .Z0_f (new_AGEMA_signal_6031), .Z1_t (new_AGEMA_signal_6032), .Z1_f (new_AGEMA_signal_6033) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS22ser_mux_inst_5_XOR2_U1 ( .A0_t (stateArray_MUX_inS22ser_mux_inst_5_Y), .A0_f (new_AGEMA_signal_6031), .A1_t (new_AGEMA_signal_6032), .A1_f (new_AGEMA_signal_6033), .B0_t (plaintext_s0_t[45]), .B0_f (plaintext_s0_f[45]), .B1_t (plaintext_s1_t[45]), .B1_f (plaintext_s1_f[45]), .Z0_t (stateArray_inS22ser[5]), .Z0_f (new_AGEMA_signal_6829), .Z1_t (new_AGEMA_signal_6830), .Z1_f (new_AGEMA_signal_6831) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS22ser_mux_inst_6_XOR1_U1 ( .A0_t (plaintext_s0_t[46]), .A0_f (plaintext_s0_f[46]), .A1_t (plaintext_s1_t[46]), .A1_f (plaintext_s1_f[46]), .B0_t (ciphertext_s0_t[14]), .B0_f (ciphertext_s0_f[14]), .B1_t (ciphertext_s1_t[14]), .B1_f (ciphertext_s1_f[14]), .Z0_t (stateArray_MUX_inS22ser_mux_inst_6_X), .Z0_f (new_AGEMA_signal_4158), .Z1_t (new_AGEMA_signal_4159), .Z1_f (new_AGEMA_signal_4160) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS22ser_mux_inst_6_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS22ser_mux_inst_6_X), .B0_f (new_AGEMA_signal_4158), .B1_t (new_AGEMA_signal_4159), .B1_f (new_AGEMA_signal_4160), .Z0_t (stateArray_MUX_inS22ser_mux_inst_6_Y), .Z0_f (new_AGEMA_signal_6034), .Z1_t (new_AGEMA_signal_6035), .Z1_f (new_AGEMA_signal_6036) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS22ser_mux_inst_6_XOR2_U1 ( .A0_t (stateArray_MUX_inS22ser_mux_inst_6_Y), .A0_f (new_AGEMA_signal_6034), .A1_t (new_AGEMA_signal_6035), .A1_f (new_AGEMA_signal_6036), .B0_t (plaintext_s0_t[46]), .B0_f (plaintext_s0_f[46]), .B1_t (plaintext_s1_t[46]), .B1_f (plaintext_s1_f[46]), .Z0_t (stateArray_inS22ser[6]), .Z0_f (new_AGEMA_signal_6832), .Z1_t (new_AGEMA_signal_6833), .Z1_f (new_AGEMA_signal_6834) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS22ser_mux_inst_7_XOR1_U1 ( .A0_t (plaintext_s0_t[47]), .A0_f (plaintext_s0_f[47]), .A1_t (plaintext_s1_t[47]), .A1_f (plaintext_s1_f[47]), .B0_t (ciphertext_s0_t[15]), .B0_f (ciphertext_s0_f[15]), .B1_t (ciphertext_s1_t[15]), .B1_f (ciphertext_s1_f[15]), .Z0_t (stateArray_MUX_inS22ser_mux_inst_7_X), .Z0_f (new_AGEMA_signal_4167), .Z1_t (new_AGEMA_signal_4168), .Z1_f (new_AGEMA_signal_4169) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS22ser_mux_inst_7_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS22ser_mux_inst_7_X), .B0_f (new_AGEMA_signal_4167), .B1_t (new_AGEMA_signal_4168), .B1_f (new_AGEMA_signal_4169), .Z0_t (stateArray_MUX_inS22ser_mux_inst_7_Y), .Z0_f (new_AGEMA_signal_6037), .Z1_t (new_AGEMA_signal_6038), .Z1_f (new_AGEMA_signal_6039) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS22ser_mux_inst_7_XOR2_U1 ( .A0_t (stateArray_MUX_inS22ser_mux_inst_7_Y), .A0_f (new_AGEMA_signal_6037), .A1_t (new_AGEMA_signal_6038), .A1_f (new_AGEMA_signal_6039), .B0_t (plaintext_s0_t[47]), .B0_f (plaintext_s0_f[47]), .B1_t (plaintext_s1_t[47]), .B1_f (plaintext_s1_f[47]), .Z0_t (stateArray_inS22ser[7]), .Z0_f (new_AGEMA_signal_6835), .Z1_t (new_AGEMA_signal_6836), .Z1_f (new_AGEMA_signal_6837) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS30_MC_mux_inst_0_XOR1_U1 ( .A0_t (ciphertext_s0_t[96]), .A0_f (ciphertext_s0_f[96]), .A1_t (ciphertext_s1_t[96]), .A1_f (ciphertext_s1_f[96]), .B0_t (StateInMC[8]), .B0_f (new_AGEMA_signal_9328), .B1_t (new_AGEMA_signal_9329), .B1_f (new_AGEMA_signal_9330), .Z0_t (stateArray_MUX_outS30_MC_mux_inst_0_X), .Z0_f (new_AGEMA_signal_9825), .Z1_t (new_AGEMA_signal_9826), .Z1_f (new_AGEMA_signal_9827) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS30_MC_mux_inst_0_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (stateArray_MUX_outS30_MC_mux_inst_0_X), .B0_f (new_AGEMA_signal_9825), .B1_t (new_AGEMA_signal_9826), .B1_f (new_AGEMA_signal_9827), .Z0_t (stateArray_MUX_outS30_MC_mux_inst_0_Y), .Z0_f (new_AGEMA_signal_10355), .Z1_t (new_AGEMA_signal_10356), .Z1_f (new_AGEMA_signal_10357) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS30_MC_mux_inst_0_XOR2_U1 ( .A0_t (stateArray_MUX_outS30_MC_mux_inst_0_Y), .A0_f (new_AGEMA_signal_10355), .A1_t (new_AGEMA_signal_10356), .A1_f (new_AGEMA_signal_10357), .B0_t (ciphertext_s0_t[96]), .B0_f (ciphertext_s0_f[96]), .B1_t (ciphertext_s1_t[96]), .B1_f (ciphertext_s1_f[96]), .Z0_t (stateArray_outS30ser_MC[0]), .Z0_f (new_AGEMA_signal_10478), .Z1_t (new_AGEMA_signal_10479), .Z1_f (new_AGEMA_signal_10480) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS30_MC_mux_inst_1_XOR1_U1 ( .A0_t (ciphertext_s0_t[97]), .A0_f (ciphertext_s0_f[97]), .A1_t (ciphertext_s1_t[97]), .A1_f (ciphertext_s1_f[97]), .B0_t (StateInMC[9]), .B0_f (new_AGEMA_signal_9849), .B1_t (new_AGEMA_signal_9850), .B1_f (new_AGEMA_signal_9851), .Z0_t (stateArray_MUX_outS30_MC_mux_inst_1_X), .Z0_f (new_AGEMA_signal_10358), .Z1_t (new_AGEMA_signal_10359), .Z1_f (new_AGEMA_signal_10360) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS30_MC_mux_inst_1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (stateArray_MUX_outS30_MC_mux_inst_1_X), .B0_f (new_AGEMA_signal_10358), .B1_t (new_AGEMA_signal_10359), .B1_f (new_AGEMA_signal_10360), .Z0_t (stateArray_MUX_outS30_MC_mux_inst_1_Y), .Z0_f (new_AGEMA_signal_10481), .Z1_t (new_AGEMA_signal_10482), .Z1_f (new_AGEMA_signal_10483) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS30_MC_mux_inst_1_XOR2_U1 ( .A0_t (stateArray_MUX_outS30_MC_mux_inst_1_Y), .A0_f (new_AGEMA_signal_10481), .A1_t (new_AGEMA_signal_10482), .A1_f (new_AGEMA_signal_10483), .B0_t (ciphertext_s0_t[97]), .B0_f (ciphertext_s0_f[97]), .B1_t (ciphertext_s1_t[97]), .B1_f (ciphertext_s1_f[97]), .Z0_t (stateArray_outS30ser_MC[1]), .Z0_f (new_AGEMA_signal_10619), .Z1_t (new_AGEMA_signal_10620), .Z1_f (new_AGEMA_signal_10621) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS30_MC_mux_inst_2_XOR1_U1 ( .A0_t (ciphertext_s0_t[98]), .A0_f (ciphertext_s0_f[98]), .A1_t (ciphertext_s1_t[98]), .A1_f (ciphertext_s1_f[98]), .B0_t (StateInMC[10]), .B0_f (new_AGEMA_signal_9334), .B1_t (new_AGEMA_signal_9335), .B1_f (new_AGEMA_signal_9336), .Z0_t (stateArray_MUX_outS30_MC_mux_inst_2_X), .Z0_f (new_AGEMA_signal_9828), .Z1_t (new_AGEMA_signal_9829), .Z1_f (new_AGEMA_signal_9830) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS30_MC_mux_inst_2_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (stateArray_MUX_outS30_MC_mux_inst_2_X), .B0_f (new_AGEMA_signal_9828), .B1_t (new_AGEMA_signal_9829), .B1_f (new_AGEMA_signal_9830), .Z0_t (stateArray_MUX_outS30_MC_mux_inst_2_Y), .Z0_f (new_AGEMA_signal_10361), .Z1_t (new_AGEMA_signal_10362), .Z1_f (new_AGEMA_signal_10363) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS30_MC_mux_inst_2_XOR2_U1 ( .A0_t (stateArray_MUX_outS30_MC_mux_inst_2_Y), .A0_f (new_AGEMA_signal_10361), .A1_t (new_AGEMA_signal_10362), .A1_f (new_AGEMA_signal_10363), .B0_t (ciphertext_s0_t[98]), .B0_f (ciphertext_s0_f[98]), .B1_t (ciphertext_s1_t[98]), .B1_f (ciphertext_s1_f[98]), .Z0_t (stateArray_outS30ser_MC[2]), .Z0_f (new_AGEMA_signal_10484), .Z1_t (new_AGEMA_signal_10485), .Z1_f (new_AGEMA_signal_10486) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS30_MC_mux_inst_3_XOR1_U1 ( .A0_t (ciphertext_s0_t[99]), .A0_f (ciphertext_s0_f[99]), .A1_t (ciphertext_s1_t[99]), .A1_f (ciphertext_s1_f[99]), .B0_t (StateInMC[11]), .B0_f (new_AGEMA_signal_9852), .B1_t (new_AGEMA_signal_9853), .B1_f (new_AGEMA_signal_9854), .Z0_t (stateArray_MUX_outS30_MC_mux_inst_3_X), .Z0_f (new_AGEMA_signal_10364), .Z1_t (new_AGEMA_signal_10365), .Z1_f (new_AGEMA_signal_10366) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS30_MC_mux_inst_3_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (stateArray_MUX_outS30_MC_mux_inst_3_X), .B0_f (new_AGEMA_signal_10364), .B1_t (new_AGEMA_signal_10365), .B1_f (new_AGEMA_signal_10366), .Z0_t (stateArray_MUX_outS30_MC_mux_inst_3_Y), .Z0_f (new_AGEMA_signal_10487), .Z1_t (new_AGEMA_signal_10488), .Z1_f (new_AGEMA_signal_10489) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS30_MC_mux_inst_3_XOR2_U1 ( .A0_t (stateArray_MUX_outS30_MC_mux_inst_3_Y), .A0_f (new_AGEMA_signal_10487), .A1_t (new_AGEMA_signal_10488), .A1_f (new_AGEMA_signal_10489), .B0_t (ciphertext_s0_t[99]), .B0_f (ciphertext_s0_f[99]), .B1_t (ciphertext_s1_t[99]), .B1_f (ciphertext_s1_f[99]), .Z0_t (stateArray_outS30ser_MC[3]), .Z0_f (new_AGEMA_signal_10622), .Z1_t (new_AGEMA_signal_10623), .Z1_f (new_AGEMA_signal_10624) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS30_MC_mux_inst_4_XOR1_U1 ( .A0_t (ciphertext_s0_t[100]), .A0_f (ciphertext_s0_f[100]), .A1_t (ciphertext_s1_t[100]), .A1_f (ciphertext_s1_f[100]), .B0_t (StateInMC[12]), .B0_f (new_AGEMA_signal_9855), .B1_t (new_AGEMA_signal_9856), .B1_f (new_AGEMA_signal_9857), .Z0_t (stateArray_MUX_outS30_MC_mux_inst_4_X), .Z0_f (new_AGEMA_signal_10367), .Z1_t (new_AGEMA_signal_10368), .Z1_f (new_AGEMA_signal_10369) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS30_MC_mux_inst_4_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (stateArray_MUX_outS30_MC_mux_inst_4_X), .B0_f (new_AGEMA_signal_10367), .B1_t (new_AGEMA_signal_10368), .B1_f (new_AGEMA_signal_10369), .Z0_t (stateArray_MUX_outS30_MC_mux_inst_4_Y), .Z0_f (new_AGEMA_signal_10490), .Z1_t (new_AGEMA_signal_10491), .Z1_f (new_AGEMA_signal_10492) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS30_MC_mux_inst_4_XOR2_U1 ( .A0_t (stateArray_MUX_outS30_MC_mux_inst_4_Y), .A0_f (new_AGEMA_signal_10490), .A1_t (new_AGEMA_signal_10491), .A1_f (new_AGEMA_signal_10492), .B0_t (ciphertext_s0_t[100]), .B0_f (ciphertext_s0_f[100]), .B1_t (ciphertext_s1_t[100]), .B1_f (ciphertext_s1_f[100]), .Z0_t (stateArray_outS30ser_MC[4]), .Z0_f (new_AGEMA_signal_10625), .Z1_t (new_AGEMA_signal_10626), .Z1_f (new_AGEMA_signal_10627) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS30_MC_mux_inst_5_XOR1_U1 ( .A0_t (ciphertext_s0_t[101]), .A0_f (ciphertext_s0_f[101]), .A1_t (ciphertext_s1_t[101]), .A1_f (ciphertext_s1_f[101]), .B0_t (StateInMC[13]), .B0_f (new_AGEMA_signal_9343), .B1_t (new_AGEMA_signal_9344), .B1_f (new_AGEMA_signal_9345), .Z0_t (stateArray_MUX_outS30_MC_mux_inst_5_X), .Z0_f (new_AGEMA_signal_9831), .Z1_t (new_AGEMA_signal_9832), .Z1_f (new_AGEMA_signal_9833) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS30_MC_mux_inst_5_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (stateArray_MUX_outS30_MC_mux_inst_5_X), .B0_f (new_AGEMA_signal_9831), .B1_t (new_AGEMA_signal_9832), .B1_f (new_AGEMA_signal_9833), .Z0_t (stateArray_MUX_outS30_MC_mux_inst_5_Y), .Z0_f (new_AGEMA_signal_10370), .Z1_t (new_AGEMA_signal_10371), .Z1_f (new_AGEMA_signal_10372) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS30_MC_mux_inst_5_XOR2_U1 ( .A0_t (stateArray_MUX_outS30_MC_mux_inst_5_Y), .A0_f (new_AGEMA_signal_10370), .A1_t (new_AGEMA_signal_10371), .A1_f (new_AGEMA_signal_10372), .B0_t (ciphertext_s0_t[101]), .B0_f (ciphertext_s0_f[101]), .B1_t (ciphertext_s1_t[101]), .B1_f (ciphertext_s1_f[101]), .Z0_t (stateArray_outS30ser_MC[5]), .Z0_f (new_AGEMA_signal_10493), .Z1_t (new_AGEMA_signal_10494), .Z1_f (new_AGEMA_signal_10495) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS30_MC_mux_inst_6_XOR1_U1 ( .A0_t (ciphertext_s0_t[102]), .A0_f (ciphertext_s0_f[102]), .A1_t (ciphertext_s1_t[102]), .A1_f (ciphertext_s1_f[102]), .B0_t (StateInMC[14]), .B0_f (new_AGEMA_signal_9346), .B1_t (new_AGEMA_signal_9347), .B1_f (new_AGEMA_signal_9348), .Z0_t (stateArray_MUX_outS30_MC_mux_inst_6_X), .Z0_f (new_AGEMA_signal_9834), .Z1_t (new_AGEMA_signal_9835), .Z1_f (new_AGEMA_signal_9836) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS30_MC_mux_inst_6_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (stateArray_MUX_outS30_MC_mux_inst_6_X), .B0_f (new_AGEMA_signal_9834), .B1_t (new_AGEMA_signal_9835), .B1_f (new_AGEMA_signal_9836), .Z0_t (stateArray_MUX_outS30_MC_mux_inst_6_Y), .Z0_f (new_AGEMA_signal_10373), .Z1_t (new_AGEMA_signal_10374), .Z1_f (new_AGEMA_signal_10375) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS30_MC_mux_inst_6_XOR2_U1 ( .A0_t (stateArray_MUX_outS30_MC_mux_inst_6_Y), .A0_f (new_AGEMA_signal_10373), .A1_t (new_AGEMA_signal_10374), .A1_f (new_AGEMA_signal_10375), .B0_t (ciphertext_s0_t[102]), .B0_f (ciphertext_s0_f[102]), .B1_t (ciphertext_s1_t[102]), .B1_f (ciphertext_s1_f[102]), .Z0_t (stateArray_outS30ser_MC[6]), .Z0_f (new_AGEMA_signal_10496), .Z1_t (new_AGEMA_signal_10497), .Z1_f (new_AGEMA_signal_10498) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS30_MC_mux_inst_7_XOR1_U1 ( .A0_t (ciphertext_s0_t[103]), .A0_f (ciphertext_s0_f[103]), .A1_t (ciphertext_s1_t[103]), .A1_f (ciphertext_s1_f[103]), .B0_t (StateInMC[15]), .B0_f (new_AGEMA_signal_9349), .B1_t (new_AGEMA_signal_9350), .B1_f (new_AGEMA_signal_9351), .Z0_t (stateArray_MUX_outS30_MC_mux_inst_7_X), .Z0_f (new_AGEMA_signal_9837), .Z1_t (new_AGEMA_signal_9838), .Z1_f (new_AGEMA_signal_9839) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS30_MC_mux_inst_7_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (stateArray_MUX_outS30_MC_mux_inst_7_X), .B0_f (new_AGEMA_signal_9837), .B1_t (new_AGEMA_signal_9838), .B1_f (new_AGEMA_signal_9839), .Z0_t (stateArray_MUX_outS30_MC_mux_inst_7_Y), .Z0_f (new_AGEMA_signal_10376), .Z1_t (new_AGEMA_signal_10377), .Z1_f (new_AGEMA_signal_10378) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_outS30_MC_mux_inst_7_XOR2_U1 ( .A0_t (stateArray_MUX_outS30_MC_mux_inst_7_Y), .A0_f (new_AGEMA_signal_10376), .A1_t (new_AGEMA_signal_10377), .A1_f (new_AGEMA_signal_10378), .B0_t (ciphertext_s0_t[103]), .B0_f (ciphertext_s0_f[103]), .B1_t (ciphertext_s1_t[103]), .B1_f (ciphertext_s1_f[103]), .Z0_t (stateArray_outS30ser_MC[7]), .Z0_f (new_AGEMA_signal_10499), .Z1_t (new_AGEMA_signal_10500), .Z1_f (new_AGEMA_signal_10501) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_0_XOR1_U1 ( .A0_t (plaintext_s0_t[8]), .A0_f (plaintext_s0_f[8]), .A1_t (plaintext_s1_t[8]), .A1_f (plaintext_s1_f[8]), .B0_t (stateArray_outS30ser_MC[0]), .B0_f (new_AGEMA_signal_10478), .B1_t (new_AGEMA_signal_10479), .B1_f (new_AGEMA_signal_10480), .Z0_t (stateArray_MUX_inS23ser_mux_inst_0_X), .Z0_f (new_AGEMA_signal_10631), .Z1_t (new_AGEMA_signal_10632), .Z1_f (new_AGEMA_signal_10633) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_0_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS23ser_mux_inst_0_X), .B0_f (new_AGEMA_signal_10631), .B1_t (new_AGEMA_signal_10632), .B1_f (new_AGEMA_signal_10633), .Z0_t (stateArray_MUX_inS23ser_mux_inst_0_Y), .Z0_f (new_AGEMA_signal_10760), .Z1_t (new_AGEMA_signal_10761), .Z1_f (new_AGEMA_signal_10762) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_0_XOR2_U1 ( .A0_t (stateArray_MUX_inS23ser_mux_inst_0_Y), .A0_f (new_AGEMA_signal_10760), .A1_t (new_AGEMA_signal_10761), .A1_f (new_AGEMA_signal_10762), .B0_t (plaintext_s0_t[8]), .B0_f (plaintext_s0_f[8]), .B1_t (plaintext_s1_t[8]), .B1_f (plaintext_s1_f[8]), .Z0_t (stateArray_inS23ser[0]), .Z0_f (new_AGEMA_signal_10877), .Z1_t (new_AGEMA_signal_10878), .Z1_f (new_AGEMA_signal_10879) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_1_XOR1_U1 ( .A0_t (plaintext_s0_t[9]), .A0_f (plaintext_s0_f[9]), .A1_t (plaintext_s1_t[9]), .A1_f (plaintext_s1_f[9]), .B0_t (stateArray_outS30ser_MC[1]), .B0_f (new_AGEMA_signal_10619), .B1_t (new_AGEMA_signal_10620), .B1_f (new_AGEMA_signal_10621), .Z0_t (stateArray_MUX_inS23ser_mux_inst_1_X), .Z0_f (new_AGEMA_signal_10766), .Z1_t (new_AGEMA_signal_10767), .Z1_f (new_AGEMA_signal_10768) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS23ser_mux_inst_1_X), .B0_f (new_AGEMA_signal_10766), .B1_t (new_AGEMA_signal_10767), .B1_f (new_AGEMA_signal_10768), .Z0_t (stateArray_MUX_inS23ser_mux_inst_1_Y), .Z0_f (new_AGEMA_signal_10880), .Z1_t (new_AGEMA_signal_10881), .Z1_f (new_AGEMA_signal_10882) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_1_XOR2_U1 ( .A0_t (stateArray_MUX_inS23ser_mux_inst_1_Y), .A0_f (new_AGEMA_signal_10880), .A1_t (new_AGEMA_signal_10881), .A1_f (new_AGEMA_signal_10882), .B0_t (plaintext_s0_t[9]), .B0_f (plaintext_s0_f[9]), .B1_t (plaintext_s1_t[9]), .B1_f (plaintext_s1_f[9]), .Z0_t (stateArray_inS23ser[1]), .Z0_f (new_AGEMA_signal_11003), .Z1_t (new_AGEMA_signal_11004), .Z1_f (new_AGEMA_signal_11005) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_2_XOR1_U1 ( .A0_t (plaintext_s0_t[10]), .A0_f (plaintext_s0_f[10]), .A1_t (plaintext_s1_t[10]), .A1_f (plaintext_s1_f[10]), .B0_t (stateArray_outS30ser_MC[2]), .B0_f (new_AGEMA_signal_10484), .B1_t (new_AGEMA_signal_10485), .B1_f (new_AGEMA_signal_10486), .Z0_t (stateArray_MUX_inS23ser_mux_inst_2_X), .Z0_f (new_AGEMA_signal_10637), .Z1_t (new_AGEMA_signal_10638), .Z1_f (new_AGEMA_signal_10639) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_2_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS23ser_mux_inst_2_X), .B0_f (new_AGEMA_signal_10637), .B1_t (new_AGEMA_signal_10638), .B1_f (new_AGEMA_signal_10639), .Z0_t (stateArray_MUX_inS23ser_mux_inst_2_Y), .Z0_f (new_AGEMA_signal_10769), .Z1_t (new_AGEMA_signal_10770), .Z1_f (new_AGEMA_signal_10771) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_2_XOR2_U1 ( .A0_t (stateArray_MUX_inS23ser_mux_inst_2_Y), .A0_f (new_AGEMA_signal_10769), .A1_t (new_AGEMA_signal_10770), .A1_f (new_AGEMA_signal_10771), .B0_t (plaintext_s0_t[10]), .B0_f (plaintext_s0_f[10]), .B1_t (plaintext_s1_t[10]), .B1_f (plaintext_s1_f[10]), .Z0_t (stateArray_inS23ser[2]), .Z0_f (new_AGEMA_signal_10883), .Z1_t (new_AGEMA_signal_10884), .Z1_f (new_AGEMA_signal_10885) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_3_XOR1_U1 ( .A0_t (plaintext_s0_t[11]), .A0_f (plaintext_s0_f[11]), .A1_t (plaintext_s1_t[11]), .A1_f (plaintext_s1_f[11]), .B0_t (stateArray_outS30ser_MC[3]), .B0_f (new_AGEMA_signal_10622), .B1_t (new_AGEMA_signal_10623), .B1_f (new_AGEMA_signal_10624), .Z0_t (stateArray_MUX_inS23ser_mux_inst_3_X), .Z0_f (new_AGEMA_signal_10775), .Z1_t (new_AGEMA_signal_10776), .Z1_f (new_AGEMA_signal_10777) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_3_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS23ser_mux_inst_3_X), .B0_f (new_AGEMA_signal_10775), .B1_t (new_AGEMA_signal_10776), .B1_f (new_AGEMA_signal_10777), .Z0_t (stateArray_MUX_inS23ser_mux_inst_3_Y), .Z0_f (new_AGEMA_signal_10886), .Z1_t (new_AGEMA_signal_10887), .Z1_f (new_AGEMA_signal_10888) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_3_XOR2_U1 ( .A0_t (stateArray_MUX_inS23ser_mux_inst_3_Y), .A0_f (new_AGEMA_signal_10886), .A1_t (new_AGEMA_signal_10887), .A1_f (new_AGEMA_signal_10888), .B0_t (plaintext_s0_t[11]), .B0_f (plaintext_s0_f[11]), .B1_t (plaintext_s1_t[11]), .B1_f (plaintext_s1_f[11]), .Z0_t (stateArray_inS23ser[3]), .Z0_f (new_AGEMA_signal_11006), .Z1_t (new_AGEMA_signal_11007), .Z1_f (new_AGEMA_signal_11008) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_4_XOR1_U1 ( .A0_t (plaintext_s0_t[12]), .A0_f (plaintext_s0_f[12]), .A1_t (plaintext_s1_t[12]), .A1_f (plaintext_s1_f[12]), .B0_t (stateArray_outS30ser_MC[4]), .B0_f (new_AGEMA_signal_10625), .B1_t (new_AGEMA_signal_10626), .B1_f (new_AGEMA_signal_10627), .Z0_t (stateArray_MUX_inS23ser_mux_inst_4_X), .Z0_f (new_AGEMA_signal_10781), .Z1_t (new_AGEMA_signal_10782), .Z1_f (new_AGEMA_signal_10783) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_4_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS23ser_mux_inst_4_X), .B0_f (new_AGEMA_signal_10781), .B1_t (new_AGEMA_signal_10782), .B1_f (new_AGEMA_signal_10783), .Z0_t (stateArray_MUX_inS23ser_mux_inst_4_Y), .Z0_f (new_AGEMA_signal_10889), .Z1_t (new_AGEMA_signal_10890), .Z1_f (new_AGEMA_signal_10891) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_4_XOR2_U1 ( .A0_t (stateArray_MUX_inS23ser_mux_inst_4_Y), .A0_f (new_AGEMA_signal_10889), .A1_t (new_AGEMA_signal_10890), .A1_f (new_AGEMA_signal_10891), .B0_t (plaintext_s0_t[12]), .B0_f (plaintext_s0_f[12]), .B1_t (plaintext_s1_t[12]), .B1_f (plaintext_s1_f[12]), .Z0_t (stateArray_inS23ser[4]), .Z0_f (new_AGEMA_signal_11009), .Z1_t (new_AGEMA_signal_11010), .Z1_f (new_AGEMA_signal_11011) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_5_XOR1_U1 ( .A0_t (plaintext_s0_t[13]), .A0_f (plaintext_s0_f[13]), .A1_t (plaintext_s1_t[13]), .A1_f (plaintext_s1_f[13]), .B0_t (stateArray_outS30ser_MC[5]), .B0_f (new_AGEMA_signal_10493), .B1_t (new_AGEMA_signal_10494), .B1_f (new_AGEMA_signal_10495), .Z0_t (stateArray_MUX_inS23ser_mux_inst_5_X), .Z0_f (new_AGEMA_signal_10643), .Z1_t (new_AGEMA_signal_10644), .Z1_f (new_AGEMA_signal_10645) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_5_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS23ser_mux_inst_5_X), .B0_f (new_AGEMA_signal_10643), .B1_t (new_AGEMA_signal_10644), .B1_f (new_AGEMA_signal_10645), .Z0_t (stateArray_MUX_inS23ser_mux_inst_5_Y), .Z0_f (new_AGEMA_signal_10784), .Z1_t (new_AGEMA_signal_10785), .Z1_f (new_AGEMA_signal_10786) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_5_XOR2_U1 ( .A0_t (stateArray_MUX_inS23ser_mux_inst_5_Y), .A0_f (new_AGEMA_signal_10784), .A1_t (new_AGEMA_signal_10785), .A1_f (new_AGEMA_signal_10786), .B0_t (plaintext_s0_t[13]), .B0_f (plaintext_s0_f[13]), .B1_t (plaintext_s1_t[13]), .B1_f (plaintext_s1_f[13]), .Z0_t (stateArray_inS23ser[5]), .Z0_f (new_AGEMA_signal_10892), .Z1_t (new_AGEMA_signal_10893), .Z1_f (new_AGEMA_signal_10894) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_6_XOR1_U1 ( .A0_t (plaintext_s0_t[14]), .A0_f (plaintext_s0_f[14]), .A1_t (plaintext_s1_t[14]), .A1_f (plaintext_s1_f[14]), .B0_t (stateArray_outS30ser_MC[6]), .B0_f (new_AGEMA_signal_10496), .B1_t (new_AGEMA_signal_10497), .B1_f (new_AGEMA_signal_10498), .Z0_t (stateArray_MUX_inS23ser_mux_inst_6_X), .Z0_f (new_AGEMA_signal_10649), .Z1_t (new_AGEMA_signal_10650), .Z1_f (new_AGEMA_signal_10651) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_6_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS23ser_mux_inst_6_X), .B0_f (new_AGEMA_signal_10649), .B1_t (new_AGEMA_signal_10650), .B1_f (new_AGEMA_signal_10651), .Z0_t (stateArray_MUX_inS23ser_mux_inst_6_Y), .Z0_f (new_AGEMA_signal_10787), .Z1_t (new_AGEMA_signal_10788), .Z1_f (new_AGEMA_signal_10789) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_6_XOR2_U1 ( .A0_t (stateArray_MUX_inS23ser_mux_inst_6_Y), .A0_f (new_AGEMA_signal_10787), .A1_t (new_AGEMA_signal_10788), .A1_f (new_AGEMA_signal_10789), .B0_t (plaintext_s0_t[14]), .B0_f (plaintext_s0_f[14]), .B1_t (plaintext_s1_t[14]), .B1_f (plaintext_s1_f[14]), .Z0_t (stateArray_inS23ser[6]), .Z0_f (new_AGEMA_signal_10895), .Z1_t (new_AGEMA_signal_10896), .Z1_f (new_AGEMA_signal_10897) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_7_XOR1_U1 ( .A0_t (plaintext_s0_t[15]), .A0_f (plaintext_s0_f[15]), .A1_t (plaintext_s1_t[15]), .A1_f (plaintext_s1_f[15]), .B0_t (stateArray_outS30ser_MC[7]), .B0_f (new_AGEMA_signal_10499), .B1_t (new_AGEMA_signal_10500), .B1_f (new_AGEMA_signal_10501), .Z0_t (stateArray_MUX_inS23ser_mux_inst_7_X), .Z0_f (new_AGEMA_signal_10655), .Z1_t (new_AGEMA_signal_10656), .Z1_f (new_AGEMA_signal_10657) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_7_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS23ser_mux_inst_7_X), .B0_f (new_AGEMA_signal_10655), .B1_t (new_AGEMA_signal_10656), .B1_f (new_AGEMA_signal_10657), .Z0_t (stateArray_MUX_inS23ser_mux_inst_7_Y), .Z0_f (new_AGEMA_signal_10790), .Z1_t (new_AGEMA_signal_10791), .Z1_f (new_AGEMA_signal_10792) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_7_XOR2_U1 ( .A0_t (stateArray_MUX_inS23ser_mux_inst_7_Y), .A0_f (new_AGEMA_signal_10790), .A1_t (new_AGEMA_signal_10791), .A1_f (new_AGEMA_signal_10792), .B0_t (plaintext_s0_t[15]), .B0_f (plaintext_s0_f[15]), .B1_t (plaintext_s1_t[15]), .B1_f (plaintext_s1_f[15]), .Z0_t (stateArray_inS23ser[7]), .Z0_f (new_AGEMA_signal_10898), .Z1_t (new_AGEMA_signal_10899), .Z1_f (new_AGEMA_signal_10900) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS30ser_mux_inst_0_XOR1_U1 ( .A0_t (plaintext_s0_t[96]), .A0_f (plaintext_s0_f[96]), .A1_t (plaintext_s1_t[96]), .A1_f (plaintext_s1_f[96]), .B0_t (ciphertext_s0_t[64]), .B0_f (ciphertext_s0_f[64]), .B1_t (ciphertext_s1_t[64]), .B1_f (ciphertext_s1_f[64]), .Z0_t (stateArray_MUX_inS30ser_mux_inst_0_X), .Z0_f (new_AGEMA_signal_4176), .Z1_t (new_AGEMA_signal_4177), .Z1_f (new_AGEMA_signal_4178) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS30ser_mux_inst_0_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS30ser_mux_inst_0_X), .B0_f (new_AGEMA_signal_4176), .B1_t (new_AGEMA_signal_4177), .B1_f (new_AGEMA_signal_4178), .Z0_t (stateArray_MUX_inS30ser_mux_inst_0_Y), .Z0_f (new_AGEMA_signal_6040), .Z1_t (new_AGEMA_signal_6041), .Z1_f (new_AGEMA_signal_6042) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS30ser_mux_inst_0_XOR2_U1 ( .A0_t (stateArray_MUX_inS30ser_mux_inst_0_Y), .A0_f (new_AGEMA_signal_6040), .A1_t (new_AGEMA_signal_6041), .A1_f (new_AGEMA_signal_6042), .B0_t (plaintext_s0_t[96]), .B0_f (plaintext_s0_f[96]), .B1_t (plaintext_s1_t[96]), .B1_f (plaintext_s1_f[96]), .Z0_t (stateArray_inS30ser[0]), .Z0_f (new_AGEMA_signal_6838), .Z1_t (new_AGEMA_signal_6839), .Z1_f (new_AGEMA_signal_6840) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS30ser_mux_inst_1_XOR1_U1 ( .A0_t (plaintext_s0_t[97]), .A0_f (plaintext_s0_f[97]), .A1_t (plaintext_s1_t[97]), .A1_f (plaintext_s1_f[97]), .B0_t (ciphertext_s0_t[65]), .B0_f (ciphertext_s0_f[65]), .B1_t (ciphertext_s1_t[65]), .B1_f (ciphertext_s1_f[65]), .Z0_t (stateArray_MUX_inS30ser_mux_inst_1_X), .Z0_f (new_AGEMA_signal_4185), .Z1_t (new_AGEMA_signal_4186), .Z1_f (new_AGEMA_signal_4187) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS30ser_mux_inst_1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS30ser_mux_inst_1_X), .B0_f (new_AGEMA_signal_4185), .B1_t (new_AGEMA_signal_4186), .B1_f (new_AGEMA_signal_4187), .Z0_t (stateArray_MUX_inS30ser_mux_inst_1_Y), .Z0_f (new_AGEMA_signal_6043), .Z1_t (new_AGEMA_signal_6044), .Z1_f (new_AGEMA_signal_6045) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS30ser_mux_inst_1_XOR2_U1 ( .A0_t (stateArray_MUX_inS30ser_mux_inst_1_Y), .A0_f (new_AGEMA_signal_6043), .A1_t (new_AGEMA_signal_6044), .A1_f (new_AGEMA_signal_6045), .B0_t (plaintext_s0_t[97]), .B0_f (plaintext_s0_f[97]), .B1_t (plaintext_s1_t[97]), .B1_f (plaintext_s1_f[97]), .Z0_t (stateArray_inS30ser[1]), .Z0_f (new_AGEMA_signal_6841), .Z1_t (new_AGEMA_signal_6842), .Z1_f (new_AGEMA_signal_6843) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS30ser_mux_inst_2_XOR1_U1 ( .A0_t (plaintext_s0_t[98]), .A0_f (plaintext_s0_f[98]), .A1_t (plaintext_s1_t[98]), .A1_f (plaintext_s1_f[98]), .B0_t (ciphertext_s0_t[66]), .B0_f (ciphertext_s0_f[66]), .B1_t (ciphertext_s1_t[66]), .B1_f (ciphertext_s1_f[66]), .Z0_t (stateArray_MUX_inS30ser_mux_inst_2_X), .Z0_f (new_AGEMA_signal_4194), .Z1_t (new_AGEMA_signal_4195), .Z1_f (new_AGEMA_signal_4196) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS30ser_mux_inst_2_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS30ser_mux_inst_2_X), .B0_f (new_AGEMA_signal_4194), .B1_t (new_AGEMA_signal_4195), .B1_f (new_AGEMA_signal_4196), .Z0_t (stateArray_MUX_inS30ser_mux_inst_2_Y), .Z0_f (new_AGEMA_signal_6046), .Z1_t (new_AGEMA_signal_6047), .Z1_f (new_AGEMA_signal_6048) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS30ser_mux_inst_2_XOR2_U1 ( .A0_t (stateArray_MUX_inS30ser_mux_inst_2_Y), .A0_f (new_AGEMA_signal_6046), .A1_t (new_AGEMA_signal_6047), .A1_f (new_AGEMA_signal_6048), .B0_t (plaintext_s0_t[98]), .B0_f (plaintext_s0_f[98]), .B1_t (plaintext_s1_t[98]), .B1_f (plaintext_s1_f[98]), .Z0_t (stateArray_inS30ser[2]), .Z0_f (new_AGEMA_signal_6844), .Z1_t (new_AGEMA_signal_6845), .Z1_f (new_AGEMA_signal_6846) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS30ser_mux_inst_3_XOR1_U1 ( .A0_t (plaintext_s0_t[99]), .A0_f (plaintext_s0_f[99]), .A1_t (plaintext_s1_t[99]), .A1_f (plaintext_s1_f[99]), .B0_t (ciphertext_s0_t[67]), .B0_f (ciphertext_s0_f[67]), .B1_t (ciphertext_s1_t[67]), .B1_f (ciphertext_s1_f[67]), .Z0_t (stateArray_MUX_inS30ser_mux_inst_3_X), .Z0_f (new_AGEMA_signal_4203), .Z1_t (new_AGEMA_signal_4204), .Z1_f (new_AGEMA_signal_4205) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS30ser_mux_inst_3_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS30ser_mux_inst_3_X), .B0_f (new_AGEMA_signal_4203), .B1_t (new_AGEMA_signal_4204), .B1_f (new_AGEMA_signal_4205), .Z0_t (stateArray_MUX_inS30ser_mux_inst_3_Y), .Z0_f (new_AGEMA_signal_6049), .Z1_t (new_AGEMA_signal_6050), .Z1_f (new_AGEMA_signal_6051) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS30ser_mux_inst_3_XOR2_U1 ( .A0_t (stateArray_MUX_inS30ser_mux_inst_3_Y), .A0_f (new_AGEMA_signal_6049), .A1_t (new_AGEMA_signal_6050), .A1_f (new_AGEMA_signal_6051), .B0_t (plaintext_s0_t[99]), .B0_f (plaintext_s0_f[99]), .B1_t (plaintext_s1_t[99]), .B1_f (plaintext_s1_f[99]), .Z0_t (stateArray_inS30ser[3]), .Z0_f (new_AGEMA_signal_6847), .Z1_t (new_AGEMA_signal_6848), .Z1_f (new_AGEMA_signal_6849) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS30ser_mux_inst_4_XOR1_U1 ( .A0_t (plaintext_s0_t[100]), .A0_f (plaintext_s0_f[100]), .A1_t (plaintext_s1_t[100]), .A1_f (plaintext_s1_f[100]), .B0_t (ciphertext_s0_t[68]), .B0_f (ciphertext_s0_f[68]), .B1_t (ciphertext_s1_t[68]), .B1_f (ciphertext_s1_f[68]), .Z0_t (stateArray_MUX_inS30ser_mux_inst_4_X), .Z0_f (new_AGEMA_signal_4212), .Z1_t (new_AGEMA_signal_4213), .Z1_f (new_AGEMA_signal_4214) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS30ser_mux_inst_4_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS30ser_mux_inst_4_X), .B0_f (new_AGEMA_signal_4212), .B1_t (new_AGEMA_signal_4213), .B1_f (new_AGEMA_signal_4214), .Z0_t (stateArray_MUX_inS30ser_mux_inst_4_Y), .Z0_f (new_AGEMA_signal_6052), .Z1_t (new_AGEMA_signal_6053), .Z1_f (new_AGEMA_signal_6054) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS30ser_mux_inst_4_XOR2_U1 ( .A0_t (stateArray_MUX_inS30ser_mux_inst_4_Y), .A0_f (new_AGEMA_signal_6052), .A1_t (new_AGEMA_signal_6053), .A1_f (new_AGEMA_signal_6054), .B0_t (plaintext_s0_t[100]), .B0_f (plaintext_s0_f[100]), .B1_t (plaintext_s1_t[100]), .B1_f (plaintext_s1_f[100]), .Z0_t (stateArray_inS30ser[4]), .Z0_f (new_AGEMA_signal_6850), .Z1_t (new_AGEMA_signal_6851), .Z1_f (new_AGEMA_signal_6852) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS30ser_mux_inst_5_XOR1_U1 ( .A0_t (plaintext_s0_t[101]), .A0_f (plaintext_s0_f[101]), .A1_t (plaintext_s1_t[101]), .A1_f (plaintext_s1_f[101]), .B0_t (ciphertext_s0_t[69]), .B0_f (ciphertext_s0_f[69]), .B1_t (ciphertext_s1_t[69]), .B1_f (ciphertext_s1_f[69]), .Z0_t (stateArray_MUX_inS30ser_mux_inst_5_X), .Z0_f (new_AGEMA_signal_4221), .Z1_t (new_AGEMA_signal_4222), .Z1_f (new_AGEMA_signal_4223) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS30ser_mux_inst_5_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS30ser_mux_inst_5_X), .B0_f (new_AGEMA_signal_4221), .B1_t (new_AGEMA_signal_4222), .B1_f (new_AGEMA_signal_4223), .Z0_t (stateArray_MUX_inS30ser_mux_inst_5_Y), .Z0_f (new_AGEMA_signal_6055), .Z1_t (new_AGEMA_signal_6056), .Z1_f (new_AGEMA_signal_6057) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS30ser_mux_inst_5_XOR2_U1 ( .A0_t (stateArray_MUX_inS30ser_mux_inst_5_Y), .A0_f (new_AGEMA_signal_6055), .A1_t (new_AGEMA_signal_6056), .A1_f (new_AGEMA_signal_6057), .B0_t (plaintext_s0_t[101]), .B0_f (plaintext_s0_f[101]), .B1_t (plaintext_s1_t[101]), .B1_f (plaintext_s1_f[101]), .Z0_t (stateArray_inS30ser[5]), .Z0_f (new_AGEMA_signal_6853), .Z1_t (new_AGEMA_signal_6854), .Z1_f (new_AGEMA_signal_6855) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS30ser_mux_inst_6_XOR1_U1 ( .A0_t (plaintext_s0_t[102]), .A0_f (plaintext_s0_f[102]), .A1_t (plaintext_s1_t[102]), .A1_f (plaintext_s1_f[102]), .B0_t (ciphertext_s0_t[70]), .B0_f (ciphertext_s0_f[70]), .B1_t (ciphertext_s1_t[70]), .B1_f (ciphertext_s1_f[70]), .Z0_t (stateArray_MUX_inS30ser_mux_inst_6_X), .Z0_f (new_AGEMA_signal_4230), .Z1_t (new_AGEMA_signal_4231), .Z1_f (new_AGEMA_signal_4232) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS30ser_mux_inst_6_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS30ser_mux_inst_6_X), .B0_f (new_AGEMA_signal_4230), .B1_t (new_AGEMA_signal_4231), .B1_f (new_AGEMA_signal_4232), .Z0_t (stateArray_MUX_inS30ser_mux_inst_6_Y), .Z0_f (new_AGEMA_signal_6058), .Z1_t (new_AGEMA_signal_6059), .Z1_f (new_AGEMA_signal_6060) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS30ser_mux_inst_6_XOR2_U1 ( .A0_t (stateArray_MUX_inS30ser_mux_inst_6_Y), .A0_f (new_AGEMA_signal_6058), .A1_t (new_AGEMA_signal_6059), .A1_f (new_AGEMA_signal_6060), .B0_t (plaintext_s0_t[102]), .B0_f (plaintext_s0_f[102]), .B1_t (plaintext_s1_t[102]), .B1_f (plaintext_s1_f[102]), .Z0_t (stateArray_inS30ser[6]), .Z0_f (new_AGEMA_signal_6856), .Z1_t (new_AGEMA_signal_6857), .Z1_f (new_AGEMA_signal_6858) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS30ser_mux_inst_7_XOR1_U1 ( .A0_t (plaintext_s0_t[103]), .A0_f (plaintext_s0_f[103]), .A1_t (plaintext_s1_t[103]), .A1_f (plaintext_s1_f[103]), .B0_t (ciphertext_s0_t[71]), .B0_f (ciphertext_s0_f[71]), .B1_t (ciphertext_s1_t[71]), .B1_f (ciphertext_s1_f[71]), .Z0_t (stateArray_MUX_inS30ser_mux_inst_7_X), .Z0_f (new_AGEMA_signal_4239), .Z1_t (new_AGEMA_signal_4240), .Z1_f (new_AGEMA_signal_4241) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS30ser_mux_inst_7_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS30ser_mux_inst_7_X), .B0_f (new_AGEMA_signal_4239), .B1_t (new_AGEMA_signal_4240), .B1_f (new_AGEMA_signal_4241), .Z0_t (stateArray_MUX_inS30ser_mux_inst_7_Y), .Z0_f (new_AGEMA_signal_6061), .Z1_t (new_AGEMA_signal_6062), .Z1_f (new_AGEMA_signal_6063) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS30ser_mux_inst_7_XOR2_U1 ( .A0_t (stateArray_MUX_inS30ser_mux_inst_7_Y), .A0_f (new_AGEMA_signal_6061), .A1_t (new_AGEMA_signal_6062), .A1_f (new_AGEMA_signal_6063), .B0_t (plaintext_s0_t[103]), .B0_f (plaintext_s0_f[103]), .B1_t (plaintext_s1_t[103]), .B1_f (plaintext_s1_f[103]), .Z0_t (stateArray_inS30ser[7]), .Z0_f (new_AGEMA_signal_6859), .Z1_t (new_AGEMA_signal_6860), .Z1_f (new_AGEMA_signal_6861) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS31ser_mux_inst_0_XOR1_U1 ( .A0_t (plaintext_s0_t[64]), .A0_f (plaintext_s0_f[64]), .A1_t (plaintext_s1_t[64]), .A1_f (plaintext_s1_f[64]), .B0_t (ciphertext_s0_t[32]), .B0_f (ciphertext_s0_f[32]), .B1_t (ciphertext_s1_t[32]), .B1_f (ciphertext_s1_f[32]), .Z0_t (stateArray_MUX_inS31ser_mux_inst_0_X), .Z0_f (new_AGEMA_signal_4248), .Z1_t (new_AGEMA_signal_4249), .Z1_f (new_AGEMA_signal_4250) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS31ser_mux_inst_0_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS31ser_mux_inst_0_X), .B0_f (new_AGEMA_signal_4248), .B1_t (new_AGEMA_signal_4249), .B1_f (new_AGEMA_signal_4250), .Z0_t (stateArray_MUX_inS31ser_mux_inst_0_Y), .Z0_f (new_AGEMA_signal_6064), .Z1_t (new_AGEMA_signal_6065), .Z1_f (new_AGEMA_signal_6066) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS31ser_mux_inst_0_XOR2_U1 ( .A0_t (stateArray_MUX_inS31ser_mux_inst_0_Y), .A0_f (new_AGEMA_signal_6064), .A1_t (new_AGEMA_signal_6065), .A1_f (new_AGEMA_signal_6066), .B0_t (plaintext_s0_t[64]), .B0_f (plaintext_s0_f[64]), .B1_t (plaintext_s1_t[64]), .B1_f (plaintext_s1_f[64]), .Z0_t (stateArray_inS31ser[0]), .Z0_f (new_AGEMA_signal_6862), .Z1_t (new_AGEMA_signal_6863), .Z1_f (new_AGEMA_signal_6864) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS31ser_mux_inst_1_XOR1_U1 ( .A0_t (plaintext_s0_t[65]), .A0_f (plaintext_s0_f[65]), .A1_t (plaintext_s1_t[65]), .A1_f (plaintext_s1_f[65]), .B0_t (ciphertext_s0_t[33]), .B0_f (ciphertext_s0_f[33]), .B1_t (ciphertext_s1_t[33]), .B1_f (ciphertext_s1_f[33]), .Z0_t (stateArray_MUX_inS31ser_mux_inst_1_X), .Z0_f (new_AGEMA_signal_4257), .Z1_t (new_AGEMA_signal_4258), .Z1_f (new_AGEMA_signal_4259) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS31ser_mux_inst_1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS31ser_mux_inst_1_X), .B0_f (new_AGEMA_signal_4257), .B1_t (new_AGEMA_signal_4258), .B1_f (new_AGEMA_signal_4259), .Z0_t (stateArray_MUX_inS31ser_mux_inst_1_Y), .Z0_f (new_AGEMA_signal_6067), .Z1_t (new_AGEMA_signal_6068), .Z1_f (new_AGEMA_signal_6069) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS31ser_mux_inst_1_XOR2_U1 ( .A0_t (stateArray_MUX_inS31ser_mux_inst_1_Y), .A0_f (new_AGEMA_signal_6067), .A1_t (new_AGEMA_signal_6068), .A1_f (new_AGEMA_signal_6069), .B0_t (plaintext_s0_t[65]), .B0_f (plaintext_s0_f[65]), .B1_t (plaintext_s1_t[65]), .B1_f (plaintext_s1_f[65]), .Z0_t (stateArray_inS31ser[1]), .Z0_f (new_AGEMA_signal_6865), .Z1_t (new_AGEMA_signal_6866), .Z1_f (new_AGEMA_signal_6867) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS31ser_mux_inst_2_XOR1_U1 ( .A0_t (plaintext_s0_t[66]), .A0_f (plaintext_s0_f[66]), .A1_t (plaintext_s1_t[66]), .A1_f (plaintext_s1_f[66]), .B0_t (ciphertext_s0_t[34]), .B0_f (ciphertext_s0_f[34]), .B1_t (ciphertext_s1_t[34]), .B1_f (ciphertext_s1_f[34]), .Z0_t (stateArray_MUX_inS31ser_mux_inst_2_X), .Z0_f (new_AGEMA_signal_4266), .Z1_t (new_AGEMA_signal_4267), .Z1_f (new_AGEMA_signal_4268) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS31ser_mux_inst_2_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS31ser_mux_inst_2_X), .B0_f (new_AGEMA_signal_4266), .B1_t (new_AGEMA_signal_4267), .B1_f (new_AGEMA_signal_4268), .Z0_t (stateArray_MUX_inS31ser_mux_inst_2_Y), .Z0_f (new_AGEMA_signal_6070), .Z1_t (new_AGEMA_signal_6071), .Z1_f (new_AGEMA_signal_6072) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS31ser_mux_inst_2_XOR2_U1 ( .A0_t (stateArray_MUX_inS31ser_mux_inst_2_Y), .A0_f (new_AGEMA_signal_6070), .A1_t (new_AGEMA_signal_6071), .A1_f (new_AGEMA_signal_6072), .B0_t (plaintext_s0_t[66]), .B0_f (plaintext_s0_f[66]), .B1_t (plaintext_s1_t[66]), .B1_f (plaintext_s1_f[66]), .Z0_t (stateArray_inS31ser[2]), .Z0_f (new_AGEMA_signal_6868), .Z1_t (new_AGEMA_signal_6869), .Z1_f (new_AGEMA_signal_6870) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS31ser_mux_inst_3_XOR1_U1 ( .A0_t (plaintext_s0_t[67]), .A0_f (plaintext_s0_f[67]), .A1_t (plaintext_s1_t[67]), .A1_f (plaintext_s1_f[67]), .B0_t (ciphertext_s0_t[35]), .B0_f (ciphertext_s0_f[35]), .B1_t (ciphertext_s1_t[35]), .B1_f (ciphertext_s1_f[35]), .Z0_t (stateArray_MUX_inS31ser_mux_inst_3_X), .Z0_f (new_AGEMA_signal_4275), .Z1_t (new_AGEMA_signal_4276), .Z1_f (new_AGEMA_signal_4277) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS31ser_mux_inst_3_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS31ser_mux_inst_3_X), .B0_f (new_AGEMA_signal_4275), .B1_t (new_AGEMA_signal_4276), .B1_f (new_AGEMA_signal_4277), .Z0_t (stateArray_MUX_inS31ser_mux_inst_3_Y), .Z0_f (new_AGEMA_signal_6073), .Z1_t (new_AGEMA_signal_6074), .Z1_f (new_AGEMA_signal_6075) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS31ser_mux_inst_3_XOR2_U1 ( .A0_t (stateArray_MUX_inS31ser_mux_inst_3_Y), .A0_f (new_AGEMA_signal_6073), .A1_t (new_AGEMA_signal_6074), .A1_f (new_AGEMA_signal_6075), .B0_t (plaintext_s0_t[67]), .B0_f (plaintext_s0_f[67]), .B1_t (plaintext_s1_t[67]), .B1_f (plaintext_s1_f[67]), .Z0_t (stateArray_inS31ser[3]), .Z0_f (new_AGEMA_signal_6871), .Z1_t (new_AGEMA_signal_6872), .Z1_f (new_AGEMA_signal_6873) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS31ser_mux_inst_4_XOR1_U1 ( .A0_t (plaintext_s0_t[68]), .A0_f (plaintext_s0_f[68]), .A1_t (plaintext_s1_t[68]), .A1_f (plaintext_s1_f[68]), .B0_t (ciphertext_s0_t[36]), .B0_f (ciphertext_s0_f[36]), .B1_t (ciphertext_s1_t[36]), .B1_f (ciphertext_s1_f[36]), .Z0_t (stateArray_MUX_inS31ser_mux_inst_4_X), .Z0_f (new_AGEMA_signal_4284), .Z1_t (new_AGEMA_signal_4285), .Z1_f (new_AGEMA_signal_4286) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS31ser_mux_inst_4_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS31ser_mux_inst_4_X), .B0_f (new_AGEMA_signal_4284), .B1_t (new_AGEMA_signal_4285), .B1_f (new_AGEMA_signal_4286), .Z0_t (stateArray_MUX_inS31ser_mux_inst_4_Y), .Z0_f (new_AGEMA_signal_6076), .Z1_t (new_AGEMA_signal_6077), .Z1_f (new_AGEMA_signal_6078) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS31ser_mux_inst_4_XOR2_U1 ( .A0_t (stateArray_MUX_inS31ser_mux_inst_4_Y), .A0_f (new_AGEMA_signal_6076), .A1_t (new_AGEMA_signal_6077), .A1_f (new_AGEMA_signal_6078), .B0_t (plaintext_s0_t[68]), .B0_f (plaintext_s0_f[68]), .B1_t (plaintext_s1_t[68]), .B1_f (plaintext_s1_f[68]), .Z0_t (stateArray_inS31ser[4]), .Z0_f (new_AGEMA_signal_6874), .Z1_t (new_AGEMA_signal_6875), .Z1_f (new_AGEMA_signal_6876) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS31ser_mux_inst_5_XOR1_U1 ( .A0_t (plaintext_s0_t[69]), .A0_f (plaintext_s0_f[69]), .A1_t (plaintext_s1_t[69]), .A1_f (plaintext_s1_f[69]), .B0_t (ciphertext_s0_t[37]), .B0_f (ciphertext_s0_f[37]), .B1_t (ciphertext_s1_t[37]), .B1_f (ciphertext_s1_f[37]), .Z0_t (stateArray_MUX_inS31ser_mux_inst_5_X), .Z0_f (new_AGEMA_signal_4293), .Z1_t (new_AGEMA_signal_4294), .Z1_f (new_AGEMA_signal_4295) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS31ser_mux_inst_5_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS31ser_mux_inst_5_X), .B0_f (new_AGEMA_signal_4293), .B1_t (new_AGEMA_signal_4294), .B1_f (new_AGEMA_signal_4295), .Z0_t (stateArray_MUX_inS31ser_mux_inst_5_Y), .Z0_f (new_AGEMA_signal_6079), .Z1_t (new_AGEMA_signal_6080), .Z1_f (new_AGEMA_signal_6081) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS31ser_mux_inst_5_XOR2_U1 ( .A0_t (stateArray_MUX_inS31ser_mux_inst_5_Y), .A0_f (new_AGEMA_signal_6079), .A1_t (new_AGEMA_signal_6080), .A1_f (new_AGEMA_signal_6081), .B0_t (plaintext_s0_t[69]), .B0_f (plaintext_s0_f[69]), .B1_t (plaintext_s1_t[69]), .B1_f (plaintext_s1_f[69]), .Z0_t (stateArray_inS31ser[5]), .Z0_f (new_AGEMA_signal_6877), .Z1_t (new_AGEMA_signal_6878), .Z1_f (new_AGEMA_signal_6879) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS31ser_mux_inst_6_XOR1_U1 ( .A0_t (plaintext_s0_t[70]), .A0_f (plaintext_s0_f[70]), .A1_t (plaintext_s1_t[70]), .A1_f (plaintext_s1_f[70]), .B0_t (ciphertext_s0_t[38]), .B0_f (ciphertext_s0_f[38]), .B1_t (ciphertext_s1_t[38]), .B1_f (ciphertext_s1_f[38]), .Z0_t (stateArray_MUX_inS31ser_mux_inst_6_X), .Z0_f (new_AGEMA_signal_4302), .Z1_t (new_AGEMA_signal_4303), .Z1_f (new_AGEMA_signal_4304) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS31ser_mux_inst_6_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS31ser_mux_inst_6_X), .B0_f (new_AGEMA_signal_4302), .B1_t (new_AGEMA_signal_4303), .B1_f (new_AGEMA_signal_4304), .Z0_t (stateArray_MUX_inS31ser_mux_inst_6_Y), .Z0_f (new_AGEMA_signal_6082), .Z1_t (new_AGEMA_signal_6083), .Z1_f (new_AGEMA_signal_6084) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS31ser_mux_inst_6_XOR2_U1 ( .A0_t (stateArray_MUX_inS31ser_mux_inst_6_Y), .A0_f (new_AGEMA_signal_6082), .A1_t (new_AGEMA_signal_6083), .A1_f (new_AGEMA_signal_6084), .B0_t (plaintext_s0_t[70]), .B0_f (plaintext_s0_f[70]), .B1_t (plaintext_s1_t[70]), .B1_f (plaintext_s1_f[70]), .Z0_t (stateArray_inS31ser[6]), .Z0_f (new_AGEMA_signal_6880), .Z1_t (new_AGEMA_signal_6881), .Z1_f (new_AGEMA_signal_6882) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS31ser_mux_inst_7_XOR1_U1 ( .A0_t (plaintext_s0_t[71]), .A0_f (plaintext_s0_f[71]), .A1_t (plaintext_s1_t[71]), .A1_f (plaintext_s1_f[71]), .B0_t (ciphertext_s0_t[39]), .B0_f (ciphertext_s0_f[39]), .B1_t (ciphertext_s1_t[39]), .B1_f (ciphertext_s1_f[39]), .Z0_t (stateArray_MUX_inS31ser_mux_inst_7_X), .Z0_f (new_AGEMA_signal_4311), .Z1_t (new_AGEMA_signal_4312), .Z1_f (new_AGEMA_signal_4313) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS31ser_mux_inst_7_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS31ser_mux_inst_7_X), .B0_f (new_AGEMA_signal_4311), .B1_t (new_AGEMA_signal_4312), .B1_f (new_AGEMA_signal_4313), .Z0_t (stateArray_MUX_inS31ser_mux_inst_7_Y), .Z0_f (new_AGEMA_signal_6085), .Z1_t (new_AGEMA_signal_6086), .Z1_f (new_AGEMA_signal_6087) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS31ser_mux_inst_7_XOR2_U1 ( .A0_t (stateArray_MUX_inS31ser_mux_inst_7_Y), .A0_f (new_AGEMA_signal_6085), .A1_t (new_AGEMA_signal_6086), .A1_f (new_AGEMA_signal_6087), .B0_t (plaintext_s0_t[71]), .B0_f (plaintext_s0_f[71]), .B1_t (plaintext_s1_t[71]), .B1_f (plaintext_s1_f[71]), .Z0_t (stateArray_inS31ser[7]), .Z0_f (new_AGEMA_signal_6883), .Z1_t (new_AGEMA_signal_6884), .Z1_f (new_AGEMA_signal_6885) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS32ser_mux_inst_0_XOR1_U1 ( .A0_t (plaintext_s0_t[32]), .A0_f (plaintext_s0_f[32]), .A1_t (plaintext_s1_t[32]), .A1_f (plaintext_s1_f[32]), .B0_t (ciphertext_s0_t[0]), .B0_f (ciphertext_s0_f[0]), .B1_t (ciphertext_s1_t[0]), .B1_f (ciphertext_s1_f[0]), .Z0_t (stateArray_MUX_inS32ser_mux_inst_0_X), .Z0_f (new_AGEMA_signal_4320), .Z1_t (new_AGEMA_signal_4321), .Z1_f (new_AGEMA_signal_4322) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS32ser_mux_inst_0_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS32ser_mux_inst_0_X), .B0_f (new_AGEMA_signal_4320), .B1_t (new_AGEMA_signal_4321), .B1_f (new_AGEMA_signal_4322), .Z0_t (stateArray_MUX_inS32ser_mux_inst_0_Y), .Z0_f (new_AGEMA_signal_6088), .Z1_t (new_AGEMA_signal_6089), .Z1_f (new_AGEMA_signal_6090) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS32ser_mux_inst_0_XOR2_U1 ( .A0_t (stateArray_MUX_inS32ser_mux_inst_0_Y), .A0_f (new_AGEMA_signal_6088), .A1_t (new_AGEMA_signal_6089), .A1_f (new_AGEMA_signal_6090), .B0_t (plaintext_s0_t[32]), .B0_f (plaintext_s0_f[32]), .B1_t (plaintext_s1_t[32]), .B1_f (plaintext_s1_f[32]), .Z0_t (stateArray_inS32ser[0]), .Z0_f (new_AGEMA_signal_6886), .Z1_t (new_AGEMA_signal_6887), .Z1_f (new_AGEMA_signal_6888) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS32ser_mux_inst_1_XOR1_U1 ( .A0_t (plaintext_s0_t[33]), .A0_f (plaintext_s0_f[33]), .A1_t (plaintext_s1_t[33]), .A1_f (plaintext_s1_f[33]), .B0_t (ciphertext_s0_t[1]), .B0_f (ciphertext_s0_f[1]), .B1_t (ciphertext_s1_t[1]), .B1_f (ciphertext_s1_f[1]), .Z0_t (stateArray_MUX_inS32ser_mux_inst_1_X), .Z0_f (new_AGEMA_signal_4329), .Z1_t (new_AGEMA_signal_4330), .Z1_f (new_AGEMA_signal_4331) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS32ser_mux_inst_1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS32ser_mux_inst_1_X), .B0_f (new_AGEMA_signal_4329), .B1_t (new_AGEMA_signal_4330), .B1_f (new_AGEMA_signal_4331), .Z0_t (stateArray_MUX_inS32ser_mux_inst_1_Y), .Z0_f (new_AGEMA_signal_6091), .Z1_t (new_AGEMA_signal_6092), .Z1_f (new_AGEMA_signal_6093) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS32ser_mux_inst_1_XOR2_U1 ( .A0_t (stateArray_MUX_inS32ser_mux_inst_1_Y), .A0_f (new_AGEMA_signal_6091), .A1_t (new_AGEMA_signal_6092), .A1_f (new_AGEMA_signal_6093), .B0_t (plaintext_s0_t[33]), .B0_f (plaintext_s0_f[33]), .B1_t (plaintext_s1_t[33]), .B1_f (plaintext_s1_f[33]), .Z0_t (stateArray_inS32ser[1]), .Z0_f (new_AGEMA_signal_6889), .Z1_t (new_AGEMA_signal_6890), .Z1_f (new_AGEMA_signal_6891) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS32ser_mux_inst_2_XOR1_U1 ( .A0_t (plaintext_s0_t[34]), .A0_f (plaintext_s0_f[34]), .A1_t (plaintext_s1_t[34]), .A1_f (plaintext_s1_f[34]), .B0_t (ciphertext_s0_t[2]), .B0_f (ciphertext_s0_f[2]), .B1_t (ciphertext_s1_t[2]), .B1_f (ciphertext_s1_f[2]), .Z0_t (stateArray_MUX_inS32ser_mux_inst_2_X), .Z0_f (new_AGEMA_signal_4338), .Z1_t (new_AGEMA_signal_4339), .Z1_f (new_AGEMA_signal_4340) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS32ser_mux_inst_2_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS32ser_mux_inst_2_X), .B0_f (new_AGEMA_signal_4338), .B1_t (new_AGEMA_signal_4339), .B1_f (new_AGEMA_signal_4340), .Z0_t (stateArray_MUX_inS32ser_mux_inst_2_Y), .Z0_f (new_AGEMA_signal_6094), .Z1_t (new_AGEMA_signal_6095), .Z1_f (new_AGEMA_signal_6096) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS32ser_mux_inst_2_XOR2_U1 ( .A0_t (stateArray_MUX_inS32ser_mux_inst_2_Y), .A0_f (new_AGEMA_signal_6094), .A1_t (new_AGEMA_signal_6095), .A1_f (new_AGEMA_signal_6096), .B0_t (plaintext_s0_t[34]), .B0_f (plaintext_s0_f[34]), .B1_t (plaintext_s1_t[34]), .B1_f (plaintext_s1_f[34]), .Z0_t (stateArray_inS32ser[2]), .Z0_f (new_AGEMA_signal_6892), .Z1_t (new_AGEMA_signal_6893), .Z1_f (new_AGEMA_signal_6894) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS32ser_mux_inst_3_XOR1_U1 ( .A0_t (plaintext_s0_t[35]), .A0_f (plaintext_s0_f[35]), .A1_t (plaintext_s1_t[35]), .A1_f (plaintext_s1_f[35]), .B0_t (ciphertext_s0_t[3]), .B0_f (ciphertext_s0_f[3]), .B1_t (ciphertext_s1_t[3]), .B1_f (ciphertext_s1_f[3]), .Z0_t (stateArray_MUX_inS32ser_mux_inst_3_X), .Z0_f (new_AGEMA_signal_4347), .Z1_t (new_AGEMA_signal_4348), .Z1_f (new_AGEMA_signal_4349) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS32ser_mux_inst_3_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS32ser_mux_inst_3_X), .B0_f (new_AGEMA_signal_4347), .B1_t (new_AGEMA_signal_4348), .B1_f (new_AGEMA_signal_4349), .Z0_t (stateArray_MUX_inS32ser_mux_inst_3_Y), .Z0_f (new_AGEMA_signal_6097), .Z1_t (new_AGEMA_signal_6098), .Z1_f (new_AGEMA_signal_6099) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS32ser_mux_inst_3_XOR2_U1 ( .A0_t (stateArray_MUX_inS32ser_mux_inst_3_Y), .A0_f (new_AGEMA_signal_6097), .A1_t (new_AGEMA_signal_6098), .A1_f (new_AGEMA_signal_6099), .B0_t (plaintext_s0_t[35]), .B0_f (plaintext_s0_f[35]), .B1_t (plaintext_s1_t[35]), .B1_f (plaintext_s1_f[35]), .Z0_t (stateArray_inS32ser[3]), .Z0_f (new_AGEMA_signal_6895), .Z1_t (new_AGEMA_signal_6896), .Z1_f (new_AGEMA_signal_6897) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS32ser_mux_inst_4_XOR1_U1 ( .A0_t (plaintext_s0_t[36]), .A0_f (plaintext_s0_f[36]), .A1_t (plaintext_s1_t[36]), .A1_f (plaintext_s1_f[36]), .B0_t (ciphertext_s0_t[4]), .B0_f (ciphertext_s0_f[4]), .B1_t (ciphertext_s1_t[4]), .B1_f (ciphertext_s1_f[4]), .Z0_t (stateArray_MUX_inS32ser_mux_inst_4_X), .Z0_f (new_AGEMA_signal_4356), .Z1_t (new_AGEMA_signal_4357), .Z1_f (new_AGEMA_signal_4358) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS32ser_mux_inst_4_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS32ser_mux_inst_4_X), .B0_f (new_AGEMA_signal_4356), .B1_t (new_AGEMA_signal_4357), .B1_f (new_AGEMA_signal_4358), .Z0_t (stateArray_MUX_inS32ser_mux_inst_4_Y), .Z0_f (new_AGEMA_signal_6100), .Z1_t (new_AGEMA_signal_6101), .Z1_f (new_AGEMA_signal_6102) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS32ser_mux_inst_4_XOR2_U1 ( .A0_t (stateArray_MUX_inS32ser_mux_inst_4_Y), .A0_f (new_AGEMA_signal_6100), .A1_t (new_AGEMA_signal_6101), .A1_f (new_AGEMA_signal_6102), .B0_t (plaintext_s0_t[36]), .B0_f (plaintext_s0_f[36]), .B1_t (plaintext_s1_t[36]), .B1_f (plaintext_s1_f[36]), .Z0_t (stateArray_inS32ser[4]), .Z0_f (new_AGEMA_signal_6898), .Z1_t (new_AGEMA_signal_6899), .Z1_f (new_AGEMA_signal_6900) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS32ser_mux_inst_5_XOR1_U1 ( .A0_t (plaintext_s0_t[37]), .A0_f (plaintext_s0_f[37]), .A1_t (plaintext_s1_t[37]), .A1_f (plaintext_s1_f[37]), .B0_t (ciphertext_s0_t[5]), .B0_f (ciphertext_s0_f[5]), .B1_t (ciphertext_s1_t[5]), .B1_f (ciphertext_s1_f[5]), .Z0_t (stateArray_MUX_inS32ser_mux_inst_5_X), .Z0_f (new_AGEMA_signal_4365), .Z1_t (new_AGEMA_signal_4366), .Z1_f (new_AGEMA_signal_4367) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS32ser_mux_inst_5_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS32ser_mux_inst_5_X), .B0_f (new_AGEMA_signal_4365), .B1_t (new_AGEMA_signal_4366), .B1_f (new_AGEMA_signal_4367), .Z0_t (stateArray_MUX_inS32ser_mux_inst_5_Y), .Z0_f (new_AGEMA_signal_6103), .Z1_t (new_AGEMA_signal_6104), .Z1_f (new_AGEMA_signal_6105) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS32ser_mux_inst_5_XOR2_U1 ( .A0_t (stateArray_MUX_inS32ser_mux_inst_5_Y), .A0_f (new_AGEMA_signal_6103), .A1_t (new_AGEMA_signal_6104), .A1_f (new_AGEMA_signal_6105), .B0_t (plaintext_s0_t[37]), .B0_f (plaintext_s0_f[37]), .B1_t (plaintext_s1_t[37]), .B1_f (plaintext_s1_f[37]), .Z0_t (stateArray_inS32ser[5]), .Z0_f (new_AGEMA_signal_6901), .Z1_t (new_AGEMA_signal_6902), .Z1_f (new_AGEMA_signal_6903) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS32ser_mux_inst_6_XOR1_U1 ( .A0_t (plaintext_s0_t[38]), .A0_f (plaintext_s0_f[38]), .A1_t (plaintext_s1_t[38]), .A1_f (plaintext_s1_f[38]), .B0_t (ciphertext_s0_t[6]), .B0_f (ciphertext_s0_f[6]), .B1_t (ciphertext_s1_t[6]), .B1_f (ciphertext_s1_f[6]), .Z0_t (stateArray_MUX_inS32ser_mux_inst_6_X), .Z0_f (new_AGEMA_signal_4374), .Z1_t (new_AGEMA_signal_4375), .Z1_f (new_AGEMA_signal_4376) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS32ser_mux_inst_6_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS32ser_mux_inst_6_X), .B0_f (new_AGEMA_signal_4374), .B1_t (new_AGEMA_signal_4375), .B1_f (new_AGEMA_signal_4376), .Z0_t (stateArray_MUX_inS32ser_mux_inst_6_Y), .Z0_f (new_AGEMA_signal_6106), .Z1_t (new_AGEMA_signal_6107), .Z1_f (new_AGEMA_signal_6108) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS32ser_mux_inst_6_XOR2_U1 ( .A0_t (stateArray_MUX_inS32ser_mux_inst_6_Y), .A0_f (new_AGEMA_signal_6106), .A1_t (new_AGEMA_signal_6107), .A1_f (new_AGEMA_signal_6108), .B0_t (plaintext_s0_t[38]), .B0_f (plaintext_s0_f[38]), .B1_t (plaintext_s1_t[38]), .B1_f (plaintext_s1_f[38]), .Z0_t (stateArray_inS32ser[6]), .Z0_f (new_AGEMA_signal_6904), .Z1_t (new_AGEMA_signal_6905), .Z1_f (new_AGEMA_signal_6906) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS32ser_mux_inst_7_XOR1_U1 ( .A0_t (plaintext_s0_t[39]), .A0_f (plaintext_s0_f[39]), .A1_t (plaintext_s1_t[39]), .A1_f (plaintext_s1_f[39]), .B0_t (ciphertext_s0_t[7]), .B0_f (ciphertext_s0_f[7]), .B1_t (ciphertext_s1_t[7]), .B1_f (ciphertext_s1_f[7]), .Z0_t (stateArray_MUX_inS32ser_mux_inst_7_X), .Z0_f (new_AGEMA_signal_4383), .Z1_t (new_AGEMA_signal_4384), .Z1_f (new_AGEMA_signal_4385) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS32ser_mux_inst_7_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS32ser_mux_inst_7_X), .B0_f (new_AGEMA_signal_4383), .B1_t (new_AGEMA_signal_4384), .B1_f (new_AGEMA_signal_4385), .Z0_t (stateArray_MUX_inS32ser_mux_inst_7_Y), .Z0_f (new_AGEMA_signal_6109), .Z1_t (new_AGEMA_signal_6110), .Z1_f (new_AGEMA_signal_6111) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS32ser_mux_inst_7_XOR2_U1 ( .A0_t (stateArray_MUX_inS32ser_mux_inst_7_Y), .A0_f (new_AGEMA_signal_6109), .A1_t (new_AGEMA_signal_6110), .A1_f (new_AGEMA_signal_6111), .B0_t (plaintext_s0_t[39]), .B0_f (plaintext_s0_f[39]), .B1_t (plaintext_s1_t[39]), .B1_f (plaintext_s1_f[39]), .Z0_t (stateArray_inS32ser[7]), .Z0_f (new_AGEMA_signal_6907), .Z1_t (new_AGEMA_signal_6908), .Z1_f (new_AGEMA_signal_6909) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_0_XOR1_U1 ( .A0_t (StateIn[0]), .A0_f (new_AGEMA_signal_11399), .A1_t (new_AGEMA_signal_11400), .A1_f (new_AGEMA_signal_11401), .B0_t (StateInMC[0]), .B0_f (new_AGEMA_signal_9304), .B1_t (new_AGEMA_signal_9305), .B1_f (new_AGEMA_signal_9306), .Z0_t (stateArray_MUX_input_MC_mux_inst_0_X), .Z0_f (new_AGEMA_signal_11468), .Z1_t (new_AGEMA_signal_11469), .Z1_f (new_AGEMA_signal_11470) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_0_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (stateArray_MUX_input_MC_mux_inst_0_X), .B0_f (new_AGEMA_signal_11468), .B1_t (new_AGEMA_signal_11469), .B1_f (new_AGEMA_signal_11470), .Z0_t (stateArray_MUX_input_MC_mux_inst_0_Y), .Z0_f (new_AGEMA_signal_11495), .Z1_t (new_AGEMA_signal_11496), .Z1_f (new_AGEMA_signal_11497) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_0_XOR2_U1 ( .A0_t (stateArray_MUX_input_MC_mux_inst_0_Y), .A0_f (new_AGEMA_signal_11495), .A1_t (new_AGEMA_signal_11496), .A1_f (new_AGEMA_signal_11497), .B0_t (StateIn[0]), .B0_f (new_AGEMA_signal_11399), .B1_t (new_AGEMA_signal_11400), .B1_f (new_AGEMA_signal_11401), .Z0_t (stateArray_input_MC[0]), .Z0_f (new_AGEMA_signal_11543), .Z1_t (new_AGEMA_signal_11544), .Z1_f (new_AGEMA_signal_11545) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_1_XOR1_U1 ( .A0_t (StateIn[1]), .A0_f (new_AGEMA_signal_11447), .A1_t (new_AGEMA_signal_11448), .A1_f (new_AGEMA_signal_11449), .B0_t (StateInMC[1]), .B0_f (new_AGEMA_signal_9840), .B1_t (new_AGEMA_signal_9841), .B1_f (new_AGEMA_signal_9842), .Z0_t (stateArray_MUX_input_MC_mux_inst_1_X), .Z0_f (new_AGEMA_signal_11498), .Z1_t (new_AGEMA_signal_11499), .Z1_f (new_AGEMA_signal_11500) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (stateArray_MUX_input_MC_mux_inst_1_X), .B0_f (new_AGEMA_signal_11498), .B1_t (new_AGEMA_signal_11499), .B1_f (new_AGEMA_signal_11500), .Z0_t (stateArray_MUX_input_MC_mux_inst_1_Y), .Z0_f (new_AGEMA_signal_11546), .Z1_t (new_AGEMA_signal_11547), .Z1_f (new_AGEMA_signal_11548) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_1_XOR2_U1 ( .A0_t (stateArray_MUX_input_MC_mux_inst_1_Y), .A0_f (new_AGEMA_signal_11546), .A1_t (new_AGEMA_signal_11547), .A1_f (new_AGEMA_signal_11548), .B0_t (StateIn[1]), .B0_f (new_AGEMA_signal_11447), .B1_t (new_AGEMA_signal_11448), .B1_f (new_AGEMA_signal_11449), .Z0_t (stateArray_input_MC[1]), .Z0_f (new_AGEMA_signal_11591), .Z1_t (new_AGEMA_signal_11592), .Z1_f (new_AGEMA_signal_11593) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_2_XOR1_U1 ( .A0_t (StateIn[2]), .A0_f (new_AGEMA_signal_11450), .A1_t (new_AGEMA_signal_11451), .A1_f (new_AGEMA_signal_11452), .B0_t (StateInMC[2]), .B0_f (new_AGEMA_signal_9310), .B1_t (new_AGEMA_signal_9311), .B1_f (new_AGEMA_signal_9312), .Z0_t (stateArray_MUX_input_MC_mux_inst_2_X), .Z0_f (new_AGEMA_signal_11501), .Z1_t (new_AGEMA_signal_11502), .Z1_f (new_AGEMA_signal_11503) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_2_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (stateArray_MUX_input_MC_mux_inst_2_X), .B0_f (new_AGEMA_signal_11501), .B1_t (new_AGEMA_signal_11502), .B1_f (new_AGEMA_signal_11503), .Z0_t (stateArray_MUX_input_MC_mux_inst_2_Y), .Z0_f (new_AGEMA_signal_11549), .Z1_t (new_AGEMA_signal_11550), .Z1_f (new_AGEMA_signal_11551) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_2_XOR2_U1 ( .A0_t (stateArray_MUX_input_MC_mux_inst_2_Y), .A0_f (new_AGEMA_signal_11549), .A1_t (new_AGEMA_signal_11550), .A1_f (new_AGEMA_signal_11551), .B0_t (StateIn[2]), .B0_f (new_AGEMA_signal_11450), .B1_t (new_AGEMA_signal_11451), .B1_f (new_AGEMA_signal_11452), .Z0_t (stateArray_input_MC[2]), .Z0_f (new_AGEMA_signal_11594), .Z1_t (new_AGEMA_signal_11595), .Z1_f (new_AGEMA_signal_11596) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_3_XOR1_U1 ( .A0_t (StateIn[3]), .A0_f (new_AGEMA_signal_11453), .A1_t (new_AGEMA_signal_11454), .A1_f (new_AGEMA_signal_11455), .B0_t (StateInMC[3]), .B0_f (new_AGEMA_signal_9843), .B1_t (new_AGEMA_signal_9844), .B1_f (new_AGEMA_signal_9845), .Z0_t (stateArray_MUX_input_MC_mux_inst_3_X), .Z0_f (new_AGEMA_signal_11504), .Z1_t (new_AGEMA_signal_11505), .Z1_f (new_AGEMA_signal_11506) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_3_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (stateArray_MUX_input_MC_mux_inst_3_X), .B0_f (new_AGEMA_signal_11504), .B1_t (new_AGEMA_signal_11505), .B1_f (new_AGEMA_signal_11506), .Z0_t (stateArray_MUX_input_MC_mux_inst_3_Y), .Z0_f (new_AGEMA_signal_11552), .Z1_t (new_AGEMA_signal_11553), .Z1_f (new_AGEMA_signal_11554) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_3_XOR2_U1 ( .A0_t (stateArray_MUX_input_MC_mux_inst_3_Y), .A0_f (new_AGEMA_signal_11552), .A1_t (new_AGEMA_signal_11553), .A1_f (new_AGEMA_signal_11554), .B0_t (StateIn[3]), .B0_f (new_AGEMA_signal_11453), .B1_t (new_AGEMA_signal_11454), .B1_f (new_AGEMA_signal_11455), .Z0_t (stateArray_input_MC[3]), .Z0_f (new_AGEMA_signal_11597), .Z1_t (new_AGEMA_signal_11598), .Z1_f (new_AGEMA_signal_11599) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_4_XOR1_U1 ( .A0_t (StateIn[4]), .A0_f (new_AGEMA_signal_11456), .A1_t (new_AGEMA_signal_11457), .A1_f (new_AGEMA_signal_11458), .B0_t (StateInMC[4]), .B0_f (new_AGEMA_signal_9846), .B1_t (new_AGEMA_signal_9847), .B1_f (new_AGEMA_signal_9848), .Z0_t (stateArray_MUX_input_MC_mux_inst_4_X), .Z0_f (new_AGEMA_signal_11507), .Z1_t (new_AGEMA_signal_11508), .Z1_f (new_AGEMA_signal_11509) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_4_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (stateArray_MUX_input_MC_mux_inst_4_X), .B0_f (new_AGEMA_signal_11507), .B1_t (new_AGEMA_signal_11508), .B1_f (new_AGEMA_signal_11509), .Z0_t (stateArray_MUX_input_MC_mux_inst_4_Y), .Z0_f (new_AGEMA_signal_11555), .Z1_t (new_AGEMA_signal_11556), .Z1_f (new_AGEMA_signal_11557) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_4_XOR2_U1 ( .A0_t (stateArray_MUX_input_MC_mux_inst_4_Y), .A0_f (new_AGEMA_signal_11555), .A1_t (new_AGEMA_signal_11556), .A1_f (new_AGEMA_signal_11557), .B0_t (StateIn[4]), .B0_f (new_AGEMA_signal_11456), .B1_t (new_AGEMA_signal_11457), .B1_f (new_AGEMA_signal_11458), .Z0_t (stateArray_input_MC[4]), .Z0_f (new_AGEMA_signal_11600), .Z1_t (new_AGEMA_signal_11601), .Z1_f (new_AGEMA_signal_11602) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_5_XOR1_U1 ( .A0_t (StateIn[5]), .A0_f (new_AGEMA_signal_11459), .A1_t (new_AGEMA_signal_11460), .A1_f (new_AGEMA_signal_11461), .B0_t (StateInMC[5]), .B0_f (new_AGEMA_signal_9319), .B1_t (new_AGEMA_signal_9320), .B1_f (new_AGEMA_signal_9321), .Z0_t (stateArray_MUX_input_MC_mux_inst_5_X), .Z0_f (new_AGEMA_signal_11510), .Z1_t (new_AGEMA_signal_11511), .Z1_f (new_AGEMA_signal_11512) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_5_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (stateArray_MUX_input_MC_mux_inst_5_X), .B0_f (new_AGEMA_signal_11510), .B1_t (new_AGEMA_signal_11511), .B1_f (new_AGEMA_signal_11512), .Z0_t (stateArray_MUX_input_MC_mux_inst_5_Y), .Z0_f (new_AGEMA_signal_11558), .Z1_t (new_AGEMA_signal_11559), .Z1_f (new_AGEMA_signal_11560) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_5_XOR2_U1 ( .A0_t (stateArray_MUX_input_MC_mux_inst_5_Y), .A0_f (new_AGEMA_signal_11558), .A1_t (new_AGEMA_signal_11559), .A1_f (new_AGEMA_signal_11560), .B0_t (StateIn[5]), .B0_f (new_AGEMA_signal_11459), .B1_t (new_AGEMA_signal_11460), .B1_f (new_AGEMA_signal_11461), .Z0_t (stateArray_input_MC[5]), .Z0_f (new_AGEMA_signal_11603), .Z1_t (new_AGEMA_signal_11604), .Z1_f (new_AGEMA_signal_11605) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_6_XOR1_U1 ( .A0_t (StateIn[6]), .A0_f (new_AGEMA_signal_11462), .A1_t (new_AGEMA_signal_11463), .A1_f (new_AGEMA_signal_11464), .B0_t (StateInMC[6]), .B0_f (new_AGEMA_signal_9322), .B1_t (new_AGEMA_signal_9323), .B1_f (new_AGEMA_signal_9324), .Z0_t (stateArray_MUX_input_MC_mux_inst_6_X), .Z0_f (new_AGEMA_signal_11513), .Z1_t (new_AGEMA_signal_11514), .Z1_f (new_AGEMA_signal_11515) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_6_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (stateArray_MUX_input_MC_mux_inst_6_X), .B0_f (new_AGEMA_signal_11513), .B1_t (new_AGEMA_signal_11514), .B1_f (new_AGEMA_signal_11515), .Z0_t (stateArray_MUX_input_MC_mux_inst_6_Y), .Z0_f (new_AGEMA_signal_11561), .Z1_t (new_AGEMA_signal_11562), .Z1_f (new_AGEMA_signal_11563) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_6_XOR2_U1 ( .A0_t (stateArray_MUX_input_MC_mux_inst_6_Y), .A0_f (new_AGEMA_signal_11561), .A1_t (new_AGEMA_signal_11562), .A1_f (new_AGEMA_signal_11563), .B0_t (StateIn[6]), .B0_f (new_AGEMA_signal_11462), .B1_t (new_AGEMA_signal_11463), .B1_f (new_AGEMA_signal_11464), .Z0_t (stateArray_input_MC[6]), .Z0_f (new_AGEMA_signal_11606), .Z1_t (new_AGEMA_signal_11607), .Z1_f (new_AGEMA_signal_11608) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_7_XOR1_U1 ( .A0_t (StateIn[7]), .A0_f (new_AGEMA_signal_11465), .A1_t (new_AGEMA_signal_11466), .A1_f (new_AGEMA_signal_11467), .B0_t (StateInMC[7]), .B0_f (new_AGEMA_signal_9325), .B1_t (new_AGEMA_signal_9326), .B1_f (new_AGEMA_signal_9327), .Z0_t (stateArray_MUX_input_MC_mux_inst_7_X), .Z0_f (new_AGEMA_signal_11516), .Z1_t (new_AGEMA_signal_11517), .Z1_f (new_AGEMA_signal_11518) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_7_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (stateArray_MUX_input_MC_mux_inst_7_X), .B0_f (new_AGEMA_signal_11516), .B1_t (new_AGEMA_signal_11517), .B1_f (new_AGEMA_signal_11518), .Z0_t (stateArray_MUX_input_MC_mux_inst_7_Y), .Z0_f (new_AGEMA_signal_11564), .Z1_t (new_AGEMA_signal_11565), .Z1_f (new_AGEMA_signal_11566) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_7_XOR2_U1 ( .A0_t (stateArray_MUX_input_MC_mux_inst_7_Y), .A0_f (new_AGEMA_signal_11564), .A1_t (new_AGEMA_signal_11565), .A1_f (new_AGEMA_signal_11566), .B0_t (StateIn[7]), .B0_f (new_AGEMA_signal_11465), .B1_t (new_AGEMA_signal_11466), .B1_f (new_AGEMA_signal_11467), .Z0_t (stateArray_input_MC[7]), .Z0_f (new_AGEMA_signal_11609), .Z1_t (new_AGEMA_signal_11610), .Z1_f (new_AGEMA_signal_11611) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_0_XOR1_U1 ( .A0_t (plaintext_s0_t[0]), .A0_f (plaintext_s0_f[0]), .A1_t (plaintext_s1_t[0]), .A1_f (plaintext_s1_f[0]), .B0_t (stateArray_input_MC[0]), .B0_f (new_AGEMA_signal_11543), .B1_t (new_AGEMA_signal_11544), .B1_f (new_AGEMA_signal_11545), .Z0_t (stateArray_MUX_inS33ser_mux_inst_0_X), .Z0_f (new_AGEMA_signal_11615), .Z1_t (new_AGEMA_signal_11616), .Z1_f (new_AGEMA_signal_11617) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_0_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS33ser_mux_inst_0_X), .B0_f (new_AGEMA_signal_11615), .B1_t (new_AGEMA_signal_11616), .B1_f (new_AGEMA_signal_11617), .Z0_t (stateArray_MUX_inS33ser_mux_inst_0_Y), .Z0_f (new_AGEMA_signal_11639), .Z1_t (new_AGEMA_signal_11640), .Z1_f (new_AGEMA_signal_11641) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_0_XOR2_U1 ( .A0_t (stateArray_MUX_inS33ser_mux_inst_0_Y), .A0_f (new_AGEMA_signal_11639), .A1_t (new_AGEMA_signal_11640), .A1_f (new_AGEMA_signal_11641), .B0_t (plaintext_s0_t[0]), .B0_f (plaintext_s0_f[0]), .B1_t (plaintext_s1_t[0]), .B1_f (plaintext_s1_f[0]), .Z0_t (stateArray_inS33ser[0]), .Z0_f (new_AGEMA_signal_11684), .Z1_t (new_AGEMA_signal_11685), .Z1_f (new_AGEMA_signal_11686) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_1_XOR1_U1 ( .A0_t (plaintext_s0_t[1]), .A0_f (plaintext_s0_f[1]), .A1_t (plaintext_s1_t[1]), .A1_f (plaintext_s1_f[1]), .B0_t (stateArray_input_MC[1]), .B0_f (new_AGEMA_signal_11591), .B1_t (new_AGEMA_signal_11592), .B1_f (new_AGEMA_signal_11593), .Z0_t (stateArray_MUX_inS33ser_mux_inst_1_X), .Z0_f (new_AGEMA_signal_11645), .Z1_t (new_AGEMA_signal_11646), .Z1_f (new_AGEMA_signal_11647) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS33ser_mux_inst_1_X), .B0_f (new_AGEMA_signal_11645), .B1_t (new_AGEMA_signal_11646), .B1_f (new_AGEMA_signal_11647), .Z0_t (stateArray_MUX_inS33ser_mux_inst_1_Y), .Z0_f (new_AGEMA_signal_11687), .Z1_t (new_AGEMA_signal_11688), .Z1_f (new_AGEMA_signal_11689) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_1_XOR2_U1 ( .A0_t (stateArray_MUX_inS33ser_mux_inst_1_Y), .A0_f (new_AGEMA_signal_11687), .A1_t (new_AGEMA_signal_11688), .A1_f (new_AGEMA_signal_11689), .B0_t (plaintext_s0_t[1]), .B0_f (plaintext_s0_f[1]), .B1_t (plaintext_s1_t[1]), .B1_f (plaintext_s1_f[1]), .Z0_t (stateArray_inS33ser[1]), .Z0_f (new_AGEMA_signal_11711), .Z1_t (new_AGEMA_signal_11712), .Z1_f (new_AGEMA_signal_11713) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_2_XOR1_U1 ( .A0_t (plaintext_s0_t[2]), .A0_f (plaintext_s0_f[2]), .A1_t (plaintext_s1_t[2]), .A1_f (plaintext_s1_f[2]), .B0_t (stateArray_input_MC[2]), .B0_f (new_AGEMA_signal_11594), .B1_t (new_AGEMA_signal_11595), .B1_f (new_AGEMA_signal_11596), .Z0_t (stateArray_MUX_inS33ser_mux_inst_2_X), .Z0_f (new_AGEMA_signal_11651), .Z1_t (new_AGEMA_signal_11652), .Z1_f (new_AGEMA_signal_11653) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_2_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS33ser_mux_inst_2_X), .B0_f (new_AGEMA_signal_11651), .B1_t (new_AGEMA_signal_11652), .B1_f (new_AGEMA_signal_11653), .Z0_t (stateArray_MUX_inS33ser_mux_inst_2_Y), .Z0_f (new_AGEMA_signal_11690), .Z1_t (new_AGEMA_signal_11691), .Z1_f (new_AGEMA_signal_11692) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_2_XOR2_U1 ( .A0_t (stateArray_MUX_inS33ser_mux_inst_2_Y), .A0_f (new_AGEMA_signal_11690), .A1_t (new_AGEMA_signal_11691), .A1_f (new_AGEMA_signal_11692), .B0_t (plaintext_s0_t[2]), .B0_f (plaintext_s0_f[2]), .B1_t (plaintext_s1_t[2]), .B1_f (plaintext_s1_f[2]), .Z0_t (stateArray_inS33ser[2]), .Z0_f (new_AGEMA_signal_11714), .Z1_t (new_AGEMA_signal_11715), .Z1_f (new_AGEMA_signal_11716) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_3_XOR1_U1 ( .A0_t (plaintext_s0_t[3]), .A0_f (plaintext_s0_f[3]), .A1_t (plaintext_s1_t[3]), .A1_f (plaintext_s1_f[3]), .B0_t (stateArray_input_MC[3]), .B0_f (new_AGEMA_signal_11597), .B1_t (new_AGEMA_signal_11598), .B1_f (new_AGEMA_signal_11599), .Z0_t (stateArray_MUX_inS33ser_mux_inst_3_X), .Z0_f (new_AGEMA_signal_11657), .Z1_t (new_AGEMA_signal_11658), .Z1_f (new_AGEMA_signal_11659) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_3_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS33ser_mux_inst_3_X), .B0_f (new_AGEMA_signal_11657), .B1_t (new_AGEMA_signal_11658), .B1_f (new_AGEMA_signal_11659), .Z0_t (stateArray_MUX_inS33ser_mux_inst_3_Y), .Z0_f (new_AGEMA_signal_11693), .Z1_t (new_AGEMA_signal_11694), .Z1_f (new_AGEMA_signal_11695) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_3_XOR2_U1 ( .A0_t (stateArray_MUX_inS33ser_mux_inst_3_Y), .A0_f (new_AGEMA_signal_11693), .A1_t (new_AGEMA_signal_11694), .A1_f (new_AGEMA_signal_11695), .B0_t (plaintext_s0_t[3]), .B0_f (plaintext_s0_f[3]), .B1_t (plaintext_s1_t[3]), .B1_f (plaintext_s1_f[3]), .Z0_t (stateArray_inS33ser[3]), .Z0_f (new_AGEMA_signal_11717), .Z1_t (new_AGEMA_signal_11718), .Z1_f (new_AGEMA_signal_11719) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_4_XOR1_U1 ( .A0_t (plaintext_s0_t[4]), .A0_f (plaintext_s0_f[4]), .A1_t (plaintext_s1_t[4]), .A1_f (plaintext_s1_f[4]), .B0_t (stateArray_input_MC[4]), .B0_f (new_AGEMA_signal_11600), .B1_t (new_AGEMA_signal_11601), .B1_f (new_AGEMA_signal_11602), .Z0_t (stateArray_MUX_inS33ser_mux_inst_4_X), .Z0_f (new_AGEMA_signal_11663), .Z1_t (new_AGEMA_signal_11664), .Z1_f (new_AGEMA_signal_11665) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_4_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS33ser_mux_inst_4_X), .B0_f (new_AGEMA_signal_11663), .B1_t (new_AGEMA_signal_11664), .B1_f (new_AGEMA_signal_11665), .Z0_t (stateArray_MUX_inS33ser_mux_inst_4_Y), .Z0_f (new_AGEMA_signal_11696), .Z1_t (new_AGEMA_signal_11697), .Z1_f (new_AGEMA_signal_11698) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_4_XOR2_U1 ( .A0_t (stateArray_MUX_inS33ser_mux_inst_4_Y), .A0_f (new_AGEMA_signal_11696), .A1_t (new_AGEMA_signal_11697), .A1_f (new_AGEMA_signal_11698), .B0_t (plaintext_s0_t[4]), .B0_f (plaintext_s0_f[4]), .B1_t (plaintext_s1_t[4]), .B1_f (plaintext_s1_f[4]), .Z0_t (stateArray_inS33ser[4]), .Z0_f (new_AGEMA_signal_11720), .Z1_t (new_AGEMA_signal_11721), .Z1_f (new_AGEMA_signal_11722) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_5_XOR1_U1 ( .A0_t (plaintext_s0_t[5]), .A0_f (plaintext_s0_f[5]), .A1_t (plaintext_s1_t[5]), .A1_f (plaintext_s1_f[5]), .B0_t (stateArray_input_MC[5]), .B0_f (new_AGEMA_signal_11603), .B1_t (new_AGEMA_signal_11604), .B1_f (new_AGEMA_signal_11605), .Z0_t (stateArray_MUX_inS33ser_mux_inst_5_X), .Z0_f (new_AGEMA_signal_11669), .Z1_t (new_AGEMA_signal_11670), .Z1_f (new_AGEMA_signal_11671) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_5_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS33ser_mux_inst_5_X), .B0_f (new_AGEMA_signal_11669), .B1_t (new_AGEMA_signal_11670), .B1_f (new_AGEMA_signal_11671), .Z0_t (stateArray_MUX_inS33ser_mux_inst_5_Y), .Z0_f (new_AGEMA_signal_11699), .Z1_t (new_AGEMA_signal_11700), .Z1_f (new_AGEMA_signal_11701) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_5_XOR2_U1 ( .A0_t (stateArray_MUX_inS33ser_mux_inst_5_Y), .A0_f (new_AGEMA_signal_11699), .A1_t (new_AGEMA_signal_11700), .A1_f (new_AGEMA_signal_11701), .B0_t (plaintext_s0_t[5]), .B0_f (plaintext_s0_f[5]), .B1_t (plaintext_s1_t[5]), .B1_f (plaintext_s1_f[5]), .Z0_t (stateArray_inS33ser[5]), .Z0_f (new_AGEMA_signal_11723), .Z1_t (new_AGEMA_signal_11724), .Z1_f (new_AGEMA_signal_11725) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_6_XOR1_U1 ( .A0_t (plaintext_s0_t[6]), .A0_f (plaintext_s0_f[6]), .A1_t (plaintext_s1_t[6]), .A1_f (plaintext_s1_f[6]), .B0_t (stateArray_input_MC[6]), .B0_f (new_AGEMA_signal_11606), .B1_t (new_AGEMA_signal_11607), .B1_f (new_AGEMA_signal_11608), .Z0_t (stateArray_MUX_inS33ser_mux_inst_6_X), .Z0_f (new_AGEMA_signal_11675), .Z1_t (new_AGEMA_signal_11676), .Z1_f (new_AGEMA_signal_11677) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_6_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS33ser_mux_inst_6_X), .B0_f (new_AGEMA_signal_11675), .B1_t (new_AGEMA_signal_11676), .B1_f (new_AGEMA_signal_11677), .Z0_t (stateArray_MUX_inS33ser_mux_inst_6_Y), .Z0_f (new_AGEMA_signal_11702), .Z1_t (new_AGEMA_signal_11703), .Z1_f (new_AGEMA_signal_11704) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_6_XOR2_U1 ( .A0_t (stateArray_MUX_inS33ser_mux_inst_6_Y), .A0_f (new_AGEMA_signal_11702), .A1_t (new_AGEMA_signal_11703), .A1_f (new_AGEMA_signal_11704), .B0_t (plaintext_s0_t[6]), .B0_f (plaintext_s0_f[6]), .B1_t (plaintext_s1_t[6]), .B1_f (plaintext_s1_f[6]), .Z0_t (stateArray_inS33ser[6]), .Z0_f (new_AGEMA_signal_11726), .Z1_t (new_AGEMA_signal_11727), .Z1_f (new_AGEMA_signal_11728) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_7_XOR1_U1 ( .A0_t (plaintext_s0_t[7]), .A0_f (plaintext_s0_f[7]), .A1_t (plaintext_s1_t[7]), .A1_f (plaintext_s1_f[7]), .B0_t (stateArray_input_MC[7]), .B0_f (new_AGEMA_signal_11609), .B1_t (new_AGEMA_signal_11610), .B1_f (new_AGEMA_signal_11611), .Z0_t (stateArray_MUX_inS33ser_mux_inst_7_X), .Z0_f (new_AGEMA_signal_11681), .Z1_t (new_AGEMA_signal_11682), .Z1_f (new_AGEMA_signal_11683) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_7_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (stateArray_MUX_inS33ser_mux_inst_7_X), .B0_f (new_AGEMA_signal_11681), .B1_t (new_AGEMA_signal_11682), .B1_f (new_AGEMA_signal_11683), .Z0_t (stateArray_MUX_inS33ser_mux_inst_7_Y), .Z0_f (new_AGEMA_signal_11705), .Z1_t (new_AGEMA_signal_11706), .Z1_f (new_AGEMA_signal_11707) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_7_XOR2_U1 ( .A0_t (stateArray_MUX_inS33ser_mux_inst_7_Y), .A0_f (new_AGEMA_signal_11705), .A1_t (new_AGEMA_signal_11706), .A1_f (new_AGEMA_signal_11707), .B0_t (plaintext_s0_t[7]), .B0_f (plaintext_s0_f[7]), .B1_t (plaintext_s1_t[7]), .B1_f (plaintext_s1_f[7]), .Z0_t (stateArray_inS33ser[7]), .Z0_f (new_AGEMA_signal_11729), .Z1_t (new_AGEMA_signal_11730), .Z1_f (new_AGEMA_signal_11731) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_0_XOR1_U1 ( .A0_t (MCout[0]), .A0_f (new_AGEMA_signal_7363), .A1_t (new_AGEMA_signal_7364), .A1_f (new_AGEMA_signal_7365), .B0_t (ciphertext_s0_t[96]), .B0_f (ciphertext_s0_f[96]), .B1_t (ciphertext_s1_t[96]), .B1_f (ciphertext_s1_f[96]), .Z0_t (MUX_StateInMC_mux_inst_0_X), .Z0_f (new_AGEMA_signal_7683), .Z1_t (new_AGEMA_signal_7684), .Z1_f (new_AGEMA_signal_7685) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_0_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_6594), .B0_t (MUX_StateInMC_mux_inst_0_X), .B0_f (new_AGEMA_signal_7683), .B1_t (new_AGEMA_signal_7684), .B1_f (new_AGEMA_signal_7685), .Z0_t (MUX_StateInMC_mux_inst_0_Y), .Z0_f (new_AGEMA_signal_8430), .Z1_t (new_AGEMA_signal_8431), .Z1_f (new_AGEMA_signal_8432) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_0_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_0_Y), .A0_f (new_AGEMA_signal_8430), .A1_t (new_AGEMA_signal_8431), .A1_f (new_AGEMA_signal_8432), .B0_t (MCout[0]), .B0_f (new_AGEMA_signal_7363), .B1_t (new_AGEMA_signal_7364), .B1_f (new_AGEMA_signal_7365), .Z0_t (StateInMC[0]), .Z0_f (new_AGEMA_signal_9304), .Z1_t (new_AGEMA_signal_9305), .Z1_f (new_AGEMA_signal_9306) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_1_XOR1_U1 ( .A0_t (MCout[1]), .A0_f (new_AGEMA_signal_8112), .A1_t (new_AGEMA_signal_8113), .A1_f (new_AGEMA_signal_8114), .B0_t (ciphertext_s0_t[97]), .B0_f (ciphertext_s0_f[97]), .B1_t (ciphertext_s1_t[97]), .B1_f (ciphertext_s1_f[97]), .Z0_t (MUX_StateInMC_mux_inst_1_X), .Z0_f (new_AGEMA_signal_8433), .Z1_t (new_AGEMA_signal_8434), .Z1_f (new_AGEMA_signal_8435) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_6594), .B0_t (MUX_StateInMC_mux_inst_1_X), .B0_f (new_AGEMA_signal_8433), .B1_t (new_AGEMA_signal_8434), .B1_f (new_AGEMA_signal_8435), .Z0_t (MUX_StateInMC_mux_inst_1_Y), .Z0_f (new_AGEMA_signal_9307), .Z1_t (new_AGEMA_signal_9308), .Z1_f (new_AGEMA_signal_9309) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_1_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_1_Y), .A0_f (new_AGEMA_signal_9307), .A1_t (new_AGEMA_signal_9308), .A1_f (new_AGEMA_signal_9309), .B0_t (MCout[1]), .B0_f (new_AGEMA_signal_8112), .B1_t (new_AGEMA_signal_8113), .B1_f (new_AGEMA_signal_8114), .Z0_t (StateInMC[1]), .Z0_f (new_AGEMA_signal_9840), .Z1_t (new_AGEMA_signal_9841), .Z1_f (new_AGEMA_signal_9842) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_2_XOR1_U1 ( .A0_t (MCout[2]), .A0_f (new_AGEMA_signal_7357), .A1_t (new_AGEMA_signal_7358), .A1_f (new_AGEMA_signal_7359), .B0_t (ciphertext_s0_t[98]), .B0_f (ciphertext_s0_f[98]), .B1_t (ciphertext_s1_t[98]), .B1_f (ciphertext_s1_f[98]), .Z0_t (MUX_StateInMC_mux_inst_2_X), .Z0_f (new_AGEMA_signal_7686), .Z1_t (new_AGEMA_signal_7687), .Z1_f (new_AGEMA_signal_7688) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_2_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_6594), .B0_t (MUX_StateInMC_mux_inst_2_X), .B0_f (new_AGEMA_signal_7686), .B1_t (new_AGEMA_signal_7687), .B1_f (new_AGEMA_signal_7688), .Z0_t (MUX_StateInMC_mux_inst_2_Y), .Z0_f (new_AGEMA_signal_8436), .Z1_t (new_AGEMA_signal_8437), .Z1_f (new_AGEMA_signal_8438) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_2_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_2_Y), .A0_f (new_AGEMA_signal_8436), .A1_t (new_AGEMA_signal_8437), .A1_f (new_AGEMA_signal_8438), .B0_t (MCout[2]), .B0_f (new_AGEMA_signal_7357), .B1_t (new_AGEMA_signal_7358), .B1_f (new_AGEMA_signal_7359), .Z0_t (StateInMC[2]), .Z0_f (new_AGEMA_signal_9310), .Z1_t (new_AGEMA_signal_9311), .Z1_f (new_AGEMA_signal_9312) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_3_XOR1_U1 ( .A0_t (MCout[3]), .A0_f (new_AGEMA_signal_8109), .A1_t (new_AGEMA_signal_8110), .A1_f (new_AGEMA_signal_8111), .B0_t (ciphertext_s0_t[99]), .B0_f (ciphertext_s0_f[99]), .B1_t (ciphertext_s1_t[99]), .B1_f (ciphertext_s1_f[99]), .Z0_t (MUX_StateInMC_mux_inst_3_X), .Z0_f (new_AGEMA_signal_8439), .Z1_t (new_AGEMA_signal_8440), .Z1_f (new_AGEMA_signal_8441) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_3_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_6594), .B0_t (MUX_StateInMC_mux_inst_3_X), .B0_f (new_AGEMA_signal_8439), .B1_t (new_AGEMA_signal_8440), .B1_f (new_AGEMA_signal_8441), .Z0_t (MUX_StateInMC_mux_inst_3_Y), .Z0_f (new_AGEMA_signal_9313), .Z1_t (new_AGEMA_signal_9314), .Z1_f (new_AGEMA_signal_9315) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_3_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_3_Y), .A0_f (new_AGEMA_signal_9313), .A1_t (new_AGEMA_signal_9314), .A1_f (new_AGEMA_signal_9315), .B0_t (MCout[3]), .B0_f (new_AGEMA_signal_8109), .B1_t (new_AGEMA_signal_8110), .B1_f (new_AGEMA_signal_8111), .Z0_t (StateInMC[3]), .Z0_f (new_AGEMA_signal_9843), .Z1_t (new_AGEMA_signal_9844), .Z1_f (new_AGEMA_signal_9845) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_4_XOR1_U1 ( .A0_t (MCout[4]), .A0_f (new_AGEMA_signal_8106), .A1_t (new_AGEMA_signal_8107), .A1_f (new_AGEMA_signal_8108), .B0_t (ciphertext_s0_t[100]), .B0_f (ciphertext_s0_f[100]), .B1_t (ciphertext_s1_t[100]), .B1_f (ciphertext_s1_f[100]), .Z0_t (MUX_StateInMC_mux_inst_4_X), .Z0_f (new_AGEMA_signal_8442), .Z1_t (new_AGEMA_signal_8443), .Z1_f (new_AGEMA_signal_8444) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_4_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_6594), .B0_t (MUX_StateInMC_mux_inst_4_X), .B0_f (new_AGEMA_signal_8442), .B1_t (new_AGEMA_signal_8443), .B1_f (new_AGEMA_signal_8444), .Z0_t (MUX_StateInMC_mux_inst_4_Y), .Z0_f (new_AGEMA_signal_9316), .Z1_t (new_AGEMA_signal_9317), .Z1_f (new_AGEMA_signal_9318) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_4_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_4_Y), .A0_f (new_AGEMA_signal_9316), .A1_t (new_AGEMA_signal_9317), .A1_f (new_AGEMA_signal_9318), .B0_t (MCout[4]), .B0_f (new_AGEMA_signal_8106), .B1_t (new_AGEMA_signal_8107), .B1_f (new_AGEMA_signal_8108), .Z0_t (StateInMC[4]), .Z0_f (new_AGEMA_signal_9846), .Z1_t (new_AGEMA_signal_9847), .Z1_f (new_AGEMA_signal_9848) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_5_XOR1_U1 ( .A0_t (MCout[5]), .A0_f (new_AGEMA_signal_7348), .A1_t (new_AGEMA_signal_7349), .A1_f (new_AGEMA_signal_7350), .B0_t (ciphertext_s0_t[101]), .B0_f (ciphertext_s0_f[101]), .B1_t (ciphertext_s1_t[101]), .B1_f (ciphertext_s1_f[101]), .Z0_t (MUX_StateInMC_mux_inst_5_X), .Z0_f (new_AGEMA_signal_7689), .Z1_t (new_AGEMA_signal_7690), .Z1_f (new_AGEMA_signal_7691) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_5_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_6594), .B0_t (MUX_StateInMC_mux_inst_5_X), .B0_f (new_AGEMA_signal_7689), .B1_t (new_AGEMA_signal_7690), .B1_f (new_AGEMA_signal_7691), .Z0_t (MUX_StateInMC_mux_inst_5_Y), .Z0_f (new_AGEMA_signal_8445), .Z1_t (new_AGEMA_signal_8446), .Z1_f (new_AGEMA_signal_8447) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_5_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_5_Y), .A0_f (new_AGEMA_signal_8445), .A1_t (new_AGEMA_signal_8446), .A1_f (new_AGEMA_signal_8447), .B0_t (MCout[5]), .B0_f (new_AGEMA_signal_7348), .B1_t (new_AGEMA_signal_7349), .B1_f (new_AGEMA_signal_7350), .Z0_t (StateInMC[5]), .Z0_f (new_AGEMA_signal_9319), .Z1_t (new_AGEMA_signal_9320), .Z1_f (new_AGEMA_signal_9321) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_6_XOR1_U1 ( .A0_t (MCout[6]), .A0_f (new_AGEMA_signal_7345), .A1_t (new_AGEMA_signal_7346), .A1_f (new_AGEMA_signal_7347), .B0_t (ciphertext_s0_t[102]), .B0_f (ciphertext_s0_f[102]), .B1_t (ciphertext_s1_t[102]), .B1_f (ciphertext_s1_f[102]), .Z0_t (MUX_StateInMC_mux_inst_6_X), .Z0_f (new_AGEMA_signal_7692), .Z1_t (new_AGEMA_signal_7693), .Z1_f (new_AGEMA_signal_7694) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_6_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_6594), .B0_t (MUX_StateInMC_mux_inst_6_X), .B0_f (new_AGEMA_signal_7692), .B1_t (new_AGEMA_signal_7693), .B1_f (new_AGEMA_signal_7694), .Z0_t (MUX_StateInMC_mux_inst_6_Y), .Z0_f (new_AGEMA_signal_8448), .Z1_t (new_AGEMA_signal_8449), .Z1_f (new_AGEMA_signal_8450) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_6_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_6_Y), .A0_f (new_AGEMA_signal_8448), .A1_t (new_AGEMA_signal_8449), .A1_f (new_AGEMA_signal_8450), .B0_t (MCout[6]), .B0_f (new_AGEMA_signal_7345), .B1_t (new_AGEMA_signal_7346), .B1_f (new_AGEMA_signal_7347), .Z0_t (StateInMC[6]), .Z0_f (new_AGEMA_signal_9322), .Z1_t (new_AGEMA_signal_9323), .Z1_f (new_AGEMA_signal_9324) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_7_XOR1_U1 ( .A0_t (MCout[7]), .A0_f (new_AGEMA_signal_7342), .A1_t (new_AGEMA_signal_7343), .A1_f (new_AGEMA_signal_7344), .B0_t (ciphertext_s0_t[103]), .B0_f (ciphertext_s0_f[103]), .B1_t (ciphertext_s1_t[103]), .B1_f (ciphertext_s1_f[103]), .Z0_t (MUX_StateInMC_mux_inst_7_X), .Z0_f (new_AGEMA_signal_7695), .Z1_t (new_AGEMA_signal_7696), .Z1_f (new_AGEMA_signal_7697) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_7_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_6594), .B0_t (MUX_StateInMC_mux_inst_7_X), .B0_f (new_AGEMA_signal_7695), .B1_t (new_AGEMA_signal_7696), .B1_f (new_AGEMA_signal_7697), .Z0_t (MUX_StateInMC_mux_inst_7_Y), .Z0_f (new_AGEMA_signal_8451), .Z1_t (new_AGEMA_signal_8452), .Z1_f (new_AGEMA_signal_8453) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_7_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_7_Y), .A0_f (new_AGEMA_signal_8451), .A1_t (new_AGEMA_signal_8452), .A1_f (new_AGEMA_signal_8453), .B0_t (MCout[7]), .B0_f (new_AGEMA_signal_7342), .B1_t (new_AGEMA_signal_7343), .B1_f (new_AGEMA_signal_7344), .Z0_t (StateInMC[7]), .Z0_f (new_AGEMA_signal_9325), .Z1_t (new_AGEMA_signal_9326), .Z1_f (new_AGEMA_signal_9327) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_8_XOR1_U1 ( .A0_t (MCout[8]), .A0_f (new_AGEMA_signal_7339), .A1_t (new_AGEMA_signal_7340), .A1_f (new_AGEMA_signal_7341), .B0_t (ciphertext_s0_t[104]), .B0_f (ciphertext_s0_f[104]), .B1_t (ciphertext_s1_t[104]), .B1_f (ciphertext_s1_f[104]), .Z0_t (MUX_StateInMC_mux_inst_8_X), .Z0_f (new_AGEMA_signal_7698), .Z1_t (new_AGEMA_signal_7699), .Z1_f (new_AGEMA_signal_7700) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_8_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_6594), .B0_t (MUX_StateInMC_mux_inst_8_X), .B0_f (new_AGEMA_signal_7698), .B1_t (new_AGEMA_signal_7699), .B1_f (new_AGEMA_signal_7700), .Z0_t (MUX_StateInMC_mux_inst_8_Y), .Z0_f (new_AGEMA_signal_8454), .Z1_t (new_AGEMA_signal_8455), .Z1_f (new_AGEMA_signal_8456) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_8_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_8_Y), .A0_f (new_AGEMA_signal_8454), .A1_t (new_AGEMA_signal_8455), .A1_f (new_AGEMA_signal_8456), .B0_t (MCout[8]), .B0_f (new_AGEMA_signal_7339), .B1_t (new_AGEMA_signal_7340), .B1_f (new_AGEMA_signal_7341), .Z0_t (StateInMC[8]), .Z0_f (new_AGEMA_signal_9328), .Z1_t (new_AGEMA_signal_9329), .Z1_f (new_AGEMA_signal_9330) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_9_XOR1_U1 ( .A0_t (MCout[9]), .A0_f (new_AGEMA_signal_8103), .A1_t (new_AGEMA_signal_8104), .A1_f (new_AGEMA_signal_8105), .B0_t (ciphertext_s0_t[105]), .B0_f (ciphertext_s0_f[105]), .B1_t (ciphertext_s1_t[105]), .B1_f (ciphertext_s1_f[105]), .Z0_t (MUX_StateInMC_mux_inst_9_X), .Z0_f (new_AGEMA_signal_8457), .Z1_t (new_AGEMA_signal_8458), .Z1_f (new_AGEMA_signal_8459) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_9_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_6594), .B0_t (MUX_StateInMC_mux_inst_9_X), .B0_f (new_AGEMA_signal_8457), .B1_t (new_AGEMA_signal_8458), .B1_f (new_AGEMA_signal_8459), .Z0_t (MUX_StateInMC_mux_inst_9_Y), .Z0_f (new_AGEMA_signal_9331), .Z1_t (new_AGEMA_signal_9332), .Z1_f (new_AGEMA_signal_9333) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_9_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_9_Y), .A0_f (new_AGEMA_signal_9331), .A1_t (new_AGEMA_signal_9332), .A1_f (new_AGEMA_signal_9333), .B0_t (MCout[9]), .B0_f (new_AGEMA_signal_8103), .B1_t (new_AGEMA_signal_8104), .B1_f (new_AGEMA_signal_8105), .Z0_t (StateInMC[9]), .Z0_f (new_AGEMA_signal_9849), .Z1_t (new_AGEMA_signal_9850), .Z1_f (new_AGEMA_signal_9851) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_10_XOR1_U1 ( .A0_t (MCout[10]), .A0_f (new_AGEMA_signal_7333), .A1_t (new_AGEMA_signal_7334), .A1_f (new_AGEMA_signal_7335), .B0_t (ciphertext_s0_t[106]), .B0_f (ciphertext_s0_f[106]), .B1_t (ciphertext_s1_t[106]), .B1_f (ciphertext_s1_f[106]), .Z0_t (MUX_StateInMC_mux_inst_10_X), .Z0_f (new_AGEMA_signal_7701), .Z1_t (new_AGEMA_signal_7702), .Z1_f (new_AGEMA_signal_7703) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_10_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_6594), .B0_t (MUX_StateInMC_mux_inst_10_X), .B0_f (new_AGEMA_signal_7701), .B1_t (new_AGEMA_signal_7702), .B1_f (new_AGEMA_signal_7703), .Z0_t (MUX_StateInMC_mux_inst_10_Y), .Z0_f (new_AGEMA_signal_8460), .Z1_t (new_AGEMA_signal_8461), .Z1_f (new_AGEMA_signal_8462) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_10_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_10_Y), .A0_f (new_AGEMA_signal_8460), .A1_t (new_AGEMA_signal_8461), .A1_f (new_AGEMA_signal_8462), .B0_t (MCout[10]), .B0_f (new_AGEMA_signal_7333), .B1_t (new_AGEMA_signal_7334), .B1_f (new_AGEMA_signal_7335), .Z0_t (StateInMC[10]), .Z0_f (new_AGEMA_signal_9334), .Z1_t (new_AGEMA_signal_9335), .Z1_f (new_AGEMA_signal_9336) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_11_XOR1_U1 ( .A0_t (MCout[11]), .A0_f (new_AGEMA_signal_8100), .A1_t (new_AGEMA_signal_8101), .A1_f (new_AGEMA_signal_8102), .B0_t (ciphertext_s0_t[107]), .B0_f (ciphertext_s0_f[107]), .B1_t (ciphertext_s1_t[107]), .B1_f (ciphertext_s1_f[107]), .Z0_t (MUX_StateInMC_mux_inst_11_X), .Z0_f (new_AGEMA_signal_8463), .Z1_t (new_AGEMA_signal_8464), .Z1_f (new_AGEMA_signal_8465) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_11_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_6594), .B0_t (MUX_StateInMC_mux_inst_11_X), .B0_f (new_AGEMA_signal_8463), .B1_t (new_AGEMA_signal_8464), .B1_f (new_AGEMA_signal_8465), .Z0_t (MUX_StateInMC_mux_inst_11_Y), .Z0_f (new_AGEMA_signal_9337), .Z1_t (new_AGEMA_signal_9338), .Z1_f (new_AGEMA_signal_9339) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_11_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_11_Y), .A0_f (new_AGEMA_signal_9337), .A1_t (new_AGEMA_signal_9338), .A1_f (new_AGEMA_signal_9339), .B0_t (MCout[11]), .B0_f (new_AGEMA_signal_8100), .B1_t (new_AGEMA_signal_8101), .B1_f (new_AGEMA_signal_8102), .Z0_t (StateInMC[11]), .Z0_f (new_AGEMA_signal_9852), .Z1_t (new_AGEMA_signal_9853), .Z1_f (new_AGEMA_signal_9854) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_12_XOR1_U1 ( .A0_t (MCout[12]), .A0_f (new_AGEMA_signal_8097), .A1_t (new_AGEMA_signal_8098), .A1_f (new_AGEMA_signal_8099), .B0_t (ciphertext_s0_t[108]), .B0_f (ciphertext_s0_f[108]), .B1_t (ciphertext_s1_t[108]), .B1_f (ciphertext_s1_f[108]), .Z0_t (MUX_StateInMC_mux_inst_12_X), .Z0_f (new_AGEMA_signal_8466), .Z1_t (new_AGEMA_signal_8467), .Z1_f (new_AGEMA_signal_8468) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_12_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_6594), .B0_t (MUX_StateInMC_mux_inst_12_X), .B0_f (new_AGEMA_signal_8466), .B1_t (new_AGEMA_signal_8467), .B1_f (new_AGEMA_signal_8468), .Z0_t (MUX_StateInMC_mux_inst_12_Y), .Z0_f (new_AGEMA_signal_9340), .Z1_t (new_AGEMA_signal_9341), .Z1_f (new_AGEMA_signal_9342) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_12_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_12_Y), .A0_f (new_AGEMA_signal_9340), .A1_t (new_AGEMA_signal_9341), .A1_f (new_AGEMA_signal_9342), .B0_t (MCout[12]), .B0_f (new_AGEMA_signal_8097), .B1_t (new_AGEMA_signal_8098), .B1_f (new_AGEMA_signal_8099), .Z0_t (StateInMC[12]), .Z0_f (new_AGEMA_signal_9855), .Z1_t (new_AGEMA_signal_9856), .Z1_f (new_AGEMA_signal_9857) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_13_XOR1_U1 ( .A0_t (MCout[13]), .A0_f (new_AGEMA_signal_7324), .A1_t (new_AGEMA_signal_7325), .A1_f (new_AGEMA_signal_7326), .B0_t (ciphertext_s0_t[109]), .B0_f (ciphertext_s0_f[109]), .B1_t (ciphertext_s1_t[109]), .B1_f (ciphertext_s1_f[109]), .Z0_t (MUX_StateInMC_mux_inst_13_X), .Z0_f (new_AGEMA_signal_7704), .Z1_t (new_AGEMA_signal_7705), .Z1_f (new_AGEMA_signal_7706) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_13_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_6594), .B0_t (MUX_StateInMC_mux_inst_13_X), .B0_f (new_AGEMA_signal_7704), .B1_t (new_AGEMA_signal_7705), .B1_f (new_AGEMA_signal_7706), .Z0_t (MUX_StateInMC_mux_inst_13_Y), .Z0_f (new_AGEMA_signal_8469), .Z1_t (new_AGEMA_signal_8470), .Z1_f (new_AGEMA_signal_8471) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_13_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_13_Y), .A0_f (new_AGEMA_signal_8469), .A1_t (new_AGEMA_signal_8470), .A1_f (new_AGEMA_signal_8471), .B0_t (MCout[13]), .B0_f (new_AGEMA_signal_7324), .B1_t (new_AGEMA_signal_7325), .B1_f (new_AGEMA_signal_7326), .Z0_t (StateInMC[13]), .Z0_f (new_AGEMA_signal_9343), .Z1_t (new_AGEMA_signal_9344), .Z1_f (new_AGEMA_signal_9345) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_14_XOR1_U1 ( .A0_t (MCout[14]), .A0_f (new_AGEMA_signal_7321), .A1_t (new_AGEMA_signal_7322), .A1_f (new_AGEMA_signal_7323), .B0_t (ciphertext_s0_t[110]), .B0_f (ciphertext_s0_f[110]), .B1_t (ciphertext_s1_t[110]), .B1_f (ciphertext_s1_f[110]), .Z0_t (MUX_StateInMC_mux_inst_14_X), .Z0_f (new_AGEMA_signal_7707), .Z1_t (new_AGEMA_signal_7708), .Z1_f (new_AGEMA_signal_7709) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_14_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_6594), .B0_t (MUX_StateInMC_mux_inst_14_X), .B0_f (new_AGEMA_signal_7707), .B1_t (new_AGEMA_signal_7708), .B1_f (new_AGEMA_signal_7709), .Z0_t (MUX_StateInMC_mux_inst_14_Y), .Z0_f (new_AGEMA_signal_8472), .Z1_t (new_AGEMA_signal_8473), .Z1_f (new_AGEMA_signal_8474) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_14_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_14_Y), .A0_f (new_AGEMA_signal_8472), .A1_t (new_AGEMA_signal_8473), .A1_f (new_AGEMA_signal_8474), .B0_t (MCout[14]), .B0_f (new_AGEMA_signal_7321), .B1_t (new_AGEMA_signal_7322), .B1_f (new_AGEMA_signal_7323), .Z0_t (StateInMC[14]), .Z0_f (new_AGEMA_signal_9346), .Z1_t (new_AGEMA_signal_9347), .Z1_f (new_AGEMA_signal_9348) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_15_XOR1_U1 ( .A0_t (MCout[15]), .A0_f (new_AGEMA_signal_7318), .A1_t (new_AGEMA_signal_7319), .A1_f (new_AGEMA_signal_7320), .B0_t (ciphertext_s0_t[111]), .B0_f (ciphertext_s0_f[111]), .B1_t (ciphertext_s1_t[111]), .B1_f (ciphertext_s1_f[111]), .Z0_t (MUX_StateInMC_mux_inst_15_X), .Z0_f (new_AGEMA_signal_7710), .Z1_t (new_AGEMA_signal_7711), .Z1_f (new_AGEMA_signal_7712) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_15_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_6594), .B0_t (MUX_StateInMC_mux_inst_15_X), .B0_f (new_AGEMA_signal_7710), .B1_t (new_AGEMA_signal_7711), .B1_f (new_AGEMA_signal_7712), .Z0_t (MUX_StateInMC_mux_inst_15_Y), .Z0_f (new_AGEMA_signal_8475), .Z1_t (new_AGEMA_signal_8476), .Z1_f (new_AGEMA_signal_8477) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_15_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_15_Y), .A0_f (new_AGEMA_signal_8475), .A1_t (new_AGEMA_signal_8476), .A1_f (new_AGEMA_signal_8477), .B0_t (MCout[15]), .B0_f (new_AGEMA_signal_7318), .B1_t (new_AGEMA_signal_7319), .B1_f (new_AGEMA_signal_7320), .Z0_t (StateInMC[15]), .Z0_f (new_AGEMA_signal_9349), .Z1_t (new_AGEMA_signal_9350), .Z1_f (new_AGEMA_signal_9351) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_16_XOR1_U1 ( .A0_t (MCout[16]), .A0_f (new_AGEMA_signal_7315), .A1_t (new_AGEMA_signal_7316), .A1_f (new_AGEMA_signal_7317), .B0_t (ciphertext_s0_t[112]), .B0_f (ciphertext_s0_f[112]), .B1_t (ciphertext_s1_t[112]), .B1_f (ciphertext_s1_f[112]), .Z0_t (MUX_StateInMC_mux_inst_16_X), .Z0_f (new_AGEMA_signal_7713), .Z1_t (new_AGEMA_signal_7714), .Z1_f (new_AGEMA_signal_7715) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_16_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_6594), .B0_t (MUX_StateInMC_mux_inst_16_X), .B0_f (new_AGEMA_signal_7713), .B1_t (new_AGEMA_signal_7714), .B1_f (new_AGEMA_signal_7715), .Z0_t (MUX_StateInMC_mux_inst_16_Y), .Z0_f (new_AGEMA_signal_8478), .Z1_t (new_AGEMA_signal_8479), .Z1_f (new_AGEMA_signal_8480) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_16_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_16_Y), .A0_f (new_AGEMA_signal_8478), .A1_t (new_AGEMA_signal_8479), .A1_f (new_AGEMA_signal_8480), .B0_t (MCout[16]), .B0_f (new_AGEMA_signal_7315), .B1_t (new_AGEMA_signal_7316), .B1_f (new_AGEMA_signal_7317), .Z0_t (StateInMC[16]), .Z0_f (new_AGEMA_signal_9352), .Z1_t (new_AGEMA_signal_9353), .Z1_f (new_AGEMA_signal_9354) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_17_XOR1_U1 ( .A0_t (MCout[17]), .A0_f (new_AGEMA_signal_8094), .A1_t (new_AGEMA_signal_8095), .A1_f (new_AGEMA_signal_8096), .B0_t (ciphertext_s0_t[113]), .B0_f (ciphertext_s0_f[113]), .B1_t (ciphertext_s1_t[113]), .B1_f (ciphertext_s1_f[113]), .Z0_t (MUX_StateInMC_mux_inst_17_X), .Z0_f (new_AGEMA_signal_8481), .Z1_t (new_AGEMA_signal_8482), .Z1_f (new_AGEMA_signal_8483) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_17_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_6594), .B0_t (MUX_StateInMC_mux_inst_17_X), .B0_f (new_AGEMA_signal_8481), .B1_t (new_AGEMA_signal_8482), .B1_f (new_AGEMA_signal_8483), .Z0_t (MUX_StateInMC_mux_inst_17_Y), .Z0_f (new_AGEMA_signal_9355), .Z1_t (new_AGEMA_signal_9356), .Z1_f (new_AGEMA_signal_9357) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_17_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_17_Y), .A0_f (new_AGEMA_signal_9355), .A1_t (new_AGEMA_signal_9356), .A1_f (new_AGEMA_signal_9357), .B0_t (MCout[17]), .B0_f (new_AGEMA_signal_8094), .B1_t (new_AGEMA_signal_8095), .B1_f (new_AGEMA_signal_8096), .Z0_t (StateInMC[17]), .Z0_f (new_AGEMA_signal_9858), .Z1_t (new_AGEMA_signal_9859), .Z1_f (new_AGEMA_signal_9860) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_18_XOR1_U1 ( .A0_t (MCout[18]), .A0_f (new_AGEMA_signal_7309), .A1_t (new_AGEMA_signal_7310), .A1_f (new_AGEMA_signal_7311), .B0_t (ciphertext_s0_t[114]), .B0_f (ciphertext_s0_f[114]), .B1_t (ciphertext_s1_t[114]), .B1_f (ciphertext_s1_f[114]), .Z0_t (MUX_StateInMC_mux_inst_18_X), .Z0_f (new_AGEMA_signal_7716), .Z1_t (new_AGEMA_signal_7717), .Z1_f (new_AGEMA_signal_7718) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_18_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_6594), .B0_t (MUX_StateInMC_mux_inst_18_X), .B0_f (new_AGEMA_signal_7716), .B1_t (new_AGEMA_signal_7717), .B1_f (new_AGEMA_signal_7718), .Z0_t (MUX_StateInMC_mux_inst_18_Y), .Z0_f (new_AGEMA_signal_8484), .Z1_t (new_AGEMA_signal_8485), .Z1_f (new_AGEMA_signal_8486) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_18_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_18_Y), .A0_f (new_AGEMA_signal_8484), .A1_t (new_AGEMA_signal_8485), .A1_f (new_AGEMA_signal_8486), .B0_t (MCout[18]), .B0_f (new_AGEMA_signal_7309), .B1_t (new_AGEMA_signal_7310), .B1_f (new_AGEMA_signal_7311), .Z0_t (StateInMC[18]), .Z0_f (new_AGEMA_signal_9358), .Z1_t (new_AGEMA_signal_9359), .Z1_f (new_AGEMA_signal_9360) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_19_XOR1_U1 ( .A0_t (MCout[19]), .A0_f (new_AGEMA_signal_8091), .A1_t (new_AGEMA_signal_8092), .A1_f (new_AGEMA_signal_8093), .B0_t (ciphertext_s0_t[115]), .B0_f (ciphertext_s0_f[115]), .B1_t (ciphertext_s1_t[115]), .B1_f (ciphertext_s1_f[115]), .Z0_t (MUX_StateInMC_mux_inst_19_X), .Z0_f (new_AGEMA_signal_8487), .Z1_t (new_AGEMA_signal_8488), .Z1_f (new_AGEMA_signal_8489) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_19_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_6594), .B0_t (MUX_StateInMC_mux_inst_19_X), .B0_f (new_AGEMA_signal_8487), .B1_t (new_AGEMA_signal_8488), .B1_f (new_AGEMA_signal_8489), .Z0_t (MUX_StateInMC_mux_inst_19_Y), .Z0_f (new_AGEMA_signal_9361), .Z1_t (new_AGEMA_signal_9362), .Z1_f (new_AGEMA_signal_9363) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_19_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_19_Y), .A0_f (new_AGEMA_signal_9361), .A1_t (new_AGEMA_signal_9362), .A1_f (new_AGEMA_signal_9363), .B0_t (MCout[19]), .B0_f (new_AGEMA_signal_8091), .B1_t (new_AGEMA_signal_8092), .B1_f (new_AGEMA_signal_8093), .Z0_t (StateInMC[19]), .Z0_f (new_AGEMA_signal_9861), .Z1_t (new_AGEMA_signal_9862), .Z1_f (new_AGEMA_signal_9863) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_20_XOR1_U1 ( .A0_t (MCout[20]), .A0_f (new_AGEMA_signal_8088), .A1_t (new_AGEMA_signal_8089), .A1_f (new_AGEMA_signal_8090), .B0_t (ciphertext_s0_t[116]), .B0_f (ciphertext_s0_f[116]), .B1_t (ciphertext_s1_t[116]), .B1_f (ciphertext_s1_f[116]), .Z0_t (MUX_StateInMC_mux_inst_20_X), .Z0_f (new_AGEMA_signal_8490), .Z1_t (new_AGEMA_signal_8491), .Z1_f (new_AGEMA_signal_8492) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_20_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_6594), .B0_t (MUX_StateInMC_mux_inst_20_X), .B0_f (new_AGEMA_signal_8490), .B1_t (new_AGEMA_signal_8491), .B1_f (new_AGEMA_signal_8492), .Z0_t (MUX_StateInMC_mux_inst_20_Y), .Z0_f (new_AGEMA_signal_9364), .Z1_t (new_AGEMA_signal_9365), .Z1_f (new_AGEMA_signal_9366) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_20_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_20_Y), .A0_f (new_AGEMA_signal_9364), .A1_t (new_AGEMA_signal_9365), .A1_f (new_AGEMA_signal_9366), .B0_t (MCout[20]), .B0_f (new_AGEMA_signal_8088), .B1_t (new_AGEMA_signal_8089), .B1_f (new_AGEMA_signal_8090), .Z0_t (StateInMC[20]), .Z0_f (new_AGEMA_signal_9864), .Z1_t (new_AGEMA_signal_9865), .Z1_f (new_AGEMA_signal_9866) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_21_XOR1_U1 ( .A0_t (MCout[21]), .A0_f (new_AGEMA_signal_7300), .A1_t (new_AGEMA_signal_7301), .A1_f (new_AGEMA_signal_7302), .B0_t (ciphertext_s0_t[117]), .B0_f (ciphertext_s0_f[117]), .B1_t (ciphertext_s1_t[117]), .B1_f (ciphertext_s1_f[117]), .Z0_t (MUX_StateInMC_mux_inst_21_X), .Z0_f (new_AGEMA_signal_7719), .Z1_t (new_AGEMA_signal_7720), .Z1_f (new_AGEMA_signal_7721) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_21_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_6594), .B0_t (MUX_StateInMC_mux_inst_21_X), .B0_f (new_AGEMA_signal_7719), .B1_t (new_AGEMA_signal_7720), .B1_f (new_AGEMA_signal_7721), .Z0_t (MUX_StateInMC_mux_inst_21_Y), .Z0_f (new_AGEMA_signal_8493), .Z1_t (new_AGEMA_signal_8494), .Z1_f (new_AGEMA_signal_8495) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_21_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_21_Y), .A0_f (new_AGEMA_signal_8493), .A1_t (new_AGEMA_signal_8494), .A1_f (new_AGEMA_signal_8495), .B0_t (MCout[21]), .B0_f (new_AGEMA_signal_7300), .B1_t (new_AGEMA_signal_7301), .B1_f (new_AGEMA_signal_7302), .Z0_t (StateInMC[21]), .Z0_f (new_AGEMA_signal_9367), .Z1_t (new_AGEMA_signal_9368), .Z1_f (new_AGEMA_signal_9369) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_22_XOR1_U1 ( .A0_t (MCout[22]), .A0_f (new_AGEMA_signal_7297), .A1_t (new_AGEMA_signal_7298), .A1_f (new_AGEMA_signal_7299), .B0_t (ciphertext_s0_t[118]), .B0_f (ciphertext_s0_f[118]), .B1_t (ciphertext_s1_t[118]), .B1_f (ciphertext_s1_f[118]), .Z0_t (MUX_StateInMC_mux_inst_22_X), .Z0_f (new_AGEMA_signal_7722), .Z1_t (new_AGEMA_signal_7723), .Z1_f (new_AGEMA_signal_7724) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_22_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_6594), .B0_t (MUX_StateInMC_mux_inst_22_X), .B0_f (new_AGEMA_signal_7722), .B1_t (new_AGEMA_signal_7723), .B1_f (new_AGEMA_signal_7724), .Z0_t (MUX_StateInMC_mux_inst_22_Y), .Z0_f (new_AGEMA_signal_8496), .Z1_t (new_AGEMA_signal_8497), .Z1_f (new_AGEMA_signal_8498) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_22_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_22_Y), .A0_f (new_AGEMA_signal_8496), .A1_t (new_AGEMA_signal_8497), .A1_f (new_AGEMA_signal_8498), .B0_t (MCout[22]), .B0_f (new_AGEMA_signal_7297), .B1_t (new_AGEMA_signal_7298), .B1_f (new_AGEMA_signal_7299), .Z0_t (StateInMC[22]), .Z0_f (new_AGEMA_signal_9370), .Z1_t (new_AGEMA_signal_9371), .Z1_f (new_AGEMA_signal_9372) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_23_XOR1_U1 ( .A0_t (MCout[23]), .A0_f (new_AGEMA_signal_7294), .A1_t (new_AGEMA_signal_7295), .A1_f (new_AGEMA_signal_7296), .B0_t (ciphertext_s0_t[119]), .B0_f (ciphertext_s0_f[119]), .B1_t (ciphertext_s1_t[119]), .B1_f (ciphertext_s1_f[119]), .Z0_t (MUX_StateInMC_mux_inst_23_X), .Z0_f (new_AGEMA_signal_7725), .Z1_t (new_AGEMA_signal_7726), .Z1_f (new_AGEMA_signal_7727) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_23_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_6594), .B0_t (MUX_StateInMC_mux_inst_23_X), .B0_f (new_AGEMA_signal_7725), .B1_t (new_AGEMA_signal_7726), .B1_f (new_AGEMA_signal_7727), .Z0_t (MUX_StateInMC_mux_inst_23_Y), .Z0_f (new_AGEMA_signal_8499), .Z1_t (new_AGEMA_signal_8500), .Z1_f (new_AGEMA_signal_8501) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_23_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_23_Y), .A0_f (new_AGEMA_signal_8499), .A1_t (new_AGEMA_signal_8500), .A1_f (new_AGEMA_signal_8501), .B0_t (MCout[23]), .B0_f (new_AGEMA_signal_7294), .B1_t (new_AGEMA_signal_7295), .B1_f (new_AGEMA_signal_7296), .Z0_t (StateInMC[23]), .Z0_f (new_AGEMA_signal_9373), .Z1_t (new_AGEMA_signal_9374), .Z1_f (new_AGEMA_signal_9375) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_24_XOR1_U1 ( .A0_t (MCout[24]), .A0_f (new_AGEMA_signal_7291), .A1_t (new_AGEMA_signal_7292), .A1_f (new_AGEMA_signal_7293), .B0_t (ciphertext_s0_t[120]), .B0_f (ciphertext_s0_f[120]), .B1_t (ciphertext_s1_t[120]), .B1_f (ciphertext_s1_f[120]), .Z0_t (MUX_StateInMC_mux_inst_24_X), .Z0_f (new_AGEMA_signal_7728), .Z1_t (new_AGEMA_signal_7729), .Z1_f (new_AGEMA_signal_7730) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_24_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_6594), .B0_t (MUX_StateInMC_mux_inst_24_X), .B0_f (new_AGEMA_signal_7728), .B1_t (new_AGEMA_signal_7729), .B1_f (new_AGEMA_signal_7730), .Z0_t (MUX_StateInMC_mux_inst_24_Y), .Z0_f (new_AGEMA_signal_8502), .Z1_t (new_AGEMA_signal_8503), .Z1_f (new_AGEMA_signal_8504) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_24_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_24_Y), .A0_f (new_AGEMA_signal_8502), .A1_t (new_AGEMA_signal_8503), .A1_f (new_AGEMA_signal_8504), .B0_t (MCout[24]), .B0_f (new_AGEMA_signal_7291), .B1_t (new_AGEMA_signal_7292), .B1_f (new_AGEMA_signal_7293), .Z0_t (StateInMC[24]), .Z0_f (new_AGEMA_signal_9376), .Z1_t (new_AGEMA_signal_9377), .Z1_f (new_AGEMA_signal_9378) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_25_XOR1_U1 ( .A0_t (MCout[25]), .A0_f (new_AGEMA_signal_8085), .A1_t (new_AGEMA_signal_8086), .A1_f (new_AGEMA_signal_8087), .B0_t (ciphertext_s0_t[121]), .B0_f (ciphertext_s0_f[121]), .B1_t (ciphertext_s1_t[121]), .B1_f (ciphertext_s1_f[121]), .Z0_t (MUX_StateInMC_mux_inst_25_X), .Z0_f (new_AGEMA_signal_8505), .Z1_t (new_AGEMA_signal_8506), .Z1_f (new_AGEMA_signal_8507) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_25_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_6594), .B0_t (MUX_StateInMC_mux_inst_25_X), .B0_f (new_AGEMA_signal_8505), .B1_t (new_AGEMA_signal_8506), .B1_f (new_AGEMA_signal_8507), .Z0_t (MUX_StateInMC_mux_inst_25_Y), .Z0_f (new_AGEMA_signal_9379), .Z1_t (new_AGEMA_signal_9380), .Z1_f (new_AGEMA_signal_9381) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_25_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_25_Y), .A0_f (new_AGEMA_signal_9379), .A1_t (new_AGEMA_signal_9380), .A1_f (new_AGEMA_signal_9381), .B0_t (MCout[25]), .B0_f (new_AGEMA_signal_8085), .B1_t (new_AGEMA_signal_8086), .B1_f (new_AGEMA_signal_8087), .Z0_t (StateInMC[25]), .Z0_f (new_AGEMA_signal_9867), .Z1_t (new_AGEMA_signal_9868), .Z1_f (new_AGEMA_signal_9869) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_26_XOR1_U1 ( .A0_t (MCout[26]), .A0_f (new_AGEMA_signal_7285), .A1_t (new_AGEMA_signal_7286), .A1_f (new_AGEMA_signal_7287), .B0_t (ciphertext_s0_t[122]), .B0_f (ciphertext_s0_f[122]), .B1_t (ciphertext_s1_t[122]), .B1_f (ciphertext_s1_f[122]), .Z0_t (MUX_StateInMC_mux_inst_26_X), .Z0_f (new_AGEMA_signal_7731), .Z1_t (new_AGEMA_signal_7732), .Z1_f (new_AGEMA_signal_7733) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_26_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_6594), .B0_t (MUX_StateInMC_mux_inst_26_X), .B0_f (new_AGEMA_signal_7731), .B1_t (new_AGEMA_signal_7732), .B1_f (new_AGEMA_signal_7733), .Z0_t (MUX_StateInMC_mux_inst_26_Y), .Z0_f (new_AGEMA_signal_8508), .Z1_t (new_AGEMA_signal_8509), .Z1_f (new_AGEMA_signal_8510) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_26_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_26_Y), .A0_f (new_AGEMA_signal_8508), .A1_t (new_AGEMA_signal_8509), .A1_f (new_AGEMA_signal_8510), .B0_t (MCout[26]), .B0_f (new_AGEMA_signal_7285), .B1_t (new_AGEMA_signal_7286), .B1_f (new_AGEMA_signal_7287), .Z0_t (StateInMC[26]), .Z0_f (new_AGEMA_signal_9382), .Z1_t (new_AGEMA_signal_9383), .Z1_f (new_AGEMA_signal_9384) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_27_XOR1_U1 ( .A0_t (MCout[27]), .A0_f (new_AGEMA_signal_8082), .A1_t (new_AGEMA_signal_8083), .A1_f (new_AGEMA_signal_8084), .B0_t (ciphertext_s0_t[123]), .B0_f (ciphertext_s0_f[123]), .B1_t (ciphertext_s1_t[123]), .B1_f (ciphertext_s1_f[123]), .Z0_t (MUX_StateInMC_mux_inst_27_X), .Z0_f (new_AGEMA_signal_8511), .Z1_t (new_AGEMA_signal_8512), .Z1_f (new_AGEMA_signal_8513) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_27_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_6594), .B0_t (MUX_StateInMC_mux_inst_27_X), .B0_f (new_AGEMA_signal_8511), .B1_t (new_AGEMA_signal_8512), .B1_f (new_AGEMA_signal_8513), .Z0_t (MUX_StateInMC_mux_inst_27_Y), .Z0_f (new_AGEMA_signal_9385), .Z1_t (new_AGEMA_signal_9386), .Z1_f (new_AGEMA_signal_9387) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_27_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_27_Y), .A0_f (new_AGEMA_signal_9385), .A1_t (new_AGEMA_signal_9386), .A1_f (new_AGEMA_signal_9387), .B0_t (MCout[27]), .B0_f (new_AGEMA_signal_8082), .B1_t (new_AGEMA_signal_8083), .B1_f (new_AGEMA_signal_8084), .Z0_t (StateInMC[27]), .Z0_f (new_AGEMA_signal_9870), .Z1_t (new_AGEMA_signal_9871), .Z1_f (new_AGEMA_signal_9872) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_28_XOR1_U1 ( .A0_t (MCout[28]), .A0_f (new_AGEMA_signal_8079), .A1_t (new_AGEMA_signal_8080), .A1_f (new_AGEMA_signal_8081), .B0_t (ciphertext_s0_t[124]), .B0_f (ciphertext_s0_f[124]), .B1_t (ciphertext_s1_t[124]), .B1_f (ciphertext_s1_f[124]), .Z0_t (MUX_StateInMC_mux_inst_28_X), .Z0_f (new_AGEMA_signal_8514), .Z1_t (new_AGEMA_signal_8515), .Z1_f (new_AGEMA_signal_8516) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_28_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_6594), .B0_t (MUX_StateInMC_mux_inst_28_X), .B0_f (new_AGEMA_signal_8514), .B1_t (new_AGEMA_signal_8515), .B1_f (new_AGEMA_signal_8516), .Z0_t (MUX_StateInMC_mux_inst_28_Y), .Z0_f (new_AGEMA_signal_9388), .Z1_t (new_AGEMA_signal_9389), .Z1_f (new_AGEMA_signal_9390) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_28_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_28_Y), .A0_f (new_AGEMA_signal_9388), .A1_t (new_AGEMA_signal_9389), .A1_f (new_AGEMA_signal_9390), .B0_t (MCout[28]), .B0_f (new_AGEMA_signal_8079), .B1_t (new_AGEMA_signal_8080), .B1_f (new_AGEMA_signal_8081), .Z0_t (StateInMC[28]), .Z0_f (new_AGEMA_signal_9873), .Z1_t (new_AGEMA_signal_9874), .Z1_f (new_AGEMA_signal_9875) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_29_XOR1_U1 ( .A0_t (MCout[29]), .A0_f (new_AGEMA_signal_7276), .A1_t (new_AGEMA_signal_7277), .A1_f (new_AGEMA_signal_7278), .B0_t (ciphertext_s0_t[125]), .B0_f (ciphertext_s0_f[125]), .B1_t (ciphertext_s1_t[125]), .B1_f (ciphertext_s1_f[125]), .Z0_t (MUX_StateInMC_mux_inst_29_X), .Z0_f (new_AGEMA_signal_7734), .Z1_t (new_AGEMA_signal_7735), .Z1_f (new_AGEMA_signal_7736) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_29_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_6594), .B0_t (MUX_StateInMC_mux_inst_29_X), .B0_f (new_AGEMA_signal_7734), .B1_t (new_AGEMA_signal_7735), .B1_f (new_AGEMA_signal_7736), .Z0_t (MUX_StateInMC_mux_inst_29_Y), .Z0_f (new_AGEMA_signal_8517), .Z1_t (new_AGEMA_signal_8518), .Z1_f (new_AGEMA_signal_8519) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_29_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_29_Y), .A0_f (new_AGEMA_signal_8517), .A1_t (new_AGEMA_signal_8518), .A1_f (new_AGEMA_signal_8519), .B0_t (MCout[29]), .B0_f (new_AGEMA_signal_7276), .B1_t (new_AGEMA_signal_7277), .B1_f (new_AGEMA_signal_7278), .Z0_t (StateInMC[29]), .Z0_f (new_AGEMA_signal_9391), .Z1_t (new_AGEMA_signal_9392), .Z1_f (new_AGEMA_signal_9393) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_30_XOR1_U1 ( .A0_t (MCout[30]), .A0_f (new_AGEMA_signal_7273), .A1_t (new_AGEMA_signal_7274), .A1_f (new_AGEMA_signal_7275), .B0_t (ciphertext_s0_t[126]), .B0_f (ciphertext_s0_f[126]), .B1_t (ciphertext_s1_t[126]), .B1_f (ciphertext_s1_f[126]), .Z0_t (MUX_StateInMC_mux_inst_30_X), .Z0_f (new_AGEMA_signal_7737), .Z1_t (new_AGEMA_signal_7738), .Z1_f (new_AGEMA_signal_7739) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_30_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_6594), .B0_t (MUX_StateInMC_mux_inst_30_X), .B0_f (new_AGEMA_signal_7737), .B1_t (new_AGEMA_signal_7738), .B1_f (new_AGEMA_signal_7739), .Z0_t (MUX_StateInMC_mux_inst_30_Y), .Z0_f (new_AGEMA_signal_8520), .Z1_t (new_AGEMA_signal_8521), .Z1_f (new_AGEMA_signal_8522) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_30_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_30_Y), .A0_f (new_AGEMA_signal_8520), .A1_t (new_AGEMA_signal_8521), .A1_f (new_AGEMA_signal_8522), .B0_t (MCout[30]), .B0_f (new_AGEMA_signal_7273), .B1_t (new_AGEMA_signal_7274), .B1_f (new_AGEMA_signal_7275), .Z0_t (StateInMC[30]), .Z0_f (new_AGEMA_signal_9394), .Z1_t (new_AGEMA_signal_9395), .Z1_f (new_AGEMA_signal_9396) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_31_XOR1_U1 ( .A0_t (MCout[31]), .A0_f (new_AGEMA_signal_7270), .A1_t (new_AGEMA_signal_7271), .A1_f (new_AGEMA_signal_7272), .B0_t (ciphertext_s0_t[127]), .B0_f (ciphertext_s0_f[127]), .B1_t (ciphertext_s1_t[127]), .B1_f (ciphertext_s1_f[127]), .Z0_t (MUX_StateInMC_mux_inst_31_X), .Z0_f (new_AGEMA_signal_7740), .Z1_t (new_AGEMA_signal_7741), .Z1_f (new_AGEMA_signal_7742) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_31_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_6594), .B0_t (MUX_StateInMC_mux_inst_31_X), .B0_f (new_AGEMA_signal_7740), .B1_t (new_AGEMA_signal_7741), .B1_f (new_AGEMA_signal_7742), .Z0_t (MUX_StateInMC_mux_inst_31_Y), .Z0_f (new_AGEMA_signal_8523), .Z1_t (new_AGEMA_signal_8524), .Z1_f (new_AGEMA_signal_8525) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_31_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_31_Y), .A0_f (new_AGEMA_signal_8523), .A1_t (new_AGEMA_signal_8524), .A1_f (new_AGEMA_signal_8525), .B0_t (MCout[31]), .B0_f (new_AGEMA_signal_7270), .B1_t (new_AGEMA_signal_7271), .B1_f (new_AGEMA_signal_7272), .Z0_t (StateInMC[31]), .Z0_f (new_AGEMA_signal_9397), .Z1_t (new_AGEMA_signal_9398), .Z1_f (new_AGEMA_signal_9399) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_U34 ( .A0_t (KeyArray_outS01ser_7_), .A0_f (new_AGEMA_signal_4386), .A1_t (new_AGEMA_signal_4387), .A1_f (new_AGEMA_signal_4388), .B0_t (keyStateIn[7]), .B0_f (new_AGEMA_signal_3495), .B1_t (new_AGEMA_signal_3496), .B1_f (new_AGEMA_signal_3497), .Z0_t (KeyArray_outS01ser_XOR_00[7]), .Z0_f (new_AGEMA_signal_4389), .Z1_t (new_AGEMA_signal_4390), .Z1_f (new_AGEMA_signal_4391) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_U33 ( .A0_t (KeyArray_outS01ser_6_), .A0_f (new_AGEMA_signal_4392), .A1_t (new_AGEMA_signal_4393), .A1_f (new_AGEMA_signal_4394), .B0_t (keyStateIn[6]), .B0_f (new_AGEMA_signal_3486), .B1_t (new_AGEMA_signal_3487), .B1_f (new_AGEMA_signal_3488), .Z0_t (KeyArray_outS01ser_XOR_00[6]), .Z0_f (new_AGEMA_signal_4395), .Z1_t (new_AGEMA_signal_4396), .Z1_f (new_AGEMA_signal_4397) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_U32 ( .A0_t (KeyArray_outS01ser_5_), .A0_f (new_AGEMA_signal_4398), .A1_t (new_AGEMA_signal_4399), .A1_f (new_AGEMA_signal_4400), .B0_t (keyStateIn[5]), .B0_f (new_AGEMA_signal_3477), .B1_t (new_AGEMA_signal_3478), .B1_f (new_AGEMA_signal_3479), .Z0_t (KeyArray_outS01ser_XOR_00[5]), .Z0_f (new_AGEMA_signal_4401), .Z1_t (new_AGEMA_signal_4402), .Z1_f (new_AGEMA_signal_4403) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_U31 ( .A0_t (KeyArray_outS01ser_4_), .A0_f (new_AGEMA_signal_4404), .A1_t (new_AGEMA_signal_4405), .A1_f (new_AGEMA_signal_4406), .B0_t (keyStateIn[4]), .B0_f (new_AGEMA_signal_3468), .B1_t (new_AGEMA_signal_3469), .B1_f (new_AGEMA_signal_3470), .Z0_t (KeyArray_outS01ser_XOR_00[4]), .Z0_f (new_AGEMA_signal_4407), .Z1_t (new_AGEMA_signal_4408), .Z1_f (new_AGEMA_signal_4409) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_U30 ( .A0_t (KeyArray_outS01ser_3_), .A0_f (new_AGEMA_signal_4410), .A1_t (new_AGEMA_signal_4411), .A1_f (new_AGEMA_signal_4412), .B0_t (keyStateIn[3]), .B0_f (new_AGEMA_signal_3459), .B1_t (new_AGEMA_signal_3460), .B1_f (new_AGEMA_signal_3461), .Z0_t (KeyArray_outS01ser_XOR_00[3]), .Z0_f (new_AGEMA_signal_4413), .Z1_t (new_AGEMA_signal_4414), .Z1_f (new_AGEMA_signal_4415) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_U29 ( .A0_t (KeyArray_outS01ser_2_), .A0_f (new_AGEMA_signal_4416), .A1_t (new_AGEMA_signal_4417), .A1_f (new_AGEMA_signal_4418), .B0_t (keyStateIn[2]), .B0_f (new_AGEMA_signal_3450), .B1_t (new_AGEMA_signal_3451), .B1_f (new_AGEMA_signal_3452), .Z0_t (KeyArray_outS01ser_XOR_00[2]), .Z0_f (new_AGEMA_signal_4419), .Z1_t (new_AGEMA_signal_4420), .Z1_f (new_AGEMA_signal_4421) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_U28 ( .A0_t (KeyArray_outS01ser_1_), .A0_f (new_AGEMA_signal_4422), .A1_t (new_AGEMA_signal_4423), .A1_f (new_AGEMA_signal_4424), .B0_t (keyStateIn[1]), .B0_f (new_AGEMA_signal_3441), .B1_t (new_AGEMA_signal_3442), .B1_f (new_AGEMA_signal_3443), .Z0_t (KeyArray_outS01ser_XOR_00[1]), .Z0_f (new_AGEMA_signal_4425), .Z1_t (new_AGEMA_signal_4426), .Z1_f (new_AGEMA_signal_4427) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_U27 ( .A0_t (KeyArray_outS01ser_0_), .A0_f (new_AGEMA_signal_4428), .A1_t (new_AGEMA_signal_4429), .A1_f (new_AGEMA_signal_4430), .B0_t (keyStateIn[0]), .B0_f (new_AGEMA_signal_3432), .B1_t (new_AGEMA_signal_3433), .B1_f (new_AGEMA_signal_3434), .Z0_t (KeyArray_outS01ser_XOR_00[0]), .Z0_f (new_AGEMA_signal_4431), .Z1_t (new_AGEMA_signal_4432), .Z1_f (new_AGEMA_signal_4433) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_U26 ( .A0_t (KeyArray_n40), .A0_f (new_AGEMA_signal_11375), .A1_t (new_AGEMA_signal_11376), .A1_f (new_AGEMA_signal_11377), .B0_t (keyStateIn[7]), .B0_f (new_AGEMA_signal_3495), .B1_t (new_AGEMA_signal_3496), .B1_f (new_AGEMA_signal_3497), .Z0_t (KeyArray_inS30par[7]), .Z0_f (new_AGEMA_signal_11423), .Z1_t (new_AGEMA_signal_11424), .Z1_f (new_AGEMA_signal_11425) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_U25 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (roundConstant[7]), .A1_f (new_AGEMA_signal_5792), .B0_t (SboxOut[7]), .B0_f (new_AGEMA_signal_11330), .B1_t (new_AGEMA_signal_11331), .B1_f (new_AGEMA_signal_11332), .Z0_t (KeyArray_n40), .Z0_f (new_AGEMA_signal_11375), .Z1_t (new_AGEMA_signal_11376), .Z1_f (new_AGEMA_signal_11377) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_U24 ( .A0_t (KeyArray_n39), .A0_f (new_AGEMA_signal_11378), .A1_t (new_AGEMA_signal_11379), .A1_f (new_AGEMA_signal_11380), .B0_t (keyStateIn[6]), .B0_f (new_AGEMA_signal_3486), .B1_t (new_AGEMA_signal_3487), .B1_f (new_AGEMA_signal_3488), .Z0_t (KeyArray_inS30par[6]), .Z0_f (new_AGEMA_signal_11426), .Z1_t (new_AGEMA_signal_11427), .Z1_f (new_AGEMA_signal_11428) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_U23 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (roundConstant[6]), .A1_f (new_AGEMA_signal_5794), .B0_t (SboxOut[6]), .B0_f (new_AGEMA_signal_11333), .B1_t (new_AGEMA_signal_11334), .B1_f (new_AGEMA_signal_11335), .Z0_t (KeyArray_n39), .Z0_f (new_AGEMA_signal_11378), .Z1_t (new_AGEMA_signal_11379), .Z1_f (new_AGEMA_signal_11380) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_U22 ( .A0_t (KeyArray_n38), .A0_f (new_AGEMA_signal_11381), .A1_t (new_AGEMA_signal_11382), .A1_f (new_AGEMA_signal_11383), .B0_t (keyStateIn[5]), .B0_f (new_AGEMA_signal_3477), .B1_t (new_AGEMA_signal_3478), .B1_f (new_AGEMA_signal_3479), .Z0_t (KeyArray_inS30par[5]), .Z0_f (new_AGEMA_signal_11429), .Z1_t (new_AGEMA_signal_11430), .Z1_f (new_AGEMA_signal_11431) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_U21 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (roundConstant[5]), .A1_f (new_AGEMA_signal_5796), .B0_t (SboxOut[5]), .B0_f (new_AGEMA_signal_11336), .B1_t (new_AGEMA_signal_11337), .B1_f (new_AGEMA_signal_11338), .Z0_t (KeyArray_n38), .Z0_f (new_AGEMA_signal_11381), .Z1_t (new_AGEMA_signal_11382), .Z1_f (new_AGEMA_signal_11383) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_U20 ( .A0_t (KeyArray_n37), .A0_f (new_AGEMA_signal_11384), .A1_t (new_AGEMA_signal_11385), .A1_f (new_AGEMA_signal_11386), .B0_t (keyStateIn[4]), .B0_f (new_AGEMA_signal_3468), .B1_t (new_AGEMA_signal_3469), .B1_f (new_AGEMA_signal_3470), .Z0_t (KeyArray_inS30par[4]), .Z0_f (new_AGEMA_signal_11432), .Z1_t (new_AGEMA_signal_11433), .Z1_f (new_AGEMA_signal_11434) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_U19 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (roundConstant[4]), .A1_f (new_AGEMA_signal_5798), .B0_t (SboxOut[4]), .B0_f (new_AGEMA_signal_11339), .B1_t (new_AGEMA_signal_11340), .B1_f (new_AGEMA_signal_11341), .Z0_t (KeyArray_n37), .Z0_f (new_AGEMA_signal_11384), .Z1_t (new_AGEMA_signal_11385), .Z1_f (new_AGEMA_signal_11386) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_U18 ( .A0_t (KeyArray_n36), .A0_f (new_AGEMA_signal_11387), .A1_t (new_AGEMA_signal_11388), .A1_f (new_AGEMA_signal_11389), .B0_t (keyStateIn[3]), .B0_f (new_AGEMA_signal_3459), .B1_t (new_AGEMA_signal_3460), .B1_f (new_AGEMA_signal_3461), .Z0_t (KeyArray_inS30par[3]), .Z0_f (new_AGEMA_signal_11435), .Z1_t (new_AGEMA_signal_11436), .Z1_f (new_AGEMA_signal_11437) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_U17 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (roundConstant[3]), .A1_f (new_AGEMA_signal_5800), .B0_t (SboxOut[3]), .B0_f (new_AGEMA_signal_11342), .B1_t (new_AGEMA_signal_11343), .B1_f (new_AGEMA_signal_11344), .Z0_t (KeyArray_n36), .Z0_f (new_AGEMA_signal_11387), .Z1_t (new_AGEMA_signal_11388), .Z1_f (new_AGEMA_signal_11389) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_U16 ( .A0_t (KeyArray_n35), .A0_f (new_AGEMA_signal_11390), .A1_t (new_AGEMA_signal_11391), .A1_f (new_AGEMA_signal_11392), .B0_t (keyStateIn[2]), .B0_f (new_AGEMA_signal_3450), .B1_t (new_AGEMA_signal_3451), .B1_f (new_AGEMA_signal_3452), .Z0_t (KeyArray_inS30par[2]), .Z0_f (new_AGEMA_signal_11438), .Z1_t (new_AGEMA_signal_11439), .Z1_f (new_AGEMA_signal_11440) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_U15 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (roundConstant[2]), .A1_f (new_AGEMA_signal_5802), .B0_t (SboxOut[2]), .B0_f (new_AGEMA_signal_11345), .B1_t (new_AGEMA_signal_11346), .B1_f (new_AGEMA_signal_11347), .Z0_t (KeyArray_n35), .Z0_f (new_AGEMA_signal_11390), .Z1_t (new_AGEMA_signal_11391), .Z1_f (new_AGEMA_signal_11392) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_U14 ( .A0_t (KeyArray_n34), .A0_f (new_AGEMA_signal_11393), .A1_t (new_AGEMA_signal_11394), .A1_f (new_AGEMA_signal_11395), .B0_t (keyStateIn[1]), .B0_f (new_AGEMA_signal_3441), .B1_t (new_AGEMA_signal_3442), .B1_f (new_AGEMA_signal_3443), .Z0_t (KeyArray_inS30par[1]), .Z0_f (new_AGEMA_signal_11441), .Z1_t (new_AGEMA_signal_11442), .Z1_f (new_AGEMA_signal_11443) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_U13 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (roundConstant[1]), .A1_f (new_AGEMA_signal_5804), .B0_t (SboxOut[1]), .B0_f (new_AGEMA_signal_11348), .B1_t (new_AGEMA_signal_11349), .B1_f (new_AGEMA_signal_11350), .Z0_t (KeyArray_n34), .Z0_f (new_AGEMA_signal_11393), .Z1_t (new_AGEMA_signal_11394), .Z1_f (new_AGEMA_signal_11395) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_U12 ( .A0_t (KeyArray_n33), .A0_f (new_AGEMA_signal_11327), .A1_t (new_AGEMA_signal_11328), .A1_f (new_AGEMA_signal_11329), .B0_t (keyStateIn[0]), .B0_f (new_AGEMA_signal_3432), .B1_t (new_AGEMA_signal_3433), .B1_f (new_AGEMA_signal_3434), .Z0_t (KeyArray_inS30par[0]), .Z0_f (new_AGEMA_signal_11396), .Z1_t (new_AGEMA_signal_11397), .Z1_f (new_AGEMA_signal_11398) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_U11 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (roundConstant[0]), .A1_f (new_AGEMA_signal_5806), .B0_t (SboxOut[0]), .B0_f (new_AGEMA_signal_11321), .B1_t (new_AGEMA_signal_11322), .B1_f (new_AGEMA_signal_11323), .Z0_t (KeyArray_n33), .Z0_f (new_AGEMA_signal_11327), .Z1_t (new_AGEMA_signal_11328), .Z1_f (new_AGEMA_signal_11329) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S00reg_gff_1_SFF_0_U3 ( .A0_t (KeyArray_S00reg_gff_1_SFF_0_n2), .A0_f (new_AGEMA_signal_11012), .A1_t (new_AGEMA_signal_11013), .A1_f (new_AGEMA_signal_11014), .B0_t (KeyArray_S00reg_gff_1_SFF_0_n1), .B0_f (new_AGEMA_signal_8526), .B1_t (new_AGEMA_signal_8527), .B1_f (new_AGEMA_signal_8528), .Z0_t (keyStateIn[0]), .Z0_f (new_AGEMA_signal_3432), .Z1_t (new_AGEMA_signal_3433), .Z1_f (new_AGEMA_signal_3434) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_0_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (keyStateIn[0]), .B0_f (new_AGEMA_signal_3432), .B1_t (new_AGEMA_signal_3433), .B1_f (new_AGEMA_signal_3434), .Z0_t (KeyArray_S00reg_gff_1_SFF_0_n1), .Z0_f (new_AGEMA_signal_8526), .Z1_t (new_AGEMA_signal_8527), .Z1_f (new_AGEMA_signal_8528) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_0_U1 ( .A0_t (KeyArray_S00reg_gff_1_SFF_0_QD), .A0_f (new_AGEMA_signal_10901), .A1_t (new_AGEMA_signal_10902), .A1_f (new_AGEMA_signal_10903), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S00reg_gff_1_SFF_0_n2), .Z0_f (new_AGEMA_signal_11012), .Z1_t (new_AGEMA_signal_11013), .Z1_f (new_AGEMA_signal_11014) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS00ser[0]), .A0_f (new_AGEMA_signal_10502), .A1_t (new_AGEMA_signal_10503), .A1_f (new_AGEMA_signal_10504), .B0_t (KeyArray_outS10ser[0]), .B0_f (new_AGEMA_signal_4581), .B1_t (new_AGEMA_signal_4582), .B1_f (new_AGEMA_signal_4583), .Z0_t (KeyArray_S00reg_gff_1_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_10658), .Z1_t (new_AGEMA_signal_10659), .Z1_f (new_AGEMA_signal_10660) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S00reg_gff_1_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_10658), .B1_t (new_AGEMA_signal_10659), .B1_f (new_AGEMA_signal_10660), .Z0_t (KeyArray_S00reg_gff_1_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_10793), .Z1_t (new_AGEMA_signal_10794), .Z1_f (new_AGEMA_signal_10795) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S00reg_gff_1_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_10793), .A1_t (new_AGEMA_signal_10794), .A1_f (new_AGEMA_signal_10795), .B0_t (KeyArray_inS00ser[0]), .B0_f (new_AGEMA_signal_10502), .B1_t (new_AGEMA_signal_10503), .B1_f (new_AGEMA_signal_10504), .Z0_t (KeyArray_S00reg_gff_1_SFF_0_QD), .Z0_f (new_AGEMA_signal_10901), .Z1_t (new_AGEMA_signal_10902), .Z1_f (new_AGEMA_signal_10903) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S00reg_gff_1_SFF_1_U3 ( .A0_t (KeyArray_S00reg_gff_1_SFF_1_n2), .A0_f (new_AGEMA_signal_11015), .A1_t (new_AGEMA_signal_11016), .A1_f (new_AGEMA_signal_11017), .B0_t (KeyArray_S00reg_gff_1_SFF_1_n1), .B0_f (new_AGEMA_signal_8529), .B1_t (new_AGEMA_signal_8530), .B1_f (new_AGEMA_signal_8531), .Z0_t (keyStateIn[1]), .Z0_f (new_AGEMA_signal_3441), .Z1_t (new_AGEMA_signal_3442), .Z1_f (new_AGEMA_signal_3443) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_1_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (keyStateIn[1]), .B0_f (new_AGEMA_signal_3441), .B1_t (new_AGEMA_signal_3442), .B1_f (new_AGEMA_signal_3443), .Z0_t (KeyArray_S00reg_gff_1_SFF_1_n1), .Z0_f (new_AGEMA_signal_8529), .Z1_t (new_AGEMA_signal_8530), .Z1_f (new_AGEMA_signal_8531) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_1_U1 ( .A0_t (KeyArray_S00reg_gff_1_SFF_1_QD), .A0_f (new_AGEMA_signal_10904), .A1_t (new_AGEMA_signal_10905), .A1_f (new_AGEMA_signal_10906), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S00reg_gff_1_SFF_1_n2), .Z0_f (new_AGEMA_signal_11015), .Z1_t (new_AGEMA_signal_11016), .Z1_f (new_AGEMA_signal_11017) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS00ser[1]), .A0_f (new_AGEMA_signal_10505), .A1_t (new_AGEMA_signal_10506), .A1_f (new_AGEMA_signal_10507), .B0_t (KeyArray_outS10ser[1]), .B0_f (new_AGEMA_signal_4590), .B1_t (new_AGEMA_signal_4591), .B1_f (new_AGEMA_signal_4592), .Z0_t (KeyArray_S00reg_gff_1_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_10661), .Z1_t (new_AGEMA_signal_10662), .Z1_f (new_AGEMA_signal_10663) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S00reg_gff_1_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_10661), .B1_t (new_AGEMA_signal_10662), .B1_f (new_AGEMA_signal_10663), .Z0_t (KeyArray_S00reg_gff_1_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_10796), .Z1_t (new_AGEMA_signal_10797), .Z1_f (new_AGEMA_signal_10798) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S00reg_gff_1_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_10796), .A1_t (new_AGEMA_signal_10797), .A1_f (new_AGEMA_signal_10798), .B0_t (KeyArray_inS00ser[1]), .B0_f (new_AGEMA_signal_10505), .B1_t (new_AGEMA_signal_10506), .B1_f (new_AGEMA_signal_10507), .Z0_t (KeyArray_S00reg_gff_1_SFF_1_QD), .Z0_f (new_AGEMA_signal_10904), .Z1_t (new_AGEMA_signal_10905), .Z1_f (new_AGEMA_signal_10906) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S00reg_gff_1_SFF_2_U3 ( .A0_t (KeyArray_S00reg_gff_1_SFF_2_n2), .A0_f (new_AGEMA_signal_11018), .A1_t (new_AGEMA_signal_11019), .A1_f (new_AGEMA_signal_11020), .B0_t (KeyArray_S00reg_gff_1_SFF_2_n1), .B0_f (new_AGEMA_signal_8532), .B1_t (new_AGEMA_signal_8533), .B1_f (new_AGEMA_signal_8534), .Z0_t (keyStateIn[2]), .Z0_f (new_AGEMA_signal_3450), .Z1_t (new_AGEMA_signal_3451), .Z1_f (new_AGEMA_signal_3452) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_2_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (keyStateIn[2]), .B0_f (new_AGEMA_signal_3450), .B1_t (new_AGEMA_signal_3451), .B1_f (new_AGEMA_signal_3452), .Z0_t (KeyArray_S00reg_gff_1_SFF_2_n1), .Z0_f (new_AGEMA_signal_8532), .Z1_t (new_AGEMA_signal_8533), .Z1_f (new_AGEMA_signal_8534) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_2_U1 ( .A0_t (KeyArray_S00reg_gff_1_SFF_2_QD), .A0_f (new_AGEMA_signal_10907), .A1_t (new_AGEMA_signal_10908), .A1_f (new_AGEMA_signal_10909), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S00reg_gff_1_SFF_2_n2), .Z0_f (new_AGEMA_signal_11018), .Z1_t (new_AGEMA_signal_11019), .Z1_f (new_AGEMA_signal_11020) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS00ser[2]), .A0_f (new_AGEMA_signal_10508), .A1_t (new_AGEMA_signal_10509), .A1_f (new_AGEMA_signal_10510), .B0_t (KeyArray_outS10ser[2]), .B0_f (new_AGEMA_signal_4599), .B1_t (new_AGEMA_signal_4600), .B1_f (new_AGEMA_signal_4601), .Z0_t (KeyArray_S00reg_gff_1_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_10664), .Z1_t (new_AGEMA_signal_10665), .Z1_f (new_AGEMA_signal_10666) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S00reg_gff_1_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_10664), .B1_t (new_AGEMA_signal_10665), .B1_f (new_AGEMA_signal_10666), .Z0_t (KeyArray_S00reg_gff_1_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_10799), .Z1_t (new_AGEMA_signal_10800), .Z1_f (new_AGEMA_signal_10801) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S00reg_gff_1_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_10799), .A1_t (new_AGEMA_signal_10800), .A1_f (new_AGEMA_signal_10801), .B0_t (KeyArray_inS00ser[2]), .B0_f (new_AGEMA_signal_10508), .B1_t (new_AGEMA_signal_10509), .B1_f (new_AGEMA_signal_10510), .Z0_t (KeyArray_S00reg_gff_1_SFF_2_QD), .Z0_f (new_AGEMA_signal_10907), .Z1_t (new_AGEMA_signal_10908), .Z1_f (new_AGEMA_signal_10909) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S00reg_gff_1_SFF_3_U3 ( .A0_t (KeyArray_S00reg_gff_1_SFF_3_n2), .A0_f (new_AGEMA_signal_11021), .A1_t (new_AGEMA_signal_11022), .A1_f (new_AGEMA_signal_11023), .B0_t (KeyArray_S00reg_gff_1_SFF_3_n1), .B0_f (new_AGEMA_signal_8535), .B1_t (new_AGEMA_signal_8536), .B1_f (new_AGEMA_signal_8537), .Z0_t (keyStateIn[3]), .Z0_f (new_AGEMA_signal_3459), .Z1_t (new_AGEMA_signal_3460), .Z1_f (new_AGEMA_signal_3461) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_3_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (keyStateIn[3]), .B0_f (new_AGEMA_signal_3459), .B1_t (new_AGEMA_signal_3460), .B1_f (new_AGEMA_signal_3461), .Z0_t (KeyArray_S00reg_gff_1_SFF_3_n1), .Z0_f (new_AGEMA_signal_8535), .Z1_t (new_AGEMA_signal_8536), .Z1_f (new_AGEMA_signal_8537) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_3_U1 ( .A0_t (KeyArray_S00reg_gff_1_SFF_3_QD), .A0_f (new_AGEMA_signal_10910), .A1_t (new_AGEMA_signal_10911), .A1_f (new_AGEMA_signal_10912), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S00reg_gff_1_SFF_3_n2), .Z0_f (new_AGEMA_signal_11021), .Z1_t (new_AGEMA_signal_11022), .Z1_f (new_AGEMA_signal_11023) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS00ser[3]), .A0_f (new_AGEMA_signal_10511), .A1_t (new_AGEMA_signal_10512), .A1_f (new_AGEMA_signal_10513), .B0_t (KeyArray_outS10ser[3]), .B0_f (new_AGEMA_signal_4608), .B1_t (new_AGEMA_signal_4609), .B1_f (new_AGEMA_signal_4610), .Z0_t (KeyArray_S00reg_gff_1_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_10667), .Z1_t (new_AGEMA_signal_10668), .Z1_f (new_AGEMA_signal_10669) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S00reg_gff_1_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_10667), .B1_t (new_AGEMA_signal_10668), .B1_f (new_AGEMA_signal_10669), .Z0_t (KeyArray_S00reg_gff_1_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_10802), .Z1_t (new_AGEMA_signal_10803), .Z1_f (new_AGEMA_signal_10804) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S00reg_gff_1_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_10802), .A1_t (new_AGEMA_signal_10803), .A1_f (new_AGEMA_signal_10804), .B0_t (KeyArray_inS00ser[3]), .B0_f (new_AGEMA_signal_10511), .B1_t (new_AGEMA_signal_10512), .B1_f (new_AGEMA_signal_10513), .Z0_t (KeyArray_S00reg_gff_1_SFF_3_QD), .Z0_f (new_AGEMA_signal_10910), .Z1_t (new_AGEMA_signal_10911), .Z1_f (new_AGEMA_signal_10912) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S00reg_gff_1_SFF_4_U3 ( .A0_t (KeyArray_S00reg_gff_1_SFF_4_n2), .A0_f (new_AGEMA_signal_11024), .A1_t (new_AGEMA_signal_11025), .A1_f (new_AGEMA_signal_11026), .B0_t (KeyArray_S00reg_gff_1_SFF_4_n1), .B0_f (new_AGEMA_signal_8538), .B1_t (new_AGEMA_signal_8539), .B1_f (new_AGEMA_signal_8540), .Z0_t (keyStateIn[4]), .Z0_f (new_AGEMA_signal_3468), .Z1_t (new_AGEMA_signal_3469), .Z1_f (new_AGEMA_signal_3470) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_4_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (keyStateIn[4]), .B0_f (new_AGEMA_signal_3468), .B1_t (new_AGEMA_signal_3469), .B1_f (new_AGEMA_signal_3470), .Z0_t (KeyArray_S00reg_gff_1_SFF_4_n1), .Z0_f (new_AGEMA_signal_8538), .Z1_t (new_AGEMA_signal_8539), .Z1_f (new_AGEMA_signal_8540) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_4_U1 ( .A0_t (KeyArray_S00reg_gff_1_SFF_4_QD), .A0_f (new_AGEMA_signal_10913), .A1_t (new_AGEMA_signal_10914), .A1_f (new_AGEMA_signal_10915), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S00reg_gff_1_SFF_4_n2), .Z0_f (new_AGEMA_signal_11024), .Z1_t (new_AGEMA_signal_11025), .Z1_f (new_AGEMA_signal_11026) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS00ser[4]), .A0_f (new_AGEMA_signal_10514), .A1_t (new_AGEMA_signal_10515), .A1_f (new_AGEMA_signal_10516), .B0_t (KeyArray_outS10ser[4]), .B0_f (new_AGEMA_signal_4617), .B1_t (new_AGEMA_signal_4618), .B1_f (new_AGEMA_signal_4619), .Z0_t (KeyArray_S00reg_gff_1_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_10670), .Z1_t (new_AGEMA_signal_10671), .Z1_f (new_AGEMA_signal_10672) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S00reg_gff_1_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_10670), .B1_t (new_AGEMA_signal_10671), .B1_f (new_AGEMA_signal_10672), .Z0_t (KeyArray_S00reg_gff_1_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_10805), .Z1_t (new_AGEMA_signal_10806), .Z1_f (new_AGEMA_signal_10807) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S00reg_gff_1_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_10805), .A1_t (new_AGEMA_signal_10806), .A1_f (new_AGEMA_signal_10807), .B0_t (KeyArray_inS00ser[4]), .B0_f (new_AGEMA_signal_10514), .B1_t (new_AGEMA_signal_10515), .B1_f (new_AGEMA_signal_10516), .Z0_t (KeyArray_S00reg_gff_1_SFF_4_QD), .Z0_f (new_AGEMA_signal_10913), .Z1_t (new_AGEMA_signal_10914), .Z1_f (new_AGEMA_signal_10915) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S00reg_gff_1_SFF_5_U3 ( .A0_t (KeyArray_S00reg_gff_1_SFF_5_n2), .A0_f (new_AGEMA_signal_11027), .A1_t (new_AGEMA_signal_11028), .A1_f (new_AGEMA_signal_11029), .B0_t (KeyArray_S00reg_gff_1_SFF_5_n1), .B0_f (new_AGEMA_signal_8541), .B1_t (new_AGEMA_signal_8542), .B1_f (new_AGEMA_signal_8543), .Z0_t (keyStateIn[5]), .Z0_f (new_AGEMA_signal_3477), .Z1_t (new_AGEMA_signal_3478), .Z1_f (new_AGEMA_signal_3479) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_5_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (keyStateIn[5]), .B0_f (new_AGEMA_signal_3477), .B1_t (new_AGEMA_signal_3478), .B1_f (new_AGEMA_signal_3479), .Z0_t (KeyArray_S00reg_gff_1_SFF_5_n1), .Z0_f (new_AGEMA_signal_8541), .Z1_t (new_AGEMA_signal_8542), .Z1_f (new_AGEMA_signal_8543) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_5_U1 ( .A0_t (KeyArray_S00reg_gff_1_SFF_5_QD), .A0_f (new_AGEMA_signal_10916), .A1_t (new_AGEMA_signal_10917), .A1_f (new_AGEMA_signal_10918), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S00reg_gff_1_SFF_5_n2), .Z0_f (new_AGEMA_signal_11027), .Z1_t (new_AGEMA_signal_11028), .Z1_f (new_AGEMA_signal_11029) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS00ser[5]), .A0_f (new_AGEMA_signal_10517), .A1_t (new_AGEMA_signal_10518), .A1_f (new_AGEMA_signal_10519), .B0_t (KeyArray_outS10ser[5]), .B0_f (new_AGEMA_signal_4626), .B1_t (new_AGEMA_signal_4627), .B1_f (new_AGEMA_signal_4628), .Z0_t (KeyArray_S00reg_gff_1_SFF_5_MUXInst_X), .Z0_f (new_AGEMA_signal_10673), .Z1_t (new_AGEMA_signal_10674), .Z1_f (new_AGEMA_signal_10675) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S00reg_gff_1_SFF_5_MUXInst_X), .B0_f (new_AGEMA_signal_10673), .B1_t (new_AGEMA_signal_10674), .B1_f (new_AGEMA_signal_10675), .Z0_t (KeyArray_S00reg_gff_1_SFF_5_MUXInst_Y), .Z0_f (new_AGEMA_signal_10808), .Z1_t (new_AGEMA_signal_10809), .Z1_f (new_AGEMA_signal_10810) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S00reg_gff_1_SFF_5_MUXInst_Y), .A0_f (new_AGEMA_signal_10808), .A1_t (new_AGEMA_signal_10809), .A1_f (new_AGEMA_signal_10810), .B0_t (KeyArray_inS00ser[5]), .B0_f (new_AGEMA_signal_10517), .B1_t (new_AGEMA_signal_10518), .B1_f (new_AGEMA_signal_10519), .Z0_t (KeyArray_S00reg_gff_1_SFF_5_QD), .Z0_f (new_AGEMA_signal_10916), .Z1_t (new_AGEMA_signal_10917), .Z1_f (new_AGEMA_signal_10918) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S00reg_gff_1_SFF_6_U3 ( .A0_t (KeyArray_S00reg_gff_1_SFF_6_n2), .A0_f (new_AGEMA_signal_11030), .A1_t (new_AGEMA_signal_11031), .A1_f (new_AGEMA_signal_11032), .B0_t (KeyArray_S00reg_gff_1_SFF_6_n1), .B0_f (new_AGEMA_signal_8544), .B1_t (new_AGEMA_signal_8545), .B1_f (new_AGEMA_signal_8546), .Z0_t (keyStateIn[6]), .Z0_f (new_AGEMA_signal_3486), .Z1_t (new_AGEMA_signal_3487), .Z1_f (new_AGEMA_signal_3488) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_6_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (keyStateIn[6]), .B0_f (new_AGEMA_signal_3486), .B1_t (new_AGEMA_signal_3487), .B1_f (new_AGEMA_signal_3488), .Z0_t (KeyArray_S00reg_gff_1_SFF_6_n1), .Z0_f (new_AGEMA_signal_8544), .Z1_t (new_AGEMA_signal_8545), .Z1_f (new_AGEMA_signal_8546) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_6_U1 ( .A0_t (KeyArray_S00reg_gff_1_SFF_6_QD), .A0_f (new_AGEMA_signal_10919), .A1_t (new_AGEMA_signal_10920), .A1_f (new_AGEMA_signal_10921), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S00reg_gff_1_SFF_6_n2), .Z0_f (new_AGEMA_signal_11030), .Z1_t (new_AGEMA_signal_11031), .Z1_f (new_AGEMA_signal_11032) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS00ser[6]), .A0_f (new_AGEMA_signal_10520), .A1_t (new_AGEMA_signal_10521), .A1_f (new_AGEMA_signal_10522), .B0_t (KeyArray_outS10ser[6]), .B0_f (new_AGEMA_signal_4635), .B1_t (new_AGEMA_signal_4636), .B1_f (new_AGEMA_signal_4637), .Z0_t (KeyArray_S00reg_gff_1_SFF_6_MUXInst_X), .Z0_f (new_AGEMA_signal_10676), .Z1_t (new_AGEMA_signal_10677), .Z1_f (new_AGEMA_signal_10678) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S00reg_gff_1_SFF_6_MUXInst_X), .B0_f (new_AGEMA_signal_10676), .B1_t (new_AGEMA_signal_10677), .B1_f (new_AGEMA_signal_10678), .Z0_t (KeyArray_S00reg_gff_1_SFF_6_MUXInst_Y), .Z0_f (new_AGEMA_signal_10811), .Z1_t (new_AGEMA_signal_10812), .Z1_f (new_AGEMA_signal_10813) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S00reg_gff_1_SFF_6_MUXInst_Y), .A0_f (new_AGEMA_signal_10811), .A1_t (new_AGEMA_signal_10812), .A1_f (new_AGEMA_signal_10813), .B0_t (KeyArray_inS00ser[6]), .B0_f (new_AGEMA_signal_10520), .B1_t (new_AGEMA_signal_10521), .B1_f (new_AGEMA_signal_10522), .Z0_t (KeyArray_S00reg_gff_1_SFF_6_QD), .Z0_f (new_AGEMA_signal_10919), .Z1_t (new_AGEMA_signal_10920), .Z1_f (new_AGEMA_signal_10921) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S00reg_gff_1_SFF_7_U3 ( .A0_t (KeyArray_S00reg_gff_1_SFF_7_n2), .A0_f (new_AGEMA_signal_11033), .A1_t (new_AGEMA_signal_11034), .A1_f (new_AGEMA_signal_11035), .B0_t (KeyArray_S00reg_gff_1_SFF_7_n1), .B0_f (new_AGEMA_signal_8547), .B1_t (new_AGEMA_signal_8548), .B1_f (new_AGEMA_signal_8549), .Z0_t (keyStateIn[7]), .Z0_f (new_AGEMA_signal_3495), .Z1_t (new_AGEMA_signal_3496), .Z1_f (new_AGEMA_signal_3497) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_7_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (keyStateIn[7]), .B0_f (new_AGEMA_signal_3495), .B1_t (new_AGEMA_signal_3496), .B1_f (new_AGEMA_signal_3497), .Z0_t (KeyArray_S00reg_gff_1_SFF_7_n1), .Z0_f (new_AGEMA_signal_8547), .Z1_t (new_AGEMA_signal_8548), .Z1_f (new_AGEMA_signal_8549) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_7_U1 ( .A0_t (KeyArray_S00reg_gff_1_SFF_7_QD), .A0_f (new_AGEMA_signal_10922), .A1_t (new_AGEMA_signal_10923), .A1_f (new_AGEMA_signal_10924), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S00reg_gff_1_SFF_7_n2), .Z0_f (new_AGEMA_signal_11033), .Z1_t (new_AGEMA_signal_11034), .Z1_f (new_AGEMA_signal_11035) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS00ser[7]), .A0_f (new_AGEMA_signal_10523), .A1_t (new_AGEMA_signal_10524), .A1_f (new_AGEMA_signal_10525), .B0_t (KeyArray_outS10ser[7]), .B0_f (new_AGEMA_signal_4644), .B1_t (new_AGEMA_signal_4645), .B1_f (new_AGEMA_signal_4646), .Z0_t (KeyArray_S00reg_gff_1_SFF_7_MUXInst_X), .Z0_f (new_AGEMA_signal_10679), .Z1_t (new_AGEMA_signal_10680), .Z1_f (new_AGEMA_signal_10681) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S00reg_gff_1_SFF_7_MUXInst_X), .B0_f (new_AGEMA_signal_10679), .B1_t (new_AGEMA_signal_10680), .B1_f (new_AGEMA_signal_10681), .Z0_t (KeyArray_S00reg_gff_1_SFF_7_MUXInst_Y), .Z0_f (new_AGEMA_signal_10814), .Z1_t (new_AGEMA_signal_10815), .Z1_f (new_AGEMA_signal_10816) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S00reg_gff_1_SFF_7_MUXInst_Y), .A0_f (new_AGEMA_signal_10814), .A1_t (new_AGEMA_signal_10815), .A1_f (new_AGEMA_signal_10816), .B0_t (KeyArray_inS00ser[7]), .B0_f (new_AGEMA_signal_10523), .B1_t (new_AGEMA_signal_10524), .B1_f (new_AGEMA_signal_10525), .Z0_t (KeyArray_S00reg_gff_1_SFF_7_QD), .Z0_f (new_AGEMA_signal_10922), .Z1_t (new_AGEMA_signal_10923), .Z1_f (new_AGEMA_signal_10924) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S01reg_gff_1_SFF_0_U3 ( .A0_t (KeyArray_S01reg_gff_1_SFF_0_n2), .A0_f (new_AGEMA_signal_9876), .A1_t (new_AGEMA_signal_9877), .A1_f (new_AGEMA_signal_9878), .B0_t (KeyArray_S01reg_gff_1_SFF_0_n1), .B0_f (new_AGEMA_signal_8550), .B1_t (new_AGEMA_signal_8551), .B1_f (new_AGEMA_signal_8552), .Z0_t (KeyArray_outS01ser_0_), .Z0_f (new_AGEMA_signal_4428), .Z1_t (new_AGEMA_signal_4429), .Z1_f (new_AGEMA_signal_4430) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_0_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS01ser_0_), .B0_f (new_AGEMA_signal_4428), .B1_t (new_AGEMA_signal_4429), .B1_f (new_AGEMA_signal_4430), .Z0_t (KeyArray_S01reg_gff_1_SFF_0_n1), .Z0_f (new_AGEMA_signal_8550), .Z1_t (new_AGEMA_signal_8551), .Z1_f (new_AGEMA_signal_8552) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_0_U1 ( .A0_t (KeyArray_S01reg_gff_1_SFF_0_QD), .A0_f (new_AGEMA_signal_9400), .A1_t (new_AGEMA_signal_9401), .A1_f (new_AGEMA_signal_9402), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S01reg_gff_1_SFF_0_n2), .Z0_f (new_AGEMA_signal_9876), .Z1_t (new_AGEMA_signal_9877), .Z1_f (new_AGEMA_signal_9878) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS01ser[0]), .A0_f (new_AGEMA_signal_6910), .A1_t (new_AGEMA_signal_6911), .A1_f (new_AGEMA_signal_6912), .B0_t (KeyArray_outS11ser[0]), .B0_f (new_AGEMA_signal_4653), .B1_t (new_AGEMA_signal_4654), .B1_f (new_AGEMA_signal_4655), .Z0_t (KeyArray_S01reg_gff_1_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_7743), .Z1_t (new_AGEMA_signal_7744), .Z1_f (new_AGEMA_signal_7745) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S01reg_gff_1_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_7743), .B1_t (new_AGEMA_signal_7744), .B1_f (new_AGEMA_signal_7745), .Z0_t (KeyArray_S01reg_gff_1_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_8553), .Z1_t (new_AGEMA_signal_8554), .Z1_f (new_AGEMA_signal_8555) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S01reg_gff_1_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_8553), .A1_t (new_AGEMA_signal_8554), .A1_f (new_AGEMA_signal_8555), .B0_t (KeyArray_inS01ser[0]), .B0_f (new_AGEMA_signal_6910), .B1_t (new_AGEMA_signal_6911), .B1_f (new_AGEMA_signal_6912), .Z0_t (KeyArray_S01reg_gff_1_SFF_0_QD), .Z0_f (new_AGEMA_signal_9400), .Z1_t (new_AGEMA_signal_9401), .Z1_f (new_AGEMA_signal_9402) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S01reg_gff_1_SFF_1_U3 ( .A0_t (KeyArray_S01reg_gff_1_SFF_1_n2), .A0_f (new_AGEMA_signal_9879), .A1_t (new_AGEMA_signal_9880), .A1_f (new_AGEMA_signal_9881), .B0_t (KeyArray_S01reg_gff_1_SFF_1_n1), .B0_f (new_AGEMA_signal_8556), .B1_t (new_AGEMA_signal_8557), .B1_f (new_AGEMA_signal_8558), .Z0_t (KeyArray_outS01ser_1_), .Z0_f (new_AGEMA_signal_4422), .Z1_t (new_AGEMA_signal_4423), .Z1_f (new_AGEMA_signal_4424) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_1_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS01ser_1_), .B0_f (new_AGEMA_signal_4422), .B1_t (new_AGEMA_signal_4423), .B1_f (new_AGEMA_signal_4424), .Z0_t (KeyArray_S01reg_gff_1_SFF_1_n1), .Z0_f (new_AGEMA_signal_8556), .Z1_t (new_AGEMA_signal_8557), .Z1_f (new_AGEMA_signal_8558) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_1_U1 ( .A0_t (KeyArray_S01reg_gff_1_SFF_1_QD), .A0_f (new_AGEMA_signal_9403), .A1_t (new_AGEMA_signal_9404), .A1_f (new_AGEMA_signal_9405), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S01reg_gff_1_SFF_1_n2), .Z0_f (new_AGEMA_signal_9879), .Z1_t (new_AGEMA_signal_9880), .Z1_f (new_AGEMA_signal_9881) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS01ser[1]), .A0_f (new_AGEMA_signal_6913), .A1_t (new_AGEMA_signal_6914), .A1_f (new_AGEMA_signal_6915), .B0_t (KeyArray_outS11ser[1]), .B0_f (new_AGEMA_signal_4662), .B1_t (new_AGEMA_signal_4663), .B1_f (new_AGEMA_signal_4664), .Z0_t (KeyArray_S01reg_gff_1_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_7746), .Z1_t (new_AGEMA_signal_7747), .Z1_f (new_AGEMA_signal_7748) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S01reg_gff_1_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_7746), .B1_t (new_AGEMA_signal_7747), .B1_f (new_AGEMA_signal_7748), .Z0_t (KeyArray_S01reg_gff_1_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_8559), .Z1_t (new_AGEMA_signal_8560), .Z1_f (new_AGEMA_signal_8561) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S01reg_gff_1_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_8559), .A1_t (new_AGEMA_signal_8560), .A1_f (new_AGEMA_signal_8561), .B0_t (KeyArray_inS01ser[1]), .B0_f (new_AGEMA_signal_6913), .B1_t (new_AGEMA_signal_6914), .B1_f (new_AGEMA_signal_6915), .Z0_t (KeyArray_S01reg_gff_1_SFF_1_QD), .Z0_f (new_AGEMA_signal_9403), .Z1_t (new_AGEMA_signal_9404), .Z1_f (new_AGEMA_signal_9405) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S01reg_gff_1_SFF_2_U3 ( .A0_t (KeyArray_S01reg_gff_1_SFF_2_n2), .A0_f (new_AGEMA_signal_9882), .A1_t (new_AGEMA_signal_9883), .A1_f (new_AGEMA_signal_9884), .B0_t (KeyArray_S01reg_gff_1_SFF_2_n1), .B0_f (new_AGEMA_signal_8562), .B1_t (new_AGEMA_signal_8563), .B1_f (new_AGEMA_signal_8564), .Z0_t (KeyArray_outS01ser_2_), .Z0_f (new_AGEMA_signal_4416), .Z1_t (new_AGEMA_signal_4417), .Z1_f (new_AGEMA_signal_4418) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_2_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS01ser_2_), .B0_f (new_AGEMA_signal_4416), .B1_t (new_AGEMA_signal_4417), .B1_f (new_AGEMA_signal_4418), .Z0_t (KeyArray_S01reg_gff_1_SFF_2_n1), .Z0_f (new_AGEMA_signal_8562), .Z1_t (new_AGEMA_signal_8563), .Z1_f (new_AGEMA_signal_8564) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_2_U1 ( .A0_t (KeyArray_S01reg_gff_1_SFF_2_QD), .A0_f (new_AGEMA_signal_9406), .A1_t (new_AGEMA_signal_9407), .A1_f (new_AGEMA_signal_9408), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S01reg_gff_1_SFF_2_n2), .Z0_f (new_AGEMA_signal_9882), .Z1_t (new_AGEMA_signal_9883), .Z1_f (new_AGEMA_signal_9884) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS01ser[2]), .A0_f (new_AGEMA_signal_6916), .A1_t (new_AGEMA_signal_6917), .A1_f (new_AGEMA_signal_6918), .B0_t (KeyArray_outS11ser[2]), .B0_f (new_AGEMA_signal_4671), .B1_t (new_AGEMA_signal_4672), .B1_f (new_AGEMA_signal_4673), .Z0_t (KeyArray_S01reg_gff_1_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_7749), .Z1_t (new_AGEMA_signal_7750), .Z1_f (new_AGEMA_signal_7751) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S01reg_gff_1_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_7749), .B1_t (new_AGEMA_signal_7750), .B1_f (new_AGEMA_signal_7751), .Z0_t (KeyArray_S01reg_gff_1_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_8565), .Z1_t (new_AGEMA_signal_8566), .Z1_f (new_AGEMA_signal_8567) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S01reg_gff_1_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_8565), .A1_t (new_AGEMA_signal_8566), .A1_f (new_AGEMA_signal_8567), .B0_t (KeyArray_inS01ser[2]), .B0_f (new_AGEMA_signal_6916), .B1_t (new_AGEMA_signal_6917), .B1_f (new_AGEMA_signal_6918), .Z0_t (KeyArray_S01reg_gff_1_SFF_2_QD), .Z0_f (new_AGEMA_signal_9406), .Z1_t (new_AGEMA_signal_9407), .Z1_f (new_AGEMA_signal_9408) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S01reg_gff_1_SFF_3_U3 ( .A0_t (KeyArray_S01reg_gff_1_SFF_3_n2), .A0_f (new_AGEMA_signal_9885), .A1_t (new_AGEMA_signal_9886), .A1_f (new_AGEMA_signal_9887), .B0_t (KeyArray_S01reg_gff_1_SFF_3_n1), .B0_f (new_AGEMA_signal_8568), .B1_t (new_AGEMA_signal_8569), .B1_f (new_AGEMA_signal_8570), .Z0_t (KeyArray_outS01ser_3_), .Z0_f (new_AGEMA_signal_4410), .Z1_t (new_AGEMA_signal_4411), .Z1_f (new_AGEMA_signal_4412) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_3_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS01ser_3_), .B0_f (new_AGEMA_signal_4410), .B1_t (new_AGEMA_signal_4411), .B1_f (new_AGEMA_signal_4412), .Z0_t (KeyArray_S01reg_gff_1_SFF_3_n1), .Z0_f (new_AGEMA_signal_8568), .Z1_t (new_AGEMA_signal_8569), .Z1_f (new_AGEMA_signal_8570) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_3_U1 ( .A0_t (KeyArray_S01reg_gff_1_SFF_3_QD), .A0_f (new_AGEMA_signal_9409), .A1_t (new_AGEMA_signal_9410), .A1_f (new_AGEMA_signal_9411), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S01reg_gff_1_SFF_3_n2), .Z0_f (new_AGEMA_signal_9885), .Z1_t (new_AGEMA_signal_9886), .Z1_f (new_AGEMA_signal_9887) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS01ser[3]), .A0_f (new_AGEMA_signal_6919), .A1_t (new_AGEMA_signal_6920), .A1_f (new_AGEMA_signal_6921), .B0_t (KeyArray_outS11ser[3]), .B0_f (new_AGEMA_signal_4680), .B1_t (new_AGEMA_signal_4681), .B1_f (new_AGEMA_signal_4682), .Z0_t (KeyArray_S01reg_gff_1_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_7752), .Z1_t (new_AGEMA_signal_7753), .Z1_f (new_AGEMA_signal_7754) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S01reg_gff_1_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_7752), .B1_t (new_AGEMA_signal_7753), .B1_f (new_AGEMA_signal_7754), .Z0_t (KeyArray_S01reg_gff_1_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_8571), .Z1_t (new_AGEMA_signal_8572), .Z1_f (new_AGEMA_signal_8573) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S01reg_gff_1_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_8571), .A1_t (new_AGEMA_signal_8572), .A1_f (new_AGEMA_signal_8573), .B0_t (KeyArray_inS01ser[3]), .B0_f (new_AGEMA_signal_6919), .B1_t (new_AGEMA_signal_6920), .B1_f (new_AGEMA_signal_6921), .Z0_t (KeyArray_S01reg_gff_1_SFF_3_QD), .Z0_f (new_AGEMA_signal_9409), .Z1_t (new_AGEMA_signal_9410), .Z1_f (new_AGEMA_signal_9411) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S01reg_gff_1_SFF_4_U3 ( .A0_t (KeyArray_S01reg_gff_1_SFF_4_n2), .A0_f (new_AGEMA_signal_9888), .A1_t (new_AGEMA_signal_9889), .A1_f (new_AGEMA_signal_9890), .B0_t (KeyArray_S01reg_gff_1_SFF_4_n1), .B0_f (new_AGEMA_signal_8574), .B1_t (new_AGEMA_signal_8575), .B1_f (new_AGEMA_signal_8576), .Z0_t (KeyArray_outS01ser_4_), .Z0_f (new_AGEMA_signal_4404), .Z1_t (new_AGEMA_signal_4405), .Z1_f (new_AGEMA_signal_4406) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_4_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS01ser_4_), .B0_f (new_AGEMA_signal_4404), .B1_t (new_AGEMA_signal_4405), .B1_f (new_AGEMA_signal_4406), .Z0_t (KeyArray_S01reg_gff_1_SFF_4_n1), .Z0_f (new_AGEMA_signal_8574), .Z1_t (new_AGEMA_signal_8575), .Z1_f (new_AGEMA_signal_8576) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_4_U1 ( .A0_t (KeyArray_S01reg_gff_1_SFF_4_QD), .A0_f (new_AGEMA_signal_9412), .A1_t (new_AGEMA_signal_9413), .A1_f (new_AGEMA_signal_9414), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S01reg_gff_1_SFF_4_n2), .Z0_f (new_AGEMA_signal_9888), .Z1_t (new_AGEMA_signal_9889), .Z1_f (new_AGEMA_signal_9890) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS01ser[4]), .A0_f (new_AGEMA_signal_6922), .A1_t (new_AGEMA_signal_6923), .A1_f (new_AGEMA_signal_6924), .B0_t (KeyArray_outS11ser[4]), .B0_f (new_AGEMA_signal_4689), .B1_t (new_AGEMA_signal_4690), .B1_f (new_AGEMA_signal_4691), .Z0_t (KeyArray_S01reg_gff_1_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_7755), .Z1_t (new_AGEMA_signal_7756), .Z1_f (new_AGEMA_signal_7757) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S01reg_gff_1_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_7755), .B1_t (new_AGEMA_signal_7756), .B1_f (new_AGEMA_signal_7757), .Z0_t (KeyArray_S01reg_gff_1_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_8577), .Z1_t (new_AGEMA_signal_8578), .Z1_f (new_AGEMA_signal_8579) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S01reg_gff_1_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_8577), .A1_t (new_AGEMA_signal_8578), .A1_f (new_AGEMA_signal_8579), .B0_t (KeyArray_inS01ser[4]), .B0_f (new_AGEMA_signal_6922), .B1_t (new_AGEMA_signal_6923), .B1_f (new_AGEMA_signal_6924), .Z0_t (KeyArray_S01reg_gff_1_SFF_4_QD), .Z0_f (new_AGEMA_signal_9412), .Z1_t (new_AGEMA_signal_9413), .Z1_f (new_AGEMA_signal_9414) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S01reg_gff_1_SFF_5_U3 ( .A0_t (KeyArray_S01reg_gff_1_SFF_5_n2), .A0_f (new_AGEMA_signal_9891), .A1_t (new_AGEMA_signal_9892), .A1_f (new_AGEMA_signal_9893), .B0_t (KeyArray_S01reg_gff_1_SFF_5_n1), .B0_f (new_AGEMA_signal_8580), .B1_t (new_AGEMA_signal_8581), .B1_f (new_AGEMA_signal_8582), .Z0_t (KeyArray_outS01ser_5_), .Z0_f (new_AGEMA_signal_4398), .Z1_t (new_AGEMA_signal_4399), .Z1_f (new_AGEMA_signal_4400) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_5_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS01ser_5_), .B0_f (new_AGEMA_signal_4398), .B1_t (new_AGEMA_signal_4399), .B1_f (new_AGEMA_signal_4400), .Z0_t (KeyArray_S01reg_gff_1_SFF_5_n1), .Z0_f (new_AGEMA_signal_8580), .Z1_t (new_AGEMA_signal_8581), .Z1_f (new_AGEMA_signal_8582) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_5_U1 ( .A0_t (KeyArray_S01reg_gff_1_SFF_5_QD), .A0_f (new_AGEMA_signal_9415), .A1_t (new_AGEMA_signal_9416), .A1_f (new_AGEMA_signal_9417), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S01reg_gff_1_SFF_5_n2), .Z0_f (new_AGEMA_signal_9891), .Z1_t (new_AGEMA_signal_9892), .Z1_f (new_AGEMA_signal_9893) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS01ser[5]), .A0_f (new_AGEMA_signal_6925), .A1_t (new_AGEMA_signal_6926), .A1_f (new_AGEMA_signal_6927), .B0_t (KeyArray_outS11ser[5]), .B0_f (new_AGEMA_signal_4698), .B1_t (new_AGEMA_signal_4699), .B1_f (new_AGEMA_signal_4700), .Z0_t (KeyArray_S01reg_gff_1_SFF_5_MUXInst_X), .Z0_f (new_AGEMA_signal_7758), .Z1_t (new_AGEMA_signal_7759), .Z1_f (new_AGEMA_signal_7760) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S01reg_gff_1_SFF_5_MUXInst_X), .B0_f (new_AGEMA_signal_7758), .B1_t (new_AGEMA_signal_7759), .B1_f (new_AGEMA_signal_7760), .Z0_t (KeyArray_S01reg_gff_1_SFF_5_MUXInst_Y), .Z0_f (new_AGEMA_signal_8583), .Z1_t (new_AGEMA_signal_8584), .Z1_f (new_AGEMA_signal_8585) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S01reg_gff_1_SFF_5_MUXInst_Y), .A0_f (new_AGEMA_signal_8583), .A1_t (new_AGEMA_signal_8584), .A1_f (new_AGEMA_signal_8585), .B0_t (KeyArray_inS01ser[5]), .B0_f (new_AGEMA_signal_6925), .B1_t (new_AGEMA_signal_6926), .B1_f (new_AGEMA_signal_6927), .Z0_t (KeyArray_S01reg_gff_1_SFF_5_QD), .Z0_f (new_AGEMA_signal_9415), .Z1_t (new_AGEMA_signal_9416), .Z1_f (new_AGEMA_signal_9417) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S01reg_gff_1_SFF_6_U3 ( .A0_t (KeyArray_S01reg_gff_1_SFF_6_n2), .A0_f (new_AGEMA_signal_9894), .A1_t (new_AGEMA_signal_9895), .A1_f (new_AGEMA_signal_9896), .B0_t (KeyArray_S01reg_gff_1_SFF_6_n1), .B0_f (new_AGEMA_signal_8586), .B1_t (new_AGEMA_signal_8587), .B1_f (new_AGEMA_signal_8588), .Z0_t (KeyArray_outS01ser_6_), .Z0_f (new_AGEMA_signal_4392), .Z1_t (new_AGEMA_signal_4393), .Z1_f (new_AGEMA_signal_4394) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_6_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS01ser_6_), .B0_f (new_AGEMA_signal_4392), .B1_t (new_AGEMA_signal_4393), .B1_f (new_AGEMA_signal_4394), .Z0_t (KeyArray_S01reg_gff_1_SFF_6_n1), .Z0_f (new_AGEMA_signal_8586), .Z1_t (new_AGEMA_signal_8587), .Z1_f (new_AGEMA_signal_8588) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_6_U1 ( .A0_t (KeyArray_S01reg_gff_1_SFF_6_QD), .A0_f (new_AGEMA_signal_9418), .A1_t (new_AGEMA_signal_9419), .A1_f (new_AGEMA_signal_9420), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S01reg_gff_1_SFF_6_n2), .Z0_f (new_AGEMA_signal_9894), .Z1_t (new_AGEMA_signal_9895), .Z1_f (new_AGEMA_signal_9896) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS01ser[6]), .A0_f (new_AGEMA_signal_6928), .A1_t (new_AGEMA_signal_6929), .A1_f (new_AGEMA_signal_6930), .B0_t (KeyArray_outS11ser[6]), .B0_f (new_AGEMA_signal_4707), .B1_t (new_AGEMA_signal_4708), .B1_f (new_AGEMA_signal_4709), .Z0_t (KeyArray_S01reg_gff_1_SFF_6_MUXInst_X), .Z0_f (new_AGEMA_signal_7761), .Z1_t (new_AGEMA_signal_7762), .Z1_f (new_AGEMA_signal_7763) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S01reg_gff_1_SFF_6_MUXInst_X), .B0_f (new_AGEMA_signal_7761), .B1_t (new_AGEMA_signal_7762), .B1_f (new_AGEMA_signal_7763), .Z0_t (KeyArray_S01reg_gff_1_SFF_6_MUXInst_Y), .Z0_f (new_AGEMA_signal_8589), .Z1_t (new_AGEMA_signal_8590), .Z1_f (new_AGEMA_signal_8591) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S01reg_gff_1_SFF_6_MUXInst_Y), .A0_f (new_AGEMA_signal_8589), .A1_t (new_AGEMA_signal_8590), .A1_f (new_AGEMA_signal_8591), .B0_t (KeyArray_inS01ser[6]), .B0_f (new_AGEMA_signal_6928), .B1_t (new_AGEMA_signal_6929), .B1_f (new_AGEMA_signal_6930), .Z0_t (KeyArray_S01reg_gff_1_SFF_6_QD), .Z0_f (new_AGEMA_signal_9418), .Z1_t (new_AGEMA_signal_9419), .Z1_f (new_AGEMA_signal_9420) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S01reg_gff_1_SFF_7_U3 ( .A0_t (KeyArray_S01reg_gff_1_SFF_7_n2), .A0_f (new_AGEMA_signal_9897), .A1_t (new_AGEMA_signal_9898), .A1_f (new_AGEMA_signal_9899), .B0_t (KeyArray_S01reg_gff_1_SFF_7_n1), .B0_f (new_AGEMA_signal_8592), .B1_t (new_AGEMA_signal_8593), .B1_f (new_AGEMA_signal_8594), .Z0_t (KeyArray_outS01ser_7_), .Z0_f (new_AGEMA_signal_4386), .Z1_t (new_AGEMA_signal_4387), .Z1_f (new_AGEMA_signal_4388) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_7_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS01ser_7_), .B0_f (new_AGEMA_signal_4386), .B1_t (new_AGEMA_signal_4387), .B1_f (new_AGEMA_signal_4388), .Z0_t (KeyArray_S01reg_gff_1_SFF_7_n1), .Z0_f (new_AGEMA_signal_8592), .Z1_t (new_AGEMA_signal_8593), .Z1_f (new_AGEMA_signal_8594) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_7_U1 ( .A0_t (KeyArray_S01reg_gff_1_SFF_7_QD), .A0_f (new_AGEMA_signal_9421), .A1_t (new_AGEMA_signal_9422), .A1_f (new_AGEMA_signal_9423), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S01reg_gff_1_SFF_7_n2), .Z0_f (new_AGEMA_signal_9897), .Z1_t (new_AGEMA_signal_9898), .Z1_f (new_AGEMA_signal_9899) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS01ser[7]), .A0_f (new_AGEMA_signal_6931), .A1_t (new_AGEMA_signal_6932), .A1_f (new_AGEMA_signal_6933), .B0_t (KeyArray_outS11ser[7]), .B0_f (new_AGEMA_signal_4716), .B1_t (new_AGEMA_signal_4717), .B1_f (new_AGEMA_signal_4718), .Z0_t (KeyArray_S01reg_gff_1_SFF_7_MUXInst_X), .Z0_f (new_AGEMA_signal_7764), .Z1_t (new_AGEMA_signal_7765), .Z1_f (new_AGEMA_signal_7766) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S01reg_gff_1_SFF_7_MUXInst_X), .B0_f (new_AGEMA_signal_7764), .B1_t (new_AGEMA_signal_7765), .B1_f (new_AGEMA_signal_7766), .Z0_t (KeyArray_S01reg_gff_1_SFF_7_MUXInst_Y), .Z0_f (new_AGEMA_signal_8595), .Z1_t (new_AGEMA_signal_8596), .Z1_f (new_AGEMA_signal_8597) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S01reg_gff_1_SFF_7_MUXInst_Y), .A0_f (new_AGEMA_signal_8595), .A1_t (new_AGEMA_signal_8596), .A1_f (new_AGEMA_signal_8597), .B0_t (KeyArray_inS01ser[7]), .B0_f (new_AGEMA_signal_6931), .B1_t (new_AGEMA_signal_6932), .B1_f (new_AGEMA_signal_6933), .Z0_t (KeyArray_S01reg_gff_1_SFF_7_QD), .Z0_f (new_AGEMA_signal_9421), .Z1_t (new_AGEMA_signal_9422), .Z1_f (new_AGEMA_signal_9423) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S02reg_gff_1_SFF_0_U3 ( .A0_t (KeyArray_S02reg_gff_1_SFF_0_n2), .A0_f (new_AGEMA_signal_9900), .A1_t (new_AGEMA_signal_9901), .A1_f (new_AGEMA_signal_9902), .B0_t (KeyArray_S02reg_gff_1_SFF_0_n1), .B0_f (new_AGEMA_signal_8598), .B1_t (new_AGEMA_signal_8599), .B1_f (new_AGEMA_signal_8600), .Z0_t (KeyArray_outS02ser[0]), .Z0_f (new_AGEMA_signal_4437), .Z1_t (new_AGEMA_signal_4438), .Z1_f (new_AGEMA_signal_4439) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_0_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS02ser[0]), .B0_f (new_AGEMA_signal_4437), .B1_t (new_AGEMA_signal_4438), .B1_f (new_AGEMA_signal_4439), .Z0_t (KeyArray_S02reg_gff_1_SFF_0_n1), .Z0_f (new_AGEMA_signal_8598), .Z1_t (new_AGEMA_signal_8599), .Z1_f (new_AGEMA_signal_8600) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_0_U1 ( .A0_t (KeyArray_S02reg_gff_1_SFF_0_QD), .A0_f (new_AGEMA_signal_9424), .A1_t (new_AGEMA_signal_9425), .A1_f (new_AGEMA_signal_9426), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S02reg_gff_1_SFF_0_n2), .Z0_f (new_AGEMA_signal_9900), .Z1_t (new_AGEMA_signal_9901), .Z1_f (new_AGEMA_signal_9902) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS02ser[0]), .A0_f (new_AGEMA_signal_6934), .A1_t (new_AGEMA_signal_6935), .A1_f (new_AGEMA_signal_6936), .B0_t (KeyArray_outS12ser[0]), .B0_f (new_AGEMA_signal_4725), .B1_t (new_AGEMA_signal_4726), .B1_f (new_AGEMA_signal_4727), .Z0_t (KeyArray_S02reg_gff_1_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_7767), .Z1_t (new_AGEMA_signal_7768), .Z1_f (new_AGEMA_signal_7769) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S02reg_gff_1_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_7767), .B1_t (new_AGEMA_signal_7768), .B1_f (new_AGEMA_signal_7769), .Z0_t (KeyArray_S02reg_gff_1_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_8601), .Z1_t (new_AGEMA_signal_8602), .Z1_f (new_AGEMA_signal_8603) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S02reg_gff_1_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_8601), .A1_t (new_AGEMA_signal_8602), .A1_f (new_AGEMA_signal_8603), .B0_t (KeyArray_inS02ser[0]), .B0_f (new_AGEMA_signal_6934), .B1_t (new_AGEMA_signal_6935), .B1_f (new_AGEMA_signal_6936), .Z0_t (KeyArray_S02reg_gff_1_SFF_0_QD), .Z0_f (new_AGEMA_signal_9424), .Z1_t (new_AGEMA_signal_9425), .Z1_f (new_AGEMA_signal_9426) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S02reg_gff_1_SFF_1_U3 ( .A0_t (KeyArray_S02reg_gff_1_SFF_1_n2), .A0_f (new_AGEMA_signal_9903), .A1_t (new_AGEMA_signal_9904), .A1_f (new_AGEMA_signal_9905), .B0_t (KeyArray_S02reg_gff_1_SFF_1_n1), .B0_f (new_AGEMA_signal_8604), .B1_t (new_AGEMA_signal_8605), .B1_f (new_AGEMA_signal_8606), .Z0_t (KeyArray_outS02ser[1]), .Z0_f (new_AGEMA_signal_4446), .Z1_t (new_AGEMA_signal_4447), .Z1_f (new_AGEMA_signal_4448) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_1_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS02ser[1]), .B0_f (new_AGEMA_signal_4446), .B1_t (new_AGEMA_signal_4447), .B1_f (new_AGEMA_signal_4448), .Z0_t (KeyArray_S02reg_gff_1_SFF_1_n1), .Z0_f (new_AGEMA_signal_8604), .Z1_t (new_AGEMA_signal_8605), .Z1_f (new_AGEMA_signal_8606) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_1_U1 ( .A0_t (KeyArray_S02reg_gff_1_SFF_1_QD), .A0_f (new_AGEMA_signal_9427), .A1_t (new_AGEMA_signal_9428), .A1_f (new_AGEMA_signal_9429), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S02reg_gff_1_SFF_1_n2), .Z0_f (new_AGEMA_signal_9903), .Z1_t (new_AGEMA_signal_9904), .Z1_f (new_AGEMA_signal_9905) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS02ser[1]), .A0_f (new_AGEMA_signal_6937), .A1_t (new_AGEMA_signal_6938), .A1_f (new_AGEMA_signal_6939), .B0_t (KeyArray_outS12ser[1]), .B0_f (new_AGEMA_signal_4734), .B1_t (new_AGEMA_signal_4735), .B1_f (new_AGEMA_signal_4736), .Z0_t (KeyArray_S02reg_gff_1_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_7770), .Z1_t (new_AGEMA_signal_7771), .Z1_f (new_AGEMA_signal_7772) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S02reg_gff_1_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_7770), .B1_t (new_AGEMA_signal_7771), .B1_f (new_AGEMA_signal_7772), .Z0_t (KeyArray_S02reg_gff_1_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_8607), .Z1_t (new_AGEMA_signal_8608), .Z1_f (new_AGEMA_signal_8609) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S02reg_gff_1_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_8607), .A1_t (new_AGEMA_signal_8608), .A1_f (new_AGEMA_signal_8609), .B0_t (KeyArray_inS02ser[1]), .B0_f (new_AGEMA_signal_6937), .B1_t (new_AGEMA_signal_6938), .B1_f (new_AGEMA_signal_6939), .Z0_t (KeyArray_S02reg_gff_1_SFF_1_QD), .Z0_f (new_AGEMA_signal_9427), .Z1_t (new_AGEMA_signal_9428), .Z1_f (new_AGEMA_signal_9429) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S02reg_gff_1_SFF_2_U3 ( .A0_t (KeyArray_S02reg_gff_1_SFF_2_n2), .A0_f (new_AGEMA_signal_9906), .A1_t (new_AGEMA_signal_9907), .A1_f (new_AGEMA_signal_9908), .B0_t (KeyArray_S02reg_gff_1_SFF_2_n1), .B0_f (new_AGEMA_signal_8610), .B1_t (new_AGEMA_signal_8611), .B1_f (new_AGEMA_signal_8612), .Z0_t (KeyArray_outS02ser[2]), .Z0_f (new_AGEMA_signal_4455), .Z1_t (new_AGEMA_signal_4456), .Z1_f (new_AGEMA_signal_4457) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_2_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS02ser[2]), .B0_f (new_AGEMA_signal_4455), .B1_t (new_AGEMA_signal_4456), .B1_f (new_AGEMA_signal_4457), .Z0_t (KeyArray_S02reg_gff_1_SFF_2_n1), .Z0_f (new_AGEMA_signal_8610), .Z1_t (new_AGEMA_signal_8611), .Z1_f (new_AGEMA_signal_8612) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_2_U1 ( .A0_t (KeyArray_S02reg_gff_1_SFF_2_QD), .A0_f (new_AGEMA_signal_9430), .A1_t (new_AGEMA_signal_9431), .A1_f (new_AGEMA_signal_9432), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S02reg_gff_1_SFF_2_n2), .Z0_f (new_AGEMA_signal_9906), .Z1_t (new_AGEMA_signal_9907), .Z1_f (new_AGEMA_signal_9908) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS02ser[2]), .A0_f (new_AGEMA_signal_6940), .A1_t (new_AGEMA_signal_6941), .A1_f (new_AGEMA_signal_6942), .B0_t (KeyArray_outS12ser[2]), .B0_f (new_AGEMA_signal_4743), .B1_t (new_AGEMA_signal_4744), .B1_f (new_AGEMA_signal_4745), .Z0_t (KeyArray_S02reg_gff_1_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_7773), .Z1_t (new_AGEMA_signal_7774), .Z1_f (new_AGEMA_signal_7775) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S02reg_gff_1_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_7773), .B1_t (new_AGEMA_signal_7774), .B1_f (new_AGEMA_signal_7775), .Z0_t (KeyArray_S02reg_gff_1_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_8613), .Z1_t (new_AGEMA_signal_8614), .Z1_f (new_AGEMA_signal_8615) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S02reg_gff_1_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_8613), .A1_t (new_AGEMA_signal_8614), .A1_f (new_AGEMA_signal_8615), .B0_t (KeyArray_inS02ser[2]), .B0_f (new_AGEMA_signal_6940), .B1_t (new_AGEMA_signal_6941), .B1_f (new_AGEMA_signal_6942), .Z0_t (KeyArray_S02reg_gff_1_SFF_2_QD), .Z0_f (new_AGEMA_signal_9430), .Z1_t (new_AGEMA_signal_9431), .Z1_f (new_AGEMA_signal_9432) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S02reg_gff_1_SFF_3_U3 ( .A0_t (KeyArray_S02reg_gff_1_SFF_3_n2), .A0_f (new_AGEMA_signal_9909), .A1_t (new_AGEMA_signal_9910), .A1_f (new_AGEMA_signal_9911), .B0_t (KeyArray_S02reg_gff_1_SFF_3_n1), .B0_f (new_AGEMA_signal_8616), .B1_t (new_AGEMA_signal_8617), .B1_f (new_AGEMA_signal_8618), .Z0_t (KeyArray_outS02ser[3]), .Z0_f (new_AGEMA_signal_4464), .Z1_t (new_AGEMA_signal_4465), .Z1_f (new_AGEMA_signal_4466) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_3_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS02ser[3]), .B0_f (new_AGEMA_signal_4464), .B1_t (new_AGEMA_signal_4465), .B1_f (new_AGEMA_signal_4466), .Z0_t (KeyArray_S02reg_gff_1_SFF_3_n1), .Z0_f (new_AGEMA_signal_8616), .Z1_t (new_AGEMA_signal_8617), .Z1_f (new_AGEMA_signal_8618) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_3_U1 ( .A0_t (KeyArray_S02reg_gff_1_SFF_3_QD), .A0_f (new_AGEMA_signal_9433), .A1_t (new_AGEMA_signal_9434), .A1_f (new_AGEMA_signal_9435), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S02reg_gff_1_SFF_3_n2), .Z0_f (new_AGEMA_signal_9909), .Z1_t (new_AGEMA_signal_9910), .Z1_f (new_AGEMA_signal_9911) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS02ser[3]), .A0_f (new_AGEMA_signal_6943), .A1_t (new_AGEMA_signal_6944), .A1_f (new_AGEMA_signal_6945), .B0_t (KeyArray_outS12ser[3]), .B0_f (new_AGEMA_signal_4752), .B1_t (new_AGEMA_signal_4753), .B1_f (new_AGEMA_signal_4754), .Z0_t (KeyArray_S02reg_gff_1_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_7776), .Z1_t (new_AGEMA_signal_7777), .Z1_f (new_AGEMA_signal_7778) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S02reg_gff_1_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_7776), .B1_t (new_AGEMA_signal_7777), .B1_f (new_AGEMA_signal_7778), .Z0_t (KeyArray_S02reg_gff_1_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_8619), .Z1_t (new_AGEMA_signal_8620), .Z1_f (new_AGEMA_signal_8621) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S02reg_gff_1_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_8619), .A1_t (new_AGEMA_signal_8620), .A1_f (new_AGEMA_signal_8621), .B0_t (KeyArray_inS02ser[3]), .B0_f (new_AGEMA_signal_6943), .B1_t (new_AGEMA_signal_6944), .B1_f (new_AGEMA_signal_6945), .Z0_t (KeyArray_S02reg_gff_1_SFF_3_QD), .Z0_f (new_AGEMA_signal_9433), .Z1_t (new_AGEMA_signal_9434), .Z1_f (new_AGEMA_signal_9435) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S02reg_gff_1_SFF_4_U3 ( .A0_t (KeyArray_S02reg_gff_1_SFF_4_n2), .A0_f (new_AGEMA_signal_9912), .A1_t (new_AGEMA_signal_9913), .A1_f (new_AGEMA_signal_9914), .B0_t (KeyArray_S02reg_gff_1_SFF_4_n1), .B0_f (new_AGEMA_signal_8622), .B1_t (new_AGEMA_signal_8623), .B1_f (new_AGEMA_signal_8624), .Z0_t (KeyArray_outS02ser[4]), .Z0_f (new_AGEMA_signal_4473), .Z1_t (new_AGEMA_signal_4474), .Z1_f (new_AGEMA_signal_4475) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_4_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS02ser[4]), .B0_f (new_AGEMA_signal_4473), .B1_t (new_AGEMA_signal_4474), .B1_f (new_AGEMA_signal_4475), .Z0_t (KeyArray_S02reg_gff_1_SFF_4_n1), .Z0_f (new_AGEMA_signal_8622), .Z1_t (new_AGEMA_signal_8623), .Z1_f (new_AGEMA_signal_8624) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_4_U1 ( .A0_t (KeyArray_S02reg_gff_1_SFF_4_QD), .A0_f (new_AGEMA_signal_9436), .A1_t (new_AGEMA_signal_9437), .A1_f (new_AGEMA_signal_9438), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S02reg_gff_1_SFF_4_n2), .Z0_f (new_AGEMA_signal_9912), .Z1_t (new_AGEMA_signal_9913), .Z1_f (new_AGEMA_signal_9914) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS02ser[4]), .A0_f (new_AGEMA_signal_6946), .A1_t (new_AGEMA_signal_6947), .A1_f (new_AGEMA_signal_6948), .B0_t (KeyArray_outS12ser[4]), .B0_f (new_AGEMA_signal_4761), .B1_t (new_AGEMA_signal_4762), .B1_f (new_AGEMA_signal_4763), .Z0_t (KeyArray_S02reg_gff_1_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_7779), .Z1_t (new_AGEMA_signal_7780), .Z1_f (new_AGEMA_signal_7781) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S02reg_gff_1_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_7779), .B1_t (new_AGEMA_signal_7780), .B1_f (new_AGEMA_signal_7781), .Z0_t (KeyArray_S02reg_gff_1_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_8625), .Z1_t (new_AGEMA_signal_8626), .Z1_f (new_AGEMA_signal_8627) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S02reg_gff_1_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_8625), .A1_t (new_AGEMA_signal_8626), .A1_f (new_AGEMA_signal_8627), .B0_t (KeyArray_inS02ser[4]), .B0_f (new_AGEMA_signal_6946), .B1_t (new_AGEMA_signal_6947), .B1_f (new_AGEMA_signal_6948), .Z0_t (KeyArray_S02reg_gff_1_SFF_4_QD), .Z0_f (new_AGEMA_signal_9436), .Z1_t (new_AGEMA_signal_9437), .Z1_f (new_AGEMA_signal_9438) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S02reg_gff_1_SFF_5_U3 ( .A0_t (KeyArray_S02reg_gff_1_SFF_5_n2), .A0_f (new_AGEMA_signal_9915), .A1_t (new_AGEMA_signal_9916), .A1_f (new_AGEMA_signal_9917), .B0_t (KeyArray_S02reg_gff_1_SFF_5_n1), .B0_f (new_AGEMA_signal_8628), .B1_t (new_AGEMA_signal_8629), .B1_f (new_AGEMA_signal_8630), .Z0_t (KeyArray_outS02ser[5]), .Z0_f (new_AGEMA_signal_4482), .Z1_t (new_AGEMA_signal_4483), .Z1_f (new_AGEMA_signal_4484) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_5_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS02ser[5]), .B0_f (new_AGEMA_signal_4482), .B1_t (new_AGEMA_signal_4483), .B1_f (new_AGEMA_signal_4484), .Z0_t (KeyArray_S02reg_gff_1_SFF_5_n1), .Z0_f (new_AGEMA_signal_8628), .Z1_t (new_AGEMA_signal_8629), .Z1_f (new_AGEMA_signal_8630) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_5_U1 ( .A0_t (KeyArray_S02reg_gff_1_SFF_5_QD), .A0_f (new_AGEMA_signal_9439), .A1_t (new_AGEMA_signal_9440), .A1_f (new_AGEMA_signal_9441), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S02reg_gff_1_SFF_5_n2), .Z0_f (new_AGEMA_signal_9915), .Z1_t (new_AGEMA_signal_9916), .Z1_f (new_AGEMA_signal_9917) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS02ser[5]), .A0_f (new_AGEMA_signal_6949), .A1_t (new_AGEMA_signal_6950), .A1_f (new_AGEMA_signal_6951), .B0_t (KeyArray_outS12ser[5]), .B0_f (new_AGEMA_signal_4770), .B1_t (new_AGEMA_signal_4771), .B1_f (new_AGEMA_signal_4772), .Z0_t (KeyArray_S02reg_gff_1_SFF_5_MUXInst_X), .Z0_f (new_AGEMA_signal_7782), .Z1_t (new_AGEMA_signal_7783), .Z1_f (new_AGEMA_signal_7784) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S02reg_gff_1_SFF_5_MUXInst_X), .B0_f (new_AGEMA_signal_7782), .B1_t (new_AGEMA_signal_7783), .B1_f (new_AGEMA_signal_7784), .Z0_t (KeyArray_S02reg_gff_1_SFF_5_MUXInst_Y), .Z0_f (new_AGEMA_signal_8631), .Z1_t (new_AGEMA_signal_8632), .Z1_f (new_AGEMA_signal_8633) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S02reg_gff_1_SFF_5_MUXInst_Y), .A0_f (new_AGEMA_signal_8631), .A1_t (new_AGEMA_signal_8632), .A1_f (new_AGEMA_signal_8633), .B0_t (KeyArray_inS02ser[5]), .B0_f (new_AGEMA_signal_6949), .B1_t (new_AGEMA_signal_6950), .B1_f (new_AGEMA_signal_6951), .Z0_t (KeyArray_S02reg_gff_1_SFF_5_QD), .Z0_f (new_AGEMA_signal_9439), .Z1_t (new_AGEMA_signal_9440), .Z1_f (new_AGEMA_signal_9441) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S02reg_gff_1_SFF_6_U3 ( .A0_t (KeyArray_S02reg_gff_1_SFF_6_n2), .A0_f (new_AGEMA_signal_9918), .A1_t (new_AGEMA_signal_9919), .A1_f (new_AGEMA_signal_9920), .B0_t (KeyArray_S02reg_gff_1_SFF_6_n1), .B0_f (new_AGEMA_signal_8634), .B1_t (new_AGEMA_signal_8635), .B1_f (new_AGEMA_signal_8636), .Z0_t (KeyArray_outS02ser[6]), .Z0_f (new_AGEMA_signal_4491), .Z1_t (new_AGEMA_signal_4492), .Z1_f (new_AGEMA_signal_4493) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_6_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS02ser[6]), .B0_f (new_AGEMA_signal_4491), .B1_t (new_AGEMA_signal_4492), .B1_f (new_AGEMA_signal_4493), .Z0_t (KeyArray_S02reg_gff_1_SFF_6_n1), .Z0_f (new_AGEMA_signal_8634), .Z1_t (new_AGEMA_signal_8635), .Z1_f (new_AGEMA_signal_8636) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_6_U1 ( .A0_t (KeyArray_S02reg_gff_1_SFF_6_QD), .A0_f (new_AGEMA_signal_9442), .A1_t (new_AGEMA_signal_9443), .A1_f (new_AGEMA_signal_9444), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S02reg_gff_1_SFF_6_n2), .Z0_f (new_AGEMA_signal_9918), .Z1_t (new_AGEMA_signal_9919), .Z1_f (new_AGEMA_signal_9920) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS02ser[6]), .A0_f (new_AGEMA_signal_6952), .A1_t (new_AGEMA_signal_6953), .A1_f (new_AGEMA_signal_6954), .B0_t (KeyArray_outS12ser[6]), .B0_f (new_AGEMA_signal_4779), .B1_t (new_AGEMA_signal_4780), .B1_f (new_AGEMA_signal_4781), .Z0_t (KeyArray_S02reg_gff_1_SFF_6_MUXInst_X), .Z0_f (new_AGEMA_signal_7785), .Z1_t (new_AGEMA_signal_7786), .Z1_f (new_AGEMA_signal_7787) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S02reg_gff_1_SFF_6_MUXInst_X), .B0_f (new_AGEMA_signal_7785), .B1_t (new_AGEMA_signal_7786), .B1_f (new_AGEMA_signal_7787), .Z0_t (KeyArray_S02reg_gff_1_SFF_6_MUXInst_Y), .Z0_f (new_AGEMA_signal_8637), .Z1_t (new_AGEMA_signal_8638), .Z1_f (new_AGEMA_signal_8639) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S02reg_gff_1_SFF_6_MUXInst_Y), .A0_f (new_AGEMA_signal_8637), .A1_t (new_AGEMA_signal_8638), .A1_f (new_AGEMA_signal_8639), .B0_t (KeyArray_inS02ser[6]), .B0_f (new_AGEMA_signal_6952), .B1_t (new_AGEMA_signal_6953), .B1_f (new_AGEMA_signal_6954), .Z0_t (KeyArray_S02reg_gff_1_SFF_6_QD), .Z0_f (new_AGEMA_signal_9442), .Z1_t (new_AGEMA_signal_9443), .Z1_f (new_AGEMA_signal_9444) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S02reg_gff_1_SFF_7_U3 ( .A0_t (KeyArray_S02reg_gff_1_SFF_7_n2), .A0_f (new_AGEMA_signal_9921), .A1_t (new_AGEMA_signal_9922), .A1_f (new_AGEMA_signal_9923), .B0_t (KeyArray_S02reg_gff_1_SFF_7_n1), .B0_f (new_AGEMA_signal_8640), .B1_t (new_AGEMA_signal_8641), .B1_f (new_AGEMA_signal_8642), .Z0_t (KeyArray_outS02ser[7]), .Z0_f (new_AGEMA_signal_4500), .Z1_t (new_AGEMA_signal_4501), .Z1_f (new_AGEMA_signal_4502) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_7_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS02ser[7]), .B0_f (new_AGEMA_signal_4500), .B1_t (new_AGEMA_signal_4501), .B1_f (new_AGEMA_signal_4502), .Z0_t (KeyArray_S02reg_gff_1_SFF_7_n1), .Z0_f (new_AGEMA_signal_8640), .Z1_t (new_AGEMA_signal_8641), .Z1_f (new_AGEMA_signal_8642) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_7_U1 ( .A0_t (KeyArray_S02reg_gff_1_SFF_7_QD), .A0_f (new_AGEMA_signal_9445), .A1_t (new_AGEMA_signal_9446), .A1_f (new_AGEMA_signal_9447), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S02reg_gff_1_SFF_7_n2), .Z0_f (new_AGEMA_signal_9921), .Z1_t (new_AGEMA_signal_9922), .Z1_f (new_AGEMA_signal_9923) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS02ser[7]), .A0_f (new_AGEMA_signal_6955), .A1_t (new_AGEMA_signal_6956), .A1_f (new_AGEMA_signal_6957), .B0_t (KeyArray_outS12ser[7]), .B0_f (new_AGEMA_signal_4788), .B1_t (new_AGEMA_signal_4789), .B1_f (new_AGEMA_signal_4790), .Z0_t (KeyArray_S02reg_gff_1_SFF_7_MUXInst_X), .Z0_f (new_AGEMA_signal_7788), .Z1_t (new_AGEMA_signal_7789), .Z1_f (new_AGEMA_signal_7790) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S02reg_gff_1_SFF_7_MUXInst_X), .B0_f (new_AGEMA_signal_7788), .B1_t (new_AGEMA_signal_7789), .B1_f (new_AGEMA_signal_7790), .Z0_t (KeyArray_S02reg_gff_1_SFF_7_MUXInst_Y), .Z0_f (new_AGEMA_signal_8643), .Z1_t (new_AGEMA_signal_8644), .Z1_f (new_AGEMA_signal_8645) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S02reg_gff_1_SFF_7_MUXInst_Y), .A0_f (new_AGEMA_signal_8643), .A1_t (new_AGEMA_signal_8644), .A1_f (new_AGEMA_signal_8645), .B0_t (KeyArray_inS02ser[7]), .B0_f (new_AGEMA_signal_6955), .B1_t (new_AGEMA_signal_6956), .B1_f (new_AGEMA_signal_6957), .Z0_t (KeyArray_S02reg_gff_1_SFF_7_QD), .Z0_f (new_AGEMA_signal_9445), .Z1_t (new_AGEMA_signal_9446), .Z1_f (new_AGEMA_signal_9447) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S03reg_gff_1_SFF_0_U3 ( .A0_t (KeyArray_S03reg_gff_1_SFF_0_n2), .A0_f (new_AGEMA_signal_9924), .A1_t (new_AGEMA_signal_9925), .A1_f (new_AGEMA_signal_9926), .B0_t (KeyArray_S03reg_gff_1_SFF_0_n1), .B0_f (new_AGEMA_signal_8646), .B1_t (new_AGEMA_signal_8647), .B1_f (new_AGEMA_signal_8648), .Z0_t (KeyArray_outS03ser[0]), .Z0_f (new_AGEMA_signal_4509), .Z1_t (new_AGEMA_signal_4510), .Z1_f (new_AGEMA_signal_4511) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_0_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS03ser[0]), .B0_f (new_AGEMA_signal_4509), .B1_t (new_AGEMA_signal_4510), .B1_f (new_AGEMA_signal_4511), .Z0_t (KeyArray_S03reg_gff_1_SFF_0_n1), .Z0_f (new_AGEMA_signal_8646), .Z1_t (new_AGEMA_signal_8647), .Z1_f (new_AGEMA_signal_8648) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_0_U1 ( .A0_t (KeyArray_S03reg_gff_1_SFF_0_QD), .A0_f (new_AGEMA_signal_9448), .A1_t (new_AGEMA_signal_9449), .A1_f (new_AGEMA_signal_9450), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S03reg_gff_1_SFF_0_n2), .Z0_f (new_AGEMA_signal_9924), .Z1_t (new_AGEMA_signal_9925), .Z1_f (new_AGEMA_signal_9926) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS03ser[0]), .A0_f (new_AGEMA_signal_6958), .A1_t (new_AGEMA_signal_6959), .A1_f (new_AGEMA_signal_6960), .B0_t (keySBIn[0]), .B0_f (new_AGEMA_signal_4797), .B1_t (new_AGEMA_signal_4798), .B1_f (new_AGEMA_signal_4799), .Z0_t (KeyArray_S03reg_gff_1_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_7791), .Z1_t (new_AGEMA_signal_7792), .Z1_f (new_AGEMA_signal_7793) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S03reg_gff_1_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_7791), .B1_t (new_AGEMA_signal_7792), .B1_f (new_AGEMA_signal_7793), .Z0_t (KeyArray_S03reg_gff_1_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_8649), .Z1_t (new_AGEMA_signal_8650), .Z1_f (new_AGEMA_signal_8651) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S03reg_gff_1_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_8649), .A1_t (new_AGEMA_signal_8650), .A1_f (new_AGEMA_signal_8651), .B0_t (KeyArray_inS03ser[0]), .B0_f (new_AGEMA_signal_6958), .B1_t (new_AGEMA_signal_6959), .B1_f (new_AGEMA_signal_6960), .Z0_t (KeyArray_S03reg_gff_1_SFF_0_QD), .Z0_f (new_AGEMA_signal_9448), .Z1_t (new_AGEMA_signal_9449), .Z1_f (new_AGEMA_signal_9450) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S03reg_gff_1_SFF_1_U3 ( .A0_t (KeyArray_S03reg_gff_1_SFF_1_n2), .A0_f (new_AGEMA_signal_9927), .A1_t (new_AGEMA_signal_9928), .A1_f (new_AGEMA_signal_9929), .B0_t (KeyArray_S03reg_gff_1_SFF_1_n1), .B0_f (new_AGEMA_signal_8652), .B1_t (new_AGEMA_signal_8653), .B1_f (new_AGEMA_signal_8654), .Z0_t (KeyArray_outS03ser[1]), .Z0_f (new_AGEMA_signal_4518), .Z1_t (new_AGEMA_signal_4519), .Z1_f (new_AGEMA_signal_4520) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_1_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS03ser[1]), .B0_f (new_AGEMA_signal_4518), .B1_t (new_AGEMA_signal_4519), .B1_f (new_AGEMA_signal_4520), .Z0_t (KeyArray_S03reg_gff_1_SFF_1_n1), .Z0_f (new_AGEMA_signal_8652), .Z1_t (new_AGEMA_signal_8653), .Z1_f (new_AGEMA_signal_8654) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_1_U1 ( .A0_t (KeyArray_S03reg_gff_1_SFF_1_QD), .A0_f (new_AGEMA_signal_9451), .A1_t (new_AGEMA_signal_9452), .A1_f (new_AGEMA_signal_9453), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S03reg_gff_1_SFF_1_n2), .Z0_f (new_AGEMA_signal_9927), .Z1_t (new_AGEMA_signal_9928), .Z1_f (new_AGEMA_signal_9929) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS03ser[1]), .A0_f (new_AGEMA_signal_6961), .A1_t (new_AGEMA_signal_6962), .A1_f (new_AGEMA_signal_6963), .B0_t (keySBIn[1]), .B0_f (new_AGEMA_signal_4806), .B1_t (new_AGEMA_signal_4807), .B1_f (new_AGEMA_signal_4808), .Z0_t (KeyArray_S03reg_gff_1_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_7794), .Z1_t (new_AGEMA_signal_7795), .Z1_f (new_AGEMA_signal_7796) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S03reg_gff_1_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_7794), .B1_t (new_AGEMA_signal_7795), .B1_f (new_AGEMA_signal_7796), .Z0_t (KeyArray_S03reg_gff_1_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_8655), .Z1_t (new_AGEMA_signal_8656), .Z1_f (new_AGEMA_signal_8657) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S03reg_gff_1_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_8655), .A1_t (new_AGEMA_signal_8656), .A1_f (new_AGEMA_signal_8657), .B0_t (KeyArray_inS03ser[1]), .B0_f (new_AGEMA_signal_6961), .B1_t (new_AGEMA_signal_6962), .B1_f (new_AGEMA_signal_6963), .Z0_t (KeyArray_S03reg_gff_1_SFF_1_QD), .Z0_f (new_AGEMA_signal_9451), .Z1_t (new_AGEMA_signal_9452), .Z1_f (new_AGEMA_signal_9453) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S03reg_gff_1_SFF_2_U3 ( .A0_t (KeyArray_S03reg_gff_1_SFF_2_n2), .A0_f (new_AGEMA_signal_9930), .A1_t (new_AGEMA_signal_9931), .A1_f (new_AGEMA_signal_9932), .B0_t (KeyArray_S03reg_gff_1_SFF_2_n1), .B0_f (new_AGEMA_signal_8658), .B1_t (new_AGEMA_signal_8659), .B1_f (new_AGEMA_signal_8660), .Z0_t (KeyArray_outS03ser[2]), .Z0_f (new_AGEMA_signal_4527), .Z1_t (new_AGEMA_signal_4528), .Z1_f (new_AGEMA_signal_4529) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_2_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS03ser[2]), .B0_f (new_AGEMA_signal_4527), .B1_t (new_AGEMA_signal_4528), .B1_f (new_AGEMA_signal_4529), .Z0_t (KeyArray_S03reg_gff_1_SFF_2_n1), .Z0_f (new_AGEMA_signal_8658), .Z1_t (new_AGEMA_signal_8659), .Z1_f (new_AGEMA_signal_8660) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_2_U1 ( .A0_t (KeyArray_S03reg_gff_1_SFF_2_QD), .A0_f (new_AGEMA_signal_9454), .A1_t (new_AGEMA_signal_9455), .A1_f (new_AGEMA_signal_9456), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S03reg_gff_1_SFF_2_n2), .Z0_f (new_AGEMA_signal_9930), .Z1_t (new_AGEMA_signal_9931), .Z1_f (new_AGEMA_signal_9932) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS03ser[2]), .A0_f (new_AGEMA_signal_6964), .A1_t (new_AGEMA_signal_6965), .A1_f (new_AGEMA_signal_6966), .B0_t (keySBIn[2]), .B0_f (new_AGEMA_signal_4815), .B1_t (new_AGEMA_signal_4816), .B1_f (new_AGEMA_signal_4817), .Z0_t (KeyArray_S03reg_gff_1_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_7797), .Z1_t (new_AGEMA_signal_7798), .Z1_f (new_AGEMA_signal_7799) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S03reg_gff_1_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_7797), .B1_t (new_AGEMA_signal_7798), .B1_f (new_AGEMA_signal_7799), .Z0_t (KeyArray_S03reg_gff_1_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_8661), .Z1_t (new_AGEMA_signal_8662), .Z1_f (new_AGEMA_signal_8663) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S03reg_gff_1_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_8661), .A1_t (new_AGEMA_signal_8662), .A1_f (new_AGEMA_signal_8663), .B0_t (KeyArray_inS03ser[2]), .B0_f (new_AGEMA_signal_6964), .B1_t (new_AGEMA_signal_6965), .B1_f (new_AGEMA_signal_6966), .Z0_t (KeyArray_S03reg_gff_1_SFF_2_QD), .Z0_f (new_AGEMA_signal_9454), .Z1_t (new_AGEMA_signal_9455), .Z1_f (new_AGEMA_signal_9456) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S03reg_gff_1_SFF_3_U3 ( .A0_t (KeyArray_S03reg_gff_1_SFF_3_n2), .A0_f (new_AGEMA_signal_9933), .A1_t (new_AGEMA_signal_9934), .A1_f (new_AGEMA_signal_9935), .B0_t (KeyArray_S03reg_gff_1_SFF_3_n1), .B0_f (new_AGEMA_signal_8664), .B1_t (new_AGEMA_signal_8665), .B1_f (new_AGEMA_signal_8666), .Z0_t (KeyArray_outS03ser[3]), .Z0_f (new_AGEMA_signal_4536), .Z1_t (new_AGEMA_signal_4537), .Z1_f (new_AGEMA_signal_4538) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_3_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS03ser[3]), .B0_f (new_AGEMA_signal_4536), .B1_t (new_AGEMA_signal_4537), .B1_f (new_AGEMA_signal_4538), .Z0_t (KeyArray_S03reg_gff_1_SFF_3_n1), .Z0_f (new_AGEMA_signal_8664), .Z1_t (new_AGEMA_signal_8665), .Z1_f (new_AGEMA_signal_8666) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_3_U1 ( .A0_t (KeyArray_S03reg_gff_1_SFF_3_QD), .A0_f (new_AGEMA_signal_9457), .A1_t (new_AGEMA_signal_9458), .A1_f (new_AGEMA_signal_9459), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S03reg_gff_1_SFF_3_n2), .Z0_f (new_AGEMA_signal_9933), .Z1_t (new_AGEMA_signal_9934), .Z1_f (new_AGEMA_signal_9935) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS03ser[3]), .A0_f (new_AGEMA_signal_6967), .A1_t (new_AGEMA_signal_6968), .A1_f (new_AGEMA_signal_6969), .B0_t (keySBIn[3]), .B0_f (new_AGEMA_signal_4824), .B1_t (new_AGEMA_signal_4825), .B1_f (new_AGEMA_signal_4826), .Z0_t (KeyArray_S03reg_gff_1_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_7800), .Z1_t (new_AGEMA_signal_7801), .Z1_f (new_AGEMA_signal_7802) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S03reg_gff_1_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_7800), .B1_t (new_AGEMA_signal_7801), .B1_f (new_AGEMA_signal_7802), .Z0_t (KeyArray_S03reg_gff_1_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_8667), .Z1_t (new_AGEMA_signal_8668), .Z1_f (new_AGEMA_signal_8669) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S03reg_gff_1_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_8667), .A1_t (new_AGEMA_signal_8668), .A1_f (new_AGEMA_signal_8669), .B0_t (KeyArray_inS03ser[3]), .B0_f (new_AGEMA_signal_6967), .B1_t (new_AGEMA_signal_6968), .B1_f (new_AGEMA_signal_6969), .Z0_t (KeyArray_S03reg_gff_1_SFF_3_QD), .Z0_f (new_AGEMA_signal_9457), .Z1_t (new_AGEMA_signal_9458), .Z1_f (new_AGEMA_signal_9459) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S03reg_gff_1_SFF_4_U3 ( .A0_t (KeyArray_S03reg_gff_1_SFF_4_n2), .A0_f (new_AGEMA_signal_9936), .A1_t (new_AGEMA_signal_9937), .A1_f (new_AGEMA_signal_9938), .B0_t (KeyArray_S03reg_gff_1_SFF_4_n1), .B0_f (new_AGEMA_signal_8670), .B1_t (new_AGEMA_signal_8671), .B1_f (new_AGEMA_signal_8672), .Z0_t (KeyArray_outS03ser[4]), .Z0_f (new_AGEMA_signal_4545), .Z1_t (new_AGEMA_signal_4546), .Z1_f (new_AGEMA_signal_4547) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_4_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS03ser[4]), .B0_f (new_AGEMA_signal_4545), .B1_t (new_AGEMA_signal_4546), .B1_f (new_AGEMA_signal_4547), .Z0_t (KeyArray_S03reg_gff_1_SFF_4_n1), .Z0_f (new_AGEMA_signal_8670), .Z1_t (new_AGEMA_signal_8671), .Z1_f (new_AGEMA_signal_8672) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_4_U1 ( .A0_t (KeyArray_S03reg_gff_1_SFF_4_QD), .A0_f (new_AGEMA_signal_9460), .A1_t (new_AGEMA_signal_9461), .A1_f (new_AGEMA_signal_9462), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S03reg_gff_1_SFF_4_n2), .Z0_f (new_AGEMA_signal_9936), .Z1_t (new_AGEMA_signal_9937), .Z1_f (new_AGEMA_signal_9938) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS03ser[4]), .A0_f (new_AGEMA_signal_6970), .A1_t (new_AGEMA_signal_6971), .A1_f (new_AGEMA_signal_6972), .B0_t (keySBIn[4]), .B0_f (new_AGEMA_signal_4833), .B1_t (new_AGEMA_signal_4834), .B1_f (new_AGEMA_signal_4835), .Z0_t (KeyArray_S03reg_gff_1_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_7803), .Z1_t (new_AGEMA_signal_7804), .Z1_f (new_AGEMA_signal_7805) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S03reg_gff_1_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_7803), .B1_t (new_AGEMA_signal_7804), .B1_f (new_AGEMA_signal_7805), .Z0_t (KeyArray_S03reg_gff_1_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_8673), .Z1_t (new_AGEMA_signal_8674), .Z1_f (new_AGEMA_signal_8675) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S03reg_gff_1_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_8673), .A1_t (new_AGEMA_signal_8674), .A1_f (new_AGEMA_signal_8675), .B0_t (KeyArray_inS03ser[4]), .B0_f (new_AGEMA_signal_6970), .B1_t (new_AGEMA_signal_6971), .B1_f (new_AGEMA_signal_6972), .Z0_t (KeyArray_S03reg_gff_1_SFF_4_QD), .Z0_f (new_AGEMA_signal_9460), .Z1_t (new_AGEMA_signal_9461), .Z1_f (new_AGEMA_signal_9462) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S03reg_gff_1_SFF_5_U3 ( .A0_t (KeyArray_S03reg_gff_1_SFF_5_n2), .A0_f (new_AGEMA_signal_9939), .A1_t (new_AGEMA_signal_9940), .A1_f (new_AGEMA_signal_9941), .B0_t (KeyArray_S03reg_gff_1_SFF_5_n1), .B0_f (new_AGEMA_signal_8676), .B1_t (new_AGEMA_signal_8677), .B1_f (new_AGEMA_signal_8678), .Z0_t (KeyArray_outS03ser[5]), .Z0_f (new_AGEMA_signal_4554), .Z1_t (new_AGEMA_signal_4555), .Z1_f (new_AGEMA_signal_4556) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_5_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS03ser[5]), .B0_f (new_AGEMA_signal_4554), .B1_t (new_AGEMA_signal_4555), .B1_f (new_AGEMA_signal_4556), .Z0_t (KeyArray_S03reg_gff_1_SFF_5_n1), .Z0_f (new_AGEMA_signal_8676), .Z1_t (new_AGEMA_signal_8677), .Z1_f (new_AGEMA_signal_8678) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_5_U1 ( .A0_t (KeyArray_S03reg_gff_1_SFF_5_QD), .A0_f (new_AGEMA_signal_9463), .A1_t (new_AGEMA_signal_9464), .A1_f (new_AGEMA_signal_9465), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S03reg_gff_1_SFF_5_n2), .Z0_f (new_AGEMA_signal_9939), .Z1_t (new_AGEMA_signal_9940), .Z1_f (new_AGEMA_signal_9941) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS03ser[5]), .A0_f (new_AGEMA_signal_6973), .A1_t (new_AGEMA_signal_6974), .A1_f (new_AGEMA_signal_6975), .B0_t (keySBIn[5]), .B0_f (new_AGEMA_signal_4842), .B1_t (new_AGEMA_signal_4843), .B1_f (new_AGEMA_signal_4844), .Z0_t (KeyArray_S03reg_gff_1_SFF_5_MUXInst_X), .Z0_f (new_AGEMA_signal_7806), .Z1_t (new_AGEMA_signal_7807), .Z1_f (new_AGEMA_signal_7808) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S03reg_gff_1_SFF_5_MUXInst_X), .B0_f (new_AGEMA_signal_7806), .B1_t (new_AGEMA_signal_7807), .B1_f (new_AGEMA_signal_7808), .Z0_t (KeyArray_S03reg_gff_1_SFF_5_MUXInst_Y), .Z0_f (new_AGEMA_signal_8679), .Z1_t (new_AGEMA_signal_8680), .Z1_f (new_AGEMA_signal_8681) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S03reg_gff_1_SFF_5_MUXInst_Y), .A0_f (new_AGEMA_signal_8679), .A1_t (new_AGEMA_signal_8680), .A1_f (new_AGEMA_signal_8681), .B0_t (KeyArray_inS03ser[5]), .B0_f (new_AGEMA_signal_6973), .B1_t (new_AGEMA_signal_6974), .B1_f (new_AGEMA_signal_6975), .Z0_t (KeyArray_S03reg_gff_1_SFF_5_QD), .Z0_f (new_AGEMA_signal_9463), .Z1_t (new_AGEMA_signal_9464), .Z1_f (new_AGEMA_signal_9465) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S03reg_gff_1_SFF_6_U3 ( .A0_t (KeyArray_S03reg_gff_1_SFF_6_n2), .A0_f (new_AGEMA_signal_9942), .A1_t (new_AGEMA_signal_9943), .A1_f (new_AGEMA_signal_9944), .B0_t (KeyArray_S03reg_gff_1_SFF_6_n1), .B0_f (new_AGEMA_signal_8682), .B1_t (new_AGEMA_signal_8683), .B1_f (new_AGEMA_signal_8684), .Z0_t (KeyArray_outS03ser[6]), .Z0_f (new_AGEMA_signal_4563), .Z1_t (new_AGEMA_signal_4564), .Z1_f (new_AGEMA_signal_4565) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_6_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS03ser[6]), .B0_f (new_AGEMA_signal_4563), .B1_t (new_AGEMA_signal_4564), .B1_f (new_AGEMA_signal_4565), .Z0_t (KeyArray_S03reg_gff_1_SFF_6_n1), .Z0_f (new_AGEMA_signal_8682), .Z1_t (new_AGEMA_signal_8683), .Z1_f (new_AGEMA_signal_8684) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_6_U1 ( .A0_t (KeyArray_S03reg_gff_1_SFF_6_QD), .A0_f (new_AGEMA_signal_9466), .A1_t (new_AGEMA_signal_9467), .A1_f (new_AGEMA_signal_9468), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S03reg_gff_1_SFF_6_n2), .Z0_f (new_AGEMA_signal_9942), .Z1_t (new_AGEMA_signal_9943), .Z1_f (new_AGEMA_signal_9944) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS03ser[6]), .A0_f (new_AGEMA_signal_6976), .A1_t (new_AGEMA_signal_6977), .A1_f (new_AGEMA_signal_6978), .B0_t (keySBIn[6]), .B0_f (new_AGEMA_signal_4851), .B1_t (new_AGEMA_signal_4852), .B1_f (new_AGEMA_signal_4853), .Z0_t (KeyArray_S03reg_gff_1_SFF_6_MUXInst_X), .Z0_f (new_AGEMA_signal_7809), .Z1_t (new_AGEMA_signal_7810), .Z1_f (new_AGEMA_signal_7811) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S03reg_gff_1_SFF_6_MUXInst_X), .B0_f (new_AGEMA_signal_7809), .B1_t (new_AGEMA_signal_7810), .B1_f (new_AGEMA_signal_7811), .Z0_t (KeyArray_S03reg_gff_1_SFF_6_MUXInst_Y), .Z0_f (new_AGEMA_signal_8685), .Z1_t (new_AGEMA_signal_8686), .Z1_f (new_AGEMA_signal_8687) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S03reg_gff_1_SFF_6_MUXInst_Y), .A0_f (new_AGEMA_signal_8685), .A1_t (new_AGEMA_signal_8686), .A1_f (new_AGEMA_signal_8687), .B0_t (KeyArray_inS03ser[6]), .B0_f (new_AGEMA_signal_6976), .B1_t (new_AGEMA_signal_6977), .B1_f (new_AGEMA_signal_6978), .Z0_t (KeyArray_S03reg_gff_1_SFF_6_QD), .Z0_f (new_AGEMA_signal_9466), .Z1_t (new_AGEMA_signal_9467), .Z1_f (new_AGEMA_signal_9468) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S03reg_gff_1_SFF_7_U3 ( .A0_t (KeyArray_S03reg_gff_1_SFF_7_n2), .A0_f (new_AGEMA_signal_9945), .A1_t (new_AGEMA_signal_9946), .A1_f (new_AGEMA_signal_9947), .B0_t (KeyArray_S03reg_gff_1_SFF_7_n1), .B0_f (new_AGEMA_signal_8688), .B1_t (new_AGEMA_signal_8689), .B1_f (new_AGEMA_signal_8690), .Z0_t (KeyArray_outS03ser[7]), .Z0_f (new_AGEMA_signal_4572), .Z1_t (new_AGEMA_signal_4573), .Z1_f (new_AGEMA_signal_4574) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_7_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS03ser[7]), .B0_f (new_AGEMA_signal_4572), .B1_t (new_AGEMA_signal_4573), .B1_f (new_AGEMA_signal_4574), .Z0_t (KeyArray_S03reg_gff_1_SFF_7_n1), .Z0_f (new_AGEMA_signal_8688), .Z1_t (new_AGEMA_signal_8689), .Z1_f (new_AGEMA_signal_8690) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_7_U1 ( .A0_t (KeyArray_S03reg_gff_1_SFF_7_QD), .A0_f (new_AGEMA_signal_9469), .A1_t (new_AGEMA_signal_9470), .A1_f (new_AGEMA_signal_9471), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S03reg_gff_1_SFF_7_n2), .Z0_f (new_AGEMA_signal_9945), .Z1_t (new_AGEMA_signal_9946), .Z1_f (new_AGEMA_signal_9947) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS03ser[7]), .A0_f (new_AGEMA_signal_6979), .A1_t (new_AGEMA_signal_6980), .A1_f (new_AGEMA_signal_6981), .B0_t (keySBIn[7]), .B0_f (new_AGEMA_signal_4860), .B1_t (new_AGEMA_signal_4861), .B1_f (new_AGEMA_signal_4862), .Z0_t (KeyArray_S03reg_gff_1_SFF_7_MUXInst_X), .Z0_f (new_AGEMA_signal_7812), .Z1_t (new_AGEMA_signal_7813), .Z1_f (new_AGEMA_signal_7814) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S03reg_gff_1_SFF_7_MUXInst_X), .B0_f (new_AGEMA_signal_7812), .B1_t (new_AGEMA_signal_7813), .B1_f (new_AGEMA_signal_7814), .Z0_t (KeyArray_S03reg_gff_1_SFF_7_MUXInst_Y), .Z0_f (new_AGEMA_signal_8691), .Z1_t (new_AGEMA_signal_8692), .Z1_f (new_AGEMA_signal_8693) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S03reg_gff_1_SFF_7_MUXInst_Y), .A0_f (new_AGEMA_signal_8691), .A1_t (new_AGEMA_signal_8692), .A1_f (new_AGEMA_signal_8693), .B0_t (KeyArray_inS03ser[7]), .B0_f (new_AGEMA_signal_6979), .B1_t (new_AGEMA_signal_6980), .B1_f (new_AGEMA_signal_6981), .Z0_t (KeyArray_S03reg_gff_1_SFF_7_QD), .Z0_f (new_AGEMA_signal_9469), .Z1_t (new_AGEMA_signal_9470), .Z1_f (new_AGEMA_signal_9471) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S10reg_gff_1_SFF_0_U3 ( .A0_t (KeyArray_S10reg_gff_1_SFF_0_n2), .A0_f (new_AGEMA_signal_9948), .A1_t (new_AGEMA_signal_9949), .A1_f (new_AGEMA_signal_9950), .B0_t (KeyArray_S10reg_gff_1_SFF_0_n1), .B0_f (new_AGEMA_signal_8694), .B1_t (new_AGEMA_signal_8695), .B1_f (new_AGEMA_signal_8696), .Z0_t (KeyArray_outS10ser[0]), .Z0_f (new_AGEMA_signal_4581), .Z1_t (new_AGEMA_signal_4582), .Z1_f (new_AGEMA_signal_4583) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_0_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS10ser[0]), .B0_f (new_AGEMA_signal_4581), .B1_t (new_AGEMA_signal_4582), .B1_f (new_AGEMA_signal_4583), .Z0_t (KeyArray_S10reg_gff_1_SFF_0_n1), .Z0_f (new_AGEMA_signal_8694), .Z1_t (new_AGEMA_signal_8695), .Z1_f (new_AGEMA_signal_8696) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_0_U1 ( .A0_t (KeyArray_S10reg_gff_1_SFF_0_QD), .A0_f (new_AGEMA_signal_9472), .A1_t (new_AGEMA_signal_9473), .A1_f (new_AGEMA_signal_9474), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S10reg_gff_1_SFF_0_n2), .Z0_f (new_AGEMA_signal_9948), .Z1_t (new_AGEMA_signal_9949), .Z1_f (new_AGEMA_signal_9950) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS10ser[0]), .A0_f (new_AGEMA_signal_6982), .A1_t (new_AGEMA_signal_6983), .A1_f (new_AGEMA_signal_6984), .B0_t (KeyArray_outS20ser[0]), .B0_f (new_AGEMA_signal_4869), .B1_t (new_AGEMA_signal_4870), .B1_f (new_AGEMA_signal_4871), .Z0_t (KeyArray_S10reg_gff_1_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_7815), .Z1_t (new_AGEMA_signal_7816), .Z1_f (new_AGEMA_signal_7817) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S10reg_gff_1_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_7815), .B1_t (new_AGEMA_signal_7816), .B1_f (new_AGEMA_signal_7817), .Z0_t (KeyArray_S10reg_gff_1_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_8697), .Z1_t (new_AGEMA_signal_8698), .Z1_f (new_AGEMA_signal_8699) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S10reg_gff_1_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_8697), .A1_t (new_AGEMA_signal_8698), .A1_f (new_AGEMA_signal_8699), .B0_t (KeyArray_inS10ser[0]), .B0_f (new_AGEMA_signal_6982), .B1_t (new_AGEMA_signal_6983), .B1_f (new_AGEMA_signal_6984), .Z0_t (KeyArray_S10reg_gff_1_SFF_0_QD), .Z0_f (new_AGEMA_signal_9472), .Z1_t (new_AGEMA_signal_9473), .Z1_f (new_AGEMA_signal_9474) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S10reg_gff_1_SFF_1_U3 ( .A0_t (KeyArray_S10reg_gff_1_SFF_1_n2), .A0_f (new_AGEMA_signal_9951), .A1_t (new_AGEMA_signal_9952), .A1_f (new_AGEMA_signal_9953), .B0_t (KeyArray_S10reg_gff_1_SFF_1_n1), .B0_f (new_AGEMA_signal_8700), .B1_t (new_AGEMA_signal_8701), .B1_f (new_AGEMA_signal_8702), .Z0_t (KeyArray_outS10ser[1]), .Z0_f (new_AGEMA_signal_4590), .Z1_t (new_AGEMA_signal_4591), .Z1_f (new_AGEMA_signal_4592) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_1_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS10ser[1]), .B0_f (new_AGEMA_signal_4590), .B1_t (new_AGEMA_signal_4591), .B1_f (new_AGEMA_signal_4592), .Z0_t (KeyArray_S10reg_gff_1_SFF_1_n1), .Z0_f (new_AGEMA_signal_8700), .Z1_t (new_AGEMA_signal_8701), .Z1_f (new_AGEMA_signal_8702) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_1_U1 ( .A0_t (KeyArray_S10reg_gff_1_SFF_1_QD), .A0_f (new_AGEMA_signal_9475), .A1_t (new_AGEMA_signal_9476), .A1_f (new_AGEMA_signal_9477), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S10reg_gff_1_SFF_1_n2), .Z0_f (new_AGEMA_signal_9951), .Z1_t (new_AGEMA_signal_9952), .Z1_f (new_AGEMA_signal_9953) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS10ser[1]), .A0_f (new_AGEMA_signal_6985), .A1_t (new_AGEMA_signal_6986), .A1_f (new_AGEMA_signal_6987), .B0_t (KeyArray_outS20ser[1]), .B0_f (new_AGEMA_signal_4878), .B1_t (new_AGEMA_signal_4879), .B1_f (new_AGEMA_signal_4880), .Z0_t (KeyArray_S10reg_gff_1_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_7818), .Z1_t (new_AGEMA_signal_7819), .Z1_f (new_AGEMA_signal_7820) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S10reg_gff_1_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_7818), .B1_t (new_AGEMA_signal_7819), .B1_f (new_AGEMA_signal_7820), .Z0_t (KeyArray_S10reg_gff_1_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_8703), .Z1_t (new_AGEMA_signal_8704), .Z1_f (new_AGEMA_signal_8705) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S10reg_gff_1_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_8703), .A1_t (new_AGEMA_signal_8704), .A1_f (new_AGEMA_signal_8705), .B0_t (KeyArray_inS10ser[1]), .B0_f (new_AGEMA_signal_6985), .B1_t (new_AGEMA_signal_6986), .B1_f (new_AGEMA_signal_6987), .Z0_t (KeyArray_S10reg_gff_1_SFF_1_QD), .Z0_f (new_AGEMA_signal_9475), .Z1_t (new_AGEMA_signal_9476), .Z1_f (new_AGEMA_signal_9477) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S10reg_gff_1_SFF_2_U3 ( .A0_t (KeyArray_S10reg_gff_1_SFF_2_n2), .A0_f (new_AGEMA_signal_9954), .A1_t (new_AGEMA_signal_9955), .A1_f (new_AGEMA_signal_9956), .B0_t (KeyArray_S10reg_gff_1_SFF_2_n1), .B0_f (new_AGEMA_signal_8706), .B1_t (new_AGEMA_signal_8707), .B1_f (new_AGEMA_signal_8708), .Z0_t (KeyArray_outS10ser[2]), .Z0_f (new_AGEMA_signal_4599), .Z1_t (new_AGEMA_signal_4600), .Z1_f (new_AGEMA_signal_4601) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_2_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS10ser[2]), .B0_f (new_AGEMA_signal_4599), .B1_t (new_AGEMA_signal_4600), .B1_f (new_AGEMA_signal_4601), .Z0_t (KeyArray_S10reg_gff_1_SFF_2_n1), .Z0_f (new_AGEMA_signal_8706), .Z1_t (new_AGEMA_signal_8707), .Z1_f (new_AGEMA_signal_8708) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_2_U1 ( .A0_t (KeyArray_S10reg_gff_1_SFF_2_QD), .A0_f (new_AGEMA_signal_9478), .A1_t (new_AGEMA_signal_9479), .A1_f (new_AGEMA_signal_9480), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S10reg_gff_1_SFF_2_n2), .Z0_f (new_AGEMA_signal_9954), .Z1_t (new_AGEMA_signal_9955), .Z1_f (new_AGEMA_signal_9956) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS10ser[2]), .A0_f (new_AGEMA_signal_6988), .A1_t (new_AGEMA_signal_6989), .A1_f (new_AGEMA_signal_6990), .B0_t (KeyArray_outS20ser[2]), .B0_f (new_AGEMA_signal_4887), .B1_t (new_AGEMA_signal_4888), .B1_f (new_AGEMA_signal_4889), .Z0_t (KeyArray_S10reg_gff_1_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_7821), .Z1_t (new_AGEMA_signal_7822), .Z1_f (new_AGEMA_signal_7823) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S10reg_gff_1_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_7821), .B1_t (new_AGEMA_signal_7822), .B1_f (new_AGEMA_signal_7823), .Z0_t (KeyArray_S10reg_gff_1_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_8709), .Z1_t (new_AGEMA_signal_8710), .Z1_f (new_AGEMA_signal_8711) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S10reg_gff_1_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_8709), .A1_t (new_AGEMA_signal_8710), .A1_f (new_AGEMA_signal_8711), .B0_t (KeyArray_inS10ser[2]), .B0_f (new_AGEMA_signal_6988), .B1_t (new_AGEMA_signal_6989), .B1_f (new_AGEMA_signal_6990), .Z0_t (KeyArray_S10reg_gff_1_SFF_2_QD), .Z0_f (new_AGEMA_signal_9478), .Z1_t (new_AGEMA_signal_9479), .Z1_f (new_AGEMA_signal_9480) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S10reg_gff_1_SFF_3_U3 ( .A0_t (KeyArray_S10reg_gff_1_SFF_3_n2), .A0_f (new_AGEMA_signal_9957), .A1_t (new_AGEMA_signal_9958), .A1_f (new_AGEMA_signal_9959), .B0_t (KeyArray_S10reg_gff_1_SFF_3_n1), .B0_f (new_AGEMA_signal_8712), .B1_t (new_AGEMA_signal_8713), .B1_f (new_AGEMA_signal_8714), .Z0_t (KeyArray_outS10ser[3]), .Z0_f (new_AGEMA_signal_4608), .Z1_t (new_AGEMA_signal_4609), .Z1_f (new_AGEMA_signal_4610) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_3_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS10ser[3]), .B0_f (new_AGEMA_signal_4608), .B1_t (new_AGEMA_signal_4609), .B1_f (new_AGEMA_signal_4610), .Z0_t (KeyArray_S10reg_gff_1_SFF_3_n1), .Z0_f (new_AGEMA_signal_8712), .Z1_t (new_AGEMA_signal_8713), .Z1_f (new_AGEMA_signal_8714) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_3_U1 ( .A0_t (KeyArray_S10reg_gff_1_SFF_3_QD), .A0_f (new_AGEMA_signal_9481), .A1_t (new_AGEMA_signal_9482), .A1_f (new_AGEMA_signal_9483), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S10reg_gff_1_SFF_3_n2), .Z0_f (new_AGEMA_signal_9957), .Z1_t (new_AGEMA_signal_9958), .Z1_f (new_AGEMA_signal_9959) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS10ser[3]), .A0_f (new_AGEMA_signal_6991), .A1_t (new_AGEMA_signal_6992), .A1_f (new_AGEMA_signal_6993), .B0_t (KeyArray_outS20ser[3]), .B0_f (new_AGEMA_signal_4896), .B1_t (new_AGEMA_signal_4897), .B1_f (new_AGEMA_signal_4898), .Z0_t (KeyArray_S10reg_gff_1_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_7824), .Z1_t (new_AGEMA_signal_7825), .Z1_f (new_AGEMA_signal_7826) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S10reg_gff_1_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_7824), .B1_t (new_AGEMA_signal_7825), .B1_f (new_AGEMA_signal_7826), .Z0_t (KeyArray_S10reg_gff_1_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_8715), .Z1_t (new_AGEMA_signal_8716), .Z1_f (new_AGEMA_signal_8717) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S10reg_gff_1_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_8715), .A1_t (new_AGEMA_signal_8716), .A1_f (new_AGEMA_signal_8717), .B0_t (KeyArray_inS10ser[3]), .B0_f (new_AGEMA_signal_6991), .B1_t (new_AGEMA_signal_6992), .B1_f (new_AGEMA_signal_6993), .Z0_t (KeyArray_S10reg_gff_1_SFF_3_QD), .Z0_f (new_AGEMA_signal_9481), .Z1_t (new_AGEMA_signal_9482), .Z1_f (new_AGEMA_signal_9483) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S10reg_gff_1_SFF_4_U3 ( .A0_t (KeyArray_S10reg_gff_1_SFF_4_n2), .A0_f (new_AGEMA_signal_9960), .A1_t (new_AGEMA_signal_9961), .A1_f (new_AGEMA_signal_9962), .B0_t (KeyArray_S10reg_gff_1_SFF_4_n1), .B0_f (new_AGEMA_signal_8718), .B1_t (new_AGEMA_signal_8719), .B1_f (new_AGEMA_signal_8720), .Z0_t (KeyArray_outS10ser[4]), .Z0_f (new_AGEMA_signal_4617), .Z1_t (new_AGEMA_signal_4618), .Z1_f (new_AGEMA_signal_4619) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_4_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS10ser[4]), .B0_f (new_AGEMA_signal_4617), .B1_t (new_AGEMA_signal_4618), .B1_f (new_AGEMA_signal_4619), .Z0_t (KeyArray_S10reg_gff_1_SFF_4_n1), .Z0_f (new_AGEMA_signal_8718), .Z1_t (new_AGEMA_signal_8719), .Z1_f (new_AGEMA_signal_8720) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_4_U1 ( .A0_t (KeyArray_S10reg_gff_1_SFF_4_QD), .A0_f (new_AGEMA_signal_9484), .A1_t (new_AGEMA_signal_9485), .A1_f (new_AGEMA_signal_9486), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S10reg_gff_1_SFF_4_n2), .Z0_f (new_AGEMA_signal_9960), .Z1_t (new_AGEMA_signal_9961), .Z1_f (new_AGEMA_signal_9962) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS10ser[4]), .A0_f (new_AGEMA_signal_6994), .A1_t (new_AGEMA_signal_6995), .A1_f (new_AGEMA_signal_6996), .B0_t (KeyArray_outS20ser[4]), .B0_f (new_AGEMA_signal_4905), .B1_t (new_AGEMA_signal_4906), .B1_f (new_AGEMA_signal_4907), .Z0_t (KeyArray_S10reg_gff_1_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_7827), .Z1_t (new_AGEMA_signal_7828), .Z1_f (new_AGEMA_signal_7829) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S10reg_gff_1_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_7827), .B1_t (new_AGEMA_signal_7828), .B1_f (new_AGEMA_signal_7829), .Z0_t (KeyArray_S10reg_gff_1_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_8721), .Z1_t (new_AGEMA_signal_8722), .Z1_f (new_AGEMA_signal_8723) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S10reg_gff_1_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_8721), .A1_t (new_AGEMA_signal_8722), .A1_f (new_AGEMA_signal_8723), .B0_t (KeyArray_inS10ser[4]), .B0_f (new_AGEMA_signal_6994), .B1_t (new_AGEMA_signal_6995), .B1_f (new_AGEMA_signal_6996), .Z0_t (KeyArray_S10reg_gff_1_SFF_4_QD), .Z0_f (new_AGEMA_signal_9484), .Z1_t (new_AGEMA_signal_9485), .Z1_f (new_AGEMA_signal_9486) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S10reg_gff_1_SFF_5_U3 ( .A0_t (KeyArray_S10reg_gff_1_SFF_5_n2), .A0_f (new_AGEMA_signal_9963), .A1_t (new_AGEMA_signal_9964), .A1_f (new_AGEMA_signal_9965), .B0_t (KeyArray_S10reg_gff_1_SFF_5_n1), .B0_f (new_AGEMA_signal_8724), .B1_t (new_AGEMA_signal_8725), .B1_f (new_AGEMA_signal_8726), .Z0_t (KeyArray_outS10ser[5]), .Z0_f (new_AGEMA_signal_4626), .Z1_t (new_AGEMA_signal_4627), .Z1_f (new_AGEMA_signal_4628) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_5_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS10ser[5]), .B0_f (new_AGEMA_signal_4626), .B1_t (new_AGEMA_signal_4627), .B1_f (new_AGEMA_signal_4628), .Z0_t (KeyArray_S10reg_gff_1_SFF_5_n1), .Z0_f (new_AGEMA_signal_8724), .Z1_t (new_AGEMA_signal_8725), .Z1_f (new_AGEMA_signal_8726) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_5_U1 ( .A0_t (KeyArray_S10reg_gff_1_SFF_5_QD), .A0_f (new_AGEMA_signal_9487), .A1_t (new_AGEMA_signal_9488), .A1_f (new_AGEMA_signal_9489), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S10reg_gff_1_SFF_5_n2), .Z0_f (new_AGEMA_signal_9963), .Z1_t (new_AGEMA_signal_9964), .Z1_f (new_AGEMA_signal_9965) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS10ser[5]), .A0_f (new_AGEMA_signal_6997), .A1_t (new_AGEMA_signal_6998), .A1_f (new_AGEMA_signal_6999), .B0_t (KeyArray_outS20ser[5]), .B0_f (new_AGEMA_signal_4914), .B1_t (new_AGEMA_signal_4915), .B1_f (new_AGEMA_signal_4916), .Z0_t (KeyArray_S10reg_gff_1_SFF_5_MUXInst_X), .Z0_f (new_AGEMA_signal_7830), .Z1_t (new_AGEMA_signal_7831), .Z1_f (new_AGEMA_signal_7832) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S10reg_gff_1_SFF_5_MUXInst_X), .B0_f (new_AGEMA_signal_7830), .B1_t (new_AGEMA_signal_7831), .B1_f (new_AGEMA_signal_7832), .Z0_t (KeyArray_S10reg_gff_1_SFF_5_MUXInst_Y), .Z0_f (new_AGEMA_signal_8727), .Z1_t (new_AGEMA_signal_8728), .Z1_f (new_AGEMA_signal_8729) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S10reg_gff_1_SFF_5_MUXInst_Y), .A0_f (new_AGEMA_signal_8727), .A1_t (new_AGEMA_signal_8728), .A1_f (new_AGEMA_signal_8729), .B0_t (KeyArray_inS10ser[5]), .B0_f (new_AGEMA_signal_6997), .B1_t (new_AGEMA_signal_6998), .B1_f (new_AGEMA_signal_6999), .Z0_t (KeyArray_S10reg_gff_1_SFF_5_QD), .Z0_f (new_AGEMA_signal_9487), .Z1_t (new_AGEMA_signal_9488), .Z1_f (new_AGEMA_signal_9489) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S10reg_gff_1_SFF_6_U3 ( .A0_t (KeyArray_S10reg_gff_1_SFF_6_n2), .A0_f (new_AGEMA_signal_9966), .A1_t (new_AGEMA_signal_9967), .A1_f (new_AGEMA_signal_9968), .B0_t (KeyArray_S10reg_gff_1_SFF_6_n1), .B0_f (new_AGEMA_signal_8730), .B1_t (new_AGEMA_signal_8731), .B1_f (new_AGEMA_signal_8732), .Z0_t (KeyArray_outS10ser[6]), .Z0_f (new_AGEMA_signal_4635), .Z1_t (new_AGEMA_signal_4636), .Z1_f (new_AGEMA_signal_4637) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_6_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS10ser[6]), .B0_f (new_AGEMA_signal_4635), .B1_t (new_AGEMA_signal_4636), .B1_f (new_AGEMA_signal_4637), .Z0_t (KeyArray_S10reg_gff_1_SFF_6_n1), .Z0_f (new_AGEMA_signal_8730), .Z1_t (new_AGEMA_signal_8731), .Z1_f (new_AGEMA_signal_8732) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_6_U1 ( .A0_t (KeyArray_S10reg_gff_1_SFF_6_QD), .A0_f (new_AGEMA_signal_9490), .A1_t (new_AGEMA_signal_9491), .A1_f (new_AGEMA_signal_9492), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S10reg_gff_1_SFF_6_n2), .Z0_f (new_AGEMA_signal_9966), .Z1_t (new_AGEMA_signal_9967), .Z1_f (new_AGEMA_signal_9968) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS10ser[6]), .A0_f (new_AGEMA_signal_7000), .A1_t (new_AGEMA_signal_7001), .A1_f (new_AGEMA_signal_7002), .B0_t (KeyArray_outS20ser[6]), .B0_f (new_AGEMA_signal_4923), .B1_t (new_AGEMA_signal_4924), .B1_f (new_AGEMA_signal_4925), .Z0_t (KeyArray_S10reg_gff_1_SFF_6_MUXInst_X), .Z0_f (new_AGEMA_signal_7833), .Z1_t (new_AGEMA_signal_7834), .Z1_f (new_AGEMA_signal_7835) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S10reg_gff_1_SFF_6_MUXInst_X), .B0_f (new_AGEMA_signal_7833), .B1_t (new_AGEMA_signal_7834), .B1_f (new_AGEMA_signal_7835), .Z0_t (KeyArray_S10reg_gff_1_SFF_6_MUXInst_Y), .Z0_f (new_AGEMA_signal_8733), .Z1_t (new_AGEMA_signal_8734), .Z1_f (new_AGEMA_signal_8735) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S10reg_gff_1_SFF_6_MUXInst_Y), .A0_f (new_AGEMA_signal_8733), .A1_t (new_AGEMA_signal_8734), .A1_f (new_AGEMA_signal_8735), .B0_t (KeyArray_inS10ser[6]), .B0_f (new_AGEMA_signal_7000), .B1_t (new_AGEMA_signal_7001), .B1_f (new_AGEMA_signal_7002), .Z0_t (KeyArray_S10reg_gff_1_SFF_6_QD), .Z0_f (new_AGEMA_signal_9490), .Z1_t (new_AGEMA_signal_9491), .Z1_f (new_AGEMA_signal_9492) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S10reg_gff_1_SFF_7_U3 ( .A0_t (KeyArray_S10reg_gff_1_SFF_7_n2), .A0_f (new_AGEMA_signal_9969), .A1_t (new_AGEMA_signal_9970), .A1_f (new_AGEMA_signal_9971), .B0_t (KeyArray_S10reg_gff_1_SFF_7_n1), .B0_f (new_AGEMA_signal_8736), .B1_t (new_AGEMA_signal_8737), .B1_f (new_AGEMA_signal_8738), .Z0_t (KeyArray_outS10ser[7]), .Z0_f (new_AGEMA_signal_4644), .Z1_t (new_AGEMA_signal_4645), .Z1_f (new_AGEMA_signal_4646) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_7_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS10ser[7]), .B0_f (new_AGEMA_signal_4644), .B1_t (new_AGEMA_signal_4645), .B1_f (new_AGEMA_signal_4646), .Z0_t (KeyArray_S10reg_gff_1_SFF_7_n1), .Z0_f (new_AGEMA_signal_8736), .Z1_t (new_AGEMA_signal_8737), .Z1_f (new_AGEMA_signal_8738) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_7_U1 ( .A0_t (KeyArray_S10reg_gff_1_SFF_7_QD), .A0_f (new_AGEMA_signal_9493), .A1_t (new_AGEMA_signal_9494), .A1_f (new_AGEMA_signal_9495), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S10reg_gff_1_SFF_7_n2), .Z0_f (new_AGEMA_signal_9969), .Z1_t (new_AGEMA_signal_9970), .Z1_f (new_AGEMA_signal_9971) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS10ser[7]), .A0_f (new_AGEMA_signal_7003), .A1_t (new_AGEMA_signal_7004), .A1_f (new_AGEMA_signal_7005), .B0_t (KeyArray_outS20ser[7]), .B0_f (new_AGEMA_signal_4932), .B1_t (new_AGEMA_signal_4933), .B1_f (new_AGEMA_signal_4934), .Z0_t (KeyArray_S10reg_gff_1_SFF_7_MUXInst_X), .Z0_f (new_AGEMA_signal_7836), .Z1_t (new_AGEMA_signal_7837), .Z1_f (new_AGEMA_signal_7838) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S10reg_gff_1_SFF_7_MUXInst_X), .B0_f (new_AGEMA_signal_7836), .B1_t (new_AGEMA_signal_7837), .B1_f (new_AGEMA_signal_7838), .Z0_t (KeyArray_S10reg_gff_1_SFF_7_MUXInst_Y), .Z0_f (new_AGEMA_signal_8739), .Z1_t (new_AGEMA_signal_8740), .Z1_f (new_AGEMA_signal_8741) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S10reg_gff_1_SFF_7_MUXInst_Y), .A0_f (new_AGEMA_signal_8739), .A1_t (new_AGEMA_signal_8740), .A1_f (new_AGEMA_signal_8741), .B0_t (KeyArray_inS10ser[7]), .B0_f (new_AGEMA_signal_7003), .B1_t (new_AGEMA_signal_7004), .B1_f (new_AGEMA_signal_7005), .Z0_t (KeyArray_S10reg_gff_1_SFF_7_QD), .Z0_f (new_AGEMA_signal_9493), .Z1_t (new_AGEMA_signal_9494), .Z1_f (new_AGEMA_signal_9495) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S11reg_gff_1_SFF_0_U3 ( .A0_t (KeyArray_S11reg_gff_1_SFF_0_n2), .A0_f (new_AGEMA_signal_9972), .A1_t (new_AGEMA_signal_9973), .A1_f (new_AGEMA_signal_9974), .B0_t (KeyArray_S11reg_gff_1_SFF_0_n1), .B0_f (new_AGEMA_signal_8742), .B1_t (new_AGEMA_signal_8743), .B1_f (new_AGEMA_signal_8744), .Z0_t (KeyArray_outS11ser[0]), .Z0_f (new_AGEMA_signal_4653), .Z1_t (new_AGEMA_signal_4654), .Z1_f (new_AGEMA_signal_4655) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_0_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS11ser[0]), .B0_f (new_AGEMA_signal_4653), .B1_t (new_AGEMA_signal_4654), .B1_f (new_AGEMA_signal_4655), .Z0_t (KeyArray_S11reg_gff_1_SFF_0_n1), .Z0_f (new_AGEMA_signal_8742), .Z1_t (new_AGEMA_signal_8743), .Z1_f (new_AGEMA_signal_8744) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_0_U1 ( .A0_t (KeyArray_S11reg_gff_1_SFF_0_QD), .A0_f (new_AGEMA_signal_9496), .A1_t (new_AGEMA_signal_9497), .A1_f (new_AGEMA_signal_9498), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S11reg_gff_1_SFF_0_n2), .Z0_f (new_AGEMA_signal_9972), .Z1_t (new_AGEMA_signal_9973), .Z1_f (new_AGEMA_signal_9974) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS11ser[0]), .A0_f (new_AGEMA_signal_7006), .A1_t (new_AGEMA_signal_7007), .A1_f (new_AGEMA_signal_7008), .B0_t (KeyArray_outS21ser[0]), .B0_f (new_AGEMA_signal_4941), .B1_t (new_AGEMA_signal_4942), .B1_f (new_AGEMA_signal_4943), .Z0_t (KeyArray_S11reg_gff_1_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_7839), .Z1_t (new_AGEMA_signal_7840), .Z1_f (new_AGEMA_signal_7841) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S11reg_gff_1_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_7839), .B1_t (new_AGEMA_signal_7840), .B1_f (new_AGEMA_signal_7841), .Z0_t (KeyArray_S11reg_gff_1_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_8745), .Z1_t (new_AGEMA_signal_8746), .Z1_f (new_AGEMA_signal_8747) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S11reg_gff_1_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_8745), .A1_t (new_AGEMA_signal_8746), .A1_f (new_AGEMA_signal_8747), .B0_t (KeyArray_inS11ser[0]), .B0_f (new_AGEMA_signal_7006), .B1_t (new_AGEMA_signal_7007), .B1_f (new_AGEMA_signal_7008), .Z0_t (KeyArray_S11reg_gff_1_SFF_0_QD), .Z0_f (new_AGEMA_signal_9496), .Z1_t (new_AGEMA_signal_9497), .Z1_f (new_AGEMA_signal_9498) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S11reg_gff_1_SFF_1_U3 ( .A0_t (KeyArray_S11reg_gff_1_SFF_1_n2), .A0_f (new_AGEMA_signal_9975), .A1_t (new_AGEMA_signal_9976), .A1_f (new_AGEMA_signal_9977), .B0_t (KeyArray_S11reg_gff_1_SFF_1_n1), .B0_f (new_AGEMA_signal_8748), .B1_t (new_AGEMA_signal_8749), .B1_f (new_AGEMA_signal_8750), .Z0_t (KeyArray_outS11ser[1]), .Z0_f (new_AGEMA_signal_4662), .Z1_t (new_AGEMA_signal_4663), .Z1_f (new_AGEMA_signal_4664) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_1_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS11ser[1]), .B0_f (new_AGEMA_signal_4662), .B1_t (new_AGEMA_signal_4663), .B1_f (new_AGEMA_signal_4664), .Z0_t (KeyArray_S11reg_gff_1_SFF_1_n1), .Z0_f (new_AGEMA_signal_8748), .Z1_t (new_AGEMA_signal_8749), .Z1_f (new_AGEMA_signal_8750) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_1_U1 ( .A0_t (KeyArray_S11reg_gff_1_SFF_1_QD), .A0_f (new_AGEMA_signal_9499), .A1_t (new_AGEMA_signal_9500), .A1_f (new_AGEMA_signal_9501), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S11reg_gff_1_SFF_1_n2), .Z0_f (new_AGEMA_signal_9975), .Z1_t (new_AGEMA_signal_9976), .Z1_f (new_AGEMA_signal_9977) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS11ser[1]), .A0_f (new_AGEMA_signal_7009), .A1_t (new_AGEMA_signal_7010), .A1_f (new_AGEMA_signal_7011), .B0_t (KeyArray_outS21ser[1]), .B0_f (new_AGEMA_signal_4950), .B1_t (new_AGEMA_signal_4951), .B1_f (new_AGEMA_signal_4952), .Z0_t (KeyArray_S11reg_gff_1_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_7842), .Z1_t (new_AGEMA_signal_7843), .Z1_f (new_AGEMA_signal_7844) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S11reg_gff_1_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_7842), .B1_t (new_AGEMA_signal_7843), .B1_f (new_AGEMA_signal_7844), .Z0_t (KeyArray_S11reg_gff_1_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_8751), .Z1_t (new_AGEMA_signal_8752), .Z1_f (new_AGEMA_signal_8753) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S11reg_gff_1_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_8751), .A1_t (new_AGEMA_signal_8752), .A1_f (new_AGEMA_signal_8753), .B0_t (KeyArray_inS11ser[1]), .B0_f (new_AGEMA_signal_7009), .B1_t (new_AGEMA_signal_7010), .B1_f (new_AGEMA_signal_7011), .Z0_t (KeyArray_S11reg_gff_1_SFF_1_QD), .Z0_f (new_AGEMA_signal_9499), .Z1_t (new_AGEMA_signal_9500), .Z1_f (new_AGEMA_signal_9501) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S11reg_gff_1_SFF_2_U3 ( .A0_t (KeyArray_S11reg_gff_1_SFF_2_n2), .A0_f (new_AGEMA_signal_9978), .A1_t (new_AGEMA_signal_9979), .A1_f (new_AGEMA_signal_9980), .B0_t (KeyArray_S11reg_gff_1_SFF_2_n1), .B0_f (new_AGEMA_signal_8754), .B1_t (new_AGEMA_signal_8755), .B1_f (new_AGEMA_signal_8756), .Z0_t (KeyArray_outS11ser[2]), .Z0_f (new_AGEMA_signal_4671), .Z1_t (new_AGEMA_signal_4672), .Z1_f (new_AGEMA_signal_4673) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_2_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS11ser[2]), .B0_f (new_AGEMA_signal_4671), .B1_t (new_AGEMA_signal_4672), .B1_f (new_AGEMA_signal_4673), .Z0_t (KeyArray_S11reg_gff_1_SFF_2_n1), .Z0_f (new_AGEMA_signal_8754), .Z1_t (new_AGEMA_signal_8755), .Z1_f (new_AGEMA_signal_8756) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_2_U1 ( .A0_t (KeyArray_S11reg_gff_1_SFF_2_QD), .A0_f (new_AGEMA_signal_9502), .A1_t (new_AGEMA_signal_9503), .A1_f (new_AGEMA_signal_9504), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S11reg_gff_1_SFF_2_n2), .Z0_f (new_AGEMA_signal_9978), .Z1_t (new_AGEMA_signal_9979), .Z1_f (new_AGEMA_signal_9980) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS11ser[2]), .A0_f (new_AGEMA_signal_7012), .A1_t (new_AGEMA_signal_7013), .A1_f (new_AGEMA_signal_7014), .B0_t (KeyArray_outS21ser[2]), .B0_f (new_AGEMA_signal_4959), .B1_t (new_AGEMA_signal_4960), .B1_f (new_AGEMA_signal_4961), .Z0_t (KeyArray_S11reg_gff_1_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_7845), .Z1_t (new_AGEMA_signal_7846), .Z1_f (new_AGEMA_signal_7847) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S11reg_gff_1_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_7845), .B1_t (new_AGEMA_signal_7846), .B1_f (new_AGEMA_signal_7847), .Z0_t (KeyArray_S11reg_gff_1_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_8757), .Z1_t (new_AGEMA_signal_8758), .Z1_f (new_AGEMA_signal_8759) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S11reg_gff_1_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_8757), .A1_t (new_AGEMA_signal_8758), .A1_f (new_AGEMA_signal_8759), .B0_t (KeyArray_inS11ser[2]), .B0_f (new_AGEMA_signal_7012), .B1_t (new_AGEMA_signal_7013), .B1_f (new_AGEMA_signal_7014), .Z0_t (KeyArray_S11reg_gff_1_SFF_2_QD), .Z0_f (new_AGEMA_signal_9502), .Z1_t (new_AGEMA_signal_9503), .Z1_f (new_AGEMA_signal_9504) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S11reg_gff_1_SFF_3_U3 ( .A0_t (KeyArray_S11reg_gff_1_SFF_3_n2), .A0_f (new_AGEMA_signal_9981), .A1_t (new_AGEMA_signal_9982), .A1_f (new_AGEMA_signal_9983), .B0_t (KeyArray_S11reg_gff_1_SFF_3_n1), .B0_f (new_AGEMA_signal_8760), .B1_t (new_AGEMA_signal_8761), .B1_f (new_AGEMA_signal_8762), .Z0_t (KeyArray_outS11ser[3]), .Z0_f (new_AGEMA_signal_4680), .Z1_t (new_AGEMA_signal_4681), .Z1_f (new_AGEMA_signal_4682) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_3_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS11ser[3]), .B0_f (new_AGEMA_signal_4680), .B1_t (new_AGEMA_signal_4681), .B1_f (new_AGEMA_signal_4682), .Z0_t (KeyArray_S11reg_gff_1_SFF_3_n1), .Z0_f (new_AGEMA_signal_8760), .Z1_t (new_AGEMA_signal_8761), .Z1_f (new_AGEMA_signal_8762) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_3_U1 ( .A0_t (KeyArray_S11reg_gff_1_SFF_3_QD), .A0_f (new_AGEMA_signal_9505), .A1_t (new_AGEMA_signal_9506), .A1_f (new_AGEMA_signal_9507), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S11reg_gff_1_SFF_3_n2), .Z0_f (new_AGEMA_signal_9981), .Z1_t (new_AGEMA_signal_9982), .Z1_f (new_AGEMA_signal_9983) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS11ser[3]), .A0_f (new_AGEMA_signal_7015), .A1_t (new_AGEMA_signal_7016), .A1_f (new_AGEMA_signal_7017), .B0_t (KeyArray_outS21ser[3]), .B0_f (new_AGEMA_signal_4968), .B1_t (new_AGEMA_signal_4969), .B1_f (new_AGEMA_signal_4970), .Z0_t (KeyArray_S11reg_gff_1_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_7848), .Z1_t (new_AGEMA_signal_7849), .Z1_f (new_AGEMA_signal_7850) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S11reg_gff_1_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_7848), .B1_t (new_AGEMA_signal_7849), .B1_f (new_AGEMA_signal_7850), .Z0_t (KeyArray_S11reg_gff_1_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_8763), .Z1_t (new_AGEMA_signal_8764), .Z1_f (new_AGEMA_signal_8765) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S11reg_gff_1_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_8763), .A1_t (new_AGEMA_signal_8764), .A1_f (new_AGEMA_signal_8765), .B0_t (KeyArray_inS11ser[3]), .B0_f (new_AGEMA_signal_7015), .B1_t (new_AGEMA_signal_7016), .B1_f (new_AGEMA_signal_7017), .Z0_t (KeyArray_S11reg_gff_1_SFF_3_QD), .Z0_f (new_AGEMA_signal_9505), .Z1_t (new_AGEMA_signal_9506), .Z1_f (new_AGEMA_signal_9507) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S11reg_gff_1_SFF_4_U3 ( .A0_t (KeyArray_S11reg_gff_1_SFF_4_n2), .A0_f (new_AGEMA_signal_9984), .A1_t (new_AGEMA_signal_9985), .A1_f (new_AGEMA_signal_9986), .B0_t (KeyArray_S11reg_gff_1_SFF_4_n1), .B0_f (new_AGEMA_signal_8766), .B1_t (new_AGEMA_signal_8767), .B1_f (new_AGEMA_signal_8768), .Z0_t (KeyArray_outS11ser[4]), .Z0_f (new_AGEMA_signal_4689), .Z1_t (new_AGEMA_signal_4690), .Z1_f (new_AGEMA_signal_4691) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_4_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS11ser[4]), .B0_f (new_AGEMA_signal_4689), .B1_t (new_AGEMA_signal_4690), .B1_f (new_AGEMA_signal_4691), .Z0_t (KeyArray_S11reg_gff_1_SFF_4_n1), .Z0_f (new_AGEMA_signal_8766), .Z1_t (new_AGEMA_signal_8767), .Z1_f (new_AGEMA_signal_8768) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_4_U1 ( .A0_t (KeyArray_S11reg_gff_1_SFF_4_QD), .A0_f (new_AGEMA_signal_9508), .A1_t (new_AGEMA_signal_9509), .A1_f (new_AGEMA_signal_9510), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S11reg_gff_1_SFF_4_n2), .Z0_f (new_AGEMA_signal_9984), .Z1_t (new_AGEMA_signal_9985), .Z1_f (new_AGEMA_signal_9986) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS11ser[4]), .A0_f (new_AGEMA_signal_7018), .A1_t (new_AGEMA_signal_7019), .A1_f (new_AGEMA_signal_7020), .B0_t (KeyArray_outS21ser[4]), .B0_f (new_AGEMA_signal_4977), .B1_t (new_AGEMA_signal_4978), .B1_f (new_AGEMA_signal_4979), .Z0_t (KeyArray_S11reg_gff_1_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_7851), .Z1_t (new_AGEMA_signal_7852), .Z1_f (new_AGEMA_signal_7853) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S11reg_gff_1_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_7851), .B1_t (new_AGEMA_signal_7852), .B1_f (new_AGEMA_signal_7853), .Z0_t (KeyArray_S11reg_gff_1_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_8769), .Z1_t (new_AGEMA_signal_8770), .Z1_f (new_AGEMA_signal_8771) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S11reg_gff_1_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_8769), .A1_t (new_AGEMA_signal_8770), .A1_f (new_AGEMA_signal_8771), .B0_t (KeyArray_inS11ser[4]), .B0_f (new_AGEMA_signal_7018), .B1_t (new_AGEMA_signal_7019), .B1_f (new_AGEMA_signal_7020), .Z0_t (KeyArray_S11reg_gff_1_SFF_4_QD), .Z0_f (new_AGEMA_signal_9508), .Z1_t (new_AGEMA_signal_9509), .Z1_f (new_AGEMA_signal_9510) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S11reg_gff_1_SFF_5_U3 ( .A0_t (KeyArray_S11reg_gff_1_SFF_5_n2), .A0_f (new_AGEMA_signal_9987), .A1_t (new_AGEMA_signal_9988), .A1_f (new_AGEMA_signal_9989), .B0_t (KeyArray_S11reg_gff_1_SFF_5_n1), .B0_f (new_AGEMA_signal_8772), .B1_t (new_AGEMA_signal_8773), .B1_f (new_AGEMA_signal_8774), .Z0_t (KeyArray_outS11ser[5]), .Z0_f (new_AGEMA_signal_4698), .Z1_t (new_AGEMA_signal_4699), .Z1_f (new_AGEMA_signal_4700) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_5_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS11ser[5]), .B0_f (new_AGEMA_signal_4698), .B1_t (new_AGEMA_signal_4699), .B1_f (new_AGEMA_signal_4700), .Z0_t (KeyArray_S11reg_gff_1_SFF_5_n1), .Z0_f (new_AGEMA_signal_8772), .Z1_t (new_AGEMA_signal_8773), .Z1_f (new_AGEMA_signal_8774) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_5_U1 ( .A0_t (KeyArray_S11reg_gff_1_SFF_5_QD), .A0_f (new_AGEMA_signal_9511), .A1_t (new_AGEMA_signal_9512), .A1_f (new_AGEMA_signal_9513), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S11reg_gff_1_SFF_5_n2), .Z0_f (new_AGEMA_signal_9987), .Z1_t (new_AGEMA_signal_9988), .Z1_f (new_AGEMA_signal_9989) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS11ser[5]), .A0_f (new_AGEMA_signal_7021), .A1_t (new_AGEMA_signal_7022), .A1_f (new_AGEMA_signal_7023), .B0_t (KeyArray_outS21ser[5]), .B0_f (new_AGEMA_signal_4986), .B1_t (new_AGEMA_signal_4987), .B1_f (new_AGEMA_signal_4988), .Z0_t (KeyArray_S11reg_gff_1_SFF_5_MUXInst_X), .Z0_f (new_AGEMA_signal_7854), .Z1_t (new_AGEMA_signal_7855), .Z1_f (new_AGEMA_signal_7856) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S11reg_gff_1_SFF_5_MUXInst_X), .B0_f (new_AGEMA_signal_7854), .B1_t (new_AGEMA_signal_7855), .B1_f (new_AGEMA_signal_7856), .Z0_t (KeyArray_S11reg_gff_1_SFF_5_MUXInst_Y), .Z0_f (new_AGEMA_signal_8775), .Z1_t (new_AGEMA_signal_8776), .Z1_f (new_AGEMA_signal_8777) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S11reg_gff_1_SFF_5_MUXInst_Y), .A0_f (new_AGEMA_signal_8775), .A1_t (new_AGEMA_signal_8776), .A1_f (new_AGEMA_signal_8777), .B0_t (KeyArray_inS11ser[5]), .B0_f (new_AGEMA_signal_7021), .B1_t (new_AGEMA_signal_7022), .B1_f (new_AGEMA_signal_7023), .Z0_t (KeyArray_S11reg_gff_1_SFF_5_QD), .Z0_f (new_AGEMA_signal_9511), .Z1_t (new_AGEMA_signal_9512), .Z1_f (new_AGEMA_signal_9513) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S11reg_gff_1_SFF_6_U3 ( .A0_t (KeyArray_S11reg_gff_1_SFF_6_n2), .A0_f (new_AGEMA_signal_9990), .A1_t (new_AGEMA_signal_9991), .A1_f (new_AGEMA_signal_9992), .B0_t (KeyArray_S11reg_gff_1_SFF_6_n1), .B0_f (new_AGEMA_signal_8778), .B1_t (new_AGEMA_signal_8779), .B1_f (new_AGEMA_signal_8780), .Z0_t (KeyArray_outS11ser[6]), .Z0_f (new_AGEMA_signal_4707), .Z1_t (new_AGEMA_signal_4708), .Z1_f (new_AGEMA_signal_4709) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_6_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS11ser[6]), .B0_f (new_AGEMA_signal_4707), .B1_t (new_AGEMA_signal_4708), .B1_f (new_AGEMA_signal_4709), .Z0_t (KeyArray_S11reg_gff_1_SFF_6_n1), .Z0_f (new_AGEMA_signal_8778), .Z1_t (new_AGEMA_signal_8779), .Z1_f (new_AGEMA_signal_8780) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_6_U1 ( .A0_t (KeyArray_S11reg_gff_1_SFF_6_QD), .A0_f (new_AGEMA_signal_9514), .A1_t (new_AGEMA_signal_9515), .A1_f (new_AGEMA_signal_9516), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S11reg_gff_1_SFF_6_n2), .Z0_f (new_AGEMA_signal_9990), .Z1_t (new_AGEMA_signal_9991), .Z1_f (new_AGEMA_signal_9992) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS11ser[6]), .A0_f (new_AGEMA_signal_7024), .A1_t (new_AGEMA_signal_7025), .A1_f (new_AGEMA_signal_7026), .B0_t (KeyArray_outS21ser[6]), .B0_f (new_AGEMA_signal_4995), .B1_t (new_AGEMA_signal_4996), .B1_f (new_AGEMA_signal_4997), .Z0_t (KeyArray_S11reg_gff_1_SFF_6_MUXInst_X), .Z0_f (new_AGEMA_signal_7857), .Z1_t (new_AGEMA_signal_7858), .Z1_f (new_AGEMA_signal_7859) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S11reg_gff_1_SFF_6_MUXInst_X), .B0_f (new_AGEMA_signal_7857), .B1_t (new_AGEMA_signal_7858), .B1_f (new_AGEMA_signal_7859), .Z0_t (KeyArray_S11reg_gff_1_SFF_6_MUXInst_Y), .Z0_f (new_AGEMA_signal_8781), .Z1_t (new_AGEMA_signal_8782), .Z1_f (new_AGEMA_signal_8783) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S11reg_gff_1_SFF_6_MUXInst_Y), .A0_f (new_AGEMA_signal_8781), .A1_t (new_AGEMA_signal_8782), .A1_f (new_AGEMA_signal_8783), .B0_t (KeyArray_inS11ser[6]), .B0_f (new_AGEMA_signal_7024), .B1_t (new_AGEMA_signal_7025), .B1_f (new_AGEMA_signal_7026), .Z0_t (KeyArray_S11reg_gff_1_SFF_6_QD), .Z0_f (new_AGEMA_signal_9514), .Z1_t (new_AGEMA_signal_9515), .Z1_f (new_AGEMA_signal_9516) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S11reg_gff_1_SFF_7_U3 ( .A0_t (KeyArray_S11reg_gff_1_SFF_7_n2), .A0_f (new_AGEMA_signal_9993), .A1_t (new_AGEMA_signal_9994), .A1_f (new_AGEMA_signal_9995), .B0_t (KeyArray_S11reg_gff_1_SFF_7_n1), .B0_f (new_AGEMA_signal_8784), .B1_t (new_AGEMA_signal_8785), .B1_f (new_AGEMA_signal_8786), .Z0_t (KeyArray_outS11ser[7]), .Z0_f (new_AGEMA_signal_4716), .Z1_t (new_AGEMA_signal_4717), .Z1_f (new_AGEMA_signal_4718) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_7_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS11ser[7]), .B0_f (new_AGEMA_signal_4716), .B1_t (new_AGEMA_signal_4717), .B1_f (new_AGEMA_signal_4718), .Z0_t (KeyArray_S11reg_gff_1_SFF_7_n1), .Z0_f (new_AGEMA_signal_8784), .Z1_t (new_AGEMA_signal_8785), .Z1_f (new_AGEMA_signal_8786) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_7_U1 ( .A0_t (KeyArray_S11reg_gff_1_SFF_7_QD), .A0_f (new_AGEMA_signal_9517), .A1_t (new_AGEMA_signal_9518), .A1_f (new_AGEMA_signal_9519), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S11reg_gff_1_SFF_7_n2), .Z0_f (new_AGEMA_signal_9993), .Z1_t (new_AGEMA_signal_9994), .Z1_f (new_AGEMA_signal_9995) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS11ser[7]), .A0_f (new_AGEMA_signal_7027), .A1_t (new_AGEMA_signal_7028), .A1_f (new_AGEMA_signal_7029), .B0_t (KeyArray_outS21ser[7]), .B0_f (new_AGEMA_signal_5004), .B1_t (new_AGEMA_signal_5005), .B1_f (new_AGEMA_signal_5006), .Z0_t (KeyArray_S11reg_gff_1_SFF_7_MUXInst_X), .Z0_f (new_AGEMA_signal_7860), .Z1_t (new_AGEMA_signal_7861), .Z1_f (new_AGEMA_signal_7862) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S11reg_gff_1_SFF_7_MUXInst_X), .B0_f (new_AGEMA_signal_7860), .B1_t (new_AGEMA_signal_7861), .B1_f (new_AGEMA_signal_7862), .Z0_t (KeyArray_S11reg_gff_1_SFF_7_MUXInst_Y), .Z0_f (new_AGEMA_signal_8787), .Z1_t (new_AGEMA_signal_8788), .Z1_f (new_AGEMA_signal_8789) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S11reg_gff_1_SFF_7_MUXInst_Y), .A0_f (new_AGEMA_signal_8787), .A1_t (new_AGEMA_signal_8788), .A1_f (new_AGEMA_signal_8789), .B0_t (KeyArray_inS11ser[7]), .B0_f (new_AGEMA_signal_7027), .B1_t (new_AGEMA_signal_7028), .B1_f (new_AGEMA_signal_7029), .Z0_t (KeyArray_S11reg_gff_1_SFF_7_QD), .Z0_f (new_AGEMA_signal_9517), .Z1_t (new_AGEMA_signal_9518), .Z1_f (new_AGEMA_signal_9519) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S12reg_gff_1_SFF_0_U3 ( .A0_t (KeyArray_S12reg_gff_1_SFF_0_n2), .A0_f (new_AGEMA_signal_9996), .A1_t (new_AGEMA_signal_9997), .A1_f (new_AGEMA_signal_9998), .B0_t (KeyArray_S12reg_gff_1_SFF_0_n1), .B0_f (new_AGEMA_signal_8790), .B1_t (new_AGEMA_signal_8791), .B1_f (new_AGEMA_signal_8792), .Z0_t (KeyArray_outS12ser[0]), .Z0_f (new_AGEMA_signal_4725), .Z1_t (new_AGEMA_signal_4726), .Z1_f (new_AGEMA_signal_4727) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_0_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS12ser[0]), .B0_f (new_AGEMA_signal_4725), .B1_t (new_AGEMA_signal_4726), .B1_f (new_AGEMA_signal_4727), .Z0_t (KeyArray_S12reg_gff_1_SFF_0_n1), .Z0_f (new_AGEMA_signal_8790), .Z1_t (new_AGEMA_signal_8791), .Z1_f (new_AGEMA_signal_8792) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_0_U1 ( .A0_t (KeyArray_S12reg_gff_1_SFF_0_QD), .A0_f (new_AGEMA_signal_9520), .A1_t (new_AGEMA_signal_9521), .A1_f (new_AGEMA_signal_9522), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S12reg_gff_1_SFF_0_n2), .Z0_f (new_AGEMA_signal_9996), .Z1_t (new_AGEMA_signal_9997), .Z1_f (new_AGEMA_signal_9998) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS12ser[0]), .A0_f (new_AGEMA_signal_7030), .A1_t (new_AGEMA_signal_7031), .A1_f (new_AGEMA_signal_7032), .B0_t (KeyArray_outS22ser[0]), .B0_f (new_AGEMA_signal_5013), .B1_t (new_AGEMA_signal_5014), .B1_f (new_AGEMA_signal_5015), .Z0_t (KeyArray_S12reg_gff_1_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_7863), .Z1_t (new_AGEMA_signal_7864), .Z1_f (new_AGEMA_signal_7865) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S12reg_gff_1_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_7863), .B1_t (new_AGEMA_signal_7864), .B1_f (new_AGEMA_signal_7865), .Z0_t (KeyArray_S12reg_gff_1_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_8793), .Z1_t (new_AGEMA_signal_8794), .Z1_f (new_AGEMA_signal_8795) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S12reg_gff_1_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_8793), .A1_t (new_AGEMA_signal_8794), .A1_f (new_AGEMA_signal_8795), .B0_t (KeyArray_inS12ser[0]), .B0_f (new_AGEMA_signal_7030), .B1_t (new_AGEMA_signal_7031), .B1_f (new_AGEMA_signal_7032), .Z0_t (KeyArray_S12reg_gff_1_SFF_0_QD), .Z0_f (new_AGEMA_signal_9520), .Z1_t (new_AGEMA_signal_9521), .Z1_f (new_AGEMA_signal_9522) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S12reg_gff_1_SFF_1_U3 ( .A0_t (KeyArray_S12reg_gff_1_SFF_1_n2), .A0_f (new_AGEMA_signal_9999), .A1_t (new_AGEMA_signal_10000), .A1_f (new_AGEMA_signal_10001), .B0_t (KeyArray_S12reg_gff_1_SFF_1_n1), .B0_f (new_AGEMA_signal_8796), .B1_t (new_AGEMA_signal_8797), .B1_f (new_AGEMA_signal_8798), .Z0_t (KeyArray_outS12ser[1]), .Z0_f (new_AGEMA_signal_4734), .Z1_t (new_AGEMA_signal_4735), .Z1_f (new_AGEMA_signal_4736) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_1_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS12ser[1]), .B0_f (new_AGEMA_signal_4734), .B1_t (new_AGEMA_signal_4735), .B1_f (new_AGEMA_signal_4736), .Z0_t (KeyArray_S12reg_gff_1_SFF_1_n1), .Z0_f (new_AGEMA_signal_8796), .Z1_t (new_AGEMA_signal_8797), .Z1_f (new_AGEMA_signal_8798) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_1_U1 ( .A0_t (KeyArray_S12reg_gff_1_SFF_1_QD), .A0_f (new_AGEMA_signal_9523), .A1_t (new_AGEMA_signal_9524), .A1_f (new_AGEMA_signal_9525), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S12reg_gff_1_SFF_1_n2), .Z0_f (new_AGEMA_signal_9999), .Z1_t (new_AGEMA_signal_10000), .Z1_f (new_AGEMA_signal_10001) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS12ser[1]), .A0_f (new_AGEMA_signal_7033), .A1_t (new_AGEMA_signal_7034), .A1_f (new_AGEMA_signal_7035), .B0_t (KeyArray_outS22ser[1]), .B0_f (new_AGEMA_signal_5022), .B1_t (new_AGEMA_signal_5023), .B1_f (new_AGEMA_signal_5024), .Z0_t (KeyArray_S12reg_gff_1_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_7866), .Z1_t (new_AGEMA_signal_7867), .Z1_f (new_AGEMA_signal_7868) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S12reg_gff_1_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_7866), .B1_t (new_AGEMA_signal_7867), .B1_f (new_AGEMA_signal_7868), .Z0_t (KeyArray_S12reg_gff_1_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_8799), .Z1_t (new_AGEMA_signal_8800), .Z1_f (new_AGEMA_signal_8801) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S12reg_gff_1_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_8799), .A1_t (new_AGEMA_signal_8800), .A1_f (new_AGEMA_signal_8801), .B0_t (KeyArray_inS12ser[1]), .B0_f (new_AGEMA_signal_7033), .B1_t (new_AGEMA_signal_7034), .B1_f (new_AGEMA_signal_7035), .Z0_t (KeyArray_S12reg_gff_1_SFF_1_QD), .Z0_f (new_AGEMA_signal_9523), .Z1_t (new_AGEMA_signal_9524), .Z1_f (new_AGEMA_signal_9525) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S12reg_gff_1_SFF_2_U3 ( .A0_t (KeyArray_S12reg_gff_1_SFF_2_n2), .A0_f (new_AGEMA_signal_10002), .A1_t (new_AGEMA_signal_10003), .A1_f (new_AGEMA_signal_10004), .B0_t (KeyArray_S12reg_gff_1_SFF_2_n1), .B0_f (new_AGEMA_signal_8802), .B1_t (new_AGEMA_signal_8803), .B1_f (new_AGEMA_signal_8804), .Z0_t (KeyArray_outS12ser[2]), .Z0_f (new_AGEMA_signal_4743), .Z1_t (new_AGEMA_signal_4744), .Z1_f (new_AGEMA_signal_4745) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_2_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS12ser[2]), .B0_f (new_AGEMA_signal_4743), .B1_t (new_AGEMA_signal_4744), .B1_f (new_AGEMA_signal_4745), .Z0_t (KeyArray_S12reg_gff_1_SFF_2_n1), .Z0_f (new_AGEMA_signal_8802), .Z1_t (new_AGEMA_signal_8803), .Z1_f (new_AGEMA_signal_8804) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_2_U1 ( .A0_t (KeyArray_S12reg_gff_1_SFF_2_QD), .A0_f (new_AGEMA_signal_9526), .A1_t (new_AGEMA_signal_9527), .A1_f (new_AGEMA_signal_9528), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S12reg_gff_1_SFF_2_n2), .Z0_f (new_AGEMA_signal_10002), .Z1_t (new_AGEMA_signal_10003), .Z1_f (new_AGEMA_signal_10004) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS12ser[2]), .A0_f (new_AGEMA_signal_7036), .A1_t (new_AGEMA_signal_7037), .A1_f (new_AGEMA_signal_7038), .B0_t (KeyArray_outS22ser[2]), .B0_f (new_AGEMA_signal_5031), .B1_t (new_AGEMA_signal_5032), .B1_f (new_AGEMA_signal_5033), .Z0_t (KeyArray_S12reg_gff_1_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_7869), .Z1_t (new_AGEMA_signal_7870), .Z1_f (new_AGEMA_signal_7871) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S12reg_gff_1_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_7869), .B1_t (new_AGEMA_signal_7870), .B1_f (new_AGEMA_signal_7871), .Z0_t (KeyArray_S12reg_gff_1_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_8805), .Z1_t (new_AGEMA_signal_8806), .Z1_f (new_AGEMA_signal_8807) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S12reg_gff_1_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_8805), .A1_t (new_AGEMA_signal_8806), .A1_f (new_AGEMA_signal_8807), .B0_t (KeyArray_inS12ser[2]), .B0_f (new_AGEMA_signal_7036), .B1_t (new_AGEMA_signal_7037), .B1_f (new_AGEMA_signal_7038), .Z0_t (KeyArray_S12reg_gff_1_SFF_2_QD), .Z0_f (new_AGEMA_signal_9526), .Z1_t (new_AGEMA_signal_9527), .Z1_f (new_AGEMA_signal_9528) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S12reg_gff_1_SFF_3_U3 ( .A0_t (KeyArray_S12reg_gff_1_SFF_3_n2), .A0_f (new_AGEMA_signal_10005), .A1_t (new_AGEMA_signal_10006), .A1_f (new_AGEMA_signal_10007), .B0_t (KeyArray_S12reg_gff_1_SFF_3_n1), .B0_f (new_AGEMA_signal_8808), .B1_t (new_AGEMA_signal_8809), .B1_f (new_AGEMA_signal_8810), .Z0_t (KeyArray_outS12ser[3]), .Z0_f (new_AGEMA_signal_4752), .Z1_t (new_AGEMA_signal_4753), .Z1_f (new_AGEMA_signal_4754) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_3_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS12ser[3]), .B0_f (new_AGEMA_signal_4752), .B1_t (new_AGEMA_signal_4753), .B1_f (new_AGEMA_signal_4754), .Z0_t (KeyArray_S12reg_gff_1_SFF_3_n1), .Z0_f (new_AGEMA_signal_8808), .Z1_t (new_AGEMA_signal_8809), .Z1_f (new_AGEMA_signal_8810) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_3_U1 ( .A0_t (KeyArray_S12reg_gff_1_SFF_3_QD), .A0_f (new_AGEMA_signal_9529), .A1_t (new_AGEMA_signal_9530), .A1_f (new_AGEMA_signal_9531), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S12reg_gff_1_SFF_3_n2), .Z0_f (new_AGEMA_signal_10005), .Z1_t (new_AGEMA_signal_10006), .Z1_f (new_AGEMA_signal_10007) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS12ser[3]), .A0_f (new_AGEMA_signal_7039), .A1_t (new_AGEMA_signal_7040), .A1_f (new_AGEMA_signal_7041), .B0_t (KeyArray_outS22ser[3]), .B0_f (new_AGEMA_signal_5040), .B1_t (new_AGEMA_signal_5041), .B1_f (new_AGEMA_signal_5042), .Z0_t (KeyArray_S12reg_gff_1_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_7872), .Z1_t (new_AGEMA_signal_7873), .Z1_f (new_AGEMA_signal_7874) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S12reg_gff_1_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_7872), .B1_t (new_AGEMA_signal_7873), .B1_f (new_AGEMA_signal_7874), .Z0_t (KeyArray_S12reg_gff_1_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_8811), .Z1_t (new_AGEMA_signal_8812), .Z1_f (new_AGEMA_signal_8813) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S12reg_gff_1_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_8811), .A1_t (new_AGEMA_signal_8812), .A1_f (new_AGEMA_signal_8813), .B0_t (KeyArray_inS12ser[3]), .B0_f (new_AGEMA_signal_7039), .B1_t (new_AGEMA_signal_7040), .B1_f (new_AGEMA_signal_7041), .Z0_t (KeyArray_S12reg_gff_1_SFF_3_QD), .Z0_f (new_AGEMA_signal_9529), .Z1_t (new_AGEMA_signal_9530), .Z1_f (new_AGEMA_signal_9531) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S12reg_gff_1_SFF_4_U3 ( .A0_t (KeyArray_S12reg_gff_1_SFF_4_n2), .A0_f (new_AGEMA_signal_10008), .A1_t (new_AGEMA_signal_10009), .A1_f (new_AGEMA_signal_10010), .B0_t (KeyArray_S12reg_gff_1_SFF_4_n1), .B0_f (new_AGEMA_signal_8814), .B1_t (new_AGEMA_signal_8815), .B1_f (new_AGEMA_signal_8816), .Z0_t (KeyArray_outS12ser[4]), .Z0_f (new_AGEMA_signal_4761), .Z1_t (new_AGEMA_signal_4762), .Z1_f (new_AGEMA_signal_4763) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_4_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS12ser[4]), .B0_f (new_AGEMA_signal_4761), .B1_t (new_AGEMA_signal_4762), .B1_f (new_AGEMA_signal_4763), .Z0_t (KeyArray_S12reg_gff_1_SFF_4_n1), .Z0_f (new_AGEMA_signal_8814), .Z1_t (new_AGEMA_signal_8815), .Z1_f (new_AGEMA_signal_8816) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_4_U1 ( .A0_t (KeyArray_S12reg_gff_1_SFF_4_QD), .A0_f (new_AGEMA_signal_9532), .A1_t (new_AGEMA_signal_9533), .A1_f (new_AGEMA_signal_9534), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S12reg_gff_1_SFF_4_n2), .Z0_f (new_AGEMA_signal_10008), .Z1_t (new_AGEMA_signal_10009), .Z1_f (new_AGEMA_signal_10010) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS12ser[4]), .A0_f (new_AGEMA_signal_7042), .A1_t (new_AGEMA_signal_7043), .A1_f (new_AGEMA_signal_7044), .B0_t (KeyArray_outS22ser[4]), .B0_f (new_AGEMA_signal_5049), .B1_t (new_AGEMA_signal_5050), .B1_f (new_AGEMA_signal_5051), .Z0_t (KeyArray_S12reg_gff_1_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_7875), .Z1_t (new_AGEMA_signal_7876), .Z1_f (new_AGEMA_signal_7877) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S12reg_gff_1_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_7875), .B1_t (new_AGEMA_signal_7876), .B1_f (new_AGEMA_signal_7877), .Z0_t (KeyArray_S12reg_gff_1_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_8817), .Z1_t (new_AGEMA_signal_8818), .Z1_f (new_AGEMA_signal_8819) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S12reg_gff_1_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_8817), .A1_t (new_AGEMA_signal_8818), .A1_f (new_AGEMA_signal_8819), .B0_t (KeyArray_inS12ser[4]), .B0_f (new_AGEMA_signal_7042), .B1_t (new_AGEMA_signal_7043), .B1_f (new_AGEMA_signal_7044), .Z0_t (KeyArray_S12reg_gff_1_SFF_4_QD), .Z0_f (new_AGEMA_signal_9532), .Z1_t (new_AGEMA_signal_9533), .Z1_f (new_AGEMA_signal_9534) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S12reg_gff_1_SFF_5_U3 ( .A0_t (KeyArray_S12reg_gff_1_SFF_5_n2), .A0_f (new_AGEMA_signal_10011), .A1_t (new_AGEMA_signal_10012), .A1_f (new_AGEMA_signal_10013), .B0_t (KeyArray_S12reg_gff_1_SFF_5_n1), .B0_f (new_AGEMA_signal_8820), .B1_t (new_AGEMA_signal_8821), .B1_f (new_AGEMA_signal_8822), .Z0_t (KeyArray_outS12ser[5]), .Z0_f (new_AGEMA_signal_4770), .Z1_t (new_AGEMA_signal_4771), .Z1_f (new_AGEMA_signal_4772) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_5_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS12ser[5]), .B0_f (new_AGEMA_signal_4770), .B1_t (new_AGEMA_signal_4771), .B1_f (new_AGEMA_signal_4772), .Z0_t (KeyArray_S12reg_gff_1_SFF_5_n1), .Z0_f (new_AGEMA_signal_8820), .Z1_t (new_AGEMA_signal_8821), .Z1_f (new_AGEMA_signal_8822) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_5_U1 ( .A0_t (KeyArray_S12reg_gff_1_SFF_5_QD), .A0_f (new_AGEMA_signal_9535), .A1_t (new_AGEMA_signal_9536), .A1_f (new_AGEMA_signal_9537), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S12reg_gff_1_SFF_5_n2), .Z0_f (new_AGEMA_signal_10011), .Z1_t (new_AGEMA_signal_10012), .Z1_f (new_AGEMA_signal_10013) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS12ser[5]), .A0_f (new_AGEMA_signal_7045), .A1_t (new_AGEMA_signal_7046), .A1_f (new_AGEMA_signal_7047), .B0_t (KeyArray_outS22ser[5]), .B0_f (new_AGEMA_signal_5058), .B1_t (new_AGEMA_signal_5059), .B1_f (new_AGEMA_signal_5060), .Z0_t (KeyArray_S12reg_gff_1_SFF_5_MUXInst_X), .Z0_f (new_AGEMA_signal_7878), .Z1_t (new_AGEMA_signal_7879), .Z1_f (new_AGEMA_signal_7880) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S12reg_gff_1_SFF_5_MUXInst_X), .B0_f (new_AGEMA_signal_7878), .B1_t (new_AGEMA_signal_7879), .B1_f (new_AGEMA_signal_7880), .Z0_t (KeyArray_S12reg_gff_1_SFF_5_MUXInst_Y), .Z0_f (new_AGEMA_signal_8823), .Z1_t (new_AGEMA_signal_8824), .Z1_f (new_AGEMA_signal_8825) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S12reg_gff_1_SFF_5_MUXInst_Y), .A0_f (new_AGEMA_signal_8823), .A1_t (new_AGEMA_signal_8824), .A1_f (new_AGEMA_signal_8825), .B0_t (KeyArray_inS12ser[5]), .B0_f (new_AGEMA_signal_7045), .B1_t (new_AGEMA_signal_7046), .B1_f (new_AGEMA_signal_7047), .Z0_t (KeyArray_S12reg_gff_1_SFF_5_QD), .Z0_f (new_AGEMA_signal_9535), .Z1_t (new_AGEMA_signal_9536), .Z1_f (new_AGEMA_signal_9537) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S12reg_gff_1_SFF_6_U3 ( .A0_t (KeyArray_S12reg_gff_1_SFF_6_n2), .A0_f (new_AGEMA_signal_10014), .A1_t (new_AGEMA_signal_10015), .A1_f (new_AGEMA_signal_10016), .B0_t (KeyArray_S12reg_gff_1_SFF_6_n1), .B0_f (new_AGEMA_signal_8826), .B1_t (new_AGEMA_signal_8827), .B1_f (new_AGEMA_signal_8828), .Z0_t (KeyArray_outS12ser[6]), .Z0_f (new_AGEMA_signal_4779), .Z1_t (new_AGEMA_signal_4780), .Z1_f (new_AGEMA_signal_4781) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_6_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS12ser[6]), .B0_f (new_AGEMA_signal_4779), .B1_t (new_AGEMA_signal_4780), .B1_f (new_AGEMA_signal_4781), .Z0_t (KeyArray_S12reg_gff_1_SFF_6_n1), .Z0_f (new_AGEMA_signal_8826), .Z1_t (new_AGEMA_signal_8827), .Z1_f (new_AGEMA_signal_8828) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_6_U1 ( .A0_t (KeyArray_S12reg_gff_1_SFF_6_QD), .A0_f (new_AGEMA_signal_9538), .A1_t (new_AGEMA_signal_9539), .A1_f (new_AGEMA_signal_9540), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S12reg_gff_1_SFF_6_n2), .Z0_f (new_AGEMA_signal_10014), .Z1_t (new_AGEMA_signal_10015), .Z1_f (new_AGEMA_signal_10016) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS12ser[6]), .A0_f (new_AGEMA_signal_7048), .A1_t (new_AGEMA_signal_7049), .A1_f (new_AGEMA_signal_7050), .B0_t (KeyArray_outS22ser[6]), .B0_f (new_AGEMA_signal_5067), .B1_t (new_AGEMA_signal_5068), .B1_f (new_AGEMA_signal_5069), .Z0_t (KeyArray_S12reg_gff_1_SFF_6_MUXInst_X), .Z0_f (new_AGEMA_signal_7881), .Z1_t (new_AGEMA_signal_7882), .Z1_f (new_AGEMA_signal_7883) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S12reg_gff_1_SFF_6_MUXInst_X), .B0_f (new_AGEMA_signal_7881), .B1_t (new_AGEMA_signal_7882), .B1_f (new_AGEMA_signal_7883), .Z0_t (KeyArray_S12reg_gff_1_SFF_6_MUXInst_Y), .Z0_f (new_AGEMA_signal_8829), .Z1_t (new_AGEMA_signal_8830), .Z1_f (new_AGEMA_signal_8831) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S12reg_gff_1_SFF_6_MUXInst_Y), .A0_f (new_AGEMA_signal_8829), .A1_t (new_AGEMA_signal_8830), .A1_f (new_AGEMA_signal_8831), .B0_t (KeyArray_inS12ser[6]), .B0_f (new_AGEMA_signal_7048), .B1_t (new_AGEMA_signal_7049), .B1_f (new_AGEMA_signal_7050), .Z0_t (KeyArray_S12reg_gff_1_SFF_6_QD), .Z0_f (new_AGEMA_signal_9538), .Z1_t (new_AGEMA_signal_9539), .Z1_f (new_AGEMA_signal_9540) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S12reg_gff_1_SFF_7_U3 ( .A0_t (KeyArray_S12reg_gff_1_SFF_7_n2), .A0_f (new_AGEMA_signal_10017), .A1_t (new_AGEMA_signal_10018), .A1_f (new_AGEMA_signal_10019), .B0_t (KeyArray_S12reg_gff_1_SFF_7_n1), .B0_f (new_AGEMA_signal_8832), .B1_t (new_AGEMA_signal_8833), .B1_f (new_AGEMA_signal_8834), .Z0_t (KeyArray_outS12ser[7]), .Z0_f (new_AGEMA_signal_4788), .Z1_t (new_AGEMA_signal_4789), .Z1_f (new_AGEMA_signal_4790) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_7_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS12ser[7]), .B0_f (new_AGEMA_signal_4788), .B1_t (new_AGEMA_signal_4789), .B1_f (new_AGEMA_signal_4790), .Z0_t (KeyArray_S12reg_gff_1_SFF_7_n1), .Z0_f (new_AGEMA_signal_8832), .Z1_t (new_AGEMA_signal_8833), .Z1_f (new_AGEMA_signal_8834) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_7_U1 ( .A0_t (KeyArray_S12reg_gff_1_SFF_7_QD), .A0_f (new_AGEMA_signal_9541), .A1_t (new_AGEMA_signal_9542), .A1_f (new_AGEMA_signal_9543), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S12reg_gff_1_SFF_7_n2), .Z0_f (new_AGEMA_signal_10017), .Z1_t (new_AGEMA_signal_10018), .Z1_f (new_AGEMA_signal_10019) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS12ser[7]), .A0_f (new_AGEMA_signal_7051), .A1_t (new_AGEMA_signal_7052), .A1_f (new_AGEMA_signal_7053), .B0_t (KeyArray_outS22ser[7]), .B0_f (new_AGEMA_signal_5076), .B1_t (new_AGEMA_signal_5077), .B1_f (new_AGEMA_signal_5078), .Z0_t (KeyArray_S12reg_gff_1_SFF_7_MUXInst_X), .Z0_f (new_AGEMA_signal_7884), .Z1_t (new_AGEMA_signal_7885), .Z1_f (new_AGEMA_signal_7886) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S12reg_gff_1_SFF_7_MUXInst_X), .B0_f (new_AGEMA_signal_7884), .B1_t (new_AGEMA_signal_7885), .B1_f (new_AGEMA_signal_7886), .Z0_t (KeyArray_S12reg_gff_1_SFF_7_MUXInst_Y), .Z0_f (new_AGEMA_signal_8835), .Z1_t (new_AGEMA_signal_8836), .Z1_f (new_AGEMA_signal_8837) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S12reg_gff_1_SFF_7_MUXInst_Y), .A0_f (new_AGEMA_signal_8835), .A1_t (new_AGEMA_signal_8836), .A1_f (new_AGEMA_signal_8837), .B0_t (KeyArray_inS12ser[7]), .B0_f (new_AGEMA_signal_7051), .B1_t (new_AGEMA_signal_7052), .B1_f (new_AGEMA_signal_7053), .Z0_t (KeyArray_S12reg_gff_1_SFF_7_QD), .Z0_f (new_AGEMA_signal_9541), .Z1_t (new_AGEMA_signal_9542), .Z1_f (new_AGEMA_signal_9543) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S13reg_gff_1_SFF_0_U3 ( .A0_t (KeyArray_S13reg_gff_1_SFF_0_n2), .A0_f (new_AGEMA_signal_10020), .A1_t (new_AGEMA_signal_10021), .A1_f (new_AGEMA_signal_10022), .B0_t (KeyArray_S13reg_gff_1_SFF_0_n1), .B0_f (new_AGEMA_signal_8838), .B1_t (new_AGEMA_signal_8839), .B1_f (new_AGEMA_signal_8840), .Z0_t (keySBIn[0]), .Z0_f (new_AGEMA_signal_4797), .Z1_t (new_AGEMA_signal_4798), .Z1_f (new_AGEMA_signal_4799) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_0_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (keySBIn[0]), .B0_f (new_AGEMA_signal_4797), .B1_t (new_AGEMA_signal_4798), .B1_f (new_AGEMA_signal_4799), .Z0_t (KeyArray_S13reg_gff_1_SFF_0_n1), .Z0_f (new_AGEMA_signal_8838), .Z1_t (new_AGEMA_signal_8839), .Z1_f (new_AGEMA_signal_8840) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_0_U1 ( .A0_t (KeyArray_S13reg_gff_1_SFF_0_QD), .A0_f (new_AGEMA_signal_9544), .A1_t (new_AGEMA_signal_9545), .A1_f (new_AGEMA_signal_9546), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S13reg_gff_1_SFF_0_n2), .Z0_f (new_AGEMA_signal_10020), .Z1_t (new_AGEMA_signal_10021), .Z1_f (new_AGEMA_signal_10022) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS13ser[0]), .A0_f (new_AGEMA_signal_7054), .A1_t (new_AGEMA_signal_7055), .A1_f (new_AGEMA_signal_7056), .B0_t (KeyArray_outS23ser[0]), .B0_f (new_AGEMA_signal_5085), .B1_t (new_AGEMA_signal_5086), .B1_f (new_AGEMA_signal_5087), .Z0_t (KeyArray_S13reg_gff_1_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_7887), .Z1_t (new_AGEMA_signal_7888), .Z1_f (new_AGEMA_signal_7889) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S13reg_gff_1_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_7887), .B1_t (new_AGEMA_signal_7888), .B1_f (new_AGEMA_signal_7889), .Z0_t (KeyArray_S13reg_gff_1_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_8841), .Z1_t (new_AGEMA_signal_8842), .Z1_f (new_AGEMA_signal_8843) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S13reg_gff_1_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_8841), .A1_t (new_AGEMA_signal_8842), .A1_f (new_AGEMA_signal_8843), .B0_t (KeyArray_inS13ser[0]), .B0_f (new_AGEMA_signal_7054), .B1_t (new_AGEMA_signal_7055), .B1_f (new_AGEMA_signal_7056), .Z0_t (KeyArray_S13reg_gff_1_SFF_0_QD), .Z0_f (new_AGEMA_signal_9544), .Z1_t (new_AGEMA_signal_9545), .Z1_f (new_AGEMA_signal_9546) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S13reg_gff_1_SFF_1_U3 ( .A0_t (KeyArray_S13reg_gff_1_SFF_1_n2), .A0_f (new_AGEMA_signal_10023), .A1_t (new_AGEMA_signal_10024), .A1_f (new_AGEMA_signal_10025), .B0_t (KeyArray_S13reg_gff_1_SFF_1_n1), .B0_f (new_AGEMA_signal_8844), .B1_t (new_AGEMA_signal_8845), .B1_f (new_AGEMA_signal_8846), .Z0_t (keySBIn[1]), .Z0_f (new_AGEMA_signal_4806), .Z1_t (new_AGEMA_signal_4807), .Z1_f (new_AGEMA_signal_4808) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_1_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (keySBIn[1]), .B0_f (new_AGEMA_signal_4806), .B1_t (new_AGEMA_signal_4807), .B1_f (new_AGEMA_signal_4808), .Z0_t (KeyArray_S13reg_gff_1_SFF_1_n1), .Z0_f (new_AGEMA_signal_8844), .Z1_t (new_AGEMA_signal_8845), .Z1_f (new_AGEMA_signal_8846) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_1_U1 ( .A0_t (KeyArray_S13reg_gff_1_SFF_1_QD), .A0_f (new_AGEMA_signal_9547), .A1_t (new_AGEMA_signal_9548), .A1_f (new_AGEMA_signal_9549), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S13reg_gff_1_SFF_1_n2), .Z0_f (new_AGEMA_signal_10023), .Z1_t (new_AGEMA_signal_10024), .Z1_f (new_AGEMA_signal_10025) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS13ser[1]), .A0_f (new_AGEMA_signal_7057), .A1_t (new_AGEMA_signal_7058), .A1_f (new_AGEMA_signal_7059), .B0_t (KeyArray_outS23ser[1]), .B0_f (new_AGEMA_signal_5094), .B1_t (new_AGEMA_signal_5095), .B1_f (new_AGEMA_signal_5096), .Z0_t (KeyArray_S13reg_gff_1_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_7890), .Z1_t (new_AGEMA_signal_7891), .Z1_f (new_AGEMA_signal_7892) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S13reg_gff_1_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_7890), .B1_t (new_AGEMA_signal_7891), .B1_f (new_AGEMA_signal_7892), .Z0_t (KeyArray_S13reg_gff_1_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_8847), .Z1_t (new_AGEMA_signal_8848), .Z1_f (new_AGEMA_signal_8849) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S13reg_gff_1_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_8847), .A1_t (new_AGEMA_signal_8848), .A1_f (new_AGEMA_signal_8849), .B0_t (KeyArray_inS13ser[1]), .B0_f (new_AGEMA_signal_7057), .B1_t (new_AGEMA_signal_7058), .B1_f (new_AGEMA_signal_7059), .Z0_t (KeyArray_S13reg_gff_1_SFF_1_QD), .Z0_f (new_AGEMA_signal_9547), .Z1_t (new_AGEMA_signal_9548), .Z1_f (new_AGEMA_signal_9549) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S13reg_gff_1_SFF_2_U3 ( .A0_t (KeyArray_S13reg_gff_1_SFF_2_n2), .A0_f (new_AGEMA_signal_10026), .A1_t (new_AGEMA_signal_10027), .A1_f (new_AGEMA_signal_10028), .B0_t (KeyArray_S13reg_gff_1_SFF_2_n1), .B0_f (new_AGEMA_signal_8850), .B1_t (new_AGEMA_signal_8851), .B1_f (new_AGEMA_signal_8852), .Z0_t (keySBIn[2]), .Z0_f (new_AGEMA_signal_4815), .Z1_t (new_AGEMA_signal_4816), .Z1_f (new_AGEMA_signal_4817) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_2_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (keySBIn[2]), .B0_f (new_AGEMA_signal_4815), .B1_t (new_AGEMA_signal_4816), .B1_f (new_AGEMA_signal_4817), .Z0_t (KeyArray_S13reg_gff_1_SFF_2_n1), .Z0_f (new_AGEMA_signal_8850), .Z1_t (new_AGEMA_signal_8851), .Z1_f (new_AGEMA_signal_8852) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_2_U1 ( .A0_t (KeyArray_S13reg_gff_1_SFF_2_QD), .A0_f (new_AGEMA_signal_9550), .A1_t (new_AGEMA_signal_9551), .A1_f (new_AGEMA_signal_9552), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S13reg_gff_1_SFF_2_n2), .Z0_f (new_AGEMA_signal_10026), .Z1_t (new_AGEMA_signal_10027), .Z1_f (new_AGEMA_signal_10028) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS13ser[2]), .A0_f (new_AGEMA_signal_7060), .A1_t (new_AGEMA_signal_7061), .A1_f (new_AGEMA_signal_7062), .B0_t (KeyArray_outS23ser[2]), .B0_f (new_AGEMA_signal_5103), .B1_t (new_AGEMA_signal_5104), .B1_f (new_AGEMA_signal_5105), .Z0_t (KeyArray_S13reg_gff_1_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_7893), .Z1_t (new_AGEMA_signal_7894), .Z1_f (new_AGEMA_signal_7895) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S13reg_gff_1_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_7893), .B1_t (new_AGEMA_signal_7894), .B1_f (new_AGEMA_signal_7895), .Z0_t (KeyArray_S13reg_gff_1_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_8853), .Z1_t (new_AGEMA_signal_8854), .Z1_f (new_AGEMA_signal_8855) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S13reg_gff_1_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_8853), .A1_t (new_AGEMA_signal_8854), .A1_f (new_AGEMA_signal_8855), .B0_t (KeyArray_inS13ser[2]), .B0_f (new_AGEMA_signal_7060), .B1_t (new_AGEMA_signal_7061), .B1_f (new_AGEMA_signal_7062), .Z0_t (KeyArray_S13reg_gff_1_SFF_2_QD), .Z0_f (new_AGEMA_signal_9550), .Z1_t (new_AGEMA_signal_9551), .Z1_f (new_AGEMA_signal_9552) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S13reg_gff_1_SFF_3_U3 ( .A0_t (KeyArray_S13reg_gff_1_SFF_3_n2), .A0_f (new_AGEMA_signal_10029), .A1_t (new_AGEMA_signal_10030), .A1_f (new_AGEMA_signal_10031), .B0_t (KeyArray_S13reg_gff_1_SFF_3_n1), .B0_f (new_AGEMA_signal_8856), .B1_t (new_AGEMA_signal_8857), .B1_f (new_AGEMA_signal_8858), .Z0_t (keySBIn[3]), .Z0_f (new_AGEMA_signal_4824), .Z1_t (new_AGEMA_signal_4825), .Z1_f (new_AGEMA_signal_4826) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_3_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (keySBIn[3]), .B0_f (new_AGEMA_signal_4824), .B1_t (new_AGEMA_signal_4825), .B1_f (new_AGEMA_signal_4826), .Z0_t (KeyArray_S13reg_gff_1_SFF_3_n1), .Z0_f (new_AGEMA_signal_8856), .Z1_t (new_AGEMA_signal_8857), .Z1_f (new_AGEMA_signal_8858) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_3_U1 ( .A0_t (KeyArray_S13reg_gff_1_SFF_3_QD), .A0_f (new_AGEMA_signal_9553), .A1_t (new_AGEMA_signal_9554), .A1_f (new_AGEMA_signal_9555), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S13reg_gff_1_SFF_3_n2), .Z0_f (new_AGEMA_signal_10029), .Z1_t (new_AGEMA_signal_10030), .Z1_f (new_AGEMA_signal_10031) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS13ser[3]), .A0_f (new_AGEMA_signal_7063), .A1_t (new_AGEMA_signal_7064), .A1_f (new_AGEMA_signal_7065), .B0_t (KeyArray_outS23ser[3]), .B0_f (new_AGEMA_signal_5112), .B1_t (new_AGEMA_signal_5113), .B1_f (new_AGEMA_signal_5114), .Z0_t (KeyArray_S13reg_gff_1_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_7896), .Z1_t (new_AGEMA_signal_7897), .Z1_f (new_AGEMA_signal_7898) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S13reg_gff_1_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_7896), .B1_t (new_AGEMA_signal_7897), .B1_f (new_AGEMA_signal_7898), .Z0_t (KeyArray_S13reg_gff_1_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_8859), .Z1_t (new_AGEMA_signal_8860), .Z1_f (new_AGEMA_signal_8861) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S13reg_gff_1_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_8859), .A1_t (new_AGEMA_signal_8860), .A1_f (new_AGEMA_signal_8861), .B0_t (KeyArray_inS13ser[3]), .B0_f (new_AGEMA_signal_7063), .B1_t (new_AGEMA_signal_7064), .B1_f (new_AGEMA_signal_7065), .Z0_t (KeyArray_S13reg_gff_1_SFF_3_QD), .Z0_f (new_AGEMA_signal_9553), .Z1_t (new_AGEMA_signal_9554), .Z1_f (new_AGEMA_signal_9555) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S13reg_gff_1_SFF_4_U3 ( .A0_t (KeyArray_S13reg_gff_1_SFF_4_n2), .A0_f (new_AGEMA_signal_10032), .A1_t (new_AGEMA_signal_10033), .A1_f (new_AGEMA_signal_10034), .B0_t (KeyArray_S13reg_gff_1_SFF_4_n1), .B0_f (new_AGEMA_signal_8862), .B1_t (new_AGEMA_signal_8863), .B1_f (new_AGEMA_signal_8864), .Z0_t (keySBIn[4]), .Z0_f (new_AGEMA_signal_4833), .Z1_t (new_AGEMA_signal_4834), .Z1_f (new_AGEMA_signal_4835) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_4_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (keySBIn[4]), .B0_f (new_AGEMA_signal_4833), .B1_t (new_AGEMA_signal_4834), .B1_f (new_AGEMA_signal_4835), .Z0_t (KeyArray_S13reg_gff_1_SFF_4_n1), .Z0_f (new_AGEMA_signal_8862), .Z1_t (new_AGEMA_signal_8863), .Z1_f (new_AGEMA_signal_8864) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_4_U1 ( .A0_t (KeyArray_S13reg_gff_1_SFF_4_QD), .A0_f (new_AGEMA_signal_9556), .A1_t (new_AGEMA_signal_9557), .A1_f (new_AGEMA_signal_9558), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S13reg_gff_1_SFF_4_n2), .Z0_f (new_AGEMA_signal_10032), .Z1_t (new_AGEMA_signal_10033), .Z1_f (new_AGEMA_signal_10034) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS13ser[4]), .A0_f (new_AGEMA_signal_7066), .A1_t (new_AGEMA_signal_7067), .A1_f (new_AGEMA_signal_7068), .B0_t (KeyArray_outS23ser[4]), .B0_f (new_AGEMA_signal_5121), .B1_t (new_AGEMA_signal_5122), .B1_f (new_AGEMA_signal_5123), .Z0_t (KeyArray_S13reg_gff_1_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_7899), .Z1_t (new_AGEMA_signal_7900), .Z1_f (new_AGEMA_signal_7901) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S13reg_gff_1_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_7899), .B1_t (new_AGEMA_signal_7900), .B1_f (new_AGEMA_signal_7901), .Z0_t (KeyArray_S13reg_gff_1_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_8865), .Z1_t (new_AGEMA_signal_8866), .Z1_f (new_AGEMA_signal_8867) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S13reg_gff_1_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_8865), .A1_t (new_AGEMA_signal_8866), .A1_f (new_AGEMA_signal_8867), .B0_t (KeyArray_inS13ser[4]), .B0_f (new_AGEMA_signal_7066), .B1_t (new_AGEMA_signal_7067), .B1_f (new_AGEMA_signal_7068), .Z0_t (KeyArray_S13reg_gff_1_SFF_4_QD), .Z0_f (new_AGEMA_signal_9556), .Z1_t (new_AGEMA_signal_9557), .Z1_f (new_AGEMA_signal_9558) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S13reg_gff_1_SFF_5_U3 ( .A0_t (KeyArray_S13reg_gff_1_SFF_5_n2), .A0_f (new_AGEMA_signal_10035), .A1_t (new_AGEMA_signal_10036), .A1_f (new_AGEMA_signal_10037), .B0_t (KeyArray_S13reg_gff_1_SFF_5_n1), .B0_f (new_AGEMA_signal_8868), .B1_t (new_AGEMA_signal_8869), .B1_f (new_AGEMA_signal_8870), .Z0_t (keySBIn[5]), .Z0_f (new_AGEMA_signal_4842), .Z1_t (new_AGEMA_signal_4843), .Z1_f (new_AGEMA_signal_4844) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_5_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (keySBIn[5]), .B0_f (new_AGEMA_signal_4842), .B1_t (new_AGEMA_signal_4843), .B1_f (new_AGEMA_signal_4844), .Z0_t (KeyArray_S13reg_gff_1_SFF_5_n1), .Z0_f (new_AGEMA_signal_8868), .Z1_t (new_AGEMA_signal_8869), .Z1_f (new_AGEMA_signal_8870) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_5_U1 ( .A0_t (KeyArray_S13reg_gff_1_SFF_5_QD), .A0_f (new_AGEMA_signal_9559), .A1_t (new_AGEMA_signal_9560), .A1_f (new_AGEMA_signal_9561), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S13reg_gff_1_SFF_5_n2), .Z0_f (new_AGEMA_signal_10035), .Z1_t (new_AGEMA_signal_10036), .Z1_f (new_AGEMA_signal_10037) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS13ser[5]), .A0_f (new_AGEMA_signal_7069), .A1_t (new_AGEMA_signal_7070), .A1_f (new_AGEMA_signal_7071), .B0_t (KeyArray_outS23ser[5]), .B0_f (new_AGEMA_signal_5130), .B1_t (new_AGEMA_signal_5131), .B1_f (new_AGEMA_signal_5132), .Z0_t (KeyArray_S13reg_gff_1_SFF_5_MUXInst_X), .Z0_f (new_AGEMA_signal_7902), .Z1_t (new_AGEMA_signal_7903), .Z1_f (new_AGEMA_signal_7904) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S13reg_gff_1_SFF_5_MUXInst_X), .B0_f (new_AGEMA_signal_7902), .B1_t (new_AGEMA_signal_7903), .B1_f (new_AGEMA_signal_7904), .Z0_t (KeyArray_S13reg_gff_1_SFF_5_MUXInst_Y), .Z0_f (new_AGEMA_signal_8871), .Z1_t (new_AGEMA_signal_8872), .Z1_f (new_AGEMA_signal_8873) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S13reg_gff_1_SFF_5_MUXInst_Y), .A0_f (new_AGEMA_signal_8871), .A1_t (new_AGEMA_signal_8872), .A1_f (new_AGEMA_signal_8873), .B0_t (KeyArray_inS13ser[5]), .B0_f (new_AGEMA_signal_7069), .B1_t (new_AGEMA_signal_7070), .B1_f (new_AGEMA_signal_7071), .Z0_t (KeyArray_S13reg_gff_1_SFF_5_QD), .Z0_f (new_AGEMA_signal_9559), .Z1_t (new_AGEMA_signal_9560), .Z1_f (new_AGEMA_signal_9561) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S13reg_gff_1_SFF_6_U3 ( .A0_t (KeyArray_S13reg_gff_1_SFF_6_n2), .A0_f (new_AGEMA_signal_10038), .A1_t (new_AGEMA_signal_10039), .A1_f (new_AGEMA_signal_10040), .B0_t (KeyArray_S13reg_gff_1_SFF_6_n1), .B0_f (new_AGEMA_signal_8874), .B1_t (new_AGEMA_signal_8875), .B1_f (new_AGEMA_signal_8876), .Z0_t (keySBIn[6]), .Z0_f (new_AGEMA_signal_4851), .Z1_t (new_AGEMA_signal_4852), .Z1_f (new_AGEMA_signal_4853) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_6_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (keySBIn[6]), .B0_f (new_AGEMA_signal_4851), .B1_t (new_AGEMA_signal_4852), .B1_f (new_AGEMA_signal_4853), .Z0_t (KeyArray_S13reg_gff_1_SFF_6_n1), .Z0_f (new_AGEMA_signal_8874), .Z1_t (new_AGEMA_signal_8875), .Z1_f (new_AGEMA_signal_8876) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_6_U1 ( .A0_t (KeyArray_S13reg_gff_1_SFF_6_QD), .A0_f (new_AGEMA_signal_9562), .A1_t (new_AGEMA_signal_9563), .A1_f (new_AGEMA_signal_9564), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S13reg_gff_1_SFF_6_n2), .Z0_f (new_AGEMA_signal_10038), .Z1_t (new_AGEMA_signal_10039), .Z1_f (new_AGEMA_signal_10040) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS13ser[6]), .A0_f (new_AGEMA_signal_7072), .A1_t (new_AGEMA_signal_7073), .A1_f (new_AGEMA_signal_7074), .B0_t (KeyArray_outS23ser[6]), .B0_f (new_AGEMA_signal_5139), .B1_t (new_AGEMA_signal_5140), .B1_f (new_AGEMA_signal_5141), .Z0_t (KeyArray_S13reg_gff_1_SFF_6_MUXInst_X), .Z0_f (new_AGEMA_signal_7905), .Z1_t (new_AGEMA_signal_7906), .Z1_f (new_AGEMA_signal_7907) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S13reg_gff_1_SFF_6_MUXInst_X), .B0_f (new_AGEMA_signal_7905), .B1_t (new_AGEMA_signal_7906), .B1_f (new_AGEMA_signal_7907), .Z0_t (KeyArray_S13reg_gff_1_SFF_6_MUXInst_Y), .Z0_f (new_AGEMA_signal_8877), .Z1_t (new_AGEMA_signal_8878), .Z1_f (new_AGEMA_signal_8879) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S13reg_gff_1_SFF_6_MUXInst_Y), .A0_f (new_AGEMA_signal_8877), .A1_t (new_AGEMA_signal_8878), .A1_f (new_AGEMA_signal_8879), .B0_t (KeyArray_inS13ser[6]), .B0_f (new_AGEMA_signal_7072), .B1_t (new_AGEMA_signal_7073), .B1_f (new_AGEMA_signal_7074), .Z0_t (KeyArray_S13reg_gff_1_SFF_6_QD), .Z0_f (new_AGEMA_signal_9562), .Z1_t (new_AGEMA_signal_9563), .Z1_f (new_AGEMA_signal_9564) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S13reg_gff_1_SFF_7_U3 ( .A0_t (KeyArray_S13reg_gff_1_SFF_7_n2), .A0_f (new_AGEMA_signal_10041), .A1_t (new_AGEMA_signal_10042), .A1_f (new_AGEMA_signal_10043), .B0_t (KeyArray_S13reg_gff_1_SFF_7_n1), .B0_f (new_AGEMA_signal_8880), .B1_t (new_AGEMA_signal_8881), .B1_f (new_AGEMA_signal_8882), .Z0_t (keySBIn[7]), .Z0_f (new_AGEMA_signal_4860), .Z1_t (new_AGEMA_signal_4861), .Z1_f (new_AGEMA_signal_4862) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_7_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (keySBIn[7]), .B0_f (new_AGEMA_signal_4860), .B1_t (new_AGEMA_signal_4861), .B1_f (new_AGEMA_signal_4862), .Z0_t (KeyArray_S13reg_gff_1_SFF_7_n1), .Z0_f (new_AGEMA_signal_8880), .Z1_t (new_AGEMA_signal_8881), .Z1_f (new_AGEMA_signal_8882) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_7_U1 ( .A0_t (KeyArray_S13reg_gff_1_SFF_7_QD), .A0_f (new_AGEMA_signal_9565), .A1_t (new_AGEMA_signal_9566), .A1_f (new_AGEMA_signal_9567), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S13reg_gff_1_SFF_7_n2), .Z0_f (new_AGEMA_signal_10041), .Z1_t (new_AGEMA_signal_10042), .Z1_f (new_AGEMA_signal_10043) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS13ser[7]), .A0_f (new_AGEMA_signal_7075), .A1_t (new_AGEMA_signal_7076), .A1_f (new_AGEMA_signal_7077), .B0_t (KeyArray_outS23ser[7]), .B0_f (new_AGEMA_signal_5148), .B1_t (new_AGEMA_signal_5149), .B1_f (new_AGEMA_signal_5150), .Z0_t (KeyArray_S13reg_gff_1_SFF_7_MUXInst_X), .Z0_f (new_AGEMA_signal_7908), .Z1_t (new_AGEMA_signal_7909), .Z1_f (new_AGEMA_signal_7910) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S13reg_gff_1_SFF_7_MUXInst_X), .B0_f (new_AGEMA_signal_7908), .B1_t (new_AGEMA_signal_7909), .B1_f (new_AGEMA_signal_7910), .Z0_t (KeyArray_S13reg_gff_1_SFF_7_MUXInst_Y), .Z0_f (new_AGEMA_signal_8883), .Z1_t (new_AGEMA_signal_8884), .Z1_f (new_AGEMA_signal_8885) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S13reg_gff_1_SFF_7_MUXInst_Y), .A0_f (new_AGEMA_signal_8883), .A1_t (new_AGEMA_signal_8884), .A1_f (new_AGEMA_signal_8885), .B0_t (KeyArray_inS13ser[7]), .B0_f (new_AGEMA_signal_7075), .B1_t (new_AGEMA_signal_7076), .B1_f (new_AGEMA_signal_7077), .Z0_t (KeyArray_S13reg_gff_1_SFF_7_QD), .Z0_f (new_AGEMA_signal_9565), .Z1_t (new_AGEMA_signal_9566), .Z1_f (new_AGEMA_signal_9567) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S20reg_gff_1_SFF_0_U3 ( .A0_t (KeyArray_S20reg_gff_1_SFF_0_n2), .A0_f (new_AGEMA_signal_10044), .A1_t (new_AGEMA_signal_10045), .A1_f (new_AGEMA_signal_10046), .B0_t (KeyArray_S20reg_gff_1_SFF_0_n1), .B0_f (new_AGEMA_signal_8886), .B1_t (new_AGEMA_signal_8887), .B1_f (new_AGEMA_signal_8888), .Z0_t (KeyArray_outS20ser[0]), .Z0_f (new_AGEMA_signal_4869), .Z1_t (new_AGEMA_signal_4870), .Z1_f (new_AGEMA_signal_4871) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_0_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS20ser[0]), .B0_f (new_AGEMA_signal_4869), .B1_t (new_AGEMA_signal_4870), .B1_f (new_AGEMA_signal_4871), .Z0_t (KeyArray_S20reg_gff_1_SFF_0_n1), .Z0_f (new_AGEMA_signal_8886), .Z1_t (new_AGEMA_signal_8887), .Z1_f (new_AGEMA_signal_8888) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_0_U1 ( .A0_t (KeyArray_S20reg_gff_1_SFF_0_QD), .A0_f (new_AGEMA_signal_9568), .A1_t (new_AGEMA_signal_9569), .A1_f (new_AGEMA_signal_9570), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S20reg_gff_1_SFF_0_n2), .Z0_f (new_AGEMA_signal_10044), .Z1_t (new_AGEMA_signal_10045), .Z1_f (new_AGEMA_signal_10046) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS20ser[0]), .A0_f (new_AGEMA_signal_7078), .A1_t (new_AGEMA_signal_7079), .A1_f (new_AGEMA_signal_7080), .B0_t (KeyArray_outS30ser[0]), .B0_f (new_AGEMA_signal_5157), .B1_t (new_AGEMA_signal_5158), .B1_f (new_AGEMA_signal_5159), .Z0_t (KeyArray_S20reg_gff_1_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_7911), .Z1_t (new_AGEMA_signal_7912), .Z1_f (new_AGEMA_signal_7913) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S20reg_gff_1_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_7911), .B1_t (new_AGEMA_signal_7912), .B1_f (new_AGEMA_signal_7913), .Z0_t (KeyArray_S20reg_gff_1_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_8889), .Z1_t (new_AGEMA_signal_8890), .Z1_f (new_AGEMA_signal_8891) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S20reg_gff_1_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_8889), .A1_t (new_AGEMA_signal_8890), .A1_f (new_AGEMA_signal_8891), .B0_t (KeyArray_inS20ser[0]), .B0_f (new_AGEMA_signal_7078), .B1_t (new_AGEMA_signal_7079), .B1_f (new_AGEMA_signal_7080), .Z0_t (KeyArray_S20reg_gff_1_SFF_0_QD), .Z0_f (new_AGEMA_signal_9568), .Z1_t (new_AGEMA_signal_9569), .Z1_f (new_AGEMA_signal_9570) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S20reg_gff_1_SFF_1_U3 ( .A0_t (KeyArray_S20reg_gff_1_SFF_1_n2), .A0_f (new_AGEMA_signal_10047), .A1_t (new_AGEMA_signal_10048), .A1_f (new_AGEMA_signal_10049), .B0_t (KeyArray_S20reg_gff_1_SFF_1_n1), .B0_f (new_AGEMA_signal_8892), .B1_t (new_AGEMA_signal_8893), .B1_f (new_AGEMA_signal_8894), .Z0_t (KeyArray_outS20ser[1]), .Z0_f (new_AGEMA_signal_4878), .Z1_t (new_AGEMA_signal_4879), .Z1_f (new_AGEMA_signal_4880) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_1_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS20ser[1]), .B0_f (new_AGEMA_signal_4878), .B1_t (new_AGEMA_signal_4879), .B1_f (new_AGEMA_signal_4880), .Z0_t (KeyArray_S20reg_gff_1_SFF_1_n1), .Z0_f (new_AGEMA_signal_8892), .Z1_t (new_AGEMA_signal_8893), .Z1_f (new_AGEMA_signal_8894) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_1_U1 ( .A0_t (KeyArray_S20reg_gff_1_SFF_1_QD), .A0_f (new_AGEMA_signal_9571), .A1_t (new_AGEMA_signal_9572), .A1_f (new_AGEMA_signal_9573), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S20reg_gff_1_SFF_1_n2), .Z0_f (new_AGEMA_signal_10047), .Z1_t (new_AGEMA_signal_10048), .Z1_f (new_AGEMA_signal_10049) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS20ser[1]), .A0_f (new_AGEMA_signal_7081), .A1_t (new_AGEMA_signal_7082), .A1_f (new_AGEMA_signal_7083), .B0_t (KeyArray_outS30ser[1]), .B0_f (new_AGEMA_signal_5166), .B1_t (new_AGEMA_signal_5167), .B1_f (new_AGEMA_signal_5168), .Z0_t (KeyArray_S20reg_gff_1_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_7914), .Z1_t (new_AGEMA_signal_7915), .Z1_f (new_AGEMA_signal_7916) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S20reg_gff_1_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_7914), .B1_t (new_AGEMA_signal_7915), .B1_f (new_AGEMA_signal_7916), .Z0_t (KeyArray_S20reg_gff_1_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_8895), .Z1_t (new_AGEMA_signal_8896), .Z1_f (new_AGEMA_signal_8897) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S20reg_gff_1_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_8895), .A1_t (new_AGEMA_signal_8896), .A1_f (new_AGEMA_signal_8897), .B0_t (KeyArray_inS20ser[1]), .B0_f (new_AGEMA_signal_7081), .B1_t (new_AGEMA_signal_7082), .B1_f (new_AGEMA_signal_7083), .Z0_t (KeyArray_S20reg_gff_1_SFF_1_QD), .Z0_f (new_AGEMA_signal_9571), .Z1_t (new_AGEMA_signal_9572), .Z1_f (new_AGEMA_signal_9573) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S20reg_gff_1_SFF_2_U3 ( .A0_t (KeyArray_S20reg_gff_1_SFF_2_n2), .A0_f (new_AGEMA_signal_10050), .A1_t (new_AGEMA_signal_10051), .A1_f (new_AGEMA_signal_10052), .B0_t (KeyArray_S20reg_gff_1_SFF_2_n1), .B0_f (new_AGEMA_signal_8898), .B1_t (new_AGEMA_signal_8899), .B1_f (new_AGEMA_signal_8900), .Z0_t (KeyArray_outS20ser[2]), .Z0_f (new_AGEMA_signal_4887), .Z1_t (new_AGEMA_signal_4888), .Z1_f (new_AGEMA_signal_4889) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_2_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS20ser[2]), .B0_f (new_AGEMA_signal_4887), .B1_t (new_AGEMA_signal_4888), .B1_f (new_AGEMA_signal_4889), .Z0_t (KeyArray_S20reg_gff_1_SFF_2_n1), .Z0_f (new_AGEMA_signal_8898), .Z1_t (new_AGEMA_signal_8899), .Z1_f (new_AGEMA_signal_8900) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_2_U1 ( .A0_t (KeyArray_S20reg_gff_1_SFF_2_QD), .A0_f (new_AGEMA_signal_9574), .A1_t (new_AGEMA_signal_9575), .A1_f (new_AGEMA_signal_9576), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S20reg_gff_1_SFF_2_n2), .Z0_f (new_AGEMA_signal_10050), .Z1_t (new_AGEMA_signal_10051), .Z1_f (new_AGEMA_signal_10052) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS20ser[2]), .A0_f (new_AGEMA_signal_7084), .A1_t (new_AGEMA_signal_7085), .A1_f (new_AGEMA_signal_7086), .B0_t (KeyArray_outS30ser[2]), .B0_f (new_AGEMA_signal_5175), .B1_t (new_AGEMA_signal_5176), .B1_f (new_AGEMA_signal_5177), .Z0_t (KeyArray_S20reg_gff_1_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_7917), .Z1_t (new_AGEMA_signal_7918), .Z1_f (new_AGEMA_signal_7919) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S20reg_gff_1_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_7917), .B1_t (new_AGEMA_signal_7918), .B1_f (new_AGEMA_signal_7919), .Z0_t (KeyArray_S20reg_gff_1_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_8901), .Z1_t (new_AGEMA_signal_8902), .Z1_f (new_AGEMA_signal_8903) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S20reg_gff_1_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_8901), .A1_t (new_AGEMA_signal_8902), .A1_f (new_AGEMA_signal_8903), .B0_t (KeyArray_inS20ser[2]), .B0_f (new_AGEMA_signal_7084), .B1_t (new_AGEMA_signal_7085), .B1_f (new_AGEMA_signal_7086), .Z0_t (KeyArray_S20reg_gff_1_SFF_2_QD), .Z0_f (new_AGEMA_signal_9574), .Z1_t (new_AGEMA_signal_9575), .Z1_f (new_AGEMA_signal_9576) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S20reg_gff_1_SFF_3_U3 ( .A0_t (KeyArray_S20reg_gff_1_SFF_3_n2), .A0_f (new_AGEMA_signal_10053), .A1_t (new_AGEMA_signal_10054), .A1_f (new_AGEMA_signal_10055), .B0_t (KeyArray_S20reg_gff_1_SFF_3_n1), .B0_f (new_AGEMA_signal_8904), .B1_t (new_AGEMA_signal_8905), .B1_f (new_AGEMA_signal_8906), .Z0_t (KeyArray_outS20ser[3]), .Z0_f (new_AGEMA_signal_4896), .Z1_t (new_AGEMA_signal_4897), .Z1_f (new_AGEMA_signal_4898) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_3_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS20ser[3]), .B0_f (new_AGEMA_signal_4896), .B1_t (new_AGEMA_signal_4897), .B1_f (new_AGEMA_signal_4898), .Z0_t (KeyArray_S20reg_gff_1_SFF_3_n1), .Z0_f (new_AGEMA_signal_8904), .Z1_t (new_AGEMA_signal_8905), .Z1_f (new_AGEMA_signal_8906) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_3_U1 ( .A0_t (KeyArray_S20reg_gff_1_SFF_3_QD), .A0_f (new_AGEMA_signal_9577), .A1_t (new_AGEMA_signal_9578), .A1_f (new_AGEMA_signal_9579), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S20reg_gff_1_SFF_3_n2), .Z0_f (new_AGEMA_signal_10053), .Z1_t (new_AGEMA_signal_10054), .Z1_f (new_AGEMA_signal_10055) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS20ser[3]), .A0_f (new_AGEMA_signal_7087), .A1_t (new_AGEMA_signal_7088), .A1_f (new_AGEMA_signal_7089), .B0_t (KeyArray_outS30ser[3]), .B0_f (new_AGEMA_signal_5184), .B1_t (new_AGEMA_signal_5185), .B1_f (new_AGEMA_signal_5186), .Z0_t (KeyArray_S20reg_gff_1_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_7920), .Z1_t (new_AGEMA_signal_7921), .Z1_f (new_AGEMA_signal_7922) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S20reg_gff_1_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_7920), .B1_t (new_AGEMA_signal_7921), .B1_f (new_AGEMA_signal_7922), .Z0_t (KeyArray_S20reg_gff_1_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_8907), .Z1_t (new_AGEMA_signal_8908), .Z1_f (new_AGEMA_signal_8909) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S20reg_gff_1_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_8907), .A1_t (new_AGEMA_signal_8908), .A1_f (new_AGEMA_signal_8909), .B0_t (KeyArray_inS20ser[3]), .B0_f (new_AGEMA_signal_7087), .B1_t (new_AGEMA_signal_7088), .B1_f (new_AGEMA_signal_7089), .Z0_t (KeyArray_S20reg_gff_1_SFF_3_QD), .Z0_f (new_AGEMA_signal_9577), .Z1_t (new_AGEMA_signal_9578), .Z1_f (new_AGEMA_signal_9579) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S20reg_gff_1_SFF_4_U3 ( .A0_t (KeyArray_S20reg_gff_1_SFF_4_n2), .A0_f (new_AGEMA_signal_10056), .A1_t (new_AGEMA_signal_10057), .A1_f (new_AGEMA_signal_10058), .B0_t (KeyArray_S20reg_gff_1_SFF_4_n1), .B0_f (new_AGEMA_signal_8910), .B1_t (new_AGEMA_signal_8911), .B1_f (new_AGEMA_signal_8912), .Z0_t (KeyArray_outS20ser[4]), .Z0_f (new_AGEMA_signal_4905), .Z1_t (new_AGEMA_signal_4906), .Z1_f (new_AGEMA_signal_4907) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_4_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS20ser[4]), .B0_f (new_AGEMA_signal_4905), .B1_t (new_AGEMA_signal_4906), .B1_f (new_AGEMA_signal_4907), .Z0_t (KeyArray_S20reg_gff_1_SFF_4_n1), .Z0_f (new_AGEMA_signal_8910), .Z1_t (new_AGEMA_signal_8911), .Z1_f (new_AGEMA_signal_8912) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_4_U1 ( .A0_t (KeyArray_S20reg_gff_1_SFF_4_QD), .A0_f (new_AGEMA_signal_9580), .A1_t (new_AGEMA_signal_9581), .A1_f (new_AGEMA_signal_9582), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S20reg_gff_1_SFF_4_n2), .Z0_f (new_AGEMA_signal_10056), .Z1_t (new_AGEMA_signal_10057), .Z1_f (new_AGEMA_signal_10058) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS20ser[4]), .A0_f (new_AGEMA_signal_7090), .A1_t (new_AGEMA_signal_7091), .A1_f (new_AGEMA_signal_7092), .B0_t (KeyArray_outS30ser[4]), .B0_f (new_AGEMA_signal_5193), .B1_t (new_AGEMA_signal_5194), .B1_f (new_AGEMA_signal_5195), .Z0_t (KeyArray_S20reg_gff_1_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_7923), .Z1_t (new_AGEMA_signal_7924), .Z1_f (new_AGEMA_signal_7925) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S20reg_gff_1_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_7923), .B1_t (new_AGEMA_signal_7924), .B1_f (new_AGEMA_signal_7925), .Z0_t (KeyArray_S20reg_gff_1_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_8913), .Z1_t (new_AGEMA_signal_8914), .Z1_f (new_AGEMA_signal_8915) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S20reg_gff_1_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_8913), .A1_t (new_AGEMA_signal_8914), .A1_f (new_AGEMA_signal_8915), .B0_t (KeyArray_inS20ser[4]), .B0_f (new_AGEMA_signal_7090), .B1_t (new_AGEMA_signal_7091), .B1_f (new_AGEMA_signal_7092), .Z0_t (KeyArray_S20reg_gff_1_SFF_4_QD), .Z0_f (new_AGEMA_signal_9580), .Z1_t (new_AGEMA_signal_9581), .Z1_f (new_AGEMA_signal_9582) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S20reg_gff_1_SFF_5_U3 ( .A0_t (KeyArray_S20reg_gff_1_SFF_5_n2), .A0_f (new_AGEMA_signal_10059), .A1_t (new_AGEMA_signal_10060), .A1_f (new_AGEMA_signal_10061), .B0_t (KeyArray_S20reg_gff_1_SFF_5_n1), .B0_f (new_AGEMA_signal_8916), .B1_t (new_AGEMA_signal_8917), .B1_f (new_AGEMA_signal_8918), .Z0_t (KeyArray_outS20ser[5]), .Z0_f (new_AGEMA_signal_4914), .Z1_t (new_AGEMA_signal_4915), .Z1_f (new_AGEMA_signal_4916) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_5_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS20ser[5]), .B0_f (new_AGEMA_signal_4914), .B1_t (new_AGEMA_signal_4915), .B1_f (new_AGEMA_signal_4916), .Z0_t (KeyArray_S20reg_gff_1_SFF_5_n1), .Z0_f (new_AGEMA_signal_8916), .Z1_t (new_AGEMA_signal_8917), .Z1_f (new_AGEMA_signal_8918) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_5_U1 ( .A0_t (KeyArray_S20reg_gff_1_SFF_5_QD), .A0_f (new_AGEMA_signal_9583), .A1_t (new_AGEMA_signal_9584), .A1_f (new_AGEMA_signal_9585), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S20reg_gff_1_SFF_5_n2), .Z0_f (new_AGEMA_signal_10059), .Z1_t (new_AGEMA_signal_10060), .Z1_f (new_AGEMA_signal_10061) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS20ser[5]), .A0_f (new_AGEMA_signal_7093), .A1_t (new_AGEMA_signal_7094), .A1_f (new_AGEMA_signal_7095), .B0_t (KeyArray_outS30ser[5]), .B0_f (new_AGEMA_signal_5202), .B1_t (new_AGEMA_signal_5203), .B1_f (new_AGEMA_signal_5204), .Z0_t (KeyArray_S20reg_gff_1_SFF_5_MUXInst_X), .Z0_f (new_AGEMA_signal_7926), .Z1_t (new_AGEMA_signal_7927), .Z1_f (new_AGEMA_signal_7928) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S20reg_gff_1_SFF_5_MUXInst_X), .B0_f (new_AGEMA_signal_7926), .B1_t (new_AGEMA_signal_7927), .B1_f (new_AGEMA_signal_7928), .Z0_t (KeyArray_S20reg_gff_1_SFF_5_MUXInst_Y), .Z0_f (new_AGEMA_signal_8919), .Z1_t (new_AGEMA_signal_8920), .Z1_f (new_AGEMA_signal_8921) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S20reg_gff_1_SFF_5_MUXInst_Y), .A0_f (new_AGEMA_signal_8919), .A1_t (new_AGEMA_signal_8920), .A1_f (new_AGEMA_signal_8921), .B0_t (KeyArray_inS20ser[5]), .B0_f (new_AGEMA_signal_7093), .B1_t (new_AGEMA_signal_7094), .B1_f (new_AGEMA_signal_7095), .Z0_t (KeyArray_S20reg_gff_1_SFF_5_QD), .Z0_f (new_AGEMA_signal_9583), .Z1_t (new_AGEMA_signal_9584), .Z1_f (new_AGEMA_signal_9585) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S20reg_gff_1_SFF_6_U3 ( .A0_t (KeyArray_S20reg_gff_1_SFF_6_n2), .A0_f (new_AGEMA_signal_10062), .A1_t (new_AGEMA_signal_10063), .A1_f (new_AGEMA_signal_10064), .B0_t (KeyArray_S20reg_gff_1_SFF_6_n1), .B0_f (new_AGEMA_signal_8922), .B1_t (new_AGEMA_signal_8923), .B1_f (new_AGEMA_signal_8924), .Z0_t (KeyArray_outS20ser[6]), .Z0_f (new_AGEMA_signal_4923), .Z1_t (new_AGEMA_signal_4924), .Z1_f (new_AGEMA_signal_4925) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_6_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS20ser[6]), .B0_f (new_AGEMA_signal_4923), .B1_t (new_AGEMA_signal_4924), .B1_f (new_AGEMA_signal_4925), .Z0_t (KeyArray_S20reg_gff_1_SFF_6_n1), .Z0_f (new_AGEMA_signal_8922), .Z1_t (new_AGEMA_signal_8923), .Z1_f (new_AGEMA_signal_8924) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_6_U1 ( .A0_t (KeyArray_S20reg_gff_1_SFF_6_QD), .A0_f (new_AGEMA_signal_9586), .A1_t (new_AGEMA_signal_9587), .A1_f (new_AGEMA_signal_9588), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S20reg_gff_1_SFF_6_n2), .Z0_f (new_AGEMA_signal_10062), .Z1_t (new_AGEMA_signal_10063), .Z1_f (new_AGEMA_signal_10064) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS20ser[6]), .A0_f (new_AGEMA_signal_7096), .A1_t (new_AGEMA_signal_7097), .A1_f (new_AGEMA_signal_7098), .B0_t (KeyArray_outS30ser[6]), .B0_f (new_AGEMA_signal_5211), .B1_t (new_AGEMA_signal_5212), .B1_f (new_AGEMA_signal_5213), .Z0_t (KeyArray_S20reg_gff_1_SFF_6_MUXInst_X), .Z0_f (new_AGEMA_signal_7929), .Z1_t (new_AGEMA_signal_7930), .Z1_f (new_AGEMA_signal_7931) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S20reg_gff_1_SFF_6_MUXInst_X), .B0_f (new_AGEMA_signal_7929), .B1_t (new_AGEMA_signal_7930), .B1_f (new_AGEMA_signal_7931), .Z0_t (KeyArray_S20reg_gff_1_SFF_6_MUXInst_Y), .Z0_f (new_AGEMA_signal_8925), .Z1_t (new_AGEMA_signal_8926), .Z1_f (new_AGEMA_signal_8927) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S20reg_gff_1_SFF_6_MUXInst_Y), .A0_f (new_AGEMA_signal_8925), .A1_t (new_AGEMA_signal_8926), .A1_f (new_AGEMA_signal_8927), .B0_t (KeyArray_inS20ser[6]), .B0_f (new_AGEMA_signal_7096), .B1_t (new_AGEMA_signal_7097), .B1_f (new_AGEMA_signal_7098), .Z0_t (KeyArray_S20reg_gff_1_SFF_6_QD), .Z0_f (new_AGEMA_signal_9586), .Z1_t (new_AGEMA_signal_9587), .Z1_f (new_AGEMA_signal_9588) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S20reg_gff_1_SFF_7_U3 ( .A0_t (KeyArray_S20reg_gff_1_SFF_7_n2), .A0_f (new_AGEMA_signal_10065), .A1_t (new_AGEMA_signal_10066), .A1_f (new_AGEMA_signal_10067), .B0_t (KeyArray_S20reg_gff_1_SFF_7_n1), .B0_f (new_AGEMA_signal_8928), .B1_t (new_AGEMA_signal_8929), .B1_f (new_AGEMA_signal_8930), .Z0_t (KeyArray_outS20ser[7]), .Z0_f (new_AGEMA_signal_4932), .Z1_t (new_AGEMA_signal_4933), .Z1_f (new_AGEMA_signal_4934) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_7_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS20ser[7]), .B0_f (new_AGEMA_signal_4932), .B1_t (new_AGEMA_signal_4933), .B1_f (new_AGEMA_signal_4934), .Z0_t (KeyArray_S20reg_gff_1_SFF_7_n1), .Z0_f (new_AGEMA_signal_8928), .Z1_t (new_AGEMA_signal_8929), .Z1_f (new_AGEMA_signal_8930) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_7_U1 ( .A0_t (KeyArray_S20reg_gff_1_SFF_7_QD), .A0_f (new_AGEMA_signal_9589), .A1_t (new_AGEMA_signal_9590), .A1_f (new_AGEMA_signal_9591), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S20reg_gff_1_SFF_7_n2), .Z0_f (new_AGEMA_signal_10065), .Z1_t (new_AGEMA_signal_10066), .Z1_f (new_AGEMA_signal_10067) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS20ser[7]), .A0_f (new_AGEMA_signal_7099), .A1_t (new_AGEMA_signal_7100), .A1_f (new_AGEMA_signal_7101), .B0_t (KeyArray_outS30ser[7]), .B0_f (new_AGEMA_signal_5220), .B1_t (new_AGEMA_signal_5221), .B1_f (new_AGEMA_signal_5222), .Z0_t (KeyArray_S20reg_gff_1_SFF_7_MUXInst_X), .Z0_f (new_AGEMA_signal_7932), .Z1_t (new_AGEMA_signal_7933), .Z1_f (new_AGEMA_signal_7934) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S20reg_gff_1_SFF_7_MUXInst_X), .B0_f (new_AGEMA_signal_7932), .B1_t (new_AGEMA_signal_7933), .B1_f (new_AGEMA_signal_7934), .Z0_t (KeyArray_S20reg_gff_1_SFF_7_MUXInst_Y), .Z0_f (new_AGEMA_signal_8931), .Z1_t (new_AGEMA_signal_8932), .Z1_f (new_AGEMA_signal_8933) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S20reg_gff_1_SFF_7_MUXInst_Y), .A0_f (new_AGEMA_signal_8931), .A1_t (new_AGEMA_signal_8932), .A1_f (new_AGEMA_signal_8933), .B0_t (KeyArray_inS20ser[7]), .B0_f (new_AGEMA_signal_7099), .B1_t (new_AGEMA_signal_7100), .B1_f (new_AGEMA_signal_7101), .Z0_t (KeyArray_S20reg_gff_1_SFF_7_QD), .Z0_f (new_AGEMA_signal_9589), .Z1_t (new_AGEMA_signal_9590), .Z1_f (new_AGEMA_signal_9591) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S21reg_gff_1_SFF_0_U3 ( .A0_t (KeyArray_S21reg_gff_1_SFF_0_n2), .A0_f (new_AGEMA_signal_10068), .A1_t (new_AGEMA_signal_10069), .A1_f (new_AGEMA_signal_10070), .B0_t (KeyArray_S21reg_gff_1_SFF_0_n1), .B0_f (new_AGEMA_signal_8934), .B1_t (new_AGEMA_signal_8935), .B1_f (new_AGEMA_signal_8936), .Z0_t (KeyArray_outS21ser[0]), .Z0_f (new_AGEMA_signal_4941), .Z1_t (new_AGEMA_signal_4942), .Z1_f (new_AGEMA_signal_4943) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_0_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS21ser[0]), .B0_f (new_AGEMA_signal_4941), .B1_t (new_AGEMA_signal_4942), .B1_f (new_AGEMA_signal_4943), .Z0_t (KeyArray_S21reg_gff_1_SFF_0_n1), .Z0_f (new_AGEMA_signal_8934), .Z1_t (new_AGEMA_signal_8935), .Z1_f (new_AGEMA_signal_8936) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_0_U1 ( .A0_t (KeyArray_S21reg_gff_1_SFF_0_QD), .A0_f (new_AGEMA_signal_9592), .A1_t (new_AGEMA_signal_9593), .A1_f (new_AGEMA_signal_9594), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S21reg_gff_1_SFF_0_n2), .Z0_f (new_AGEMA_signal_10068), .Z1_t (new_AGEMA_signal_10069), .Z1_f (new_AGEMA_signal_10070) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS21ser[0]), .A0_f (new_AGEMA_signal_7102), .A1_t (new_AGEMA_signal_7103), .A1_f (new_AGEMA_signal_7104), .B0_t (KeyArray_outS31ser[0]), .B0_f (new_AGEMA_signal_5229), .B1_t (new_AGEMA_signal_5230), .B1_f (new_AGEMA_signal_5231), .Z0_t (KeyArray_S21reg_gff_1_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_7935), .Z1_t (new_AGEMA_signal_7936), .Z1_f (new_AGEMA_signal_7937) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S21reg_gff_1_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_7935), .B1_t (new_AGEMA_signal_7936), .B1_f (new_AGEMA_signal_7937), .Z0_t (KeyArray_S21reg_gff_1_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_8937), .Z1_t (new_AGEMA_signal_8938), .Z1_f (new_AGEMA_signal_8939) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S21reg_gff_1_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_8937), .A1_t (new_AGEMA_signal_8938), .A1_f (new_AGEMA_signal_8939), .B0_t (KeyArray_inS21ser[0]), .B0_f (new_AGEMA_signal_7102), .B1_t (new_AGEMA_signal_7103), .B1_f (new_AGEMA_signal_7104), .Z0_t (KeyArray_S21reg_gff_1_SFF_0_QD), .Z0_f (new_AGEMA_signal_9592), .Z1_t (new_AGEMA_signal_9593), .Z1_f (new_AGEMA_signal_9594) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S21reg_gff_1_SFF_1_U3 ( .A0_t (KeyArray_S21reg_gff_1_SFF_1_n2), .A0_f (new_AGEMA_signal_10071), .A1_t (new_AGEMA_signal_10072), .A1_f (new_AGEMA_signal_10073), .B0_t (KeyArray_S21reg_gff_1_SFF_1_n1), .B0_f (new_AGEMA_signal_8940), .B1_t (new_AGEMA_signal_8941), .B1_f (new_AGEMA_signal_8942), .Z0_t (KeyArray_outS21ser[1]), .Z0_f (new_AGEMA_signal_4950), .Z1_t (new_AGEMA_signal_4951), .Z1_f (new_AGEMA_signal_4952) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_1_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS21ser[1]), .B0_f (new_AGEMA_signal_4950), .B1_t (new_AGEMA_signal_4951), .B1_f (new_AGEMA_signal_4952), .Z0_t (KeyArray_S21reg_gff_1_SFF_1_n1), .Z0_f (new_AGEMA_signal_8940), .Z1_t (new_AGEMA_signal_8941), .Z1_f (new_AGEMA_signal_8942) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_1_U1 ( .A0_t (KeyArray_S21reg_gff_1_SFF_1_QD), .A0_f (new_AGEMA_signal_9595), .A1_t (new_AGEMA_signal_9596), .A1_f (new_AGEMA_signal_9597), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S21reg_gff_1_SFF_1_n2), .Z0_f (new_AGEMA_signal_10071), .Z1_t (new_AGEMA_signal_10072), .Z1_f (new_AGEMA_signal_10073) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS21ser[1]), .A0_f (new_AGEMA_signal_7105), .A1_t (new_AGEMA_signal_7106), .A1_f (new_AGEMA_signal_7107), .B0_t (KeyArray_outS31ser[1]), .B0_f (new_AGEMA_signal_5238), .B1_t (new_AGEMA_signal_5239), .B1_f (new_AGEMA_signal_5240), .Z0_t (KeyArray_S21reg_gff_1_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_7938), .Z1_t (new_AGEMA_signal_7939), .Z1_f (new_AGEMA_signal_7940) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S21reg_gff_1_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_7938), .B1_t (new_AGEMA_signal_7939), .B1_f (new_AGEMA_signal_7940), .Z0_t (KeyArray_S21reg_gff_1_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_8943), .Z1_t (new_AGEMA_signal_8944), .Z1_f (new_AGEMA_signal_8945) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S21reg_gff_1_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_8943), .A1_t (new_AGEMA_signal_8944), .A1_f (new_AGEMA_signal_8945), .B0_t (KeyArray_inS21ser[1]), .B0_f (new_AGEMA_signal_7105), .B1_t (new_AGEMA_signal_7106), .B1_f (new_AGEMA_signal_7107), .Z0_t (KeyArray_S21reg_gff_1_SFF_1_QD), .Z0_f (new_AGEMA_signal_9595), .Z1_t (new_AGEMA_signal_9596), .Z1_f (new_AGEMA_signal_9597) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S21reg_gff_1_SFF_2_U3 ( .A0_t (KeyArray_S21reg_gff_1_SFF_2_n2), .A0_f (new_AGEMA_signal_10074), .A1_t (new_AGEMA_signal_10075), .A1_f (new_AGEMA_signal_10076), .B0_t (KeyArray_S21reg_gff_1_SFF_2_n1), .B0_f (new_AGEMA_signal_8946), .B1_t (new_AGEMA_signal_8947), .B1_f (new_AGEMA_signal_8948), .Z0_t (KeyArray_outS21ser[2]), .Z0_f (new_AGEMA_signal_4959), .Z1_t (new_AGEMA_signal_4960), .Z1_f (new_AGEMA_signal_4961) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_2_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS21ser[2]), .B0_f (new_AGEMA_signal_4959), .B1_t (new_AGEMA_signal_4960), .B1_f (new_AGEMA_signal_4961), .Z0_t (KeyArray_S21reg_gff_1_SFF_2_n1), .Z0_f (new_AGEMA_signal_8946), .Z1_t (new_AGEMA_signal_8947), .Z1_f (new_AGEMA_signal_8948) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_2_U1 ( .A0_t (KeyArray_S21reg_gff_1_SFF_2_QD), .A0_f (new_AGEMA_signal_9598), .A1_t (new_AGEMA_signal_9599), .A1_f (new_AGEMA_signal_9600), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S21reg_gff_1_SFF_2_n2), .Z0_f (new_AGEMA_signal_10074), .Z1_t (new_AGEMA_signal_10075), .Z1_f (new_AGEMA_signal_10076) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS21ser[2]), .A0_f (new_AGEMA_signal_7108), .A1_t (new_AGEMA_signal_7109), .A1_f (new_AGEMA_signal_7110), .B0_t (KeyArray_outS31ser[2]), .B0_f (new_AGEMA_signal_5247), .B1_t (new_AGEMA_signal_5248), .B1_f (new_AGEMA_signal_5249), .Z0_t (KeyArray_S21reg_gff_1_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_7941), .Z1_t (new_AGEMA_signal_7942), .Z1_f (new_AGEMA_signal_7943) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S21reg_gff_1_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_7941), .B1_t (new_AGEMA_signal_7942), .B1_f (new_AGEMA_signal_7943), .Z0_t (KeyArray_S21reg_gff_1_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_8949), .Z1_t (new_AGEMA_signal_8950), .Z1_f (new_AGEMA_signal_8951) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S21reg_gff_1_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_8949), .A1_t (new_AGEMA_signal_8950), .A1_f (new_AGEMA_signal_8951), .B0_t (KeyArray_inS21ser[2]), .B0_f (new_AGEMA_signal_7108), .B1_t (new_AGEMA_signal_7109), .B1_f (new_AGEMA_signal_7110), .Z0_t (KeyArray_S21reg_gff_1_SFF_2_QD), .Z0_f (new_AGEMA_signal_9598), .Z1_t (new_AGEMA_signal_9599), .Z1_f (new_AGEMA_signal_9600) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S21reg_gff_1_SFF_3_U3 ( .A0_t (KeyArray_S21reg_gff_1_SFF_3_n2), .A0_f (new_AGEMA_signal_10077), .A1_t (new_AGEMA_signal_10078), .A1_f (new_AGEMA_signal_10079), .B0_t (KeyArray_S21reg_gff_1_SFF_3_n1), .B0_f (new_AGEMA_signal_8952), .B1_t (new_AGEMA_signal_8953), .B1_f (new_AGEMA_signal_8954), .Z0_t (KeyArray_outS21ser[3]), .Z0_f (new_AGEMA_signal_4968), .Z1_t (new_AGEMA_signal_4969), .Z1_f (new_AGEMA_signal_4970) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_3_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS21ser[3]), .B0_f (new_AGEMA_signal_4968), .B1_t (new_AGEMA_signal_4969), .B1_f (new_AGEMA_signal_4970), .Z0_t (KeyArray_S21reg_gff_1_SFF_3_n1), .Z0_f (new_AGEMA_signal_8952), .Z1_t (new_AGEMA_signal_8953), .Z1_f (new_AGEMA_signal_8954) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_3_U1 ( .A0_t (KeyArray_S21reg_gff_1_SFF_3_QD), .A0_f (new_AGEMA_signal_9601), .A1_t (new_AGEMA_signal_9602), .A1_f (new_AGEMA_signal_9603), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S21reg_gff_1_SFF_3_n2), .Z0_f (new_AGEMA_signal_10077), .Z1_t (new_AGEMA_signal_10078), .Z1_f (new_AGEMA_signal_10079) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS21ser[3]), .A0_f (new_AGEMA_signal_7111), .A1_t (new_AGEMA_signal_7112), .A1_f (new_AGEMA_signal_7113), .B0_t (KeyArray_outS31ser[3]), .B0_f (new_AGEMA_signal_5256), .B1_t (new_AGEMA_signal_5257), .B1_f (new_AGEMA_signal_5258), .Z0_t (KeyArray_S21reg_gff_1_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_7944), .Z1_t (new_AGEMA_signal_7945), .Z1_f (new_AGEMA_signal_7946) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S21reg_gff_1_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_7944), .B1_t (new_AGEMA_signal_7945), .B1_f (new_AGEMA_signal_7946), .Z0_t (KeyArray_S21reg_gff_1_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_8955), .Z1_t (new_AGEMA_signal_8956), .Z1_f (new_AGEMA_signal_8957) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S21reg_gff_1_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_8955), .A1_t (new_AGEMA_signal_8956), .A1_f (new_AGEMA_signal_8957), .B0_t (KeyArray_inS21ser[3]), .B0_f (new_AGEMA_signal_7111), .B1_t (new_AGEMA_signal_7112), .B1_f (new_AGEMA_signal_7113), .Z0_t (KeyArray_S21reg_gff_1_SFF_3_QD), .Z0_f (new_AGEMA_signal_9601), .Z1_t (new_AGEMA_signal_9602), .Z1_f (new_AGEMA_signal_9603) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S21reg_gff_1_SFF_4_U3 ( .A0_t (KeyArray_S21reg_gff_1_SFF_4_n2), .A0_f (new_AGEMA_signal_10080), .A1_t (new_AGEMA_signal_10081), .A1_f (new_AGEMA_signal_10082), .B0_t (KeyArray_S21reg_gff_1_SFF_4_n1), .B0_f (new_AGEMA_signal_8958), .B1_t (new_AGEMA_signal_8959), .B1_f (new_AGEMA_signal_8960), .Z0_t (KeyArray_outS21ser[4]), .Z0_f (new_AGEMA_signal_4977), .Z1_t (new_AGEMA_signal_4978), .Z1_f (new_AGEMA_signal_4979) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_4_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS21ser[4]), .B0_f (new_AGEMA_signal_4977), .B1_t (new_AGEMA_signal_4978), .B1_f (new_AGEMA_signal_4979), .Z0_t (KeyArray_S21reg_gff_1_SFF_4_n1), .Z0_f (new_AGEMA_signal_8958), .Z1_t (new_AGEMA_signal_8959), .Z1_f (new_AGEMA_signal_8960) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_4_U1 ( .A0_t (KeyArray_S21reg_gff_1_SFF_4_QD), .A0_f (new_AGEMA_signal_9604), .A1_t (new_AGEMA_signal_9605), .A1_f (new_AGEMA_signal_9606), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S21reg_gff_1_SFF_4_n2), .Z0_f (new_AGEMA_signal_10080), .Z1_t (new_AGEMA_signal_10081), .Z1_f (new_AGEMA_signal_10082) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS21ser[4]), .A0_f (new_AGEMA_signal_7114), .A1_t (new_AGEMA_signal_7115), .A1_f (new_AGEMA_signal_7116), .B0_t (KeyArray_outS31ser[4]), .B0_f (new_AGEMA_signal_5265), .B1_t (new_AGEMA_signal_5266), .B1_f (new_AGEMA_signal_5267), .Z0_t (KeyArray_S21reg_gff_1_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_7947), .Z1_t (new_AGEMA_signal_7948), .Z1_f (new_AGEMA_signal_7949) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S21reg_gff_1_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_7947), .B1_t (new_AGEMA_signal_7948), .B1_f (new_AGEMA_signal_7949), .Z0_t (KeyArray_S21reg_gff_1_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_8961), .Z1_t (new_AGEMA_signal_8962), .Z1_f (new_AGEMA_signal_8963) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S21reg_gff_1_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_8961), .A1_t (new_AGEMA_signal_8962), .A1_f (new_AGEMA_signal_8963), .B0_t (KeyArray_inS21ser[4]), .B0_f (new_AGEMA_signal_7114), .B1_t (new_AGEMA_signal_7115), .B1_f (new_AGEMA_signal_7116), .Z0_t (KeyArray_S21reg_gff_1_SFF_4_QD), .Z0_f (new_AGEMA_signal_9604), .Z1_t (new_AGEMA_signal_9605), .Z1_f (new_AGEMA_signal_9606) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S21reg_gff_1_SFF_5_U3 ( .A0_t (KeyArray_S21reg_gff_1_SFF_5_n2), .A0_f (new_AGEMA_signal_10083), .A1_t (new_AGEMA_signal_10084), .A1_f (new_AGEMA_signal_10085), .B0_t (KeyArray_S21reg_gff_1_SFF_5_n1), .B0_f (new_AGEMA_signal_8964), .B1_t (new_AGEMA_signal_8965), .B1_f (new_AGEMA_signal_8966), .Z0_t (KeyArray_outS21ser[5]), .Z0_f (new_AGEMA_signal_4986), .Z1_t (new_AGEMA_signal_4987), .Z1_f (new_AGEMA_signal_4988) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_5_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS21ser[5]), .B0_f (new_AGEMA_signal_4986), .B1_t (new_AGEMA_signal_4987), .B1_f (new_AGEMA_signal_4988), .Z0_t (KeyArray_S21reg_gff_1_SFF_5_n1), .Z0_f (new_AGEMA_signal_8964), .Z1_t (new_AGEMA_signal_8965), .Z1_f (new_AGEMA_signal_8966) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_5_U1 ( .A0_t (KeyArray_S21reg_gff_1_SFF_5_QD), .A0_f (new_AGEMA_signal_9607), .A1_t (new_AGEMA_signal_9608), .A1_f (new_AGEMA_signal_9609), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S21reg_gff_1_SFF_5_n2), .Z0_f (new_AGEMA_signal_10083), .Z1_t (new_AGEMA_signal_10084), .Z1_f (new_AGEMA_signal_10085) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS21ser[5]), .A0_f (new_AGEMA_signal_7117), .A1_t (new_AGEMA_signal_7118), .A1_f (new_AGEMA_signal_7119), .B0_t (KeyArray_outS31ser[5]), .B0_f (new_AGEMA_signal_5274), .B1_t (new_AGEMA_signal_5275), .B1_f (new_AGEMA_signal_5276), .Z0_t (KeyArray_S21reg_gff_1_SFF_5_MUXInst_X), .Z0_f (new_AGEMA_signal_7950), .Z1_t (new_AGEMA_signal_7951), .Z1_f (new_AGEMA_signal_7952) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S21reg_gff_1_SFF_5_MUXInst_X), .B0_f (new_AGEMA_signal_7950), .B1_t (new_AGEMA_signal_7951), .B1_f (new_AGEMA_signal_7952), .Z0_t (KeyArray_S21reg_gff_1_SFF_5_MUXInst_Y), .Z0_f (new_AGEMA_signal_8967), .Z1_t (new_AGEMA_signal_8968), .Z1_f (new_AGEMA_signal_8969) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S21reg_gff_1_SFF_5_MUXInst_Y), .A0_f (new_AGEMA_signal_8967), .A1_t (new_AGEMA_signal_8968), .A1_f (new_AGEMA_signal_8969), .B0_t (KeyArray_inS21ser[5]), .B0_f (new_AGEMA_signal_7117), .B1_t (new_AGEMA_signal_7118), .B1_f (new_AGEMA_signal_7119), .Z0_t (KeyArray_S21reg_gff_1_SFF_5_QD), .Z0_f (new_AGEMA_signal_9607), .Z1_t (new_AGEMA_signal_9608), .Z1_f (new_AGEMA_signal_9609) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S21reg_gff_1_SFF_6_U3 ( .A0_t (KeyArray_S21reg_gff_1_SFF_6_n2), .A0_f (new_AGEMA_signal_10086), .A1_t (new_AGEMA_signal_10087), .A1_f (new_AGEMA_signal_10088), .B0_t (KeyArray_S21reg_gff_1_SFF_6_n1), .B0_f (new_AGEMA_signal_8970), .B1_t (new_AGEMA_signal_8971), .B1_f (new_AGEMA_signal_8972), .Z0_t (KeyArray_outS21ser[6]), .Z0_f (new_AGEMA_signal_4995), .Z1_t (new_AGEMA_signal_4996), .Z1_f (new_AGEMA_signal_4997) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_6_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS21ser[6]), .B0_f (new_AGEMA_signal_4995), .B1_t (new_AGEMA_signal_4996), .B1_f (new_AGEMA_signal_4997), .Z0_t (KeyArray_S21reg_gff_1_SFF_6_n1), .Z0_f (new_AGEMA_signal_8970), .Z1_t (new_AGEMA_signal_8971), .Z1_f (new_AGEMA_signal_8972) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_6_U1 ( .A0_t (KeyArray_S21reg_gff_1_SFF_6_QD), .A0_f (new_AGEMA_signal_9610), .A1_t (new_AGEMA_signal_9611), .A1_f (new_AGEMA_signal_9612), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S21reg_gff_1_SFF_6_n2), .Z0_f (new_AGEMA_signal_10086), .Z1_t (new_AGEMA_signal_10087), .Z1_f (new_AGEMA_signal_10088) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS21ser[6]), .A0_f (new_AGEMA_signal_7120), .A1_t (new_AGEMA_signal_7121), .A1_f (new_AGEMA_signal_7122), .B0_t (KeyArray_outS31ser[6]), .B0_f (new_AGEMA_signal_5283), .B1_t (new_AGEMA_signal_5284), .B1_f (new_AGEMA_signal_5285), .Z0_t (KeyArray_S21reg_gff_1_SFF_6_MUXInst_X), .Z0_f (new_AGEMA_signal_7953), .Z1_t (new_AGEMA_signal_7954), .Z1_f (new_AGEMA_signal_7955) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S21reg_gff_1_SFF_6_MUXInst_X), .B0_f (new_AGEMA_signal_7953), .B1_t (new_AGEMA_signal_7954), .B1_f (new_AGEMA_signal_7955), .Z0_t (KeyArray_S21reg_gff_1_SFF_6_MUXInst_Y), .Z0_f (new_AGEMA_signal_8973), .Z1_t (new_AGEMA_signal_8974), .Z1_f (new_AGEMA_signal_8975) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S21reg_gff_1_SFF_6_MUXInst_Y), .A0_f (new_AGEMA_signal_8973), .A1_t (new_AGEMA_signal_8974), .A1_f (new_AGEMA_signal_8975), .B0_t (KeyArray_inS21ser[6]), .B0_f (new_AGEMA_signal_7120), .B1_t (new_AGEMA_signal_7121), .B1_f (new_AGEMA_signal_7122), .Z0_t (KeyArray_S21reg_gff_1_SFF_6_QD), .Z0_f (new_AGEMA_signal_9610), .Z1_t (new_AGEMA_signal_9611), .Z1_f (new_AGEMA_signal_9612) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S21reg_gff_1_SFF_7_U3 ( .A0_t (KeyArray_S21reg_gff_1_SFF_7_n2), .A0_f (new_AGEMA_signal_10089), .A1_t (new_AGEMA_signal_10090), .A1_f (new_AGEMA_signal_10091), .B0_t (KeyArray_S21reg_gff_1_SFF_7_n1), .B0_f (new_AGEMA_signal_8976), .B1_t (new_AGEMA_signal_8977), .B1_f (new_AGEMA_signal_8978), .Z0_t (KeyArray_outS21ser[7]), .Z0_f (new_AGEMA_signal_5004), .Z1_t (new_AGEMA_signal_5005), .Z1_f (new_AGEMA_signal_5006) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_7_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS21ser[7]), .B0_f (new_AGEMA_signal_5004), .B1_t (new_AGEMA_signal_5005), .B1_f (new_AGEMA_signal_5006), .Z0_t (KeyArray_S21reg_gff_1_SFF_7_n1), .Z0_f (new_AGEMA_signal_8976), .Z1_t (new_AGEMA_signal_8977), .Z1_f (new_AGEMA_signal_8978) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_7_U1 ( .A0_t (KeyArray_S21reg_gff_1_SFF_7_QD), .A0_f (new_AGEMA_signal_9613), .A1_t (new_AGEMA_signal_9614), .A1_f (new_AGEMA_signal_9615), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S21reg_gff_1_SFF_7_n2), .Z0_f (new_AGEMA_signal_10089), .Z1_t (new_AGEMA_signal_10090), .Z1_f (new_AGEMA_signal_10091) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS21ser[7]), .A0_f (new_AGEMA_signal_7123), .A1_t (new_AGEMA_signal_7124), .A1_f (new_AGEMA_signal_7125), .B0_t (KeyArray_outS31ser[7]), .B0_f (new_AGEMA_signal_5292), .B1_t (new_AGEMA_signal_5293), .B1_f (new_AGEMA_signal_5294), .Z0_t (KeyArray_S21reg_gff_1_SFF_7_MUXInst_X), .Z0_f (new_AGEMA_signal_7956), .Z1_t (new_AGEMA_signal_7957), .Z1_f (new_AGEMA_signal_7958) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S21reg_gff_1_SFF_7_MUXInst_X), .B0_f (new_AGEMA_signal_7956), .B1_t (new_AGEMA_signal_7957), .B1_f (new_AGEMA_signal_7958), .Z0_t (KeyArray_S21reg_gff_1_SFF_7_MUXInst_Y), .Z0_f (new_AGEMA_signal_8979), .Z1_t (new_AGEMA_signal_8980), .Z1_f (new_AGEMA_signal_8981) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S21reg_gff_1_SFF_7_MUXInst_Y), .A0_f (new_AGEMA_signal_8979), .A1_t (new_AGEMA_signal_8980), .A1_f (new_AGEMA_signal_8981), .B0_t (KeyArray_inS21ser[7]), .B0_f (new_AGEMA_signal_7123), .B1_t (new_AGEMA_signal_7124), .B1_f (new_AGEMA_signal_7125), .Z0_t (KeyArray_S21reg_gff_1_SFF_7_QD), .Z0_f (new_AGEMA_signal_9613), .Z1_t (new_AGEMA_signal_9614), .Z1_f (new_AGEMA_signal_9615) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S22reg_gff_1_SFF_0_U3 ( .A0_t (KeyArray_S22reg_gff_1_SFF_0_n2), .A0_f (new_AGEMA_signal_10092), .A1_t (new_AGEMA_signal_10093), .A1_f (new_AGEMA_signal_10094), .B0_t (KeyArray_S22reg_gff_1_SFF_0_n1), .B0_f (new_AGEMA_signal_8982), .B1_t (new_AGEMA_signal_8983), .B1_f (new_AGEMA_signal_8984), .Z0_t (KeyArray_outS22ser[0]), .Z0_f (new_AGEMA_signal_5013), .Z1_t (new_AGEMA_signal_5014), .Z1_f (new_AGEMA_signal_5015) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_0_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS22ser[0]), .B0_f (new_AGEMA_signal_5013), .B1_t (new_AGEMA_signal_5014), .B1_f (new_AGEMA_signal_5015), .Z0_t (KeyArray_S22reg_gff_1_SFF_0_n1), .Z0_f (new_AGEMA_signal_8982), .Z1_t (new_AGEMA_signal_8983), .Z1_f (new_AGEMA_signal_8984) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_0_U1 ( .A0_t (KeyArray_S22reg_gff_1_SFF_0_QD), .A0_f (new_AGEMA_signal_9616), .A1_t (new_AGEMA_signal_9617), .A1_f (new_AGEMA_signal_9618), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S22reg_gff_1_SFF_0_n2), .Z0_f (new_AGEMA_signal_10092), .Z1_t (new_AGEMA_signal_10093), .Z1_f (new_AGEMA_signal_10094) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS22ser[0]), .A0_f (new_AGEMA_signal_7126), .A1_t (new_AGEMA_signal_7127), .A1_f (new_AGEMA_signal_7128), .B0_t (KeyArray_outS32ser[0]), .B0_f (new_AGEMA_signal_5301), .B1_t (new_AGEMA_signal_5302), .B1_f (new_AGEMA_signal_5303), .Z0_t (KeyArray_S22reg_gff_1_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_7959), .Z1_t (new_AGEMA_signal_7960), .Z1_f (new_AGEMA_signal_7961) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S22reg_gff_1_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_7959), .B1_t (new_AGEMA_signal_7960), .B1_f (new_AGEMA_signal_7961), .Z0_t (KeyArray_S22reg_gff_1_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_8985), .Z1_t (new_AGEMA_signal_8986), .Z1_f (new_AGEMA_signal_8987) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S22reg_gff_1_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_8985), .A1_t (new_AGEMA_signal_8986), .A1_f (new_AGEMA_signal_8987), .B0_t (KeyArray_inS22ser[0]), .B0_f (new_AGEMA_signal_7126), .B1_t (new_AGEMA_signal_7127), .B1_f (new_AGEMA_signal_7128), .Z0_t (KeyArray_S22reg_gff_1_SFF_0_QD), .Z0_f (new_AGEMA_signal_9616), .Z1_t (new_AGEMA_signal_9617), .Z1_f (new_AGEMA_signal_9618) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S22reg_gff_1_SFF_1_U3 ( .A0_t (KeyArray_S22reg_gff_1_SFF_1_n2), .A0_f (new_AGEMA_signal_10095), .A1_t (new_AGEMA_signal_10096), .A1_f (new_AGEMA_signal_10097), .B0_t (KeyArray_S22reg_gff_1_SFF_1_n1), .B0_f (new_AGEMA_signal_8988), .B1_t (new_AGEMA_signal_8989), .B1_f (new_AGEMA_signal_8990), .Z0_t (KeyArray_outS22ser[1]), .Z0_f (new_AGEMA_signal_5022), .Z1_t (new_AGEMA_signal_5023), .Z1_f (new_AGEMA_signal_5024) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_1_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS22ser[1]), .B0_f (new_AGEMA_signal_5022), .B1_t (new_AGEMA_signal_5023), .B1_f (new_AGEMA_signal_5024), .Z0_t (KeyArray_S22reg_gff_1_SFF_1_n1), .Z0_f (new_AGEMA_signal_8988), .Z1_t (new_AGEMA_signal_8989), .Z1_f (new_AGEMA_signal_8990) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_1_U1 ( .A0_t (KeyArray_S22reg_gff_1_SFF_1_QD), .A0_f (new_AGEMA_signal_9619), .A1_t (new_AGEMA_signal_9620), .A1_f (new_AGEMA_signal_9621), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S22reg_gff_1_SFF_1_n2), .Z0_f (new_AGEMA_signal_10095), .Z1_t (new_AGEMA_signal_10096), .Z1_f (new_AGEMA_signal_10097) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS22ser[1]), .A0_f (new_AGEMA_signal_7129), .A1_t (new_AGEMA_signal_7130), .A1_f (new_AGEMA_signal_7131), .B0_t (KeyArray_outS32ser[1]), .B0_f (new_AGEMA_signal_5310), .B1_t (new_AGEMA_signal_5311), .B1_f (new_AGEMA_signal_5312), .Z0_t (KeyArray_S22reg_gff_1_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_7962), .Z1_t (new_AGEMA_signal_7963), .Z1_f (new_AGEMA_signal_7964) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S22reg_gff_1_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_7962), .B1_t (new_AGEMA_signal_7963), .B1_f (new_AGEMA_signal_7964), .Z0_t (KeyArray_S22reg_gff_1_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_8991), .Z1_t (new_AGEMA_signal_8992), .Z1_f (new_AGEMA_signal_8993) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S22reg_gff_1_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_8991), .A1_t (new_AGEMA_signal_8992), .A1_f (new_AGEMA_signal_8993), .B0_t (KeyArray_inS22ser[1]), .B0_f (new_AGEMA_signal_7129), .B1_t (new_AGEMA_signal_7130), .B1_f (new_AGEMA_signal_7131), .Z0_t (KeyArray_S22reg_gff_1_SFF_1_QD), .Z0_f (new_AGEMA_signal_9619), .Z1_t (new_AGEMA_signal_9620), .Z1_f (new_AGEMA_signal_9621) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S22reg_gff_1_SFF_2_U3 ( .A0_t (KeyArray_S22reg_gff_1_SFF_2_n2), .A0_f (new_AGEMA_signal_10098), .A1_t (new_AGEMA_signal_10099), .A1_f (new_AGEMA_signal_10100), .B0_t (KeyArray_S22reg_gff_1_SFF_2_n1), .B0_f (new_AGEMA_signal_8994), .B1_t (new_AGEMA_signal_8995), .B1_f (new_AGEMA_signal_8996), .Z0_t (KeyArray_outS22ser[2]), .Z0_f (new_AGEMA_signal_5031), .Z1_t (new_AGEMA_signal_5032), .Z1_f (new_AGEMA_signal_5033) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_2_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS22ser[2]), .B0_f (new_AGEMA_signal_5031), .B1_t (new_AGEMA_signal_5032), .B1_f (new_AGEMA_signal_5033), .Z0_t (KeyArray_S22reg_gff_1_SFF_2_n1), .Z0_f (new_AGEMA_signal_8994), .Z1_t (new_AGEMA_signal_8995), .Z1_f (new_AGEMA_signal_8996) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_2_U1 ( .A0_t (KeyArray_S22reg_gff_1_SFF_2_QD), .A0_f (new_AGEMA_signal_9622), .A1_t (new_AGEMA_signal_9623), .A1_f (new_AGEMA_signal_9624), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S22reg_gff_1_SFF_2_n2), .Z0_f (new_AGEMA_signal_10098), .Z1_t (new_AGEMA_signal_10099), .Z1_f (new_AGEMA_signal_10100) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS22ser[2]), .A0_f (new_AGEMA_signal_7132), .A1_t (new_AGEMA_signal_7133), .A1_f (new_AGEMA_signal_7134), .B0_t (KeyArray_outS32ser[2]), .B0_f (new_AGEMA_signal_5319), .B1_t (new_AGEMA_signal_5320), .B1_f (new_AGEMA_signal_5321), .Z0_t (KeyArray_S22reg_gff_1_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_7965), .Z1_t (new_AGEMA_signal_7966), .Z1_f (new_AGEMA_signal_7967) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S22reg_gff_1_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_7965), .B1_t (new_AGEMA_signal_7966), .B1_f (new_AGEMA_signal_7967), .Z0_t (KeyArray_S22reg_gff_1_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_8997), .Z1_t (new_AGEMA_signal_8998), .Z1_f (new_AGEMA_signal_8999) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S22reg_gff_1_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_8997), .A1_t (new_AGEMA_signal_8998), .A1_f (new_AGEMA_signal_8999), .B0_t (KeyArray_inS22ser[2]), .B0_f (new_AGEMA_signal_7132), .B1_t (new_AGEMA_signal_7133), .B1_f (new_AGEMA_signal_7134), .Z0_t (KeyArray_S22reg_gff_1_SFF_2_QD), .Z0_f (new_AGEMA_signal_9622), .Z1_t (new_AGEMA_signal_9623), .Z1_f (new_AGEMA_signal_9624) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S22reg_gff_1_SFF_3_U3 ( .A0_t (KeyArray_S22reg_gff_1_SFF_3_n2), .A0_f (new_AGEMA_signal_10101), .A1_t (new_AGEMA_signal_10102), .A1_f (new_AGEMA_signal_10103), .B0_t (KeyArray_S22reg_gff_1_SFF_3_n1), .B0_f (new_AGEMA_signal_9000), .B1_t (new_AGEMA_signal_9001), .B1_f (new_AGEMA_signal_9002), .Z0_t (KeyArray_outS22ser[3]), .Z0_f (new_AGEMA_signal_5040), .Z1_t (new_AGEMA_signal_5041), .Z1_f (new_AGEMA_signal_5042) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_3_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS22ser[3]), .B0_f (new_AGEMA_signal_5040), .B1_t (new_AGEMA_signal_5041), .B1_f (new_AGEMA_signal_5042), .Z0_t (KeyArray_S22reg_gff_1_SFF_3_n1), .Z0_f (new_AGEMA_signal_9000), .Z1_t (new_AGEMA_signal_9001), .Z1_f (new_AGEMA_signal_9002) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_3_U1 ( .A0_t (KeyArray_S22reg_gff_1_SFF_3_QD), .A0_f (new_AGEMA_signal_9625), .A1_t (new_AGEMA_signal_9626), .A1_f (new_AGEMA_signal_9627), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S22reg_gff_1_SFF_3_n2), .Z0_f (new_AGEMA_signal_10101), .Z1_t (new_AGEMA_signal_10102), .Z1_f (new_AGEMA_signal_10103) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS22ser[3]), .A0_f (new_AGEMA_signal_7135), .A1_t (new_AGEMA_signal_7136), .A1_f (new_AGEMA_signal_7137), .B0_t (KeyArray_outS32ser[3]), .B0_f (new_AGEMA_signal_5328), .B1_t (new_AGEMA_signal_5329), .B1_f (new_AGEMA_signal_5330), .Z0_t (KeyArray_S22reg_gff_1_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_7968), .Z1_t (new_AGEMA_signal_7969), .Z1_f (new_AGEMA_signal_7970) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S22reg_gff_1_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_7968), .B1_t (new_AGEMA_signal_7969), .B1_f (new_AGEMA_signal_7970), .Z0_t (KeyArray_S22reg_gff_1_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_9003), .Z1_t (new_AGEMA_signal_9004), .Z1_f (new_AGEMA_signal_9005) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S22reg_gff_1_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_9003), .A1_t (new_AGEMA_signal_9004), .A1_f (new_AGEMA_signal_9005), .B0_t (KeyArray_inS22ser[3]), .B0_f (new_AGEMA_signal_7135), .B1_t (new_AGEMA_signal_7136), .B1_f (new_AGEMA_signal_7137), .Z0_t (KeyArray_S22reg_gff_1_SFF_3_QD), .Z0_f (new_AGEMA_signal_9625), .Z1_t (new_AGEMA_signal_9626), .Z1_f (new_AGEMA_signal_9627) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S22reg_gff_1_SFF_4_U3 ( .A0_t (KeyArray_S22reg_gff_1_SFF_4_n2), .A0_f (new_AGEMA_signal_10104), .A1_t (new_AGEMA_signal_10105), .A1_f (new_AGEMA_signal_10106), .B0_t (KeyArray_S22reg_gff_1_SFF_4_n1), .B0_f (new_AGEMA_signal_9006), .B1_t (new_AGEMA_signal_9007), .B1_f (new_AGEMA_signal_9008), .Z0_t (KeyArray_outS22ser[4]), .Z0_f (new_AGEMA_signal_5049), .Z1_t (new_AGEMA_signal_5050), .Z1_f (new_AGEMA_signal_5051) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_4_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS22ser[4]), .B0_f (new_AGEMA_signal_5049), .B1_t (new_AGEMA_signal_5050), .B1_f (new_AGEMA_signal_5051), .Z0_t (KeyArray_S22reg_gff_1_SFF_4_n1), .Z0_f (new_AGEMA_signal_9006), .Z1_t (new_AGEMA_signal_9007), .Z1_f (new_AGEMA_signal_9008) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_4_U1 ( .A0_t (KeyArray_S22reg_gff_1_SFF_4_QD), .A0_f (new_AGEMA_signal_9628), .A1_t (new_AGEMA_signal_9629), .A1_f (new_AGEMA_signal_9630), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S22reg_gff_1_SFF_4_n2), .Z0_f (new_AGEMA_signal_10104), .Z1_t (new_AGEMA_signal_10105), .Z1_f (new_AGEMA_signal_10106) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS22ser[4]), .A0_f (new_AGEMA_signal_7138), .A1_t (new_AGEMA_signal_7139), .A1_f (new_AGEMA_signal_7140), .B0_t (KeyArray_outS32ser[4]), .B0_f (new_AGEMA_signal_5337), .B1_t (new_AGEMA_signal_5338), .B1_f (new_AGEMA_signal_5339), .Z0_t (KeyArray_S22reg_gff_1_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_7971), .Z1_t (new_AGEMA_signal_7972), .Z1_f (new_AGEMA_signal_7973) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S22reg_gff_1_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_7971), .B1_t (new_AGEMA_signal_7972), .B1_f (new_AGEMA_signal_7973), .Z0_t (KeyArray_S22reg_gff_1_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_9009), .Z1_t (new_AGEMA_signal_9010), .Z1_f (new_AGEMA_signal_9011) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S22reg_gff_1_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_9009), .A1_t (new_AGEMA_signal_9010), .A1_f (new_AGEMA_signal_9011), .B0_t (KeyArray_inS22ser[4]), .B0_f (new_AGEMA_signal_7138), .B1_t (new_AGEMA_signal_7139), .B1_f (new_AGEMA_signal_7140), .Z0_t (KeyArray_S22reg_gff_1_SFF_4_QD), .Z0_f (new_AGEMA_signal_9628), .Z1_t (new_AGEMA_signal_9629), .Z1_f (new_AGEMA_signal_9630) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S22reg_gff_1_SFF_5_U3 ( .A0_t (KeyArray_S22reg_gff_1_SFF_5_n2), .A0_f (new_AGEMA_signal_10107), .A1_t (new_AGEMA_signal_10108), .A1_f (new_AGEMA_signal_10109), .B0_t (KeyArray_S22reg_gff_1_SFF_5_n1), .B0_f (new_AGEMA_signal_9012), .B1_t (new_AGEMA_signal_9013), .B1_f (new_AGEMA_signal_9014), .Z0_t (KeyArray_outS22ser[5]), .Z0_f (new_AGEMA_signal_5058), .Z1_t (new_AGEMA_signal_5059), .Z1_f (new_AGEMA_signal_5060) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_5_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS22ser[5]), .B0_f (new_AGEMA_signal_5058), .B1_t (new_AGEMA_signal_5059), .B1_f (new_AGEMA_signal_5060), .Z0_t (KeyArray_S22reg_gff_1_SFF_5_n1), .Z0_f (new_AGEMA_signal_9012), .Z1_t (new_AGEMA_signal_9013), .Z1_f (new_AGEMA_signal_9014) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_5_U1 ( .A0_t (KeyArray_S22reg_gff_1_SFF_5_QD), .A0_f (new_AGEMA_signal_9631), .A1_t (new_AGEMA_signal_9632), .A1_f (new_AGEMA_signal_9633), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S22reg_gff_1_SFF_5_n2), .Z0_f (new_AGEMA_signal_10107), .Z1_t (new_AGEMA_signal_10108), .Z1_f (new_AGEMA_signal_10109) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS22ser[5]), .A0_f (new_AGEMA_signal_7141), .A1_t (new_AGEMA_signal_7142), .A1_f (new_AGEMA_signal_7143), .B0_t (KeyArray_outS32ser[5]), .B0_f (new_AGEMA_signal_5346), .B1_t (new_AGEMA_signal_5347), .B1_f (new_AGEMA_signal_5348), .Z0_t (KeyArray_S22reg_gff_1_SFF_5_MUXInst_X), .Z0_f (new_AGEMA_signal_7974), .Z1_t (new_AGEMA_signal_7975), .Z1_f (new_AGEMA_signal_7976) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S22reg_gff_1_SFF_5_MUXInst_X), .B0_f (new_AGEMA_signal_7974), .B1_t (new_AGEMA_signal_7975), .B1_f (new_AGEMA_signal_7976), .Z0_t (KeyArray_S22reg_gff_1_SFF_5_MUXInst_Y), .Z0_f (new_AGEMA_signal_9015), .Z1_t (new_AGEMA_signal_9016), .Z1_f (new_AGEMA_signal_9017) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S22reg_gff_1_SFF_5_MUXInst_Y), .A0_f (new_AGEMA_signal_9015), .A1_t (new_AGEMA_signal_9016), .A1_f (new_AGEMA_signal_9017), .B0_t (KeyArray_inS22ser[5]), .B0_f (new_AGEMA_signal_7141), .B1_t (new_AGEMA_signal_7142), .B1_f (new_AGEMA_signal_7143), .Z0_t (KeyArray_S22reg_gff_1_SFF_5_QD), .Z0_f (new_AGEMA_signal_9631), .Z1_t (new_AGEMA_signal_9632), .Z1_f (new_AGEMA_signal_9633) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S22reg_gff_1_SFF_6_U3 ( .A0_t (KeyArray_S22reg_gff_1_SFF_6_n2), .A0_f (new_AGEMA_signal_10110), .A1_t (new_AGEMA_signal_10111), .A1_f (new_AGEMA_signal_10112), .B0_t (KeyArray_S22reg_gff_1_SFF_6_n1), .B0_f (new_AGEMA_signal_9018), .B1_t (new_AGEMA_signal_9019), .B1_f (new_AGEMA_signal_9020), .Z0_t (KeyArray_outS22ser[6]), .Z0_f (new_AGEMA_signal_5067), .Z1_t (new_AGEMA_signal_5068), .Z1_f (new_AGEMA_signal_5069) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_6_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS22ser[6]), .B0_f (new_AGEMA_signal_5067), .B1_t (new_AGEMA_signal_5068), .B1_f (new_AGEMA_signal_5069), .Z0_t (KeyArray_S22reg_gff_1_SFF_6_n1), .Z0_f (new_AGEMA_signal_9018), .Z1_t (new_AGEMA_signal_9019), .Z1_f (new_AGEMA_signal_9020) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_6_U1 ( .A0_t (KeyArray_S22reg_gff_1_SFF_6_QD), .A0_f (new_AGEMA_signal_9634), .A1_t (new_AGEMA_signal_9635), .A1_f (new_AGEMA_signal_9636), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S22reg_gff_1_SFF_6_n2), .Z0_f (new_AGEMA_signal_10110), .Z1_t (new_AGEMA_signal_10111), .Z1_f (new_AGEMA_signal_10112) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS22ser[6]), .A0_f (new_AGEMA_signal_7144), .A1_t (new_AGEMA_signal_7145), .A1_f (new_AGEMA_signal_7146), .B0_t (KeyArray_outS32ser[6]), .B0_f (new_AGEMA_signal_5355), .B1_t (new_AGEMA_signal_5356), .B1_f (new_AGEMA_signal_5357), .Z0_t (KeyArray_S22reg_gff_1_SFF_6_MUXInst_X), .Z0_f (new_AGEMA_signal_7977), .Z1_t (new_AGEMA_signal_7978), .Z1_f (new_AGEMA_signal_7979) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S22reg_gff_1_SFF_6_MUXInst_X), .B0_f (new_AGEMA_signal_7977), .B1_t (new_AGEMA_signal_7978), .B1_f (new_AGEMA_signal_7979), .Z0_t (KeyArray_S22reg_gff_1_SFF_6_MUXInst_Y), .Z0_f (new_AGEMA_signal_9021), .Z1_t (new_AGEMA_signal_9022), .Z1_f (new_AGEMA_signal_9023) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S22reg_gff_1_SFF_6_MUXInst_Y), .A0_f (new_AGEMA_signal_9021), .A1_t (new_AGEMA_signal_9022), .A1_f (new_AGEMA_signal_9023), .B0_t (KeyArray_inS22ser[6]), .B0_f (new_AGEMA_signal_7144), .B1_t (new_AGEMA_signal_7145), .B1_f (new_AGEMA_signal_7146), .Z0_t (KeyArray_S22reg_gff_1_SFF_6_QD), .Z0_f (new_AGEMA_signal_9634), .Z1_t (new_AGEMA_signal_9635), .Z1_f (new_AGEMA_signal_9636) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S22reg_gff_1_SFF_7_U3 ( .A0_t (KeyArray_S22reg_gff_1_SFF_7_n2), .A0_f (new_AGEMA_signal_10113), .A1_t (new_AGEMA_signal_10114), .A1_f (new_AGEMA_signal_10115), .B0_t (KeyArray_S22reg_gff_1_SFF_7_n1), .B0_f (new_AGEMA_signal_9024), .B1_t (new_AGEMA_signal_9025), .B1_f (new_AGEMA_signal_9026), .Z0_t (KeyArray_outS22ser[7]), .Z0_f (new_AGEMA_signal_5076), .Z1_t (new_AGEMA_signal_5077), .Z1_f (new_AGEMA_signal_5078) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_7_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS22ser[7]), .B0_f (new_AGEMA_signal_5076), .B1_t (new_AGEMA_signal_5077), .B1_f (new_AGEMA_signal_5078), .Z0_t (KeyArray_S22reg_gff_1_SFF_7_n1), .Z0_f (new_AGEMA_signal_9024), .Z1_t (new_AGEMA_signal_9025), .Z1_f (new_AGEMA_signal_9026) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_7_U1 ( .A0_t (KeyArray_S22reg_gff_1_SFF_7_QD), .A0_f (new_AGEMA_signal_9637), .A1_t (new_AGEMA_signal_9638), .A1_f (new_AGEMA_signal_9639), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S22reg_gff_1_SFF_7_n2), .Z0_f (new_AGEMA_signal_10113), .Z1_t (new_AGEMA_signal_10114), .Z1_f (new_AGEMA_signal_10115) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS22ser[7]), .A0_f (new_AGEMA_signal_7147), .A1_t (new_AGEMA_signal_7148), .A1_f (new_AGEMA_signal_7149), .B0_t (KeyArray_outS32ser[7]), .B0_f (new_AGEMA_signal_5364), .B1_t (new_AGEMA_signal_5365), .B1_f (new_AGEMA_signal_5366), .Z0_t (KeyArray_S22reg_gff_1_SFF_7_MUXInst_X), .Z0_f (new_AGEMA_signal_7980), .Z1_t (new_AGEMA_signal_7981), .Z1_f (new_AGEMA_signal_7982) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S22reg_gff_1_SFF_7_MUXInst_X), .B0_f (new_AGEMA_signal_7980), .B1_t (new_AGEMA_signal_7981), .B1_f (new_AGEMA_signal_7982), .Z0_t (KeyArray_S22reg_gff_1_SFF_7_MUXInst_Y), .Z0_f (new_AGEMA_signal_9027), .Z1_t (new_AGEMA_signal_9028), .Z1_f (new_AGEMA_signal_9029) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S22reg_gff_1_SFF_7_MUXInst_Y), .A0_f (new_AGEMA_signal_9027), .A1_t (new_AGEMA_signal_9028), .A1_f (new_AGEMA_signal_9029), .B0_t (KeyArray_inS22ser[7]), .B0_f (new_AGEMA_signal_7147), .B1_t (new_AGEMA_signal_7148), .B1_f (new_AGEMA_signal_7149), .Z0_t (KeyArray_S22reg_gff_1_SFF_7_QD), .Z0_f (new_AGEMA_signal_9637), .Z1_t (new_AGEMA_signal_9638), .Z1_f (new_AGEMA_signal_9639) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S23reg_gff_1_SFF_0_U3 ( .A0_t (KeyArray_S23reg_gff_1_SFF_0_n2), .A0_f (new_AGEMA_signal_10116), .A1_t (new_AGEMA_signal_10117), .A1_f (new_AGEMA_signal_10118), .B0_t (KeyArray_S23reg_gff_1_SFF_0_n1), .B0_f (new_AGEMA_signal_9030), .B1_t (new_AGEMA_signal_9031), .B1_f (new_AGEMA_signal_9032), .Z0_t (KeyArray_outS23ser[0]), .Z0_f (new_AGEMA_signal_5085), .Z1_t (new_AGEMA_signal_5086), .Z1_f (new_AGEMA_signal_5087) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_0_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS23ser[0]), .B0_f (new_AGEMA_signal_5085), .B1_t (new_AGEMA_signal_5086), .B1_f (new_AGEMA_signal_5087), .Z0_t (KeyArray_S23reg_gff_1_SFF_0_n1), .Z0_f (new_AGEMA_signal_9030), .Z1_t (new_AGEMA_signal_9031), .Z1_f (new_AGEMA_signal_9032) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_0_U1 ( .A0_t (KeyArray_S23reg_gff_1_SFF_0_QD), .A0_f (new_AGEMA_signal_9640), .A1_t (new_AGEMA_signal_9641), .A1_f (new_AGEMA_signal_9642), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S23reg_gff_1_SFF_0_n2), .Z0_f (new_AGEMA_signal_10116), .Z1_t (new_AGEMA_signal_10117), .Z1_f (new_AGEMA_signal_10118) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS23ser[0]), .A0_f (new_AGEMA_signal_7150), .A1_t (new_AGEMA_signal_7151), .A1_f (new_AGEMA_signal_7152), .B0_t (KeyArray_outS33ser[0]), .B0_f (new_AGEMA_signal_5373), .B1_t (new_AGEMA_signal_5374), .B1_f (new_AGEMA_signal_5375), .Z0_t (KeyArray_S23reg_gff_1_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_7983), .Z1_t (new_AGEMA_signal_7984), .Z1_f (new_AGEMA_signal_7985) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S23reg_gff_1_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_7983), .B1_t (new_AGEMA_signal_7984), .B1_f (new_AGEMA_signal_7985), .Z0_t (KeyArray_S23reg_gff_1_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_9033), .Z1_t (new_AGEMA_signal_9034), .Z1_f (new_AGEMA_signal_9035) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S23reg_gff_1_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_9033), .A1_t (new_AGEMA_signal_9034), .A1_f (new_AGEMA_signal_9035), .B0_t (KeyArray_inS23ser[0]), .B0_f (new_AGEMA_signal_7150), .B1_t (new_AGEMA_signal_7151), .B1_f (new_AGEMA_signal_7152), .Z0_t (KeyArray_S23reg_gff_1_SFF_0_QD), .Z0_f (new_AGEMA_signal_9640), .Z1_t (new_AGEMA_signal_9641), .Z1_f (new_AGEMA_signal_9642) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S23reg_gff_1_SFF_1_U3 ( .A0_t (KeyArray_S23reg_gff_1_SFF_1_n2), .A0_f (new_AGEMA_signal_10119), .A1_t (new_AGEMA_signal_10120), .A1_f (new_AGEMA_signal_10121), .B0_t (KeyArray_S23reg_gff_1_SFF_1_n1), .B0_f (new_AGEMA_signal_9036), .B1_t (new_AGEMA_signal_9037), .B1_f (new_AGEMA_signal_9038), .Z0_t (KeyArray_outS23ser[1]), .Z0_f (new_AGEMA_signal_5094), .Z1_t (new_AGEMA_signal_5095), .Z1_f (new_AGEMA_signal_5096) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_1_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS23ser[1]), .B0_f (new_AGEMA_signal_5094), .B1_t (new_AGEMA_signal_5095), .B1_f (new_AGEMA_signal_5096), .Z0_t (KeyArray_S23reg_gff_1_SFF_1_n1), .Z0_f (new_AGEMA_signal_9036), .Z1_t (new_AGEMA_signal_9037), .Z1_f (new_AGEMA_signal_9038) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_1_U1 ( .A0_t (KeyArray_S23reg_gff_1_SFF_1_QD), .A0_f (new_AGEMA_signal_9643), .A1_t (new_AGEMA_signal_9644), .A1_f (new_AGEMA_signal_9645), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S23reg_gff_1_SFF_1_n2), .Z0_f (new_AGEMA_signal_10119), .Z1_t (new_AGEMA_signal_10120), .Z1_f (new_AGEMA_signal_10121) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS23ser[1]), .A0_f (new_AGEMA_signal_7153), .A1_t (new_AGEMA_signal_7154), .A1_f (new_AGEMA_signal_7155), .B0_t (KeyArray_outS33ser[1]), .B0_f (new_AGEMA_signal_5382), .B1_t (new_AGEMA_signal_5383), .B1_f (new_AGEMA_signal_5384), .Z0_t (KeyArray_S23reg_gff_1_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_7986), .Z1_t (new_AGEMA_signal_7987), .Z1_f (new_AGEMA_signal_7988) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S23reg_gff_1_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_7986), .B1_t (new_AGEMA_signal_7987), .B1_f (new_AGEMA_signal_7988), .Z0_t (KeyArray_S23reg_gff_1_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_9039), .Z1_t (new_AGEMA_signal_9040), .Z1_f (new_AGEMA_signal_9041) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S23reg_gff_1_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_9039), .A1_t (new_AGEMA_signal_9040), .A1_f (new_AGEMA_signal_9041), .B0_t (KeyArray_inS23ser[1]), .B0_f (new_AGEMA_signal_7153), .B1_t (new_AGEMA_signal_7154), .B1_f (new_AGEMA_signal_7155), .Z0_t (KeyArray_S23reg_gff_1_SFF_1_QD), .Z0_f (new_AGEMA_signal_9643), .Z1_t (new_AGEMA_signal_9644), .Z1_f (new_AGEMA_signal_9645) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S23reg_gff_1_SFF_2_U3 ( .A0_t (KeyArray_S23reg_gff_1_SFF_2_n2), .A0_f (new_AGEMA_signal_10122), .A1_t (new_AGEMA_signal_10123), .A1_f (new_AGEMA_signal_10124), .B0_t (KeyArray_S23reg_gff_1_SFF_2_n1), .B0_f (new_AGEMA_signal_9042), .B1_t (new_AGEMA_signal_9043), .B1_f (new_AGEMA_signal_9044), .Z0_t (KeyArray_outS23ser[2]), .Z0_f (new_AGEMA_signal_5103), .Z1_t (new_AGEMA_signal_5104), .Z1_f (new_AGEMA_signal_5105) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_2_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS23ser[2]), .B0_f (new_AGEMA_signal_5103), .B1_t (new_AGEMA_signal_5104), .B1_f (new_AGEMA_signal_5105), .Z0_t (KeyArray_S23reg_gff_1_SFF_2_n1), .Z0_f (new_AGEMA_signal_9042), .Z1_t (new_AGEMA_signal_9043), .Z1_f (new_AGEMA_signal_9044) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_2_U1 ( .A0_t (KeyArray_S23reg_gff_1_SFF_2_QD), .A0_f (new_AGEMA_signal_9646), .A1_t (new_AGEMA_signal_9647), .A1_f (new_AGEMA_signal_9648), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S23reg_gff_1_SFF_2_n2), .Z0_f (new_AGEMA_signal_10122), .Z1_t (new_AGEMA_signal_10123), .Z1_f (new_AGEMA_signal_10124) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS23ser[2]), .A0_f (new_AGEMA_signal_7156), .A1_t (new_AGEMA_signal_7157), .A1_f (new_AGEMA_signal_7158), .B0_t (KeyArray_outS33ser[2]), .B0_f (new_AGEMA_signal_5391), .B1_t (new_AGEMA_signal_5392), .B1_f (new_AGEMA_signal_5393), .Z0_t (KeyArray_S23reg_gff_1_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_7989), .Z1_t (new_AGEMA_signal_7990), .Z1_f (new_AGEMA_signal_7991) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S23reg_gff_1_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_7989), .B1_t (new_AGEMA_signal_7990), .B1_f (new_AGEMA_signal_7991), .Z0_t (KeyArray_S23reg_gff_1_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_9045), .Z1_t (new_AGEMA_signal_9046), .Z1_f (new_AGEMA_signal_9047) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S23reg_gff_1_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_9045), .A1_t (new_AGEMA_signal_9046), .A1_f (new_AGEMA_signal_9047), .B0_t (KeyArray_inS23ser[2]), .B0_f (new_AGEMA_signal_7156), .B1_t (new_AGEMA_signal_7157), .B1_f (new_AGEMA_signal_7158), .Z0_t (KeyArray_S23reg_gff_1_SFF_2_QD), .Z0_f (new_AGEMA_signal_9646), .Z1_t (new_AGEMA_signal_9647), .Z1_f (new_AGEMA_signal_9648) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S23reg_gff_1_SFF_3_U3 ( .A0_t (KeyArray_S23reg_gff_1_SFF_3_n2), .A0_f (new_AGEMA_signal_10125), .A1_t (new_AGEMA_signal_10126), .A1_f (new_AGEMA_signal_10127), .B0_t (KeyArray_S23reg_gff_1_SFF_3_n1), .B0_f (new_AGEMA_signal_9048), .B1_t (new_AGEMA_signal_9049), .B1_f (new_AGEMA_signal_9050), .Z0_t (KeyArray_outS23ser[3]), .Z0_f (new_AGEMA_signal_5112), .Z1_t (new_AGEMA_signal_5113), .Z1_f (new_AGEMA_signal_5114) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_3_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS23ser[3]), .B0_f (new_AGEMA_signal_5112), .B1_t (new_AGEMA_signal_5113), .B1_f (new_AGEMA_signal_5114), .Z0_t (KeyArray_S23reg_gff_1_SFF_3_n1), .Z0_f (new_AGEMA_signal_9048), .Z1_t (new_AGEMA_signal_9049), .Z1_f (new_AGEMA_signal_9050) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_3_U1 ( .A0_t (KeyArray_S23reg_gff_1_SFF_3_QD), .A0_f (new_AGEMA_signal_9649), .A1_t (new_AGEMA_signal_9650), .A1_f (new_AGEMA_signal_9651), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S23reg_gff_1_SFF_3_n2), .Z0_f (new_AGEMA_signal_10125), .Z1_t (new_AGEMA_signal_10126), .Z1_f (new_AGEMA_signal_10127) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS23ser[3]), .A0_f (new_AGEMA_signal_7159), .A1_t (new_AGEMA_signal_7160), .A1_f (new_AGEMA_signal_7161), .B0_t (KeyArray_outS33ser[3]), .B0_f (new_AGEMA_signal_5400), .B1_t (new_AGEMA_signal_5401), .B1_f (new_AGEMA_signal_5402), .Z0_t (KeyArray_S23reg_gff_1_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_7992), .Z1_t (new_AGEMA_signal_7993), .Z1_f (new_AGEMA_signal_7994) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S23reg_gff_1_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_7992), .B1_t (new_AGEMA_signal_7993), .B1_f (new_AGEMA_signal_7994), .Z0_t (KeyArray_S23reg_gff_1_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_9051), .Z1_t (new_AGEMA_signal_9052), .Z1_f (new_AGEMA_signal_9053) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S23reg_gff_1_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_9051), .A1_t (new_AGEMA_signal_9052), .A1_f (new_AGEMA_signal_9053), .B0_t (KeyArray_inS23ser[3]), .B0_f (new_AGEMA_signal_7159), .B1_t (new_AGEMA_signal_7160), .B1_f (new_AGEMA_signal_7161), .Z0_t (KeyArray_S23reg_gff_1_SFF_3_QD), .Z0_f (new_AGEMA_signal_9649), .Z1_t (new_AGEMA_signal_9650), .Z1_f (new_AGEMA_signal_9651) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S23reg_gff_1_SFF_4_U3 ( .A0_t (KeyArray_S23reg_gff_1_SFF_4_n2), .A0_f (new_AGEMA_signal_10128), .A1_t (new_AGEMA_signal_10129), .A1_f (new_AGEMA_signal_10130), .B0_t (KeyArray_S23reg_gff_1_SFF_4_n1), .B0_f (new_AGEMA_signal_9054), .B1_t (new_AGEMA_signal_9055), .B1_f (new_AGEMA_signal_9056), .Z0_t (KeyArray_outS23ser[4]), .Z0_f (new_AGEMA_signal_5121), .Z1_t (new_AGEMA_signal_5122), .Z1_f (new_AGEMA_signal_5123) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_4_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS23ser[4]), .B0_f (new_AGEMA_signal_5121), .B1_t (new_AGEMA_signal_5122), .B1_f (new_AGEMA_signal_5123), .Z0_t (KeyArray_S23reg_gff_1_SFF_4_n1), .Z0_f (new_AGEMA_signal_9054), .Z1_t (new_AGEMA_signal_9055), .Z1_f (new_AGEMA_signal_9056) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_4_U1 ( .A0_t (KeyArray_S23reg_gff_1_SFF_4_QD), .A0_f (new_AGEMA_signal_9652), .A1_t (new_AGEMA_signal_9653), .A1_f (new_AGEMA_signal_9654), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S23reg_gff_1_SFF_4_n2), .Z0_f (new_AGEMA_signal_10128), .Z1_t (new_AGEMA_signal_10129), .Z1_f (new_AGEMA_signal_10130) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS23ser[4]), .A0_f (new_AGEMA_signal_7162), .A1_t (new_AGEMA_signal_7163), .A1_f (new_AGEMA_signal_7164), .B0_t (KeyArray_outS33ser[4]), .B0_f (new_AGEMA_signal_5409), .B1_t (new_AGEMA_signal_5410), .B1_f (new_AGEMA_signal_5411), .Z0_t (KeyArray_S23reg_gff_1_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_7995), .Z1_t (new_AGEMA_signal_7996), .Z1_f (new_AGEMA_signal_7997) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S23reg_gff_1_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_7995), .B1_t (new_AGEMA_signal_7996), .B1_f (new_AGEMA_signal_7997), .Z0_t (KeyArray_S23reg_gff_1_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_9057), .Z1_t (new_AGEMA_signal_9058), .Z1_f (new_AGEMA_signal_9059) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S23reg_gff_1_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_9057), .A1_t (new_AGEMA_signal_9058), .A1_f (new_AGEMA_signal_9059), .B0_t (KeyArray_inS23ser[4]), .B0_f (new_AGEMA_signal_7162), .B1_t (new_AGEMA_signal_7163), .B1_f (new_AGEMA_signal_7164), .Z0_t (KeyArray_S23reg_gff_1_SFF_4_QD), .Z0_f (new_AGEMA_signal_9652), .Z1_t (new_AGEMA_signal_9653), .Z1_f (new_AGEMA_signal_9654) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S23reg_gff_1_SFF_5_U3 ( .A0_t (KeyArray_S23reg_gff_1_SFF_5_n2), .A0_f (new_AGEMA_signal_10131), .A1_t (new_AGEMA_signal_10132), .A1_f (new_AGEMA_signal_10133), .B0_t (KeyArray_S23reg_gff_1_SFF_5_n1), .B0_f (new_AGEMA_signal_9060), .B1_t (new_AGEMA_signal_9061), .B1_f (new_AGEMA_signal_9062), .Z0_t (KeyArray_outS23ser[5]), .Z0_f (new_AGEMA_signal_5130), .Z1_t (new_AGEMA_signal_5131), .Z1_f (new_AGEMA_signal_5132) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_5_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS23ser[5]), .B0_f (new_AGEMA_signal_5130), .B1_t (new_AGEMA_signal_5131), .B1_f (new_AGEMA_signal_5132), .Z0_t (KeyArray_S23reg_gff_1_SFF_5_n1), .Z0_f (new_AGEMA_signal_9060), .Z1_t (new_AGEMA_signal_9061), .Z1_f (new_AGEMA_signal_9062) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_5_U1 ( .A0_t (KeyArray_S23reg_gff_1_SFF_5_QD), .A0_f (new_AGEMA_signal_9655), .A1_t (new_AGEMA_signal_9656), .A1_f (new_AGEMA_signal_9657), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S23reg_gff_1_SFF_5_n2), .Z0_f (new_AGEMA_signal_10131), .Z1_t (new_AGEMA_signal_10132), .Z1_f (new_AGEMA_signal_10133) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS23ser[5]), .A0_f (new_AGEMA_signal_7165), .A1_t (new_AGEMA_signal_7166), .A1_f (new_AGEMA_signal_7167), .B0_t (KeyArray_outS33ser[5]), .B0_f (new_AGEMA_signal_5418), .B1_t (new_AGEMA_signal_5419), .B1_f (new_AGEMA_signal_5420), .Z0_t (KeyArray_S23reg_gff_1_SFF_5_MUXInst_X), .Z0_f (new_AGEMA_signal_7998), .Z1_t (new_AGEMA_signal_7999), .Z1_f (new_AGEMA_signal_8000) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S23reg_gff_1_SFF_5_MUXInst_X), .B0_f (new_AGEMA_signal_7998), .B1_t (new_AGEMA_signal_7999), .B1_f (new_AGEMA_signal_8000), .Z0_t (KeyArray_S23reg_gff_1_SFF_5_MUXInst_Y), .Z0_f (new_AGEMA_signal_9063), .Z1_t (new_AGEMA_signal_9064), .Z1_f (new_AGEMA_signal_9065) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S23reg_gff_1_SFF_5_MUXInst_Y), .A0_f (new_AGEMA_signal_9063), .A1_t (new_AGEMA_signal_9064), .A1_f (new_AGEMA_signal_9065), .B0_t (KeyArray_inS23ser[5]), .B0_f (new_AGEMA_signal_7165), .B1_t (new_AGEMA_signal_7166), .B1_f (new_AGEMA_signal_7167), .Z0_t (KeyArray_S23reg_gff_1_SFF_5_QD), .Z0_f (new_AGEMA_signal_9655), .Z1_t (new_AGEMA_signal_9656), .Z1_f (new_AGEMA_signal_9657) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S23reg_gff_1_SFF_6_U3 ( .A0_t (KeyArray_S23reg_gff_1_SFF_6_n2), .A0_f (new_AGEMA_signal_10134), .A1_t (new_AGEMA_signal_10135), .A1_f (new_AGEMA_signal_10136), .B0_t (KeyArray_S23reg_gff_1_SFF_6_n1), .B0_f (new_AGEMA_signal_9066), .B1_t (new_AGEMA_signal_9067), .B1_f (new_AGEMA_signal_9068), .Z0_t (KeyArray_outS23ser[6]), .Z0_f (new_AGEMA_signal_5139), .Z1_t (new_AGEMA_signal_5140), .Z1_f (new_AGEMA_signal_5141) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_6_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS23ser[6]), .B0_f (new_AGEMA_signal_5139), .B1_t (new_AGEMA_signal_5140), .B1_f (new_AGEMA_signal_5141), .Z0_t (KeyArray_S23reg_gff_1_SFF_6_n1), .Z0_f (new_AGEMA_signal_9066), .Z1_t (new_AGEMA_signal_9067), .Z1_f (new_AGEMA_signal_9068) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_6_U1 ( .A0_t (KeyArray_S23reg_gff_1_SFF_6_QD), .A0_f (new_AGEMA_signal_9658), .A1_t (new_AGEMA_signal_9659), .A1_f (new_AGEMA_signal_9660), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S23reg_gff_1_SFF_6_n2), .Z0_f (new_AGEMA_signal_10134), .Z1_t (new_AGEMA_signal_10135), .Z1_f (new_AGEMA_signal_10136) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS23ser[6]), .A0_f (new_AGEMA_signal_7168), .A1_t (new_AGEMA_signal_7169), .A1_f (new_AGEMA_signal_7170), .B0_t (KeyArray_outS33ser[6]), .B0_f (new_AGEMA_signal_5427), .B1_t (new_AGEMA_signal_5428), .B1_f (new_AGEMA_signal_5429), .Z0_t (KeyArray_S23reg_gff_1_SFF_6_MUXInst_X), .Z0_f (new_AGEMA_signal_8001), .Z1_t (new_AGEMA_signal_8002), .Z1_f (new_AGEMA_signal_8003) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S23reg_gff_1_SFF_6_MUXInst_X), .B0_f (new_AGEMA_signal_8001), .B1_t (new_AGEMA_signal_8002), .B1_f (new_AGEMA_signal_8003), .Z0_t (KeyArray_S23reg_gff_1_SFF_6_MUXInst_Y), .Z0_f (new_AGEMA_signal_9069), .Z1_t (new_AGEMA_signal_9070), .Z1_f (new_AGEMA_signal_9071) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S23reg_gff_1_SFF_6_MUXInst_Y), .A0_f (new_AGEMA_signal_9069), .A1_t (new_AGEMA_signal_9070), .A1_f (new_AGEMA_signal_9071), .B0_t (KeyArray_inS23ser[6]), .B0_f (new_AGEMA_signal_7168), .B1_t (new_AGEMA_signal_7169), .B1_f (new_AGEMA_signal_7170), .Z0_t (KeyArray_S23reg_gff_1_SFF_6_QD), .Z0_f (new_AGEMA_signal_9658), .Z1_t (new_AGEMA_signal_9659), .Z1_f (new_AGEMA_signal_9660) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S23reg_gff_1_SFF_7_U3 ( .A0_t (KeyArray_S23reg_gff_1_SFF_7_n2), .A0_f (new_AGEMA_signal_10137), .A1_t (new_AGEMA_signal_10138), .A1_f (new_AGEMA_signal_10139), .B0_t (KeyArray_S23reg_gff_1_SFF_7_n1), .B0_f (new_AGEMA_signal_9072), .B1_t (new_AGEMA_signal_9073), .B1_f (new_AGEMA_signal_9074), .Z0_t (KeyArray_outS23ser[7]), .Z0_f (new_AGEMA_signal_5148), .Z1_t (new_AGEMA_signal_5149), .Z1_f (new_AGEMA_signal_5150) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_7_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS23ser[7]), .B0_f (new_AGEMA_signal_5148), .B1_t (new_AGEMA_signal_5149), .B1_f (new_AGEMA_signal_5150), .Z0_t (KeyArray_S23reg_gff_1_SFF_7_n1), .Z0_f (new_AGEMA_signal_9072), .Z1_t (new_AGEMA_signal_9073), .Z1_f (new_AGEMA_signal_9074) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_7_U1 ( .A0_t (KeyArray_S23reg_gff_1_SFF_7_QD), .A0_f (new_AGEMA_signal_9661), .A1_t (new_AGEMA_signal_9662), .A1_f (new_AGEMA_signal_9663), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S23reg_gff_1_SFF_7_n2), .Z0_f (new_AGEMA_signal_10137), .Z1_t (new_AGEMA_signal_10138), .Z1_f (new_AGEMA_signal_10139) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS23ser[7]), .A0_f (new_AGEMA_signal_7171), .A1_t (new_AGEMA_signal_7172), .A1_f (new_AGEMA_signal_7173), .B0_t (KeyArray_outS33ser[7]), .B0_f (new_AGEMA_signal_5436), .B1_t (new_AGEMA_signal_5437), .B1_f (new_AGEMA_signal_5438), .Z0_t (KeyArray_S23reg_gff_1_SFF_7_MUXInst_X), .Z0_f (new_AGEMA_signal_8004), .Z1_t (new_AGEMA_signal_8005), .Z1_f (new_AGEMA_signal_8006) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S23reg_gff_1_SFF_7_MUXInst_X), .B0_f (new_AGEMA_signal_8004), .B1_t (new_AGEMA_signal_8005), .B1_f (new_AGEMA_signal_8006), .Z0_t (KeyArray_S23reg_gff_1_SFF_7_MUXInst_Y), .Z0_f (new_AGEMA_signal_9075), .Z1_t (new_AGEMA_signal_9076), .Z1_f (new_AGEMA_signal_9077) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S23reg_gff_1_SFF_7_MUXInst_Y), .A0_f (new_AGEMA_signal_9075), .A1_t (new_AGEMA_signal_9076), .A1_f (new_AGEMA_signal_9077), .B0_t (KeyArray_inS23ser[7]), .B0_f (new_AGEMA_signal_7171), .B1_t (new_AGEMA_signal_7172), .B1_f (new_AGEMA_signal_7173), .Z0_t (KeyArray_S23reg_gff_1_SFF_7_QD), .Z0_f (new_AGEMA_signal_9661), .Z1_t (new_AGEMA_signal_9662), .Z1_f (new_AGEMA_signal_9663) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S30reg_gff_1_SFF_0_U3 ( .A0_t (KeyArray_S30reg_gff_1_SFF_0_n2), .A0_f (new_AGEMA_signal_11567), .A1_t (new_AGEMA_signal_11568), .A1_f (new_AGEMA_signal_11569), .B0_t (KeyArray_S30reg_gff_1_SFF_0_n1), .B0_f (new_AGEMA_signal_9078), .B1_t (new_AGEMA_signal_9079), .B1_f (new_AGEMA_signal_9080), .Z0_t (KeyArray_outS30ser[0]), .Z0_f (new_AGEMA_signal_5157), .Z1_t (new_AGEMA_signal_5158), .Z1_f (new_AGEMA_signal_5159) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_0_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS30ser[0]), .B0_f (new_AGEMA_signal_5157), .B1_t (new_AGEMA_signal_5158), .B1_f (new_AGEMA_signal_5159), .Z0_t (KeyArray_S30reg_gff_1_SFF_0_n1), .Z0_f (new_AGEMA_signal_9078), .Z1_t (new_AGEMA_signal_9079), .Z1_f (new_AGEMA_signal_9080) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_0_U1 ( .A0_t (KeyArray_S30reg_gff_1_SFF_0_QD), .A0_f (new_AGEMA_signal_11519), .A1_t (new_AGEMA_signal_11520), .A1_f (new_AGEMA_signal_11521), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S30reg_gff_1_SFF_0_n2), .Z0_f (new_AGEMA_signal_11567), .Z1_t (new_AGEMA_signal_11568), .Z1_f (new_AGEMA_signal_11569) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS30ser[0]), .A0_f (new_AGEMA_signal_7174), .A1_t (new_AGEMA_signal_7175), .A1_f (new_AGEMA_signal_7176), .B0_t (KeyArray_inS30par[0]), .B0_f (new_AGEMA_signal_11396), .B1_t (new_AGEMA_signal_11397), .B1_f (new_AGEMA_signal_11398), .Z0_t (KeyArray_S30reg_gff_1_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_11444), .Z1_t (new_AGEMA_signal_11445), .Z1_f (new_AGEMA_signal_11446) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S30reg_gff_1_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_11444), .B1_t (new_AGEMA_signal_11445), .B1_f (new_AGEMA_signal_11446), .Z0_t (KeyArray_S30reg_gff_1_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_11471), .Z1_t (new_AGEMA_signal_11472), .Z1_f (new_AGEMA_signal_11473) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S30reg_gff_1_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_11471), .A1_t (new_AGEMA_signal_11472), .A1_f (new_AGEMA_signal_11473), .B0_t (KeyArray_inS30ser[0]), .B0_f (new_AGEMA_signal_7174), .B1_t (new_AGEMA_signal_7175), .B1_f (new_AGEMA_signal_7176), .Z0_t (KeyArray_S30reg_gff_1_SFF_0_QD), .Z0_f (new_AGEMA_signal_11519), .Z1_t (new_AGEMA_signal_11520), .Z1_f (new_AGEMA_signal_11521) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S30reg_gff_1_SFF_1_U3 ( .A0_t (KeyArray_S30reg_gff_1_SFF_1_n2), .A0_f (new_AGEMA_signal_11618), .A1_t (new_AGEMA_signal_11619), .A1_f (new_AGEMA_signal_11620), .B0_t (KeyArray_S30reg_gff_1_SFF_1_n1), .B0_f (new_AGEMA_signal_9081), .B1_t (new_AGEMA_signal_9082), .B1_f (new_AGEMA_signal_9083), .Z0_t (KeyArray_outS30ser[1]), .Z0_f (new_AGEMA_signal_5166), .Z1_t (new_AGEMA_signal_5167), .Z1_f (new_AGEMA_signal_5168) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_1_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS30ser[1]), .B0_f (new_AGEMA_signal_5166), .B1_t (new_AGEMA_signal_5167), .B1_f (new_AGEMA_signal_5168), .Z0_t (KeyArray_S30reg_gff_1_SFF_1_n1), .Z0_f (new_AGEMA_signal_9081), .Z1_t (new_AGEMA_signal_9082), .Z1_f (new_AGEMA_signal_9083) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_1_U1 ( .A0_t (KeyArray_S30reg_gff_1_SFF_1_QD), .A0_f (new_AGEMA_signal_11570), .A1_t (new_AGEMA_signal_11571), .A1_f (new_AGEMA_signal_11572), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S30reg_gff_1_SFF_1_n2), .Z0_f (new_AGEMA_signal_11618), .Z1_t (new_AGEMA_signal_11619), .Z1_f (new_AGEMA_signal_11620) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS30ser[1]), .A0_f (new_AGEMA_signal_7177), .A1_t (new_AGEMA_signal_7178), .A1_f (new_AGEMA_signal_7179), .B0_t (KeyArray_inS30par[1]), .B0_f (new_AGEMA_signal_11441), .B1_t (new_AGEMA_signal_11442), .B1_f (new_AGEMA_signal_11443), .Z0_t (KeyArray_S30reg_gff_1_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_11474), .Z1_t (new_AGEMA_signal_11475), .Z1_f (new_AGEMA_signal_11476) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S30reg_gff_1_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_11474), .B1_t (new_AGEMA_signal_11475), .B1_f (new_AGEMA_signal_11476), .Z0_t (KeyArray_S30reg_gff_1_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_11522), .Z1_t (new_AGEMA_signal_11523), .Z1_f (new_AGEMA_signal_11524) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S30reg_gff_1_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_11522), .A1_t (new_AGEMA_signal_11523), .A1_f (new_AGEMA_signal_11524), .B0_t (KeyArray_inS30ser[1]), .B0_f (new_AGEMA_signal_7177), .B1_t (new_AGEMA_signal_7178), .B1_f (new_AGEMA_signal_7179), .Z0_t (KeyArray_S30reg_gff_1_SFF_1_QD), .Z0_f (new_AGEMA_signal_11570), .Z1_t (new_AGEMA_signal_11571), .Z1_f (new_AGEMA_signal_11572) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S30reg_gff_1_SFF_2_U3 ( .A0_t (KeyArray_S30reg_gff_1_SFF_2_n2), .A0_f (new_AGEMA_signal_11621), .A1_t (new_AGEMA_signal_11622), .A1_f (new_AGEMA_signal_11623), .B0_t (KeyArray_S30reg_gff_1_SFF_2_n1), .B0_f (new_AGEMA_signal_9084), .B1_t (new_AGEMA_signal_9085), .B1_f (new_AGEMA_signal_9086), .Z0_t (KeyArray_outS30ser[2]), .Z0_f (new_AGEMA_signal_5175), .Z1_t (new_AGEMA_signal_5176), .Z1_f (new_AGEMA_signal_5177) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_2_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS30ser[2]), .B0_f (new_AGEMA_signal_5175), .B1_t (new_AGEMA_signal_5176), .B1_f (new_AGEMA_signal_5177), .Z0_t (KeyArray_S30reg_gff_1_SFF_2_n1), .Z0_f (new_AGEMA_signal_9084), .Z1_t (new_AGEMA_signal_9085), .Z1_f (new_AGEMA_signal_9086) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_2_U1 ( .A0_t (KeyArray_S30reg_gff_1_SFF_2_QD), .A0_f (new_AGEMA_signal_11573), .A1_t (new_AGEMA_signal_11574), .A1_f (new_AGEMA_signal_11575), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S30reg_gff_1_SFF_2_n2), .Z0_f (new_AGEMA_signal_11621), .Z1_t (new_AGEMA_signal_11622), .Z1_f (new_AGEMA_signal_11623) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS30ser[2]), .A0_f (new_AGEMA_signal_7180), .A1_t (new_AGEMA_signal_7181), .A1_f (new_AGEMA_signal_7182), .B0_t (KeyArray_inS30par[2]), .B0_f (new_AGEMA_signal_11438), .B1_t (new_AGEMA_signal_11439), .B1_f (new_AGEMA_signal_11440), .Z0_t (KeyArray_S30reg_gff_1_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_11477), .Z1_t (new_AGEMA_signal_11478), .Z1_f (new_AGEMA_signal_11479) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S30reg_gff_1_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_11477), .B1_t (new_AGEMA_signal_11478), .B1_f (new_AGEMA_signal_11479), .Z0_t (KeyArray_S30reg_gff_1_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_11525), .Z1_t (new_AGEMA_signal_11526), .Z1_f (new_AGEMA_signal_11527) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S30reg_gff_1_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_11525), .A1_t (new_AGEMA_signal_11526), .A1_f (new_AGEMA_signal_11527), .B0_t (KeyArray_inS30ser[2]), .B0_f (new_AGEMA_signal_7180), .B1_t (new_AGEMA_signal_7181), .B1_f (new_AGEMA_signal_7182), .Z0_t (KeyArray_S30reg_gff_1_SFF_2_QD), .Z0_f (new_AGEMA_signal_11573), .Z1_t (new_AGEMA_signal_11574), .Z1_f (new_AGEMA_signal_11575) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S30reg_gff_1_SFF_3_U3 ( .A0_t (KeyArray_S30reg_gff_1_SFF_3_n2), .A0_f (new_AGEMA_signal_11624), .A1_t (new_AGEMA_signal_11625), .A1_f (new_AGEMA_signal_11626), .B0_t (KeyArray_S30reg_gff_1_SFF_3_n1), .B0_f (new_AGEMA_signal_9087), .B1_t (new_AGEMA_signal_9088), .B1_f (new_AGEMA_signal_9089), .Z0_t (KeyArray_outS30ser[3]), .Z0_f (new_AGEMA_signal_5184), .Z1_t (new_AGEMA_signal_5185), .Z1_f (new_AGEMA_signal_5186) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_3_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS30ser[3]), .B0_f (new_AGEMA_signal_5184), .B1_t (new_AGEMA_signal_5185), .B1_f (new_AGEMA_signal_5186), .Z0_t (KeyArray_S30reg_gff_1_SFF_3_n1), .Z0_f (new_AGEMA_signal_9087), .Z1_t (new_AGEMA_signal_9088), .Z1_f (new_AGEMA_signal_9089) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_3_U1 ( .A0_t (KeyArray_S30reg_gff_1_SFF_3_QD), .A0_f (new_AGEMA_signal_11576), .A1_t (new_AGEMA_signal_11577), .A1_f (new_AGEMA_signal_11578), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S30reg_gff_1_SFF_3_n2), .Z0_f (new_AGEMA_signal_11624), .Z1_t (new_AGEMA_signal_11625), .Z1_f (new_AGEMA_signal_11626) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS30ser[3]), .A0_f (new_AGEMA_signal_7183), .A1_t (new_AGEMA_signal_7184), .A1_f (new_AGEMA_signal_7185), .B0_t (KeyArray_inS30par[3]), .B0_f (new_AGEMA_signal_11435), .B1_t (new_AGEMA_signal_11436), .B1_f (new_AGEMA_signal_11437), .Z0_t (KeyArray_S30reg_gff_1_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_11480), .Z1_t (new_AGEMA_signal_11481), .Z1_f (new_AGEMA_signal_11482) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S30reg_gff_1_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_11480), .B1_t (new_AGEMA_signal_11481), .B1_f (new_AGEMA_signal_11482), .Z0_t (KeyArray_S30reg_gff_1_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_11528), .Z1_t (new_AGEMA_signal_11529), .Z1_f (new_AGEMA_signal_11530) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S30reg_gff_1_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_11528), .A1_t (new_AGEMA_signal_11529), .A1_f (new_AGEMA_signal_11530), .B0_t (KeyArray_inS30ser[3]), .B0_f (new_AGEMA_signal_7183), .B1_t (new_AGEMA_signal_7184), .B1_f (new_AGEMA_signal_7185), .Z0_t (KeyArray_S30reg_gff_1_SFF_3_QD), .Z0_f (new_AGEMA_signal_11576), .Z1_t (new_AGEMA_signal_11577), .Z1_f (new_AGEMA_signal_11578) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S30reg_gff_1_SFF_4_U3 ( .A0_t (KeyArray_S30reg_gff_1_SFF_4_n2), .A0_f (new_AGEMA_signal_11627), .A1_t (new_AGEMA_signal_11628), .A1_f (new_AGEMA_signal_11629), .B0_t (KeyArray_S30reg_gff_1_SFF_4_n1), .B0_f (new_AGEMA_signal_9090), .B1_t (new_AGEMA_signal_9091), .B1_f (new_AGEMA_signal_9092), .Z0_t (KeyArray_outS30ser[4]), .Z0_f (new_AGEMA_signal_5193), .Z1_t (new_AGEMA_signal_5194), .Z1_f (new_AGEMA_signal_5195) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_4_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS30ser[4]), .B0_f (new_AGEMA_signal_5193), .B1_t (new_AGEMA_signal_5194), .B1_f (new_AGEMA_signal_5195), .Z0_t (KeyArray_S30reg_gff_1_SFF_4_n1), .Z0_f (new_AGEMA_signal_9090), .Z1_t (new_AGEMA_signal_9091), .Z1_f (new_AGEMA_signal_9092) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_4_U1 ( .A0_t (KeyArray_S30reg_gff_1_SFF_4_QD), .A0_f (new_AGEMA_signal_11579), .A1_t (new_AGEMA_signal_11580), .A1_f (new_AGEMA_signal_11581), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S30reg_gff_1_SFF_4_n2), .Z0_f (new_AGEMA_signal_11627), .Z1_t (new_AGEMA_signal_11628), .Z1_f (new_AGEMA_signal_11629) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS30ser[4]), .A0_f (new_AGEMA_signal_7186), .A1_t (new_AGEMA_signal_7187), .A1_f (new_AGEMA_signal_7188), .B0_t (KeyArray_inS30par[4]), .B0_f (new_AGEMA_signal_11432), .B1_t (new_AGEMA_signal_11433), .B1_f (new_AGEMA_signal_11434), .Z0_t (KeyArray_S30reg_gff_1_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_11483), .Z1_t (new_AGEMA_signal_11484), .Z1_f (new_AGEMA_signal_11485) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S30reg_gff_1_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_11483), .B1_t (new_AGEMA_signal_11484), .B1_f (new_AGEMA_signal_11485), .Z0_t (KeyArray_S30reg_gff_1_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_11531), .Z1_t (new_AGEMA_signal_11532), .Z1_f (new_AGEMA_signal_11533) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S30reg_gff_1_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_11531), .A1_t (new_AGEMA_signal_11532), .A1_f (new_AGEMA_signal_11533), .B0_t (KeyArray_inS30ser[4]), .B0_f (new_AGEMA_signal_7186), .B1_t (new_AGEMA_signal_7187), .B1_f (new_AGEMA_signal_7188), .Z0_t (KeyArray_S30reg_gff_1_SFF_4_QD), .Z0_f (new_AGEMA_signal_11579), .Z1_t (new_AGEMA_signal_11580), .Z1_f (new_AGEMA_signal_11581) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S30reg_gff_1_SFF_5_U3 ( .A0_t (KeyArray_S30reg_gff_1_SFF_5_n2), .A0_f (new_AGEMA_signal_11630), .A1_t (new_AGEMA_signal_11631), .A1_f (new_AGEMA_signal_11632), .B0_t (KeyArray_S30reg_gff_1_SFF_5_n1), .B0_f (new_AGEMA_signal_9093), .B1_t (new_AGEMA_signal_9094), .B1_f (new_AGEMA_signal_9095), .Z0_t (KeyArray_outS30ser[5]), .Z0_f (new_AGEMA_signal_5202), .Z1_t (new_AGEMA_signal_5203), .Z1_f (new_AGEMA_signal_5204) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_5_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS30ser[5]), .B0_f (new_AGEMA_signal_5202), .B1_t (new_AGEMA_signal_5203), .B1_f (new_AGEMA_signal_5204), .Z0_t (KeyArray_S30reg_gff_1_SFF_5_n1), .Z0_f (new_AGEMA_signal_9093), .Z1_t (new_AGEMA_signal_9094), .Z1_f (new_AGEMA_signal_9095) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_5_U1 ( .A0_t (KeyArray_S30reg_gff_1_SFF_5_QD), .A0_f (new_AGEMA_signal_11582), .A1_t (new_AGEMA_signal_11583), .A1_f (new_AGEMA_signal_11584), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S30reg_gff_1_SFF_5_n2), .Z0_f (new_AGEMA_signal_11630), .Z1_t (new_AGEMA_signal_11631), .Z1_f (new_AGEMA_signal_11632) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS30ser[5]), .A0_f (new_AGEMA_signal_7189), .A1_t (new_AGEMA_signal_7190), .A1_f (new_AGEMA_signal_7191), .B0_t (KeyArray_inS30par[5]), .B0_f (new_AGEMA_signal_11429), .B1_t (new_AGEMA_signal_11430), .B1_f (new_AGEMA_signal_11431), .Z0_t (KeyArray_S30reg_gff_1_SFF_5_MUXInst_X), .Z0_f (new_AGEMA_signal_11486), .Z1_t (new_AGEMA_signal_11487), .Z1_f (new_AGEMA_signal_11488) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S30reg_gff_1_SFF_5_MUXInst_X), .B0_f (new_AGEMA_signal_11486), .B1_t (new_AGEMA_signal_11487), .B1_f (new_AGEMA_signal_11488), .Z0_t (KeyArray_S30reg_gff_1_SFF_5_MUXInst_Y), .Z0_f (new_AGEMA_signal_11534), .Z1_t (new_AGEMA_signal_11535), .Z1_f (new_AGEMA_signal_11536) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S30reg_gff_1_SFF_5_MUXInst_Y), .A0_f (new_AGEMA_signal_11534), .A1_t (new_AGEMA_signal_11535), .A1_f (new_AGEMA_signal_11536), .B0_t (KeyArray_inS30ser[5]), .B0_f (new_AGEMA_signal_7189), .B1_t (new_AGEMA_signal_7190), .B1_f (new_AGEMA_signal_7191), .Z0_t (KeyArray_S30reg_gff_1_SFF_5_QD), .Z0_f (new_AGEMA_signal_11582), .Z1_t (new_AGEMA_signal_11583), .Z1_f (new_AGEMA_signal_11584) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S30reg_gff_1_SFF_6_U3 ( .A0_t (KeyArray_S30reg_gff_1_SFF_6_n2), .A0_f (new_AGEMA_signal_11633), .A1_t (new_AGEMA_signal_11634), .A1_f (new_AGEMA_signal_11635), .B0_t (KeyArray_S30reg_gff_1_SFF_6_n1), .B0_f (new_AGEMA_signal_9096), .B1_t (new_AGEMA_signal_9097), .B1_f (new_AGEMA_signal_9098), .Z0_t (KeyArray_outS30ser[6]), .Z0_f (new_AGEMA_signal_5211), .Z1_t (new_AGEMA_signal_5212), .Z1_f (new_AGEMA_signal_5213) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_6_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS30ser[6]), .B0_f (new_AGEMA_signal_5211), .B1_t (new_AGEMA_signal_5212), .B1_f (new_AGEMA_signal_5213), .Z0_t (KeyArray_S30reg_gff_1_SFF_6_n1), .Z0_f (new_AGEMA_signal_9096), .Z1_t (new_AGEMA_signal_9097), .Z1_f (new_AGEMA_signal_9098) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_6_U1 ( .A0_t (KeyArray_S30reg_gff_1_SFF_6_QD), .A0_f (new_AGEMA_signal_11585), .A1_t (new_AGEMA_signal_11586), .A1_f (new_AGEMA_signal_11587), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S30reg_gff_1_SFF_6_n2), .Z0_f (new_AGEMA_signal_11633), .Z1_t (new_AGEMA_signal_11634), .Z1_f (new_AGEMA_signal_11635) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS30ser[6]), .A0_f (new_AGEMA_signal_7192), .A1_t (new_AGEMA_signal_7193), .A1_f (new_AGEMA_signal_7194), .B0_t (KeyArray_inS30par[6]), .B0_f (new_AGEMA_signal_11426), .B1_t (new_AGEMA_signal_11427), .B1_f (new_AGEMA_signal_11428), .Z0_t (KeyArray_S30reg_gff_1_SFF_6_MUXInst_X), .Z0_f (new_AGEMA_signal_11489), .Z1_t (new_AGEMA_signal_11490), .Z1_f (new_AGEMA_signal_11491) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S30reg_gff_1_SFF_6_MUXInst_X), .B0_f (new_AGEMA_signal_11489), .B1_t (new_AGEMA_signal_11490), .B1_f (new_AGEMA_signal_11491), .Z0_t (KeyArray_S30reg_gff_1_SFF_6_MUXInst_Y), .Z0_f (new_AGEMA_signal_11537), .Z1_t (new_AGEMA_signal_11538), .Z1_f (new_AGEMA_signal_11539) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S30reg_gff_1_SFF_6_MUXInst_Y), .A0_f (new_AGEMA_signal_11537), .A1_t (new_AGEMA_signal_11538), .A1_f (new_AGEMA_signal_11539), .B0_t (KeyArray_inS30ser[6]), .B0_f (new_AGEMA_signal_7192), .B1_t (new_AGEMA_signal_7193), .B1_f (new_AGEMA_signal_7194), .Z0_t (KeyArray_S30reg_gff_1_SFF_6_QD), .Z0_f (new_AGEMA_signal_11585), .Z1_t (new_AGEMA_signal_11586), .Z1_f (new_AGEMA_signal_11587) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S30reg_gff_1_SFF_7_U3 ( .A0_t (KeyArray_S30reg_gff_1_SFF_7_n2), .A0_f (new_AGEMA_signal_11636), .A1_t (new_AGEMA_signal_11637), .A1_f (new_AGEMA_signal_11638), .B0_t (KeyArray_S30reg_gff_1_SFF_7_n1), .B0_f (new_AGEMA_signal_9099), .B1_t (new_AGEMA_signal_9100), .B1_f (new_AGEMA_signal_9101), .Z0_t (KeyArray_outS30ser[7]), .Z0_f (new_AGEMA_signal_5220), .Z1_t (new_AGEMA_signal_5221), .Z1_f (new_AGEMA_signal_5222) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_7_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS30ser[7]), .B0_f (new_AGEMA_signal_5220), .B1_t (new_AGEMA_signal_5221), .B1_f (new_AGEMA_signal_5222), .Z0_t (KeyArray_S30reg_gff_1_SFF_7_n1), .Z0_f (new_AGEMA_signal_9099), .Z1_t (new_AGEMA_signal_9100), .Z1_f (new_AGEMA_signal_9101) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_7_U1 ( .A0_t (KeyArray_S30reg_gff_1_SFF_7_QD), .A0_f (new_AGEMA_signal_11588), .A1_t (new_AGEMA_signal_11589), .A1_f (new_AGEMA_signal_11590), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S30reg_gff_1_SFF_7_n2), .Z0_f (new_AGEMA_signal_11636), .Z1_t (new_AGEMA_signal_11637), .Z1_f (new_AGEMA_signal_11638) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS30ser[7]), .A0_f (new_AGEMA_signal_7195), .A1_t (new_AGEMA_signal_7196), .A1_f (new_AGEMA_signal_7197), .B0_t (KeyArray_inS30par[7]), .B0_f (new_AGEMA_signal_11423), .B1_t (new_AGEMA_signal_11424), .B1_f (new_AGEMA_signal_11425), .Z0_t (KeyArray_S30reg_gff_1_SFF_7_MUXInst_X), .Z0_f (new_AGEMA_signal_11492), .Z1_t (new_AGEMA_signal_11493), .Z1_f (new_AGEMA_signal_11494) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S30reg_gff_1_SFF_7_MUXInst_X), .B0_f (new_AGEMA_signal_11492), .B1_t (new_AGEMA_signal_11493), .B1_f (new_AGEMA_signal_11494), .Z0_t (KeyArray_S30reg_gff_1_SFF_7_MUXInst_Y), .Z0_f (new_AGEMA_signal_11540), .Z1_t (new_AGEMA_signal_11541), .Z1_f (new_AGEMA_signal_11542) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S30reg_gff_1_SFF_7_MUXInst_Y), .A0_f (new_AGEMA_signal_11540), .A1_t (new_AGEMA_signal_11541), .A1_f (new_AGEMA_signal_11542), .B0_t (KeyArray_inS30ser[7]), .B0_f (new_AGEMA_signal_7195), .B1_t (new_AGEMA_signal_7196), .B1_f (new_AGEMA_signal_7197), .Z0_t (KeyArray_S30reg_gff_1_SFF_7_QD), .Z0_f (new_AGEMA_signal_11588), .Z1_t (new_AGEMA_signal_11589), .Z1_f (new_AGEMA_signal_11590) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S31reg_gff_1_SFF_0_U3 ( .A0_t (KeyArray_S31reg_gff_1_SFF_0_n2), .A0_f (new_AGEMA_signal_10140), .A1_t (new_AGEMA_signal_10141), .A1_f (new_AGEMA_signal_10142), .B0_t (KeyArray_S31reg_gff_1_SFF_0_n1), .B0_f (new_AGEMA_signal_9102), .B1_t (new_AGEMA_signal_9103), .B1_f (new_AGEMA_signal_9104), .Z0_t (KeyArray_outS31ser[0]), .Z0_f (new_AGEMA_signal_5229), .Z1_t (new_AGEMA_signal_5230), .Z1_f (new_AGEMA_signal_5231) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_0_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS31ser[0]), .B0_f (new_AGEMA_signal_5229), .B1_t (new_AGEMA_signal_5230), .B1_f (new_AGEMA_signal_5231), .Z0_t (KeyArray_S31reg_gff_1_SFF_0_n1), .Z0_f (new_AGEMA_signal_9102), .Z1_t (new_AGEMA_signal_9103), .Z1_f (new_AGEMA_signal_9104) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_0_U1 ( .A0_t (KeyArray_S31reg_gff_1_SFF_0_QD), .A0_f (new_AGEMA_signal_9664), .A1_t (new_AGEMA_signal_9665), .A1_f (new_AGEMA_signal_9666), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S31reg_gff_1_SFF_0_n2), .Z0_f (new_AGEMA_signal_10140), .Z1_t (new_AGEMA_signal_10141), .Z1_f (new_AGEMA_signal_10142) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS31ser[0]), .A0_f (new_AGEMA_signal_7198), .A1_t (new_AGEMA_signal_7199), .A1_f (new_AGEMA_signal_7200), .B0_t (KeyArray_outS01ser_0_), .B0_f (new_AGEMA_signal_4428), .B1_t (new_AGEMA_signal_4429), .B1_f (new_AGEMA_signal_4430), .Z0_t (KeyArray_S31reg_gff_1_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_8007), .Z1_t (new_AGEMA_signal_8008), .Z1_f (new_AGEMA_signal_8009) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S31reg_gff_1_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_8007), .B1_t (new_AGEMA_signal_8008), .B1_f (new_AGEMA_signal_8009), .Z0_t (KeyArray_S31reg_gff_1_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_9105), .Z1_t (new_AGEMA_signal_9106), .Z1_f (new_AGEMA_signal_9107) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S31reg_gff_1_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_9105), .A1_t (new_AGEMA_signal_9106), .A1_f (new_AGEMA_signal_9107), .B0_t (KeyArray_inS31ser[0]), .B0_f (new_AGEMA_signal_7198), .B1_t (new_AGEMA_signal_7199), .B1_f (new_AGEMA_signal_7200), .Z0_t (KeyArray_S31reg_gff_1_SFF_0_QD), .Z0_f (new_AGEMA_signal_9664), .Z1_t (new_AGEMA_signal_9665), .Z1_f (new_AGEMA_signal_9666) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S31reg_gff_1_SFF_1_U3 ( .A0_t (KeyArray_S31reg_gff_1_SFF_1_n2), .A0_f (new_AGEMA_signal_10143), .A1_t (new_AGEMA_signal_10144), .A1_f (new_AGEMA_signal_10145), .B0_t (KeyArray_S31reg_gff_1_SFF_1_n1), .B0_f (new_AGEMA_signal_9108), .B1_t (new_AGEMA_signal_9109), .B1_f (new_AGEMA_signal_9110), .Z0_t (KeyArray_outS31ser[1]), .Z0_f (new_AGEMA_signal_5238), .Z1_t (new_AGEMA_signal_5239), .Z1_f (new_AGEMA_signal_5240) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_1_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS31ser[1]), .B0_f (new_AGEMA_signal_5238), .B1_t (new_AGEMA_signal_5239), .B1_f (new_AGEMA_signal_5240), .Z0_t (KeyArray_S31reg_gff_1_SFF_1_n1), .Z0_f (new_AGEMA_signal_9108), .Z1_t (new_AGEMA_signal_9109), .Z1_f (new_AGEMA_signal_9110) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_1_U1 ( .A0_t (KeyArray_S31reg_gff_1_SFF_1_QD), .A0_f (new_AGEMA_signal_9667), .A1_t (new_AGEMA_signal_9668), .A1_f (new_AGEMA_signal_9669), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S31reg_gff_1_SFF_1_n2), .Z0_f (new_AGEMA_signal_10143), .Z1_t (new_AGEMA_signal_10144), .Z1_f (new_AGEMA_signal_10145) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS31ser[1]), .A0_f (new_AGEMA_signal_7201), .A1_t (new_AGEMA_signal_7202), .A1_f (new_AGEMA_signal_7203), .B0_t (KeyArray_outS01ser_1_), .B0_f (new_AGEMA_signal_4422), .B1_t (new_AGEMA_signal_4423), .B1_f (new_AGEMA_signal_4424), .Z0_t (KeyArray_S31reg_gff_1_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_8010), .Z1_t (new_AGEMA_signal_8011), .Z1_f (new_AGEMA_signal_8012) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S31reg_gff_1_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_8010), .B1_t (new_AGEMA_signal_8011), .B1_f (new_AGEMA_signal_8012), .Z0_t (KeyArray_S31reg_gff_1_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_9111), .Z1_t (new_AGEMA_signal_9112), .Z1_f (new_AGEMA_signal_9113) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S31reg_gff_1_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_9111), .A1_t (new_AGEMA_signal_9112), .A1_f (new_AGEMA_signal_9113), .B0_t (KeyArray_inS31ser[1]), .B0_f (new_AGEMA_signal_7201), .B1_t (new_AGEMA_signal_7202), .B1_f (new_AGEMA_signal_7203), .Z0_t (KeyArray_S31reg_gff_1_SFF_1_QD), .Z0_f (new_AGEMA_signal_9667), .Z1_t (new_AGEMA_signal_9668), .Z1_f (new_AGEMA_signal_9669) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S31reg_gff_1_SFF_2_U3 ( .A0_t (KeyArray_S31reg_gff_1_SFF_2_n2), .A0_f (new_AGEMA_signal_10146), .A1_t (new_AGEMA_signal_10147), .A1_f (new_AGEMA_signal_10148), .B0_t (KeyArray_S31reg_gff_1_SFF_2_n1), .B0_f (new_AGEMA_signal_9114), .B1_t (new_AGEMA_signal_9115), .B1_f (new_AGEMA_signal_9116), .Z0_t (KeyArray_outS31ser[2]), .Z0_f (new_AGEMA_signal_5247), .Z1_t (new_AGEMA_signal_5248), .Z1_f (new_AGEMA_signal_5249) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_2_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS31ser[2]), .B0_f (new_AGEMA_signal_5247), .B1_t (new_AGEMA_signal_5248), .B1_f (new_AGEMA_signal_5249), .Z0_t (KeyArray_S31reg_gff_1_SFF_2_n1), .Z0_f (new_AGEMA_signal_9114), .Z1_t (new_AGEMA_signal_9115), .Z1_f (new_AGEMA_signal_9116) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_2_U1 ( .A0_t (KeyArray_S31reg_gff_1_SFF_2_QD), .A0_f (new_AGEMA_signal_9670), .A1_t (new_AGEMA_signal_9671), .A1_f (new_AGEMA_signal_9672), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S31reg_gff_1_SFF_2_n2), .Z0_f (new_AGEMA_signal_10146), .Z1_t (new_AGEMA_signal_10147), .Z1_f (new_AGEMA_signal_10148) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS31ser[2]), .A0_f (new_AGEMA_signal_7204), .A1_t (new_AGEMA_signal_7205), .A1_f (new_AGEMA_signal_7206), .B0_t (KeyArray_outS01ser_2_), .B0_f (new_AGEMA_signal_4416), .B1_t (new_AGEMA_signal_4417), .B1_f (new_AGEMA_signal_4418), .Z0_t (KeyArray_S31reg_gff_1_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_8013), .Z1_t (new_AGEMA_signal_8014), .Z1_f (new_AGEMA_signal_8015) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S31reg_gff_1_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_8013), .B1_t (new_AGEMA_signal_8014), .B1_f (new_AGEMA_signal_8015), .Z0_t (KeyArray_S31reg_gff_1_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_9117), .Z1_t (new_AGEMA_signal_9118), .Z1_f (new_AGEMA_signal_9119) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S31reg_gff_1_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_9117), .A1_t (new_AGEMA_signal_9118), .A1_f (new_AGEMA_signal_9119), .B0_t (KeyArray_inS31ser[2]), .B0_f (new_AGEMA_signal_7204), .B1_t (new_AGEMA_signal_7205), .B1_f (new_AGEMA_signal_7206), .Z0_t (KeyArray_S31reg_gff_1_SFF_2_QD), .Z0_f (new_AGEMA_signal_9670), .Z1_t (new_AGEMA_signal_9671), .Z1_f (new_AGEMA_signal_9672) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S31reg_gff_1_SFF_3_U3 ( .A0_t (KeyArray_S31reg_gff_1_SFF_3_n2), .A0_f (new_AGEMA_signal_10149), .A1_t (new_AGEMA_signal_10150), .A1_f (new_AGEMA_signal_10151), .B0_t (KeyArray_S31reg_gff_1_SFF_3_n1), .B0_f (new_AGEMA_signal_9120), .B1_t (new_AGEMA_signal_9121), .B1_f (new_AGEMA_signal_9122), .Z0_t (KeyArray_outS31ser[3]), .Z0_f (new_AGEMA_signal_5256), .Z1_t (new_AGEMA_signal_5257), .Z1_f (new_AGEMA_signal_5258) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_3_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS31ser[3]), .B0_f (new_AGEMA_signal_5256), .B1_t (new_AGEMA_signal_5257), .B1_f (new_AGEMA_signal_5258), .Z0_t (KeyArray_S31reg_gff_1_SFF_3_n1), .Z0_f (new_AGEMA_signal_9120), .Z1_t (new_AGEMA_signal_9121), .Z1_f (new_AGEMA_signal_9122) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_3_U1 ( .A0_t (KeyArray_S31reg_gff_1_SFF_3_QD), .A0_f (new_AGEMA_signal_9673), .A1_t (new_AGEMA_signal_9674), .A1_f (new_AGEMA_signal_9675), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S31reg_gff_1_SFF_3_n2), .Z0_f (new_AGEMA_signal_10149), .Z1_t (new_AGEMA_signal_10150), .Z1_f (new_AGEMA_signal_10151) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS31ser[3]), .A0_f (new_AGEMA_signal_7207), .A1_t (new_AGEMA_signal_7208), .A1_f (new_AGEMA_signal_7209), .B0_t (KeyArray_outS01ser_3_), .B0_f (new_AGEMA_signal_4410), .B1_t (new_AGEMA_signal_4411), .B1_f (new_AGEMA_signal_4412), .Z0_t (KeyArray_S31reg_gff_1_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_8016), .Z1_t (new_AGEMA_signal_8017), .Z1_f (new_AGEMA_signal_8018) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S31reg_gff_1_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_8016), .B1_t (new_AGEMA_signal_8017), .B1_f (new_AGEMA_signal_8018), .Z0_t (KeyArray_S31reg_gff_1_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_9123), .Z1_t (new_AGEMA_signal_9124), .Z1_f (new_AGEMA_signal_9125) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S31reg_gff_1_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_9123), .A1_t (new_AGEMA_signal_9124), .A1_f (new_AGEMA_signal_9125), .B0_t (KeyArray_inS31ser[3]), .B0_f (new_AGEMA_signal_7207), .B1_t (new_AGEMA_signal_7208), .B1_f (new_AGEMA_signal_7209), .Z0_t (KeyArray_S31reg_gff_1_SFF_3_QD), .Z0_f (new_AGEMA_signal_9673), .Z1_t (new_AGEMA_signal_9674), .Z1_f (new_AGEMA_signal_9675) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S31reg_gff_1_SFF_4_U3 ( .A0_t (KeyArray_S31reg_gff_1_SFF_4_n2), .A0_f (new_AGEMA_signal_10152), .A1_t (new_AGEMA_signal_10153), .A1_f (new_AGEMA_signal_10154), .B0_t (KeyArray_S31reg_gff_1_SFF_4_n1), .B0_f (new_AGEMA_signal_9126), .B1_t (new_AGEMA_signal_9127), .B1_f (new_AGEMA_signal_9128), .Z0_t (KeyArray_outS31ser[4]), .Z0_f (new_AGEMA_signal_5265), .Z1_t (new_AGEMA_signal_5266), .Z1_f (new_AGEMA_signal_5267) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_4_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS31ser[4]), .B0_f (new_AGEMA_signal_5265), .B1_t (new_AGEMA_signal_5266), .B1_f (new_AGEMA_signal_5267), .Z0_t (KeyArray_S31reg_gff_1_SFF_4_n1), .Z0_f (new_AGEMA_signal_9126), .Z1_t (new_AGEMA_signal_9127), .Z1_f (new_AGEMA_signal_9128) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_4_U1 ( .A0_t (KeyArray_S31reg_gff_1_SFF_4_QD), .A0_f (new_AGEMA_signal_9676), .A1_t (new_AGEMA_signal_9677), .A1_f (new_AGEMA_signal_9678), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S31reg_gff_1_SFF_4_n2), .Z0_f (new_AGEMA_signal_10152), .Z1_t (new_AGEMA_signal_10153), .Z1_f (new_AGEMA_signal_10154) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS31ser[4]), .A0_f (new_AGEMA_signal_7210), .A1_t (new_AGEMA_signal_7211), .A1_f (new_AGEMA_signal_7212), .B0_t (KeyArray_outS01ser_4_), .B0_f (new_AGEMA_signal_4404), .B1_t (new_AGEMA_signal_4405), .B1_f (new_AGEMA_signal_4406), .Z0_t (KeyArray_S31reg_gff_1_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_8019), .Z1_t (new_AGEMA_signal_8020), .Z1_f (new_AGEMA_signal_8021) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S31reg_gff_1_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_8019), .B1_t (new_AGEMA_signal_8020), .B1_f (new_AGEMA_signal_8021), .Z0_t (KeyArray_S31reg_gff_1_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_9129), .Z1_t (new_AGEMA_signal_9130), .Z1_f (new_AGEMA_signal_9131) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S31reg_gff_1_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_9129), .A1_t (new_AGEMA_signal_9130), .A1_f (new_AGEMA_signal_9131), .B0_t (KeyArray_inS31ser[4]), .B0_f (new_AGEMA_signal_7210), .B1_t (new_AGEMA_signal_7211), .B1_f (new_AGEMA_signal_7212), .Z0_t (KeyArray_S31reg_gff_1_SFF_4_QD), .Z0_f (new_AGEMA_signal_9676), .Z1_t (new_AGEMA_signal_9677), .Z1_f (new_AGEMA_signal_9678) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S31reg_gff_1_SFF_5_U3 ( .A0_t (KeyArray_S31reg_gff_1_SFF_5_n2), .A0_f (new_AGEMA_signal_10155), .A1_t (new_AGEMA_signal_10156), .A1_f (new_AGEMA_signal_10157), .B0_t (KeyArray_S31reg_gff_1_SFF_5_n1), .B0_f (new_AGEMA_signal_9132), .B1_t (new_AGEMA_signal_9133), .B1_f (new_AGEMA_signal_9134), .Z0_t (KeyArray_outS31ser[5]), .Z0_f (new_AGEMA_signal_5274), .Z1_t (new_AGEMA_signal_5275), .Z1_f (new_AGEMA_signal_5276) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_5_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS31ser[5]), .B0_f (new_AGEMA_signal_5274), .B1_t (new_AGEMA_signal_5275), .B1_f (new_AGEMA_signal_5276), .Z0_t (KeyArray_S31reg_gff_1_SFF_5_n1), .Z0_f (new_AGEMA_signal_9132), .Z1_t (new_AGEMA_signal_9133), .Z1_f (new_AGEMA_signal_9134) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_5_U1 ( .A0_t (KeyArray_S31reg_gff_1_SFF_5_QD), .A0_f (new_AGEMA_signal_9679), .A1_t (new_AGEMA_signal_9680), .A1_f (new_AGEMA_signal_9681), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S31reg_gff_1_SFF_5_n2), .Z0_f (new_AGEMA_signal_10155), .Z1_t (new_AGEMA_signal_10156), .Z1_f (new_AGEMA_signal_10157) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS31ser[5]), .A0_f (new_AGEMA_signal_7213), .A1_t (new_AGEMA_signal_7214), .A1_f (new_AGEMA_signal_7215), .B0_t (KeyArray_outS01ser_5_), .B0_f (new_AGEMA_signal_4398), .B1_t (new_AGEMA_signal_4399), .B1_f (new_AGEMA_signal_4400), .Z0_t (KeyArray_S31reg_gff_1_SFF_5_MUXInst_X), .Z0_f (new_AGEMA_signal_8022), .Z1_t (new_AGEMA_signal_8023), .Z1_f (new_AGEMA_signal_8024) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S31reg_gff_1_SFF_5_MUXInst_X), .B0_f (new_AGEMA_signal_8022), .B1_t (new_AGEMA_signal_8023), .B1_f (new_AGEMA_signal_8024), .Z0_t (KeyArray_S31reg_gff_1_SFF_5_MUXInst_Y), .Z0_f (new_AGEMA_signal_9135), .Z1_t (new_AGEMA_signal_9136), .Z1_f (new_AGEMA_signal_9137) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S31reg_gff_1_SFF_5_MUXInst_Y), .A0_f (new_AGEMA_signal_9135), .A1_t (new_AGEMA_signal_9136), .A1_f (new_AGEMA_signal_9137), .B0_t (KeyArray_inS31ser[5]), .B0_f (new_AGEMA_signal_7213), .B1_t (new_AGEMA_signal_7214), .B1_f (new_AGEMA_signal_7215), .Z0_t (KeyArray_S31reg_gff_1_SFF_5_QD), .Z0_f (new_AGEMA_signal_9679), .Z1_t (new_AGEMA_signal_9680), .Z1_f (new_AGEMA_signal_9681) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S31reg_gff_1_SFF_6_U3 ( .A0_t (KeyArray_S31reg_gff_1_SFF_6_n2), .A0_f (new_AGEMA_signal_10158), .A1_t (new_AGEMA_signal_10159), .A1_f (new_AGEMA_signal_10160), .B0_t (KeyArray_S31reg_gff_1_SFF_6_n1), .B0_f (new_AGEMA_signal_9138), .B1_t (new_AGEMA_signal_9139), .B1_f (new_AGEMA_signal_9140), .Z0_t (KeyArray_outS31ser[6]), .Z0_f (new_AGEMA_signal_5283), .Z1_t (new_AGEMA_signal_5284), .Z1_f (new_AGEMA_signal_5285) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_6_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS31ser[6]), .B0_f (new_AGEMA_signal_5283), .B1_t (new_AGEMA_signal_5284), .B1_f (new_AGEMA_signal_5285), .Z0_t (KeyArray_S31reg_gff_1_SFF_6_n1), .Z0_f (new_AGEMA_signal_9138), .Z1_t (new_AGEMA_signal_9139), .Z1_f (new_AGEMA_signal_9140) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_6_U1 ( .A0_t (KeyArray_S31reg_gff_1_SFF_6_QD), .A0_f (new_AGEMA_signal_9682), .A1_t (new_AGEMA_signal_9683), .A1_f (new_AGEMA_signal_9684), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S31reg_gff_1_SFF_6_n2), .Z0_f (new_AGEMA_signal_10158), .Z1_t (new_AGEMA_signal_10159), .Z1_f (new_AGEMA_signal_10160) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS31ser[6]), .A0_f (new_AGEMA_signal_7216), .A1_t (new_AGEMA_signal_7217), .A1_f (new_AGEMA_signal_7218), .B0_t (KeyArray_outS01ser_6_), .B0_f (new_AGEMA_signal_4392), .B1_t (new_AGEMA_signal_4393), .B1_f (new_AGEMA_signal_4394), .Z0_t (KeyArray_S31reg_gff_1_SFF_6_MUXInst_X), .Z0_f (new_AGEMA_signal_8025), .Z1_t (new_AGEMA_signal_8026), .Z1_f (new_AGEMA_signal_8027) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S31reg_gff_1_SFF_6_MUXInst_X), .B0_f (new_AGEMA_signal_8025), .B1_t (new_AGEMA_signal_8026), .B1_f (new_AGEMA_signal_8027), .Z0_t (KeyArray_S31reg_gff_1_SFF_6_MUXInst_Y), .Z0_f (new_AGEMA_signal_9141), .Z1_t (new_AGEMA_signal_9142), .Z1_f (new_AGEMA_signal_9143) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S31reg_gff_1_SFF_6_MUXInst_Y), .A0_f (new_AGEMA_signal_9141), .A1_t (new_AGEMA_signal_9142), .A1_f (new_AGEMA_signal_9143), .B0_t (KeyArray_inS31ser[6]), .B0_f (new_AGEMA_signal_7216), .B1_t (new_AGEMA_signal_7217), .B1_f (new_AGEMA_signal_7218), .Z0_t (KeyArray_S31reg_gff_1_SFF_6_QD), .Z0_f (new_AGEMA_signal_9682), .Z1_t (new_AGEMA_signal_9683), .Z1_f (new_AGEMA_signal_9684) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S31reg_gff_1_SFF_7_U3 ( .A0_t (KeyArray_S31reg_gff_1_SFF_7_n2), .A0_f (new_AGEMA_signal_10161), .A1_t (new_AGEMA_signal_10162), .A1_f (new_AGEMA_signal_10163), .B0_t (KeyArray_S31reg_gff_1_SFF_7_n1), .B0_f (new_AGEMA_signal_9144), .B1_t (new_AGEMA_signal_9145), .B1_f (new_AGEMA_signal_9146), .Z0_t (KeyArray_outS31ser[7]), .Z0_f (new_AGEMA_signal_5292), .Z1_t (new_AGEMA_signal_5293), .Z1_f (new_AGEMA_signal_5294) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_7_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS31ser[7]), .B0_f (new_AGEMA_signal_5292), .B1_t (new_AGEMA_signal_5293), .B1_f (new_AGEMA_signal_5294), .Z0_t (KeyArray_S31reg_gff_1_SFF_7_n1), .Z0_f (new_AGEMA_signal_9144), .Z1_t (new_AGEMA_signal_9145), .Z1_f (new_AGEMA_signal_9146) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_7_U1 ( .A0_t (KeyArray_S31reg_gff_1_SFF_7_QD), .A0_f (new_AGEMA_signal_9685), .A1_t (new_AGEMA_signal_9686), .A1_f (new_AGEMA_signal_9687), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S31reg_gff_1_SFF_7_n2), .Z0_f (new_AGEMA_signal_10161), .Z1_t (new_AGEMA_signal_10162), .Z1_f (new_AGEMA_signal_10163) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS31ser[7]), .A0_f (new_AGEMA_signal_7219), .A1_t (new_AGEMA_signal_7220), .A1_f (new_AGEMA_signal_7221), .B0_t (KeyArray_outS01ser_7_), .B0_f (new_AGEMA_signal_4386), .B1_t (new_AGEMA_signal_4387), .B1_f (new_AGEMA_signal_4388), .Z0_t (KeyArray_S31reg_gff_1_SFF_7_MUXInst_X), .Z0_f (new_AGEMA_signal_8028), .Z1_t (new_AGEMA_signal_8029), .Z1_f (new_AGEMA_signal_8030) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S31reg_gff_1_SFF_7_MUXInst_X), .B0_f (new_AGEMA_signal_8028), .B1_t (new_AGEMA_signal_8029), .B1_f (new_AGEMA_signal_8030), .Z0_t (KeyArray_S31reg_gff_1_SFF_7_MUXInst_Y), .Z0_f (new_AGEMA_signal_9147), .Z1_t (new_AGEMA_signal_9148), .Z1_f (new_AGEMA_signal_9149) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S31reg_gff_1_SFF_7_MUXInst_Y), .A0_f (new_AGEMA_signal_9147), .A1_t (new_AGEMA_signal_9148), .A1_f (new_AGEMA_signal_9149), .B0_t (KeyArray_inS31ser[7]), .B0_f (new_AGEMA_signal_7219), .B1_t (new_AGEMA_signal_7220), .B1_f (new_AGEMA_signal_7221), .Z0_t (KeyArray_S31reg_gff_1_SFF_7_QD), .Z0_f (new_AGEMA_signal_9685), .Z1_t (new_AGEMA_signal_9686), .Z1_f (new_AGEMA_signal_9687) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S32reg_gff_1_SFF_0_U3 ( .A0_t (KeyArray_S32reg_gff_1_SFF_0_n2), .A0_f (new_AGEMA_signal_10164), .A1_t (new_AGEMA_signal_10165), .A1_f (new_AGEMA_signal_10166), .B0_t (KeyArray_S32reg_gff_1_SFF_0_n1), .B0_f (new_AGEMA_signal_9150), .B1_t (new_AGEMA_signal_9151), .B1_f (new_AGEMA_signal_9152), .Z0_t (KeyArray_outS32ser[0]), .Z0_f (new_AGEMA_signal_5301), .Z1_t (new_AGEMA_signal_5302), .Z1_f (new_AGEMA_signal_5303) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_0_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS32ser[0]), .B0_f (new_AGEMA_signal_5301), .B1_t (new_AGEMA_signal_5302), .B1_f (new_AGEMA_signal_5303), .Z0_t (KeyArray_S32reg_gff_1_SFF_0_n1), .Z0_f (new_AGEMA_signal_9150), .Z1_t (new_AGEMA_signal_9151), .Z1_f (new_AGEMA_signal_9152) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_0_U1 ( .A0_t (KeyArray_S32reg_gff_1_SFF_0_QD), .A0_f (new_AGEMA_signal_9688), .A1_t (new_AGEMA_signal_9689), .A1_f (new_AGEMA_signal_9690), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S32reg_gff_1_SFF_0_n2), .Z0_f (new_AGEMA_signal_10164), .Z1_t (new_AGEMA_signal_10165), .Z1_f (new_AGEMA_signal_10166) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS32ser[0]), .A0_f (new_AGEMA_signal_7222), .A1_t (new_AGEMA_signal_7223), .A1_f (new_AGEMA_signal_7224), .B0_t (KeyArray_outS02ser[0]), .B0_f (new_AGEMA_signal_4437), .B1_t (new_AGEMA_signal_4438), .B1_f (new_AGEMA_signal_4439), .Z0_t (KeyArray_S32reg_gff_1_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_8031), .Z1_t (new_AGEMA_signal_8032), .Z1_f (new_AGEMA_signal_8033) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S32reg_gff_1_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_8031), .B1_t (new_AGEMA_signal_8032), .B1_f (new_AGEMA_signal_8033), .Z0_t (KeyArray_S32reg_gff_1_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_9153), .Z1_t (new_AGEMA_signal_9154), .Z1_f (new_AGEMA_signal_9155) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S32reg_gff_1_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_9153), .A1_t (new_AGEMA_signal_9154), .A1_f (new_AGEMA_signal_9155), .B0_t (KeyArray_inS32ser[0]), .B0_f (new_AGEMA_signal_7222), .B1_t (new_AGEMA_signal_7223), .B1_f (new_AGEMA_signal_7224), .Z0_t (KeyArray_S32reg_gff_1_SFF_0_QD), .Z0_f (new_AGEMA_signal_9688), .Z1_t (new_AGEMA_signal_9689), .Z1_f (new_AGEMA_signal_9690) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S32reg_gff_1_SFF_1_U3 ( .A0_t (KeyArray_S32reg_gff_1_SFF_1_n2), .A0_f (new_AGEMA_signal_10167), .A1_t (new_AGEMA_signal_10168), .A1_f (new_AGEMA_signal_10169), .B0_t (KeyArray_S32reg_gff_1_SFF_1_n1), .B0_f (new_AGEMA_signal_9156), .B1_t (new_AGEMA_signal_9157), .B1_f (new_AGEMA_signal_9158), .Z0_t (KeyArray_outS32ser[1]), .Z0_f (new_AGEMA_signal_5310), .Z1_t (new_AGEMA_signal_5311), .Z1_f (new_AGEMA_signal_5312) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_1_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS32ser[1]), .B0_f (new_AGEMA_signal_5310), .B1_t (new_AGEMA_signal_5311), .B1_f (new_AGEMA_signal_5312), .Z0_t (KeyArray_S32reg_gff_1_SFF_1_n1), .Z0_f (new_AGEMA_signal_9156), .Z1_t (new_AGEMA_signal_9157), .Z1_f (new_AGEMA_signal_9158) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_1_U1 ( .A0_t (KeyArray_S32reg_gff_1_SFF_1_QD), .A0_f (new_AGEMA_signal_9691), .A1_t (new_AGEMA_signal_9692), .A1_f (new_AGEMA_signal_9693), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S32reg_gff_1_SFF_1_n2), .Z0_f (new_AGEMA_signal_10167), .Z1_t (new_AGEMA_signal_10168), .Z1_f (new_AGEMA_signal_10169) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS32ser[1]), .A0_f (new_AGEMA_signal_7225), .A1_t (new_AGEMA_signal_7226), .A1_f (new_AGEMA_signal_7227), .B0_t (KeyArray_outS02ser[1]), .B0_f (new_AGEMA_signal_4446), .B1_t (new_AGEMA_signal_4447), .B1_f (new_AGEMA_signal_4448), .Z0_t (KeyArray_S32reg_gff_1_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_8034), .Z1_t (new_AGEMA_signal_8035), .Z1_f (new_AGEMA_signal_8036) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S32reg_gff_1_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_8034), .B1_t (new_AGEMA_signal_8035), .B1_f (new_AGEMA_signal_8036), .Z0_t (KeyArray_S32reg_gff_1_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_9159), .Z1_t (new_AGEMA_signal_9160), .Z1_f (new_AGEMA_signal_9161) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S32reg_gff_1_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_9159), .A1_t (new_AGEMA_signal_9160), .A1_f (new_AGEMA_signal_9161), .B0_t (KeyArray_inS32ser[1]), .B0_f (new_AGEMA_signal_7225), .B1_t (new_AGEMA_signal_7226), .B1_f (new_AGEMA_signal_7227), .Z0_t (KeyArray_S32reg_gff_1_SFF_1_QD), .Z0_f (new_AGEMA_signal_9691), .Z1_t (new_AGEMA_signal_9692), .Z1_f (new_AGEMA_signal_9693) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S32reg_gff_1_SFF_2_U3 ( .A0_t (KeyArray_S32reg_gff_1_SFF_2_n2), .A0_f (new_AGEMA_signal_10170), .A1_t (new_AGEMA_signal_10171), .A1_f (new_AGEMA_signal_10172), .B0_t (KeyArray_S32reg_gff_1_SFF_2_n1), .B0_f (new_AGEMA_signal_9162), .B1_t (new_AGEMA_signal_9163), .B1_f (new_AGEMA_signal_9164), .Z0_t (KeyArray_outS32ser[2]), .Z0_f (new_AGEMA_signal_5319), .Z1_t (new_AGEMA_signal_5320), .Z1_f (new_AGEMA_signal_5321) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_2_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS32ser[2]), .B0_f (new_AGEMA_signal_5319), .B1_t (new_AGEMA_signal_5320), .B1_f (new_AGEMA_signal_5321), .Z0_t (KeyArray_S32reg_gff_1_SFF_2_n1), .Z0_f (new_AGEMA_signal_9162), .Z1_t (new_AGEMA_signal_9163), .Z1_f (new_AGEMA_signal_9164) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_2_U1 ( .A0_t (KeyArray_S32reg_gff_1_SFF_2_QD), .A0_f (new_AGEMA_signal_9694), .A1_t (new_AGEMA_signal_9695), .A1_f (new_AGEMA_signal_9696), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S32reg_gff_1_SFF_2_n2), .Z0_f (new_AGEMA_signal_10170), .Z1_t (new_AGEMA_signal_10171), .Z1_f (new_AGEMA_signal_10172) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS32ser[2]), .A0_f (new_AGEMA_signal_7228), .A1_t (new_AGEMA_signal_7229), .A1_f (new_AGEMA_signal_7230), .B0_t (KeyArray_outS02ser[2]), .B0_f (new_AGEMA_signal_4455), .B1_t (new_AGEMA_signal_4456), .B1_f (new_AGEMA_signal_4457), .Z0_t (KeyArray_S32reg_gff_1_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_8037), .Z1_t (new_AGEMA_signal_8038), .Z1_f (new_AGEMA_signal_8039) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S32reg_gff_1_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_8037), .B1_t (new_AGEMA_signal_8038), .B1_f (new_AGEMA_signal_8039), .Z0_t (KeyArray_S32reg_gff_1_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_9165), .Z1_t (new_AGEMA_signal_9166), .Z1_f (new_AGEMA_signal_9167) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S32reg_gff_1_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_9165), .A1_t (new_AGEMA_signal_9166), .A1_f (new_AGEMA_signal_9167), .B0_t (KeyArray_inS32ser[2]), .B0_f (new_AGEMA_signal_7228), .B1_t (new_AGEMA_signal_7229), .B1_f (new_AGEMA_signal_7230), .Z0_t (KeyArray_S32reg_gff_1_SFF_2_QD), .Z0_f (new_AGEMA_signal_9694), .Z1_t (new_AGEMA_signal_9695), .Z1_f (new_AGEMA_signal_9696) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S32reg_gff_1_SFF_3_U3 ( .A0_t (KeyArray_S32reg_gff_1_SFF_3_n2), .A0_f (new_AGEMA_signal_10173), .A1_t (new_AGEMA_signal_10174), .A1_f (new_AGEMA_signal_10175), .B0_t (KeyArray_S32reg_gff_1_SFF_3_n1), .B0_f (new_AGEMA_signal_9168), .B1_t (new_AGEMA_signal_9169), .B1_f (new_AGEMA_signal_9170), .Z0_t (KeyArray_outS32ser[3]), .Z0_f (new_AGEMA_signal_5328), .Z1_t (new_AGEMA_signal_5329), .Z1_f (new_AGEMA_signal_5330) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_3_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS32ser[3]), .B0_f (new_AGEMA_signal_5328), .B1_t (new_AGEMA_signal_5329), .B1_f (new_AGEMA_signal_5330), .Z0_t (KeyArray_S32reg_gff_1_SFF_3_n1), .Z0_f (new_AGEMA_signal_9168), .Z1_t (new_AGEMA_signal_9169), .Z1_f (new_AGEMA_signal_9170) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_3_U1 ( .A0_t (KeyArray_S32reg_gff_1_SFF_3_QD), .A0_f (new_AGEMA_signal_9697), .A1_t (new_AGEMA_signal_9698), .A1_f (new_AGEMA_signal_9699), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S32reg_gff_1_SFF_3_n2), .Z0_f (new_AGEMA_signal_10173), .Z1_t (new_AGEMA_signal_10174), .Z1_f (new_AGEMA_signal_10175) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS32ser[3]), .A0_f (new_AGEMA_signal_7231), .A1_t (new_AGEMA_signal_7232), .A1_f (new_AGEMA_signal_7233), .B0_t (KeyArray_outS02ser[3]), .B0_f (new_AGEMA_signal_4464), .B1_t (new_AGEMA_signal_4465), .B1_f (new_AGEMA_signal_4466), .Z0_t (KeyArray_S32reg_gff_1_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_8040), .Z1_t (new_AGEMA_signal_8041), .Z1_f (new_AGEMA_signal_8042) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S32reg_gff_1_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_8040), .B1_t (new_AGEMA_signal_8041), .B1_f (new_AGEMA_signal_8042), .Z0_t (KeyArray_S32reg_gff_1_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_9171), .Z1_t (new_AGEMA_signal_9172), .Z1_f (new_AGEMA_signal_9173) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S32reg_gff_1_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_9171), .A1_t (new_AGEMA_signal_9172), .A1_f (new_AGEMA_signal_9173), .B0_t (KeyArray_inS32ser[3]), .B0_f (new_AGEMA_signal_7231), .B1_t (new_AGEMA_signal_7232), .B1_f (new_AGEMA_signal_7233), .Z0_t (KeyArray_S32reg_gff_1_SFF_3_QD), .Z0_f (new_AGEMA_signal_9697), .Z1_t (new_AGEMA_signal_9698), .Z1_f (new_AGEMA_signal_9699) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S32reg_gff_1_SFF_4_U3 ( .A0_t (KeyArray_S32reg_gff_1_SFF_4_n2), .A0_f (new_AGEMA_signal_10176), .A1_t (new_AGEMA_signal_10177), .A1_f (new_AGEMA_signal_10178), .B0_t (KeyArray_S32reg_gff_1_SFF_4_n1), .B0_f (new_AGEMA_signal_9174), .B1_t (new_AGEMA_signal_9175), .B1_f (new_AGEMA_signal_9176), .Z0_t (KeyArray_outS32ser[4]), .Z0_f (new_AGEMA_signal_5337), .Z1_t (new_AGEMA_signal_5338), .Z1_f (new_AGEMA_signal_5339) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_4_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS32ser[4]), .B0_f (new_AGEMA_signal_5337), .B1_t (new_AGEMA_signal_5338), .B1_f (new_AGEMA_signal_5339), .Z0_t (KeyArray_S32reg_gff_1_SFF_4_n1), .Z0_f (new_AGEMA_signal_9174), .Z1_t (new_AGEMA_signal_9175), .Z1_f (new_AGEMA_signal_9176) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_4_U1 ( .A0_t (KeyArray_S32reg_gff_1_SFF_4_QD), .A0_f (new_AGEMA_signal_9700), .A1_t (new_AGEMA_signal_9701), .A1_f (new_AGEMA_signal_9702), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S32reg_gff_1_SFF_4_n2), .Z0_f (new_AGEMA_signal_10176), .Z1_t (new_AGEMA_signal_10177), .Z1_f (new_AGEMA_signal_10178) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS32ser[4]), .A0_f (new_AGEMA_signal_7234), .A1_t (new_AGEMA_signal_7235), .A1_f (new_AGEMA_signal_7236), .B0_t (KeyArray_outS02ser[4]), .B0_f (new_AGEMA_signal_4473), .B1_t (new_AGEMA_signal_4474), .B1_f (new_AGEMA_signal_4475), .Z0_t (KeyArray_S32reg_gff_1_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_8043), .Z1_t (new_AGEMA_signal_8044), .Z1_f (new_AGEMA_signal_8045) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S32reg_gff_1_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_8043), .B1_t (new_AGEMA_signal_8044), .B1_f (new_AGEMA_signal_8045), .Z0_t (KeyArray_S32reg_gff_1_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_9177), .Z1_t (new_AGEMA_signal_9178), .Z1_f (new_AGEMA_signal_9179) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S32reg_gff_1_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_9177), .A1_t (new_AGEMA_signal_9178), .A1_f (new_AGEMA_signal_9179), .B0_t (KeyArray_inS32ser[4]), .B0_f (new_AGEMA_signal_7234), .B1_t (new_AGEMA_signal_7235), .B1_f (new_AGEMA_signal_7236), .Z0_t (KeyArray_S32reg_gff_1_SFF_4_QD), .Z0_f (new_AGEMA_signal_9700), .Z1_t (new_AGEMA_signal_9701), .Z1_f (new_AGEMA_signal_9702) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S32reg_gff_1_SFF_5_U3 ( .A0_t (KeyArray_S32reg_gff_1_SFF_5_n2), .A0_f (new_AGEMA_signal_10179), .A1_t (new_AGEMA_signal_10180), .A1_f (new_AGEMA_signal_10181), .B0_t (KeyArray_S32reg_gff_1_SFF_5_n1), .B0_f (new_AGEMA_signal_9180), .B1_t (new_AGEMA_signal_9181), .B1_f (new_AGEMA_signal_9182), .Z0_t (KeyArray_outS32ser[5]), .Z0_f (new_AGEMA_signal_5346), .Z1_t (new_AGEMA_signal_5347), .Z1_f (new_AGEMA_signal_5348) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_5_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS32ser[5]), .B0_f (new_AGEMA_signal_5346), .B1_t (new_AGEMA_signal_5347), .B1_f (new_AGEMA_signal_5348), .Z0_t (KeyArray_S32reg_gff_1_SFF_5_n1), .Z0_f (new_AGEMA_signal_9180), .Z1_t (new_AGEMA_signal_9181), .Z1_f (new_AGEMA_signal_9182) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_5_U1 ( .A0_t (KeyArray_S32reg_gff_1_SFF_5_QD), .A0_f (new_AGEMA_signal_9703), .A1_t (new_AGEMA_signal_9704), .A1_f (new_AGEMA_signal_9705), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S32reg_gff_1_SFF_5_n2), .Z0_f (new_AGEMA_signal_10179), .Z1_t (new_AGEMA_signal_10180), .Z1_f (new_AGEMA_signal_10181) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS32ser[5]), .A0_f (new_AGEMA_signal_7237), .A1_t (new_AGEMA_signal_7238), .A1_f (new_AGEMA_signal_7239), .B0_t (KeyArray_outS02ser[5]), .B0_f (new_AGEMA_signal_4482), .B1_t (new_AGEMA_signal_4483), .B1_f (new_AGEMA_signal_4484), .Z0_t (KeyArray_S32reg_gff_1_SFF_5_MUXInst_X), .Z0_f (new_AGEMA_signal_8046), .Z1_t (new_AGEMA_signal_8047), .Z1_f (new_AGEMA_signal_8048) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S32reg_gff_1_SFF_5_MUXInst_X), .B0_f (new_AGEMA_signal_8046), .B1_t (new_AGEMA_signal_8047), .B1_f (new_AGEMA_signal_8048), .Z0_t (KeyArray_S32reg_gff_1_SFF_5_MUXInst_Y), .Z0_f (new_AGEMA_signal_9183), .Z1_t (new_AGEMA_signal_9184), .Z1_f (new_AGEMA_signal_9185) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S32reg_gff_1_SFF_5_MUXInst_Y), .A0_f (new_AGEMA_signal_9183), .A1_t (new_AGEMA_signal_9184), .A1_f (new_AGEMA_signal_9185), .B0_t (KeyArray_inS32ser[5]), .B0_f (new_AGEMA_signal_7237), .B1_t (new_AGEMA_signal_7238), .B1_f (new_AGEMA_signal_7239), .Z0_t (KeyArray_S32reg_gff_1_SFF_5_QD), .Z0_f (new_AGEMA_signal_9703), .Z1_t (new_AGEMA_signal_9704), .Z1_f (new_AGEMA_signal_9705) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S32reg_gff_1_SFF_6_U3 ( .A0_t (KeyArray_S32reg_gff_1_SFF_6_n2), .A0_f (new_AGEMA_signal_10182), .A1_t (new_AGEMA_signal_10183), .A1_f (new_AGEMA_signal_10184), .B0_t (KeyArray_S32reg_gff_1_SFF_6_n1), .B0_f (new_AGEMA_signal_9186), .B1_t (new_AGEMA_signal_9187), .B1_f (new_AGEMA_signal_9188), .Z0_t (KeyArray_outS32ser[6]), .Z0_f (new_AGEMA_signal_5355), .Z1_t (new_AGEMA_signal_5356), .Z1_f (new_AGEMA_signal_5357) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_6_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS32ser[6]), .B0_f (new_AGEMA_signal_5355), .B1_t (new_AGEMA_signal_5356), .B1_f (new_AGEMA_signal_5357), .Z0_t (KeyArray_S32reg_gff_1_SFF_6_n1), .Z0_f (new_AGEMA_signal_9186), .Z1_t (new_AGEMA_signal_9187), .Z1_f (new_AGEMA_signal_9188) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_6_U1 ( .A0_t (KeyArray_S32reg_gff_1_SFF_6_QD), .A0_f (new_AGEMA_signal_9706), .A1_t (new_AGEMA_signal_9707), .A1_f (new_AGEMA_signal_9708), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S32reg_gff_1_SFF_6_n2), .Z0_f (new_AGEMA_signal_10182), .Z1_t (new_AGEMA_signal_10183), .Z1_f (new_AGEMA_signal_10184) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS32ser[6]), .A0_f (new_AGEMA_signal_7240), .A1_t (new_AGEMA_signal_7241), .A1_f (new_AGEMA_signal_7242), .B0_t (KeyArray_outS02ser[6]), .B0_f (new_AGEMA_signal_4491), .B1_t (new_AGEMA_signal_4492), .B1_f (new_AGEMA_signal_4493), .Z0_t (KeyArray_S32reg_gff_1_SFF_6_MUXInst_X), .Z0_f (new_AGEMA_signal_8049), .Z1_t (new_AGEMA_signal_8050), .Z1_f (new_AGEMA_signal_8051) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S32reg_gff_1_SFF_6_MUXInst_X), .B0_f (new_AGEMA_signal_8049), .B1_t (new_AGEMA_signal_8050), .B1_f (new_AGEMA_signal_8051), .Z0_t (KeyArray_S32reg_gff_1_SFF_6_MUXInst_Y), .Z0_f (new_AGEMA_signal_9189), .Z1_t (new_AGEMA_signal_9190), .Z1_f (new_AGEMA_signal_9191) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S32reg_gff_1_SFF_6_MUXInst_Y), .A0_f (new_AGEMA_signal_9189), .A1_t (new_AGEMA_signal_9190), .A1_f (new_AGEMA_signal_9191), .B0_t (KeyArray_inS32ser[6]), .B0_f (new_AGEMA_signal_7240), .B1_t (new_AGEMA_signal_7241), .B1_f (new_AGEMA_signal_7242), .Z0_t (KeyArray_S32reg_gff_1_SFF_6_QD), .Z0_f (new_AGEMA_signal_9706), .Z1_t (new_AGEMA_signal_9707), .Z1_f (new_AGEMA_signal_9708) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S32reg_gff_1_SFF_7_U3 ( .A0_t (KeyArray_S32reg_gff_1_SFF_7_n2), .A0_f (new_AGEMA_signal_10185), .A1_t (new_AGEMA_signal_10186), .A1_f (new_AGEMA_signal_10187), .B0_t (KeyArray_S32reg_gff_1_SFF_7_n1), .B0_f (new_AGEMA_signal_9192), .B1_t (new_AGEMA_signal_9193), .B1_f (new_AGEMA_signal_9194), .Z0_t (KeyArray_outS32ser[7]), .Z0_f (new_AGEMA_signal_5364), .Z1_t (new_AGEMA_signal_5365), .Z1_f (new_AGEMA_signal_5366) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_7_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS32ser[7]), .B0_f (new_AGEMA_signal_5364), .B1_t (new_AGEMA_signal_5365), .B1_f (new_AGEMA_signal_5366), .Z0_t (KeyArray_S32reg_gff_1_SFF_7_n1), .Z0_f (new_AGEMA_signal_9192), .Z1_t (new_AGEMA_signal_9193), .Z1_f (new_AGEMA_signal_9194) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_7_U1 ( .A0_t (KeyArray_S32reg_gff_1_SFF_7_QD), .A0_f (new_AGEMA_signal_9709), .A1_t (new_AGEMA_signal_9710), .A1_f (new_AGEMA_signal_9711), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S32reg_gff_1_SFF_7_n2), .Z0_f (new_AGEMA_signal_10185), .Z1_t (new_AGEMA_signal_10186), .Z1_f (new_AGEMA_signal_10187) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS32ser[7]), .A0_f (new_AGEMA_signal_7243), .A1_t (new_AGEMA_signal_7244), .A1_f (new_AGEMA_signal_7245), .B0_t (KeyArray_outS02ser[7]), .B0_f (new_AGEMA_signal_4500), .B1_t (new_AGEMA_signal_4501), .B1_f (new_AGEMA_signal_4502), .Z0_t (KeyArray_S32reg_gff_1_SFF_7_MUXInst_X), .Z0_f (new_AGEMA_signal_8052), .Z1_t (new_AGEMA_signal_8053), .Z1_f (new_AGEMA_signal_8054) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S32reg_gff_1_SFF_7_MUXInst_X), .B0_f (new_AGEMA_signal_8052), .B1_t (new_AGEMA_signal_8053), .B1_f (new_AGEMA_signal_8054), .Z0_t (KeyArray_S32reg_gff_1_SFF_7_MUXInst_Y), .Z0_f (new_AGEMA_signal_9195), .Z1_t (new_AGEMA_signal_9196), .Z1_f (new_AGEMA_signal_9197) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S32reg_gff_1_SFF_7_MUXInst_Y), .A0_f (new_AGEMA_signal_9195), .A1_t (new_AGEMA_signal_9196), .A1_f (new_AGEMA_signal_9197), .B0_t (KeyArray_inS32ser[7]), .B0_f (new_AGEMA_signal_7243), .B1_t (new_AGEMA_signal_7244), .B1_f (new_AGEMA_signal_7245), .Z0_t (KeyArray_S32reg_gff_1_SFF_7_QD), .Z0_f (new_AGEMA_signal_9709), .Z1_t (new_AGEMA_signal_9710), .Z1_f (new_AGEMA_signal_9711) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S33reg_gff_1_SFF_0_U3 ( .A0_t (KeyArray_S33reg_gff_1_SFF_0_n2), .A0_f (new_AGEMA_signal_10188), .A1_t (new_AGEMA_signal_10189), .A1_f (new_AGEMA_signal_10190), .B0_t (KeyArray_S33reg_gff_1_SFF_0_n1), .B0_f (new_AGEMA_signal_9198), .B1_t (new_AGEMA_signal_9199), .B1_f (new_AGEMA_signal_9200), .Z0_t (KeyArray_outS33ser[0]), .Z0_f (new_AGEMA_signal_5373), .Z1_t (new_AGEMA_signal_5374), .Z1_f (new_AGEMA_signal_5375) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_0_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS33ser[0]), .B0_f (new_AGEMA_signal_5373), .B1_t (new_AGEMA_signal_5374), .B1_f (new_AGEMA_signal_5375), .Z0_t (KeyArray_S33reg_gff_1_SFF_0_n1), .Z0_f (new_AGEMA_signal_9198), .Z1_t (new_AGEMA_signal_9199), .Z1_f (new_AGEMA_signal_9200) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_0_U1 ( .A0_t (KeyArray_S33reg_gff_1_SFF_0_QD), .A0_f (new_AGEMA_signal_9712), .A1_t (new_AGEMA_signal_9713), .A1_f (new_AGEMA_signal_9714), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S33reg_gff_1_SFF_0_n2), .Z0_f (new_AGEMA_signal_10188), .Z1_t (new_AGEMA_signal_10189), .Z1_f (new_AGEMA_signal_10190) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS33ser[0]), .A0_f (new_AGEMA_signal_7246), .A1_t (new_AGEMA_signal_7247), .A1_f (new_AGEMA_signal_7248), .B0_t (KeyArray_outS03ser[0]), .B0_f (new_AGEMA_signal_4509), .B1_t (new_AGEMA_signal_4510), .B1_f (new_AGEMA_signal_4511), .Z0_t (KeyArray_S33reg_gff_1_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_8055), .Z1_t (new_AGEMA_signal_8056), .Z1_f (new_AGEMA_signal_8057) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S33reg_gff_1_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_8055), .B1_t (new_AGEMA_signal_8056), .B1_f (new_AGEMA_signal_8057), .Z0_t (KeyArray_S33reg_gff_1_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_9201), .Z1_t (new_AGEMA_signal_9202), .Z1_f (new_AGEMA_signal_9203) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S33reg_gff_1_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_9201), .A1_t (new_AGEMA_signal_9202), .A1_f (new_AGEMA_signal_9203), .B0_t (KeyArray_inS33ser[0]), .B0_f (new_AGEMA_signal_7246), .B1_t (new_AGEMA_signal_7247), .B1_f (new_AGEMA_signal_7248), .Z0_t (KeyArray_S33reg_gff_1_SFF_0_QD), .Z0_f (new_AGEMA_signal_9712), .Z1_t (new_AGEMA_signal_9713), .Z1_f (new_AGEMA_signal_9714) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S33reg_gff_1_SFF_1_U3 ( .A0_t (KeyArray_S33reg_gff_1_SFF_1_n2), .A0_f (new_AGEMA_signal_10191), .A1_t (new_AGEMA_signal_10192), .A1_f (new_AGEMA_signal_10193), .B0_t (KeyArray_S33reg_gff_1_SFF_1_n1), .B0_f (new_AGEMA_signal_9204), .B1_t (new_AGEMA_signal_9205), .B1_f (new_AGEMA_signal_9206), .Z0_t (KeyArray_outS33ser[1]), .Z0_f (new_AGEMA_signal_5382), .Z1_t (new_AGEMA_signal_5383), .Z1_f (new_AGEMA_signal_5384) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_1_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS33ser[1]), .B0_f (new_AGEMA_signal_5382), .B1_t (new_AGEMA_signal_5383), .B1_f (new_AGEMA_signal_5384), .Z0_t (KeyArray_S33reg_gff_1_SFF_1_n1), .Z0_f (new_AGEMA_signal_9204), .Z1_t (new_AGEMA_signal_9205), .Z1_f (new_AGEMA_signal_9206) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_1_U1 ( .A0_t (KeyArray_S33reg_gff_1_SFF_1_QD), .A0_f (new_AGEMA_signal_9715), .A1_t (new_AGEMA_signal_9716), .A1_f (new_AGEMA_signal_9717), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S33reg_gff_1_SFF_1_n2), .Z0_f (new_AGEMA_signal_10191), .Z1_t (new_AGEMA_signal_10192), .Z1_f (new_AGEMA_signal_10193) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS33ser[1]), .A0_f (new_AGEMA_signal_7249), .A1_t (new_AGEMA_signal_7250), .A1_f (new_AGEMA_signal_7251), .B0_t (KeyArray_outS03ser[1]), .B0_f (new_AGEMA_signal_4518), .B1_t (new_AGEMA_signal_4519), .B1_f (new_AGEMA_signal_4520), .Z0_t (KeyArray_S33reg_gff_1_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_8058), .Z1_t (new_AGEMA_signal_8059), .Z1_f (new_AGEMA_signal_8060) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S33reg_gff_1_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_8058), .B1_t (new_AGEMA_signal_8059), .B1_f (new_AGEMA_signal_8060), .Z0_t (KeyArray_S33reg_gff_1_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_9207), .Z1_t (new_AGEMA_signal_9208), .Z1_f (new_AGEMA_signal_9209) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S33reg_gff_1_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_9207), .A1_t (new_AGEMA_signal_9208), .A1_f (new_AGEMA_signal_9209), .B0_t (KeyArray_inS33ser[1]), .B0_f (new_AGEMA_signal_7249), .B1_t (new_AGEMA_signal_7250), .B1_f (new_AGEMA_signal_7251), .Z0_t (KeyArray_S33reg_gff_1_SFF_1_QD), .Z0_f (new_AGEMA_signal_9715), .Z1_t (new_AGEMA_signal_9716), .Z1_f (new_AGEMA_signal_9717) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S33reg_gff_1_SFF_2_U3 ( .A0_t (KeyArray_S33reg_gff_1_SFF_2_n2), .A0_f (new_AGEMA_signal_10194), .A1_t (new_AGEMA_signal_10195), .A1_f (new_AGEMA_signal_10196), .B0_t (KeyArray_S33reg_gff_1_SFF_2_n1), .B0_f (new_AGEMA_signal_9210), .B1_t (new_AGEMA_signal_9211), .B1_f (new_AGEMA_signal_9212), .Z0_t (KeyArray_outS33ser[2]), .Z0_f (new_AGEMA_signal_5391), .Z1_t (new_AGEMA_signal_5392), .Z1_f (new_AGEMA_signal_5393) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_2_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS33ser[2]), .B0_f (new_AGEMA_signal_5391), .B1_t (new_AGEMA_signal_5392), .B1_f (new_AGEMA_signal_5393), .Z0_t (KeyArray_S33reg_gff_1_SFF_2_n1), .Z0_f (new_AGEMA_signal_9210), .Z1_t (new_AGEMA_signal_9211), .Z1_f (new_AGEMA_signal_9212) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_2_U1 ( .A0_t (KeyArray_S33reg_gff_1_SFF_2_QD), .A0_f (new_AGEMA_signal_9718), .A1_t (new_AGEMA_signal_9719), .A1_f (new_AGEMA_signal_9720), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S33reg_gff_1_SFF_2_n2), .Z0_f (new_AGEMA_signal_10194), .Z1_t (new_AGEMA_signal_10195), .Z1_f (new_AGEMA_signal_10196) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS33ser[2]), .A0_f (new_AGEMA_signal_7252), .A1_t (new_AGEMA_signal_7253), .A1_f (new_AGEMA_signal_7254), .B0_t (KeyArray_outS03ser[2]), .B0_f (new_AGEMA_signal_4527), .B1_t (new_AGEMA_signal_4528), .B1_f (new_AGEMA_signal_4529), .Z0_t (KeyArray_S33reg_gff_1_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_8061), .Z1_t (new_AGEMA_signal_8062), .Z1_f (new_AGEMA_signal_8063) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S33reg_gff_1_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_8061), .B1_t (new_AGEMA_signal_8062), .B1_f (new_AGEMA_signal_8063), .Z0_t (KeyArray_S33reg_gff_1_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_9213), .Z1_t (new_AGEMA_signal_9214), .Z1_f (new_AGEMA_signal_9215) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S33reg_gff_1_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_9213), .A1_t (new_AGEMA_signal_9214), .A1_f (new_AGEMA_signal_9215), .B0_t (KeyArray_inS33ser[2]), .B0_f (new_AGEMA_signal_7252), .B1_t (new_AGEMA_signal_7253), .B1_f (new_AGEMA_signal_7254), .Z0_t (KeyArray_S33reg_gff_1_SFF_2_QD), .Z0_f (new_AGEMA_signal_9718), .Z1_t (new_AGEMA_signal_9719), .Z1_f (new_AGEMA_signal_9720) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S33reg_gff_1_SFF_3_U3 ( .A0_t (KeyArray_S33reg_gff_1_SFF_3_n2), .A0_f (new_AGEMA_signal_10197), .A1_t (new_AGEMA_signal_10198), .A1_f (new_AGEMA_signal_10199), .B0_t (KeyArray_S33reg_gff_1_SFF_3_n1), .B0_f (new_AGEMA_signal_9216), .B1_t (new_AGEMA_signal_9217), .B1_f (new_AGEMA_signal_9218), .Z0_t (KeyArray_outS33ser[3]), .Z0_f (new_AGEMA_signal_5400), .Z1_t (new_AGEMA_signal_5401), .Z1_f (new_AGEMA_signal_5402) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_3_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS33ser[3]), .B0_f (new_AGEMA_signal_5400), .B1_t (new_AGEMA_signal_5401), .B1_f (new_AGEMA_signal_5402), .Z0_t (KeyArray_S33reg_gff_1_SFF_3_n1), .Z0_f (new_AGEMA_signal_9216), .Z1_t (new_AGEMA_signal_9217), .Z1_f (new_AGEMA_signal_9218) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_3_U1 ( .A0_t (KeyArray_S33reg_gff_1_SFF_3_QD), .A0_f (new_AGEMA_signal_9721), .A1_t (new_AGEMA_signal_9722), .A1_f (new_AGEMA_signal_9723), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S33reg_gff_1_SFF_3_n2), .Z0_f (new_AGEMA_signal_10197), .Z1_t (new_AGEMA_signal_10198), .Z1_f (new_AGEMA_signal_10199) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS33ser[3]), .A0_f (new_AGEMA_signal_7255), .A1_t (new_AGEMA_signal_7256), .A1_f (new_AGEMA_signal_7257), .B0_t (KeyArray_outS03ser[3]), .B0_f (new_AGEMA_signal_4536), .B1_t (new_AGEMA_signal_4537), .B1_f (new_AGEMA_signal_4538), .Z0_t (KeyArray_S33reg_gff_1_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_8064), .Z1_t (new_AGEMA_signal_8065), .Z1_f (new_AGEMA_signal_8066) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S33reg_gff_1_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_8064), .B1_t (new_AGEMA_signal_8065), .B1_f (new_AGEMA_signal_8066), .Z0_t (KeyArray_S33reg_gff_1_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_9219), .Z1_t (new_AGEMA_signal_9220), .Z1_f (new_AGEMA_signal_9221) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S33reg_gff_1_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_9219), .A1_t (new_AGEMA_signal_9220), .A1_f (new_AGEMA_signal_9221), .B0_t (KeyArray_inS33ser[3]), .B0_f (new_AGEMA_signal_7255), .B1_t (new_AGEMA_signal_7256), .B1_f (new_AGEMA_signal_7257), .Z0_t (KeyArray_S33reg_gff_1_SFF_3_QD), .Z0_f (new_AGEMA_signal_9721), .Z1_t (new_AGEMA_signal_9722), .Z1_f (new_AGEMA_signal_9723) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S33reg_gff_1_SFF_4_U3 ( .A0_t (KeyArray_S33reg_gff_1_SFF_4_n2), .A0_f (new_AGEMA_signal_10200), .A1_t (new_AGEMA_signal_10201), .A1_f (new_AGEMA_signal_10202), .B0_t (KeyArray_S33reg_gff_1_SFF_4_n1), .B0_f (new_AGEMA_signal_9222), .B1_t (new_AGEMA_signal_9223), .B1_f (new_AGEMA_signal_9224), .Z0_t (KeyArray_outS33ser[4]), .Z0_f (new_AGEMA_signal_5409), .Z1_t (new_AGEMA_signal_5410), .Z1_f (new_AGEMA_signal_5411) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_4_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS33ser[4]), .B0_f (new_AGEMA_signal_5409), .B1_t (new_AGEMA_signal_5410), .B1_f (new_AGEMA_signal_5411), .Z0_t (KeyArray_S33reg_gff_1_SFF_4_n1), .Z0_f (new_AGEMA_signal_9222), .Z1_t (new_AGEMA_signal_9223), .Z1_f (new_AGEMA_signal_9224) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_4_U1 ( .A0_t (KeyArray_S33reg_gff_1_SFF_4_QD), .A0_f (new_AGEMA_signal_9724), .A1_t (new_AGEMA_signal_9725), .A1_f (new_AGEMA_signal_9726), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S33reg_gff_1_SFF_4_n2), .Z0_f (new_AGEMA_signal_10200), .Z1_t (new_AGEMA_signal_10201), .Z1_f (new_AGEMA_signal_10202) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS33ser[4]), .A0_f (new_AGEMA_signal_7258), .A1_t (new_AGEMA_signal_7259), .A1_f (new_AGEMA_signal_7260), .B0_t (KeyArray_outS03ser[4]), .B0_f (new_AGEMA_signal_4545), .B1_t (new_AGEMA_signal_4546), .B1_f (new_AGEMA_signal_4547), .Z0_t (KeyArray_S33reg_gff_1_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_8067), .Z1_t (new_AGEMA_signal_8068), .Z1_f (new_AGEMA_signal_8069) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S33reg_gff_1_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_8067), .B1_t (new_AGEMA_signal_8068), .B1_f (new_AGEMA_signal_8069), .Z0_t (KeyArray_S33reg_gff_1_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_9225), .Z1_t (new_AGEMA_signal_9226), .Z1_f (new_AGEMA_signal_9227) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S33reg_gff_1_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_9225), .A1_t (new_AGEMA_signal_9226), .A1_f (new_AGEMA_signal_9227), .B0_t (KeyArray_inS33ser[4]), .B0_f (new_AGEMA_signal_7258), .B1_t (new_AGEMA_signal_7259), .B1_f (new_AGEMA_signal_7260), .Z0_t (KeyArray_S33reg_gff_1_SFF_4_QD), .Z0_f (new_AGEMA_signal_9724), .Z1_t (new_AGEMA_signal_9725), .Z1_f (new_AGEMA_signal_9726) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S33reg_gff_1_SFF_5_U3 ( .A0_t (KeyArray_S33reg_gff_1_SFF_5_n2), .A0_f (new_AGEMA_signal_10203), .A1_t (new_AGEMA_signal_10204), .A1_f (new_AGEMA_signal_10205), .B0_t (KeyArray_S33reg_gff_1_SFF_5_n1), .B0_f (new_AGEMA_signal_9228), .B1_t (new_AGEMA_signal_9229), .B1_f (new_AGEMA_signal_9230), .Z0_t (KeyArray_outS33ser[5]), .Z0_f (new_AGEMA_signal_5418), .Z1_t (new_AGEMA_signal_5419), .Z1_f (new_AGEMA_signal_5420) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_5_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS33ser[5]), .B0_f (new_AGEMA_signal_5418), .B1_t (new_AGEMA_signal_5419), .B1_f (new_AGEMA_signal_5420), .Z0_t (KeyArray_S33reg_gff_1_SFF_5_n1), .Z0_f (new_AGEMA_signal_9228), .Z1_t (new_AGEMA_signal_9229), .Z1_f (new_AGEMA_signal_9230) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_5_U1 ( .A0_t (KeyArray_S33reg_gff_1_SFF_5_QD), .A0_f (new_AGEMA_signal_9727), .A1_t (new_AGEMA_signal_9728), .A1_f (new_AGEMA_signal_9729), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S33reg_gff_1_SFF_5_n2), .Z0_f (new_AGEMA_signal_10203), .Z1_t (new_AGEMA_signal_10204), .Z1_f (new_AGEMA_signal_10205) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS33ser[5]), .A0_f (new_AGEMA_signal_7261), .A1_t (new_AGEMA_signal_7262), .A1_f (new_AGEMA_signal_7263), .B0_t (KeyArray_outS03ser[5]), .B0_f (new_AGEMA_signal_4554), .B1_t (new_AGEMA_signal_4555), .B1_f (new_AGEMA_signal_4556), .Z0_t (KeyArray_S33reg_gff_1_SFF_5_MUXInst_X), .Z0_f (new_AGEMA_signal_8070), .Z1_t (new_AGEMA_signal_8071), .Z1_f (new_AGEMA_signal_8072) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S33reg_gff_1_SFF_5_MUXInst_X), .B0_f (new_AGEMA_signal_8070), .B1_t (new_AGEMA_signal_8071), .B1_f (new_AGEMA_signal_8072), .Z0_t (KeyArray_S33reg_gff_1_SFF_5_MUXInst_Y), .Z0_f (new_AGEMA_signal_9231), .Z1_t (new_AGEMA_signal_9232), .Z1_f (new_AGEMA_signal_9233) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S33reg_gff_1_SFF_5_MUXInst_Y), .A0_f (new_AGEMA_signal_9231), .A1_t (new_AGEMA_signal_9232), .A1_f (new_AGEMA_signal_9233), .B0_t (KeyArray_inS33ser[5]), .B0_f (new_AGEMA_signal_7261), .B1_t (new_AGEMA_signal_7262), .B1_f (new_AGEMA_signal_7263), .Z0_t (KeyArray_S33reg_gff_1_SFF_5_QD), .Z0_f (new_AGEMA_signal_9727), .Z1_t (new_AGEMA_signal_9728), .Z1_f (new_AGEMA_signal_9729) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S33reg_gff_1_SFF_6_U3 ( .A0_t (KeyArray_S33reg_gff_1_SFF_6_n2), .A0_f (new_AGEMA_signal_10206), .A1_t (new_AGEMA_signal_10207), .A1_f (new_AGEMA_signal_10208), .B0_t (KeyArray_S33reg_gff_1_SFF_6_n1), .B0_f (new_AGEMA_signal_9234), .B1_t (new_AGEMA_signal_9235), .B1_f (new_AGEMA_signal_9236), .Z0_t (KeyArray_outS33ser[6]), .Z0_f (new_AGEMA_signal_5427), .Z1_t (new_AGEMA_signal_5428), .Z1_f (new_AGEMA_signal_5429) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_6_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS33ser[6]), .B0_f (new_AGEMA_signal_5427), .B1_t (new_AGEMA_signal_5428), .B1_f (new_AGEMA_signal_5429), .Z0_t (KeyArray_S33reg_gff_1_SFF_6_n1), .Z0_f (new_AGEMA_signal_9234), .Z1_t (new_AGEMA_signal_9235), .Z1_f (new_AGEMA_signal_9236) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_6_U1 ( .A0_t (KeyArray_S33reg_gff_1_SFF_6_QD), .A0_f (new_AGEMA_signal_9730), .A1_t (new_AGEMA_signal_9731), .A1_f (new_AGEMA_signal_9732), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S33reg_gff_1_SFF_6_n2), .Z0_f (new_AGEMA_signal_10206), .Z1_t (new_AGEMA_signal_10207), .Z1_f (new_AGEMA_signal_10208) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS33ser[6]), .A0_f (new_AGEMA_signal_7264), .A1_t (new_AGEMA_signal_7265), .A1_f (new_AGEMA_signal_7266), .B0_t (KeyArray_outS03ser[6]), .B0_f (new_AGEMA_signal_4563), .B1_t (new_AGEMA_signal_4564), .B1_f (new_AGEMA_signal_4565), .Z0_t (KeyArray_S33reg_gff_1_SFF_6_MUXInst_X), .Z0_f (new_AGEMA_signal_8073), .Z1_t (new_AGEMA_signal_8074), .Z1_f (new_AGEMA_signal_8075) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S33reg_gff_1_SFF_6_MUXInst_X), .B0_f (new_AGEMA_signal_8073), .B1_t (new_AGEMA_signal_8074), .B1_f (new_AGEMA_signal_8075), .Z0_t (KeyArray_S33reg_gff_1_SFF_6_MUXInst_Y), .Z0_f (new_AGEMA_signal_9237), .Z1_t (new_AGEMA_signal_9238), .Z1_f (new_AGEMA_signal_9239) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S33reg_gff_1_SFF_6_MUXInst_Y), .A0_f (new_AGEMA_signal_9237), .A1_t (new_AGEMA_signal_9238), .A1_f (new_AGEMA_signal_9239), .B0_t (KeyArray_inS33ser[6]), .B0_f (new_AGEMA_signal_7264), .B1_t (new_AGEMA_signal_7265), .B1_f (new_AGEMA_signal_7266), .Z0_t (KeyArray_S33reg_gff_1_SFF_6_QD), .Z0_f (new_AGEMA_signal_9730), .Z1_t (new_AGEMA_signal_9731), .Z1_f (new_AGEMA_signal_9732) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S33reg_gff_1_SFF_7_U3 ( .A0_t (KeyArray_S33reg_gff_1_SFF_7_n2), .A0_f (new_AGEMA_signal_10209), .A1_t (new_AGEMA_signal_10210), .A1_f (new_AGEMA_signal_10211), .B0_t (KeyArray_S33reg_gff_1_SFF_7_n1), .B0_f (new_AGEMA_signal_9240), .B1_t (new_AGEMA_signal_9241), .B1_f (new_AGEMA_signal_9242), .Z0_t (KeyArray_outS33ser[7]), .Z0_f (new_AGEMA_signal_5436), .Z1_t (new_AGEMA_signal_5437), .Z1_f (new_AGEMA_signal_5438) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_7_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n9), .A1_f (new_AGEMA_signal_7394), .B0_t (KeyArray_outS33ser[7]), .B0_f (new_AGEMA_signal_5436), .B1_t (new_AGEMA_signal_5437), .B1_f (new_AGEMA_signal_5438), .Z0_t (KeyArray_S33reg_gff_1_SFF_7_n1), .Z0_f (new_AGEMA_signal_9240), .Z1_t (new_AGEMA_signal_9241), .Z1_f (new_AGEMA_signal_9242) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_7_U1 ( .A0_t (KeyArray_S33reg_gff_1_SFF_7_QD), .A0_f (new_AGEMA_signal_9733), .A1_t (new_AGEMA_signal_9734), .A1_f (new_AGEMA_signal_9735), .B0_t (1'b0), .B0_f (1'b1), .B1_t (ctrl_n9), .B1_f (new_AGEMA_signal_7394), .Z0_t (KeyArray_S33reg_gff_1_SFF_7_n2), .Z0_f (new_AGEMA_signal_10209), .Z1_t (new_AGEMA_signal_10210), .Z1_f (new_AGEMA_signal_10211) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS33ser[7]), .A0_f (new_AGEMA_signal_7267), .A1_t (new_AGEMA_signal_7268), .A1_f (new_AGEMA_signal_7269), .B0_t (KeyArray_outS03ser[7]), .B0_f (new_AGEMA_signal_4572), .B1_t (new_AGEMA_signal_4573), .B1_f (new_AGEMA_signal_4574), .Z0_t (KeyArray_S33reg_gff_1_SFF_7_MUXInst_X), .Z0_f (new_AGEMA_signal_8076), .Z1_t (new_AGEMA_signal_8077), .Z1_f (new_AGEMA_signal_8078) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (KeyArray_S33reg_gff_1_SFF_7_MUXInst_X), .B0_f (new_AGEMA_signal_8076), .B1_t (new_AGEMA_signal_8077), .B1_f (new_AGEMA_signal_8078), .Z0_t (KeyArray_S33reg_gff_1_SFF_7_MUXInst_Y), .Z0_f (new_AGEMA_signal_9243), .Z1_t (new_AGEMA_signal_9244), .Z1_f (new_AGEMA_signal_9245) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S33reg_gff_1_SFF_7_MUXInst_Y), .A0_f (new_AGEMA_signal_9243), .A1_t (new_AGEMA_signal_9244), .A1_f (new_AGEMA_signal_9245), .B0_t (KeyArray_inS33ser[7]), .B0_f (new_AGEMA_signal_7267), .B1_t (new_AGEMA_signal_7268), .B1_f (new_AGEMA_signal_7269), .Z0_t (KeyArray_S33reg_gff_1_SFF_7_QD), .Z0_f (new_AGEMA_signal_9733), .Z1_t (new_AGEMA_signal_9734), .Z1_f (new_AGEMA_signal_9735) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_selXOR_mux_inst_0_XOR1_U1 ( .A0_t (KeyArray_outS01ser_0_), .A0_f (new_AGEMA_signal_4428), .A1_t (new_AGEMA_signal_4429), .A1_f (new_AGEMA_signal_4430), .B0_t (KeyArray_outS01ser_XOR_00[0]), .B0_f (new_AGEMA_signal_4431), .B1_t (new_AGEMA_signal_4432), .B1_f (new_AGEMA_signal_4433), .Z0_t (KeyArray_MUX_selXOR_mux_inst_0_X), .Z0_f (new_AGEMA_signal_6112), .Z1_t (new_AGEMA_signal_6113), .Z1_f (new_AGEMA_signal_6114) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_selXOR_mux_inst_0_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intselXOR), .A1_f (new_AGEMA_signal_7391), .B0_t (KeyArray_MUX_selXOR_mux_inst_0_X), .B0_f (new_AGEMA_signal_6112), .B1_t (new_AGEMA_signal_6113), .B1_f (new_AGEMA_signal_6114), .Z0_t (KeyArray_MUX_selXOR_mux_inst_0_Y), .Z0_f (new_AGEMA_signal_9246), .Z1_t (new_AGEMA_signal_9247), .Z1_f (new_AGEMA_signal_9248) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_selXOR_mux_inst_0_XOR2_U1 ( .A0_t (KeyArray_MUX_selXOR_mux_inst_0_Y), .A0_f (new_AGEMA_signal_9246), .A1_t (new_AGEMA_signal_9247), .A1_f (new_AGEMA_signal_9248), .B0_t (KeyArray_outS01ser_0_), .B0_f (new_AGEMA_signal_4428), .B1_t (new_AGEMA_signal_4429), .B1_f (new_AGEMA_signal_4430), .Z0_t (KeyArray_outS01ser_p[0]), .Z0_f (new_AGEMA_signal_9736), .Z1_t (new_AGEMA_signal_9737), .Z1_f (new_AGEMA_signal_9738) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_selXOR_mux_inst_1_XOR1_U1 ( .A0_t (KeyArray_outS01ser_1_), .A0_f (new_AGEMA_signal_4422), .A1_t (new_AGEMA_signal_4423), .A1_f (new_AGEMA_signal_4424), .B0_t (KeyArray_outS01ser_XOR_00[1]), .B0_f (new_AGEMA_signal_4425), .B1_t (new_AGEMA_signal_4426), .B1_f (new_AGEMA_signal_4427), .Z0_t (KeyArray_MUX_selXOR_mux_inst_1_X), .Z0_f (new_AGEMA_signal_6115), .Z1_t (new_AGEMA_signal_6116), .Z1_f (new_AGEMA_signal_6117) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_selXOR_mux_inst_1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intselXOR), .A1_f (new_AGEMA_signal_7391), .B0_t (KeyArray_MUX_selXOR_mux_inst_1_X), .B0_f (new_AGEMA_signal_6115), .B1_t (new_AGEMA_signal_6116), .B1_f (new_AGEMA_signal_6117), .Z0_t (KeyArray_MUX_selXOR_mux_inst_1_Y), .Z0_f (new_AGEMA_signal_9249), .Z1_t (new_AGEMA_signal_9250), .Z1_f (new_AGEMA_signal_9251) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_selXOR_mux_inst_1_XOR2_U1 ( .A0_t (KeyArray_MUX_selXOR_mux_inst_1_Y), .A0_f (new_AGEMA_signal_9249), .A1_t (new_AGEMA_signal_9250), .A1_f (new_AGEMA_signal_9251), .B0_t (KeyArray_outS01ser_1_), .B0_f (new_AGEMA_signal_4422), .B1_t (new_AGEMA_signal_4423), .B1_f (new_AGEMA_signal_4424), .Z0_t (KeyArray_outS01ser_p[1]), .Z0_f (new_AGEMA_signal_9739), .Z1_t (new_AGEMA_signal_9740), .Z1_f (new_AGEMA_signal_9741) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_selXOR_mux_inst_2_XOR1_U1 ( .A0_t (KeyArray_outS01ser_2_), .A0_f (new_AGEMA_signal_4416), .A1_t (new_AGEMA_signal_4417), .A1_f (new_AGEMA_signal_4418), .B0_t (KeyArray_outS01ser_XOR_00[2]), .B0_f (new_AGEMA_signal_4419), .B1_t (new_AGEMA_signal_4420), .B1_f (new_AGEMA_signal_4421), .Z0_t (KeyArray_MUX_selXOR_mux_inst_2_X), .Z0_f (new_AGEMA_signal_6118), .Z1_t (new_AGEMA_signal_6119), .Z1_f (new_AGEMA_signal_6120) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_selXOR_mux_inst_2_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intselXOR), .A1_f (new_AGEMA_signal_7391), .B0_t (KeyArray_MUX_selXOR_mux_inst_2_X), .B0_f (new_AGEMA_signal_6118), .B1_t (new_AGEMA_signal_6119), .B1_f (new_AGEMA_signal_6120), .Z0_t (KeyArray_MUX_selXOR_mux_inst_2_Y), .Z0_f (new_AGEMA_signal_9252), .Z1_t (new_AGEMA_signal_9253), .Z1_f (new_AGEMA_signal_9254) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_selXOR_mux_inst_2_XOR2_U1 ( .A0_t (KeyArray_MUX_selXOR_mux_inst_2_Y), .A0_f (new_AGEMA_signal_9252), .A1_t (new_AGEMA_signal_9253), .A1_f (new_AGEMA_signal_9254), .B0_t (KeyArray_outS01ser_2_), .B0_f (new_AGEMA_signal_4416), .B1_t (new_AGEMA_signal_4417), .B1_f (new_AGEMA_signal_4418), .Z0_t (KeyArray_outS01ser_p[2]), .Z0_f (new_AGEMA_signal_9742), .Z1_t (new_AGEMA_signal_9743), .Z1_f (new_AGEMA_signal_9744) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_selXOR_mux_inst_3_XOR1_U1 ( .A0_t (KeyArray_outS01ser_3_), .A0_f (new_AGEMA_signal_4410), .A1_t (new_AGEMA_signal_4411), .A1_f (new_AGEMA_signal_4412), .B0_t (KeyArray_outS01ser_XOR_00[3]), .B0_f (new_AGEMA_signal_4413), .B1_t (new_AGEMA_signal_4414), .B1_f (new_AGEMA_signal_4415), .Z0_t (KeyArray_MUX_selXOR_mux_inst_3_X), .Z0_f (new_AGEMA_signal_6121), .Z1_t (new_AGEMA_signal_6122), .Z1_f (new_AGEMA_signal_6123) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_selXOR_mux_inst_3_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intselXOR), .A1_f (new_AGEMA_signal_7391), .B0_t (KeyArray_MUX_selXOR_mux_inst_3_X), .B0_f (new_AGEMA_signal_6121), .B1_t (new_AGEMA_signal_6122), .B1_f (new_AGEMA_signal_6123), .Z0_t (KeyArray_MUX_selXOR_mux_inst_3_Y), .Z0_f (new_AGEMA_signal_9255), .Z1_t (new_AGEMA_signal_9256), .Z1_f (new_AGEMA_signal_9257) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_selXOR_mux_inst_3_XOR2_U1 ( .A0_t (KeyArray_MUX_selXOR_mux_inst_3_Y), .A0_f (new_AGEMA_signal_9255), .A1_t (new_AGEMA_signal_9256), .A1_f (new_AGEMA_signal_9257), .B0_t (KeyArray_outS01ser_3_), .B0_f (new_AGEMA_signal_4410), .B1_t (new_AGEMA_signal_4411), .B1_f (new_AGEMA_signal_4412), .Z0_t (KeyArray_outS01ser_p[3]), .Z0_f (new_AGEMA_signal_9745), .Z1_t (new_AGEMA_signal_9746), .Z1_f (new_AGEMA_signal_9747) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_selXOR_mux_inst_4_XOR1_U1 ( .A0_t (KeyArray_outS01ser_4_), .A0_f (new_AGEMA_signal_4404), .A1_t (new_AGEMA_signal_4405), .A1_f (new_AGEMA_signal_4406), .B0_t (KeyArray_outS01ser_XOR_00[4]), .B0_f (new_AGEMA_signal_4407), .B1_t (new_AGEMA_signal_4408), .B1_f (new_AGEMA_signal_4409), .Z0_t (KeyArray_MUX_selXOR_mux_inst_4_X), .Z0_f (new_AGEMA_signal_6124), .Z1_t (new_AGEMA_signal_6125), .Z1_f (new_AGEMA_signal_6126) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_selXOR_mux_inst_4_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intselXOR), .A1_f (new_AGEMA_signal_7391), .B0_t (KeyArray_MUX_selXOR_mux_inst_4_X), .B0_f (new_AGEMA_signal_6124), .B1_t (new_AGEMA_signal_6125), .B1_f (new_AGEMA_signal_6126), .Z0_t (KeyArray_MUX_selXOR_mux_inst_4_Y), .Z0_f (new_AGEMA_signal_9258), .Z1_t (new_AGEMA_signal_9259), .Z1_f (new_AGEMA_signal_9260) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_selXOR_mux_inst_4_XOR2_U1 ( .A0_t (KeyArray_MUX_selXOR_mux_inst_4_Y), .A0_f (new_AGEMA_signal_9258), .A1_t (new_AGEMA_signal_9259), .A1_f (new_AGEMA_signal_9260), .B0_t (KeyArray_outS01ser_4_), .B0_f (new_AGEMA_signal_4404), .B1_t (new_AGEMA_signal_4405), .B1_f (new_AGEMA_signal_4406), .Z0_t (KeyArray_outS01ser_p[4]), .Z0_f (new_AGEMA_signal_9748), .Z1_t (new_AGEMA_signal_9749), .Z1_f (new_AGEMA_signal_9750) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_selXOR_mux_inst_5_XOR1_U1 ( .A0_t (KeyArray_outS01ser_5_), .A0_f (new_AGEMA_signal_4398), .A1_t (new_AGEMA_signal_4399), .A1_f (new_AGEMA_signal_4400), .B0_t (KeyArray_outS01ser_XOR_00[5]), .B0_f (new_AGEMA_signal_4401), .B1_t (new_AGEMA_signal_4402), .B1_f (new_AGEMA_signal_4403), .Z0_t (KeyArray_MUX_selXOR_mux_inst_5_X), .Z0_f (new_AGEMA_signal_6127), .Z1_t (new_AGEMA_signal_6128), .Z1_f (new_AGEMA_signal_6129) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_selXOR_mux_inst_5_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intselXOR), .A1_f (new_AGEMA_signal_7391), .B0_t (KeyArray_MUX_selXOR_mux_inst_5_X), .B0_f (new_AGEMA_signal_6127), .B1_t (new_AGEMA_signal_6128), .B1_f (new_AGEMA_signal_6129), .Z0_t (KeyArray_MUX_selXOR_mux_inst_5_Y), .Z0_f (new_AGEMA_signal_9261), .Z1_t (new_AGEMA_signal_9262), .Z1_f (new_AGEMA_signal_9263) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_selXOR_mux_inst_5_XOR2_U1 ( .A0_t (KeyArray_MUX_selXOR_mux_inst_5_Y), .A0_f (new_AGEMA_signal_9261), .A1_t (new_AGEMA_signal_9262), .A1_f (new_AGEMA_signal_9263), .B0_t (KeyArray_outS01ser_5_), .B0_f (new_AGEMA_signal_4398), .B1_t (new_AGEMA_signal_4399), .B1_f (new_AGEMA_signal_4400), .Z0_t (KeyArray_outS01ser_p[5]), .Z0_f (new_AGEMA_signal_9751), .Z1_t (new_AGEMA_signal_9752), .Z1_f (new_AGEMA_signal_9753) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_selXOR_mux_inst_6_XOR1_U1 ( .A0_t (KeyArray_outS01ser_6_), .A0_f (new_AGEMA_signal_4392), .A1_t (new_AGEMA_signal_4393), .A1_f (new_AGEMA_signal_4394), .B0_t (KeyArray_outS01ser_XOR_00[6]), .B0_f (new_AGEMA_signal_4395), .B1_t (new_AGEMA_signal_4396), .B1_f (new_AGEMA_signal_4397), .Z0_t (KeyArray_MUX_selXOR_mux_inst_6_X), .Z0_f (new_AGEMA_signal_6130), .Z1_t (new_AGEMA_signal_6131), .Z1_f (new_AGEMA_signal_6132) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_selXOR_mux_inst_6_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intselXOR), .A1_f (new_AGEMA_signal_7391), .B0_t (KeyArray_MUX_selXOR_mux_inst_6_X), .B0_f (new_AGEMA_signal_6130), .B1_t (new_AGEMA_signal_6131), .B1_f (new_AGEMA_signal_6132), .Z0_t (KeyArray_MUX_selXOR_mux_inst_6_Y), .Z0_f (new_AGEMA_signal_9264), .Z1_t (new_AGEMA_signal_9265), .Z1_f (new_AGEMA_signal_9266) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_selXOR_mux_inst_6_XOR2_U1 ( .A0_t (KeyArray_MUX_selXOR_mux_inst_6_Y), .A0_f (new_AGEMA_signal_9264), .A1_t (new_AGEMA_signal_9265), .A1_f (new_AGEMA_signal_9266), .B0_t (KeyArray_outS01ser_6_), .B0_f (new_AGEMA_signal_4392), .B1_t (new_AGEMA_signal_4393), .B1_f (new_AGEMA_signal_4394), .Z0_t (KeyArray_outS01ser_p[6]), .Z0_f (new_AGEMA_signal_9754), .Z1_t (new_AGEMA_signal_9755), .Z1_f (new_AGEMA_signal_9756) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_selXOR_mux_inst_7_XOR1_U1 ( .A0_t (KeyArray_outS01ser_7_), .A0_f (new_AGEMA_signal_4386), .A1_t (new_AGEMA_signal_4387), .A1_f (new_AGEMA_signal_4388), .B0_t (KeyArray_outS01ser_XOR_00[7]), .B0_f (new_AGEMA_signal_4389), .B1_t (new_AGEMA_signal_4390), .B1_f (new_AGEMA_signal_4391), .Z0_t (KeyArray_MUX_selXOR_mux_inst_7_X), .Z0_f (new_AGEMA_signal_6133), .Z1_t (new_AGEMA_signal_6134), .Z1_f (new_AGEMA_signal_6135) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_selXOR_mux_inst_7_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intselXOR), .A1_f (new_AGEMA_signal_7391), .B0_t (KeyArray_MUX_selXOR_mux_inst_7_X), .B0_f (new_AGEMA_signal_6133), .B1_t (new_AGEMA_signal_6134), .B1_f (new_AGEMA_signal_6135), .Z0_t (KeyArray_MUX_selXOR_mux_inst_7_Y), .Z0_f (new_AGEMA_signal_9267), .Z1_t (new_AGEMA_signal_9268), .Z1_f (new_AGEMA_signal_9269) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_selXOR_mux_inst_7_XOR2_U1 ( .A0_t (KeyArray_MUX_selXOR_mux_inst_7_Y), .A0_f (new_AGEMA_signal_9267), .A1_t (new_AGEMA_signal_9268), .A1_f (new_AGEMA_signal_9269), .B0_t (KeyArray_outS01ser_7_), .B0_f (new_AGEMA_signal_4386), .B1_t (new_AGEMA_signal_4387), .B1_f (new_AGEMA_signal_4388), .Z0_t (KeyArray_outS01ser_p[7]), .Z0_f (new_AGEMA_signal_9757), .Z1_t (new_AGEMA_signal_9758), .Z1_f (new_AGEMA_signal_9759) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_0_XOR1_U1 ( .A0_t (key_s0_t[120]), .A0_f (key_s0_f[120]), .A1_t (key_s1_t[120]), .A1_f (key_s1_f[120]), .B0_t (KeyArray_outS01ser_p[0]), .B0_f (new_AGEMA_signal_9736), .B1_t (new_AGEMA_signal_9737), .B1_f (new_AGEMA_signal_9738), .Z0_t (KeyArray_MUX_inS00ser_mux_inst_0_X), .Z0_f (new_AGEMA_signal_10215), .Z1_t (new_AGEMA_signal_10216), .Z1_f (new_AGEMA_signal_10217) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_0_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS00ser_mux_inst_0_X), .B0_f (new_AGEMA_signal_10215), .B1_t (new_AGEMA_signal_10216), .B1_f (new_AGEMA_signal_10217), .Z0_t (KeyArray_MUX_inS00ser_mux_inst_0_Y), .Z0_f (new_AGEMA_signal_10379), .Z1_t (new_AGEMA_signal_10380), .Z1_f (new_AGEMA_signal_10381) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_0_XOR2_U1 ( .A0_t (KeyArray_MUX_inS00ser_mux_inst_0_Y), .A0_f (new_AGEMA_signal_10379), .A1_t (new_AGEMA_signal_10380), .A1_f (new_AGEMA_signal_10381), .B0_t (key_s0_t[120]), .B0_f (key_s0_f[120]), .B1_t (key_s1_t[120]), .B1_f (key_s1_f[120]), .Z0_t (KeyArray_inS00ser[0]), .Z0_f (new_AGEMA_signal_10502), .Z1_t (new_AGEMA_signal_10503), .Z1_f (new_AGEMA_signal_10504) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_1_XOR1_U1 ( .A0_t (key_s0_t[121]), .A0_f (key_s0_f[121]), .A1_t (key_s1_t[121]), .A1_f (key_s1_f[121]), .B0_t (KeyArray_outS01ser_p[1]), .B0_f (new_AGEMA_signal_9739), .B1_t (new_AGEMA_signal_9740), .B1_f (new_AGEMA_signal_9741), .Z0_t (KeyArray_MUX_inS00ser_mux_inst_1_X), .Z0_f (new_AGEMA_signal_10221), .Z1_t (new_AGEMA_signal_10222), .Z1_f (new_AGEMA_signal_10223) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS00ser_mux_inst_1_X), .B0_f (new_AGEMA_signal_10221), .B1_t (new_AGEMA_signal_10222), .B1_f (new_AGEMA_signal_10223), .Z0_t (KeyArray_MUX_inS00ser_mux_inst_1_Y), .Z0_f (new_AGEMA_signal_10382), .Z1_t (new_AGEMA_signal_10383), .Z1_f (new_AGEMA_signal_10384) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_1_XOR2_U1 ( .A0_t (KeyArray_MUX_inS00ser_mux_inst_1_Y), .A0_f (new_AGEMA_signal_10382), .A1_t (new_AGEMA_signal_10383), .A1_f (new_AGEMA_signal_10384), .B0_t (key_s0_t[121]), .B0_f (key_s0_f[121]), .B1_t (key_s1_t[121]), .B1_f (key_s1_f[121]), .Z0_t (KeyArray_inS00ser[1]), .Z0_f (new_AGEMA_signal_10505), .Z1_t (new_AGEMA_signal_10506), .Z1_f (new_AGEMA_signal_10507) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_2_XOR1_U1 ( .A0_t (key_s0_t[122]), .A0_f (key_s0_f[122]), .A1_t (key_s1_t[122]), .A1_f (key_s1_f[122]), .B0_t (KeyArray_outS01ser_p[2]), .B0_f (new_AGEMA_signal_9742), .B1_t (new_AGEMA_signal_9743), .B1_f (new_AGEMA_signal_9744), .Z0_t (KeyArray_MUX_inS00ser_mux_inst_2_X), .Z0_f (new_AGEMA_signal_10227), .Z1_t (new_AGEMA_signal_10228), .Z1_f (new_AGEMA_signal_10229) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_2_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS00ser_mux_inst_2_X), .B0_f (new_AGEMA_signal_10227), .B1_t (new_AGEMA_signal_10228), .B1_f (new_AGEMA_signal_10229), .Z0_t (KeyArray_MUX_inS00ser_mux_inst_2_Y), .Z0_f (new_AGEMA_signal_10385), .Z1_t (new_AGEMA_signal_10386), .Z1_f (new_AGEMA_signal_10387) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_2_XOR2_U1 ( .A0_t (KeyArray_MUX_inS00ser_mux_inst_2_Y), .A0_f (new_AGEMA_signal_10385), .A1_t (new_AGEMA_signal_10386), .A1_f (new_AGEMA_signal_10387), .B0_t (key_s0_t[122]), .B0_f (key_s0_f[122]), .B1_t (key_s1_t[122]), .B1_f (key_s1_f[122]), .Z0_t (KeyArray_inS00ser[2]), .Z0_f (new_AGEMA_signal_10508), .Z1_t (new_AGEMA_signal_10509), .Z1_f (new_AGEMA_signal_10510) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_3_XOR1_U1 ( .A0_t (key_s0_t[123]), .A0_f (key_s0_f[123]), .A1_t (key_s1_t[123]), .A1_f (key_s1_f[123]), .B0_t (KeyArray_outS01ser_p[3]), .B0_f (new_AGEMA_signal_9745), .B1_t (new_AGEMA_signal_9746), .B1_f (new_AGEMA_signal_9747), .Z0_t (KeyArray_MUX_inS00ser_mux_inst_3_X), .Z0_f (new_AGEMA_signal_10233), .Z1_t (new_AGEMA_signal_10234), .Z1_f (new_AGEMA_signal_10235) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_3_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS00ser_mux_inst_3_X), .B0_f (new_AGEMA_signal_10233), .B1_t (new_AGEMA_signal_10234), .B1_f (new_AGEMA_signal_10235), .Z0_t (KeyArray_MUX_inS00ser_mux_inst_3_Y), .Z0_f (new_AGEMA_signal_10388), .Z1_t (new_AGEMA_signal_10389), .Z1_f (new_AGEMA_signal_10390) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_3_XOR2_U1 ( .A0_t (KeyArray_MUX_inS00ser_mux_inst_3_Y), .A0_f (new_AGEMA_signal_10388), .A1_t (new_AGEMA_signal_10389), .A1_f (new_AGEMA_signal_10390), .B0_t (key_s0_t[123]), .B0_f (key_s0_f[123]), .B1_t (key_s1_t[123]), .B1_f (key_s1_f[123]), .Z0_t (KeyArray_inS00ser[3]), .Z0_f (new_AGEMA_signal_10511), .Z1_t (new_AGEMA_signal_10512), .Z1_f (new_AGEMA_signal_10513) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_4_XOR1_U1 ( .A0_t (key_s0_t[124]), .A0_f (key_s0_f[124]), .A1_t (key_s1_t[124]), .A1_f (key_s1_f[124]), .B0_t (KeyArray_outS01ser_p[4]), .B0_f (new_AGEMA_signal_9748), .B1_t (new_AGEMA_signal_9749), .B1_f (new_AGEMA_signal_9750), .Z0_t (KeyArray_MUX_inS00ser_mux_inst_4_X), .Z0_f (new_AGEMA_signal_10239), .Z1_t (new_AGEMA_signal_10240), .Z1_f (new_AGEMA_signal_10241) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_4_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS00ser_mux_inst_4_X), .B0_f (new_AGEMA_signal_10239), .B1_t (new_AGEMA_signal_10240), .B1_f (new_AGEMA_signal_10241), .Z0_t (KeyArray_MUX_inS00ser_mux_inst_4_Y), .Z0_f (new_AGEMA_signal_10391), .Z1_t (new_AGEMA_signal_10392), .Z1_f (new_AGEMA_signal_10393) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_4_XOR2_U1 ( .A0_t (KeyArray_MUX_inS00ser_mux_inst_4_Y), .A0_f (new_AGEMA_signal_10391), .A1_t (new_AGEMA_signal_10392), .A1_f (new_AGEMA_signal_10393), .B0_t (key_s0_t[124]), .B0_f (key_s0_f[124]), .B1_t (key_s1_t[124]), .B1_f (key_s1_f[124]), .Z0_t (KeyArray_inS00ser[4]), .Z0_f (new_AGEMA_signal_10514), .Z1_t (new_AGEMA_signal_10515), .Z1_f (new_AGEMA_signal_10516) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_5_XOR1_U1 ( .A0_t (key_s0_t[125]), .A0_f (key_s0_f[125]), .A1_t (key_s1_t[125]), .A1_f (key_s1_f[125]), .B0_t (KeyArray_outS01ser_p[5]), .B0_f (new_AGEMA_signal_9751), .B1_t (new_AGEMA_signal_9752), .B1_f (new_AGEMA_signal_9753), .Z0_t (KeyArray_MUX_inS00ser_mux_inst_5_X), .Z0_f (new_AGEMA_signal_10245), .Z1_t (new_AGEMA_signal_10246), .Z1_f (new_AGEMA_signal_10247) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_5_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS00ser_mux_inst_5_X), .B0_f (new_AGEMA_signal_10245), .B1_t (new_AGEMA_signal_10246), .B1_f (new_AGEMA_signal_10247), .Z0_t (KeyArray_MUX_inS00ser_mux_inst_5_Y), .Z0_f (new_AGEMA_signal_10394), .Z1_t (new_AGEMA_signal_10395), .Z1_f (new_AGEMA_signal_10396) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_5_XOR2_U1 ( .A0_t (KeyArray_MUX_inS00ser_mux_inst_5_Y), .A0_f (new_AGEMA_signal_10394), .A1_t (new_AGEMA_signal_10395), .A1_f (new_AGEMA_signal_10396), .B0_t (key_s0_t[125]), .B0_f (key_s0_f[125]), .B1_t (key_s1_t[125]), .B1_f (key_s1_f[125]), .Z0_t (KeyArray_inS00ser[5]), .Z0_f (new_AGEMA_signal_10517), .Z1_t (new_AGEMA_signal_10518), .Z1_f (new_AGEMA_signal_10519) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_6_XOR1_U1 ( .A0_t (key_s0_t[126]), .A0_f (key_s0_f[126]), .A1_t (key_s1_t[126]), .A1_f (key_s1_f[126]), .B0_t (KeyArray_outS01ser_p[6]), .B0_f (new_AGEMA_signal_9754), .B1_t (new_AGEMA_signal_9755), .B1_f (new_AGEMA_signal_9756), .Z0_t (KeyArray_MUX_inS00ser_mux_inst_6_X), .Z0_f (new_AGEMA_signal_10251), .Z1_t (new_AGEMA_signal_10252), .Z1_f (new_AGEMA_signal_10253) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_6_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS00ser_mux_inst_6_X), .B0_f (new_AGEMA_signal_10251), .B1_t (new_AGEMA_signal_10252), .B1_f (new_AGEMA_signal_10253), .Z0_t (KeyArray_MUX_inS00ser_mux_inst_6_Y), .Z0_f (new_AGEMA_signal_10397), .Z1_t (new_AGEMA_signal_10398), .Z1_f (new_AGEMA_signal_10399) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_6_XOR2_U1 ( .A0_t (KeyArray_MUX_inS00ser_mux_inst_6_Y), .A0_f (new_AGEMA_signal_10397), .A1_t (new_AGEMA_signal_10398), .A1_f (new_AGEMA_signal_10399), .B0_t (key_s0_t[126]), .B0_f (key_s0_f[126]), .B1_t (key_s1_t[126]), .B1_f (key_s1_f[126]), .Z0_t (KeyArray_inS00ser[6]), .Z0_f (new_AGEMA_signal_10520), .Z1_t (new_AGEMA_signal_10521), .Z1_f (new_AGEMA_signal_10522) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_7_XOR1_U1 ( .A0_t (key_s0_t[127]), .A0_f (key_s0_f[127]), .A1_t (key_s1_t[127]), .A1_f (key_s1_f[127]), .B0_t (KeyArray_outS01ser_p[7]), .B0_f (new_AGEMA_signal_9757), .B1_t (new_AGEMA_signal_9758), .B1_f (new_AGEMA_signal_9759), .Z0_t (KeyArray_MUX_inS00ser_mux_inst_7_X), .Z0_f (new_AGEMA_signal_10257), .Z1_t (new_AGEMA_signal_10258), .Z1_f (new_AGEMA_signal_10259) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_7_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS00ser_mux_inst_7_X), .B0_f (new_AGEMA_signal_10257), .B1_t (new_AGEMA_signal_10258), .B1_f (new_AGEMA_signal_10259), .Z0_t (KeyArray_MUX_inS00ser_mux_inst_7_Y), .Z0_f (new_AGEMA_signal_10400), .Z1_t (new_AGEMA_signal_10401), .Z1_f (new_AGEMA_signal_10402) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_7_XOR2_U1 ( .A0_t (KeyArray_MUX_inS00ser_mux_inst_7_Y), .A0_f (new_AGEMA_signal_10400), .A1_t (new_AGEMA_signal_10401), .A1_f (new_AGEMA_signal_10402), .B0_t (key_s0_t[127]), .B0_f (key_s0_f[127]), .B1_t (key_s1_t[127]), .B1_f (key_s1_f[127]), .Z0_t (KeyArray_inS00ser[7]), .Z0_f (new_AGEMA_signal_10523), .Z1_t (new_AGEMA_signal_10524), .Z1_f (new_AGEMA_signal_10525) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS01ser_mux_inst_0_XOR1_U1 ( .A0_t (key_s0_t[88]), .A0_f (key_s0_f[88]), .A1_t (key_s1_t[88]), .A1_f (key_s1_f[88]), .B0_t (KeyArray_outS02ser[0]), .B0_f (new_AGEMA_signal_4437), .B1_t (new_AGEMA_signal_4438), .B1_f (new_AGEMA_signal_4439), .Z0_t (KeyArray_MUX_inS01ser_mux_inst_0_X), .Z0_f (new_AGEMA_signal_4440), .Z1_t (new_AGEMA_signal_4441), .Z1_f (new_AGEMA_signal_4442) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS01ser_mux_inst_0_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS01ser_mux_inst_0_X), .B0_f (new_AGEMA_signal_4440), .B1_t (new_AGEMA_signal_4441), .B1_f (new_AGEMA_signal_4442), .Z0_t (KeyArray_MUX_inS01ser_mux_inst_0_Y), .Z0_f (new_AGEMA_signal_6136), .Z1_t (new_AGEMA_signal_6137), .Z1_f (new_AGEMA_signal_6138) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS01ser_mux_inst_0_XOR2_U1 ( .A0_t (KeyArray_MUX_inS01ser_mux_inst_0_Y), .A0_f (new_AGEMA_signal_6136), .A1_t (new_AGEMA_signal_6137), .A1_f (new_AGEMA_signal_6138), .B0_t (key_s0_t[88]), .B0_f (key_s0_f[88]), .B1_t (key_s1_t[88]), .B1_f (key_s1_f[88]), .Z0_t (KeyArray_inS01ser[0]), .Z0_f (new_AGEMA_signal_6910), .Z1_t (new_AGEMA_signal_6911), .Z1_f (new_AGEMA_signal_6912) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS01ser_mux_inst_1_XOR1_U1 ( .A0_t (key_s0_t[89]), .A0_f (key_s0_f[89]), .A1_t (key_s1_t[89]), .A1_f (key_s1_f[89]), .B0_t (KeyArray_outS02ser[1]), .B0_f (new_AGEMA_signal_4446), .B1_t (new_AGEMA_signal_4447), .B1_f (new_AGEMA_signal_4448), .Z0_t (KeyArray_MUX_inS01ser_mux_inst_1_X), .Z0_f (new_AGEMA_signal_4449), .Z1_t (new_AGEMA_signal_4450), .Z1_f (new_AGEMA_signal_4451) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS01ser_mux_inst_1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS01ser_mux_inst_1_X), .B0_f (new_AGEMA_signal_4449), .B1_t (new_AGEMA_signal_4450), .B1_f (new_AGEMA_signal_4451), .Z0_t (KeyArray_MUX_inS01ser_mux_inst_1_Y), .Z0_f (new_AGEMA_signal_6139), .Z1_t (new_AGEMA_signal_6140), .Z1_f (new_AGEMA_signal_6141) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS01ser_mux_inst_1_XOR2_U1 ( .A0_t (KeyArray_MUX_inS01ser_mux_inst_1_Y), .A0_f (new_AGEMA_signal_6139), .A1_t (new_AGEMA_signal_6140), .A1_f (new_AGEMA_signal_6141), .B0_t (key_s0_t[89]), .B0_f (key_s0_f[89]), .B1_t (key_s1_t[89]), .B1_f (key_s1_f[89]), .Z0_t (KeyArray_inS01ser[1]), .Z0_f (new_AGEMA_signal_6913), .Z1_t (new_AGEMA_signal_6914), .Z1_f (new_AGEMA_signal_6915) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS01ser_mux_inst_2_XOR1_U1 ( .A0_t (key_s0_t[90]), .A0_f (key_s0_f[90]), .A1_t (key_s1_t[90]), .A1_f (key_s1_f[90]), .B0_t (KeyArray_outS02ser[2]), .B0_f (new_AGEMA_signal_4455), .B1_t (new_AGEMA_signal_4456), .B1_f (new_AGEMA_signal_4457), .Z0_t (KeyArray_MUX_inS01ser_mux_inst_2_X), .Z0_f (new_AGEMA_signal_4458), .Z1_t (new_AGEMA_signal_4459), .Z1_f (new_AGEMA_signal_4460) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS01ser_mux_inst_2_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS01ser_mux_inst_2_X), .B0_f (new_AGEMA_signal_4458), .B1_t (new_AGEMA_signal_4459), .B1_f (new_AGEMA_signal_4460), .Z0_t (KeyArray_MUX_inS01ser_mux_inst_2_Y), .Z0_f (new_AGEMA_signal_6142), .Z1_t (new_AGEMA_signal_6143), .Z1_f (new_AGEMA_signal_6144) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS01ser_mux_inst_2_XOR2_U1 ( .A0_t (KeyArray_MUX_inS01ser_mux_inst_2_Y), .A0_f (new_AGEMA_signal_6142), .A1_t (new_AGEMA_signal_6143), .A1_f (new_AGEMA_signal_6144), .B0_t (key_s0_t[90]), .B0_f (key_s0_f[90]), .B1_t (key_s1_t[90]), .B1_f (key_s1_f[90]), .Z0_t (KeyArray_inS01ser[2]), .Z0_f (new_AGEMA_signal_6916), .Z1_t (new_AGEMA_signal_6917), .Z1_f (new_AGEMA_signal_6918) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS01ser_mux_inst_3_XOR1_U1 ( .A0_t (key_s0_t[91]), .A0_f (key_s0_f[91]), .A1_t (key_s1_t[91]), .A1_f (key_s1_f[91]), .B0_t (KeyArray_outS02ser[3]), .B0_f (new_AGEMA_signal_4464), .B1_t (new_AGEMA_signal_4465), .B1_f (new_AGEMA_signal_4466), .Z0_t (KeyArray_MUX_inS01ser_mux_inst_3_X), .Z0_f (new_AGEMA_signal_4467), .Z1_t (new_AGEMA_signal_4468), .Z1_f (new_AGEMA_signal_4469) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS01ser_mux_inst_3_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS01ser_mux_inst_3_X), .B0_f (new_AGEMA_signal_4467), .B1_t (new_AGEMA_signal_4468), .B1_f (new_AGEMA_signal_4469), .Z0_t (KeyArray_MUX_inS01ser_mux_inst_3_Y), .Z0_f (new_AGEMA_signal_6145), .Z1_t (new_AGEMA_signal_6146), .Z1_f (new_AGEMA_signal_6147) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS01ser_mux_inst_3_XOR2_U1 ( .A0_t (KeyArray_MUX_inS01ser_mux_inst_3_Y), .A0_f (new_AGEMA_signal_6145), .A1_t (new_AGEMA_signal_6146), .A1_f (new_AGEMA_signal_6147), .B0_t (key_s0_t[91]), .B0_f (key_s0_f[91]), .B1_t (key_s1_t[91]), .B1_f (key_s1_f[91]), .Z0_t (KeyArray_inS01ser[3]), .Z0_f (new_AGEMA_signal_6919), .Z1_t (new_AGEMA_signal_6920), .Z1_f (new_AGEMA_signal_6921) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS01ser_mux_inst_4_XOR1_U1 ( .A0_t (key_s0_t[92]), .A0_f (key_s0_f[92]), .A1_t (key_s1_t[92]), .A1_f (key_s1_f[92]), .B0_t (KeyArray_outS02ser[4]), .B0_f (new_AGEMA_signal_4473), .B1_t (new_AGEMA_signal_4474), .B1_f (new_AGEMA_signal_4475), .Z0_t (KeyArray_MUX_inS01ser_mux_inst_4_X), .Z0_f (new_AGEMA_signal_4476), .Z1_t (new_AGEMA_signal_4477), .Z1_f (new_AGEMA_signal_4478) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS01ser_mux_inst_4_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS01ser_mux_inst_4_X), .B0_f (new_AGEMA_signal_4476), .B1_t (new_AGEMA_signal_4477), .B1_f (new_AGEMA_signal_4478), .Z0_t (KeyArray_MUX_inS01ser_mux_inst_4_Y), .Z0_f (new_AGEMA_signal_6148), .Z1_t (new_AGEMA_signal_6149), .Z1_f (new_AGEMA_signal_6150) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS01ser_mux_inst_4_XOR2_U1 ( .A0_t (KeyArray_MUX_inS01ser_mux_inst_4_Y), .A0_f (new_AGEMA_signal_6148), .A1_t (new_AGEMA_signal_6149), .A1_f (new_AGEMA_signal_6150), .B0_t (key_s0_t[92]), .B0_f (key_s0_f[92]), .B1_t (key_s1_t[92]), .B1_f (key_s1_f[92]), .Z0_t (KeyArray_inS01ser[4]), .Z0_f (new_AGEMA_signal_6922), .Z1_t (new_AGEMA_signal_6923), .Z1_f (new_AGEMA_signal_6924) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS01ser_mux_inst_5_XOR1_U1 ( .A0_t (key_s0_t[93]), .A0_f (key_s0_f[93]), .A1_t (key_s1_t[93]), .A1_f (key_s1_f[93]), .B0_t (KeyArray_outS02ser[5]), .B0_f (new_AGEMA_signal_4482), .B1_t (new_AGEMA_signal_4483), .B1_f (new_AGEMA_signal_4484), .Z0_t (KeyArray_MUX_inS01ser_mux_inst_5_X), .Z0_f (new_AGEMA_signal_4485), .Z1_t (new_AGEMA_signal_4486), .Z1_f (new_AGEMA_signal_4487) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS01ser_mux_inst_5_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS01ser_mux_inst_5_X), .B0_f (new_AGEMA_signal_4485), .B1_t (new_AGEMA_signal_4486), .B1_f (new_AGEMA_signal_4487), .Z0_t (KeyArray_MUX_inS01ser_mux_inst_5_Y), .Z0_f (new_AGEMA_signal_6151), .Z1_t (new_AGEMA_signal_6152), .Z1_f (new_AGEMA_signal_6153) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS01ser_mux_inst_5_XOR2_U1 ( .A0_t (KeyArray_MUX_inS01ser_mux_inst_5_Y), .A0_f (new_AGEMA_signal_6151), .A1_t (new_AGEMA_signal_6152), .A1_f (new_AGEMA_signal_6153), .B0_t (key_s0_t[93]), .B0_f (key_s0_f[93]), .B1_t (key_s1_t[93]), .B1_f (key_s1_f[93]), .Z0_t (KeyArray_inS01ser[5]), .Z0_f (new_AGEMA_signal_6925), .Z1_t (new_AGEMA_signal_6926), .Z1_f (new_AGEMA_signal_6927) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS01ser_mux_inst_6_XOR1_U1 ( .A0_t (key_s0_t[94]), .A0_f (key_s0_f[94]), .A1_t (key_s1_t[94]), .A1_f (key_s1_f[94]), .B0_t (KeyArray_outS02ser[6]), .B0_f (new_AGEMA_signal_4491), .B1_t (new_AGEMA_signal_4492), .B1_f (new_AGEMA_signal_4493), .Z0_t (KeyArray_MUX_inS01ser_mux_inst_6_X), .Z0_f (new_AGEMA_signal_4494), .Z1_t (new_AGEMA_signal_4495), .Z1_f (new_AGEMA_signal_4496) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS01ser_mux_inst_6_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS01ser_mux_inst_6_X), .B0_f (new_AGEMA_signal_4494), .B1_t (new_AGEMA_signal_4495), .B1_f (new_AGEMA_signal_4496), .Z0_t (KeyArray_MUX_inS01ser_mux_inst_6_Y), .Z0_f (new_AGEMA_signal_6154), .Z1_t (new_AGEMA_signal_6155), .Z1_f (new_AGEMA_signal_6156) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS01ser_mux_inst_6_XOR2_U1 ( .A0_t (KeyArray_MUX_inS01ser_mux_inst_6_Y), .A0_f (new_AGEMA_signal_6154), .A1_t (new_AGEMA_signal_6155), .A1_f (new_AGEMA_signal_6156), .B0_t (key_s0_t[94]), .B0_f (key_s0_f[94]), .B1_t (key_s1_t[94]), .B1_f (key_s1_f[94]), .Z0_t (KeyArray_inS01ser[6]), .Z0_f (new_AGEMA_signal_6928), .Z1_t (new_AGEMA_signal_6929), .Z1_f (new_AGEMA_signal_6930) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS01ser_mux_inst_7_XOR1_U1 ( .A0_t (key_s0_t[95]), .A0_f (key_s0_f[95]), .A1_t (key_s1_t[95]), .A1_f (key_s1_f[95]), .B0_t (KeyArray_outS02ser[7]), .B0_f (new_AGEMA_signal_4500), .B1_t (new_AGEMA_signal_4501), .B1_f (new_AGEMA_signal_4502), .Z0_t (KeyArray_MUX_inS01ser_mux_inst_7_X), .Z0_f (new_AGEMA_signal_4503), .Z1_t (new_AGEMA_signal_4504), .Z1_f (new_AGEMA_signal_4505) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS01ser_mux_inst_7_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS01ser_mux_inst_7_X), .B0_f (new_AGEMA_signal_4503), .B1_t (new_AGEMA_signal_4504), .B1_f (new_AGEMA_signal_4505), .Z0_t (KeyArray_MUX_inS01ser_mux_inst_7_Y), .Z0_f (new_AGEMA_signal_6157), .Z1_t (new_AGEMA_signal_6158), .Z1_f (new_AGEMA_signal_6159) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS01ser_mux_inst_7_XOR2_U1 ( .A0_t (KeyArray_MUX_inS01ser_mux_inst_7_Y), .A0_f (new_AGEMA_signal_6157), .A1_t (new_AGEMA_signal_6158), .A1_f (new_AGEMA_signal_6159), .B0_t (key_s0_t[95]), .B0_f (key_s0_f[95]), .B1_t (key_s1_t[95]), .B1_f (key_s1_f[95]), .Z0_t (KeyArray_inS01ser[7]), .Z0_f (new_AGEMA_signal_6931), .Z1_t (new_AGEMA_signal_6932), .Z1_f (new_AGEMA_signal_6933) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS02ser_mux_inst_0_XOR1_U1 ( .A0_t (key_s0_t[56]), .A0_f (key_s0_f[56]), .A1_t (key_s1_t[56]), .A1_f (key_s1_f[56]), .B0_t (KeyArray_outS03ser[0]), .B0_f (new_AGEMA_signal_4509), .B1_t (new_AGEMA_signal_4510), .B1_f (new_AGEMA_signal_4511), .Z0_t (KeyArray_MUX_inS02ser_mux_inst_0_X), .Z0_f (new_AGEMA_signal_4512), .Z1_t (new_AGEMA_signal_4513), .Z1_f (new_AGEMA_signal_4514) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS02ser_mux_inst_0_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS02ser_mux_inst_0_X), .B0_f (new_AGEMA_signal_4512), .B1_t (new_AGEMA_signal_4513), .B1_f (new_AGEMA_signal_4514), .Z0_t (KeyArray_MUX_inS02ser_mux_inst_0_Y), .Z0_f (new_AGEMA_signal_6160), .Z1_t (new_AGEMA_signal_6161), .Z1_f (new_AGEMA_signal_6162) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS02ser_mux_inst_0_XOR2_U1 ( .A0_t (KeyArray_MUX_inS02ser_mux_inst_0_Y), .A0_f (new_AGEMA_signal_6160), .A1_t (new_AGEMA_signal_6161), .A1_f (new_AGEMA_signal_6162), .B0_t (key_s0_t[56]), .B0_f (key_s0_f[56]), .B1_t (key_s1_t[56]), .B1_f (key_s1_f[56]), .Z0_t (KeyArray_inS02ser[0]), .Z0_f (new_AGEMA_signal_6934), .Z1_t (new_AGEMA_signal_6935), .Z1_f (new_AGEMA_signal_6936) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS02ser_mux_inst_1_XOR1_U1 ( .A0_t (key_s0_t[57]), .A0_f (key_s0_f[57]), .A1_t (key_s1_t[57]), .A1_f (key_s1_f[57]), .B0_t (KeyArray_outS03ser[1]), .B0_f (new_AGEMA_signal_4518), .B1_t (new_AGEMA_signal_4519), .B1_f (new_AGEMA_signal_4520), .Z0_t (KeyArray_MUX_inS02ser_mux_inst_1_X), .Z0_f (new_AGEMA_signal_4521), .Z1_t (new_AGEMA_signal_4522), .Z1_f (new_AGEMA_signal_4523) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS02ser_mux_inst_1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS02ser_mux_inst_1_X), .B0_f (new_AGEMA_signal_4521), .B1_t (new_AGEMA_signal_4522), .B1_f (new_AGEMA_signal_4523), .Z0_t (KeyArray_MUX_inS02ser_mux_inst_1_Y), .Z0_f (new_AGEMA_signal_6163), .Z1_t (new_AGEMA_signal_6164), .Z1_f (new_AGEMA_signal_6165) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS02ser_mux_inst_1_XOR2_U1 ( .A0_t (KeyArray_MUX_inS02ser_mux_inst_1_Y), .A0_f (new_AGEMA_signal_6163), .A1_t (new_AGEMA_signal_6164), .A1_f (new_AGEMA_signal_6165), .B0_t (key_s0_t[57]), .B0_f (key_s0_f[57]), .B1_t (key_s1_t[57]), .B1_f (key_s1_f[57]), .Z0_t (KeyArray_inS02ser[1]), .Z0_f (new_AGEMA_signal_6937), .Z1_t (new_AGEMA_signal_6938), .Z1_f (new_AGEMA_signal_6939) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS02ser_mux_inst_2_XOR1_U1 ( .A0_t (key_s0_t[58]), .A0_f (key_s0_f[58]), .A1_t (key_s1_t[58]), .A1_f (key_s1_f[58]), .B0_t (KeyArray_outS03ser[2]), .B0_f (new_AGEMA_signal_4527), .B1_t (new_AGEMA_signal_4528), .B1_f (new_AGEMA_signal_4529), .Z0_t (KeyArray_MUX_inS02ser_mux_inst_2_X), .Z0_f (new_AGEMA_signal_4530), .Z1_t (new_AGEMA_signal_4531), .Z1_f (new_AGEMA_signal_4532) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS02ser_mux_inst_2_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS02ser_mux_inst_2_X), .B0_f (new_AGEMA_signal_4530), .B1_t (new_AGEMA_signal_4531), .B1_f (new_AGEMA_signal_4532), .Z0_t (KeyArray_MUX_inS02ser_mux_inst_2_Y), .Z0_f (new_AGEMA_signal_6166), .Z1_t (new_AGEMA_signal_6167), .Z1_f (new_AGEMA_signal_6168) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS02ser_mux_inst_2_XOR2_U1 ( .A0_t (KeyArray_MUX_inS02ser_mux_inst_2_Y), .A0_f (new_AGEMA_signal_6166), .A1_t (new_AGEMA_signal_6167), .A1_f (new_AGEMA_signal_6168), .B0_t (key_s0_t[58]), .B0_f (key_s0_f[58]), .B1_t (key_s1_t[58]), .B1_f (key_s1_f[58]), .Z0_t (KeyArray_inS02ser[2]), .Z0_f (new_AGEMA_signal_6940), .Z1_t (new_AGEMA_signal_6941), .Z1_f (new_AGEMA_signal_6942) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS02ser_mux_inst_3_XOR1_U1 ( .A0_t (key_s0_t[59]), .A0_f (key_s0_f[59]), .A1_t (key_s1_t[59]), .A1_f (key_s1_f[59]), .B0_t (KeyArray_outS03ser[3]), .B0_f (new_AGEMA_signal_4536), .B1_t (new_AGEMA_signal_4537), .B1_f (new_AGEMA_signal_4538), .Z0_t (KeyArray_MUX_inS02ser_mux_inst_3_X), .Z0_f (new_AGEMA_signal_4539), .Z1_t (new_AGEMA_signal_4540), .Z1_f (new_AGEMA_signal_4541) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS02ser_mux_inst_3_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS02ser_mux_inst_3_X), .B0_f (new_AGEMA_signal_4539), .B1_t (new_AGEMA_signal_4540), .B1_f (new_AGEMA_signal_4541), .Z0_t (KeyArray_MUX_inS02ser_mux_inst_3_Y), .Z0_f (new_AGEMA_signal_6169), .Z1_t (new_AGEMA_signal_6170), .Z1_f (new_AGEMA_signal_6171) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS02ser_mux_inst_3_XOR2_U1 ( .A0_t (KeyArray_MUX_inS02ser_mux_inst_3_Y), .A0_f (new_AGEMA_signal_6169), .A1_t (new_AGEMA_signal_6170), .A1_f (new_AGEMA_signal_6171), .B0_t (key_s0_t[59]), .B0_f (key_s0_f[59]), .B1_t (key_s1_t[59]), .B1_f (key_s1_f[59]), .Z0_t (KeyArray_inS02ser[3]), .Z0_f (new_AGEMA_signal_6943), .Z1_t (new_AGEMA_signal_6944), .Z1_f (new_AGEMA_signal_6945) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS02ser_mux_inst_4_XOR1_U1 ( .A0_t (key_s0_t[60]), .A0_f (key_s0_f[60]), .A1_t (key_s1_t[60]), .A1_f (key_s1_f[60]), .B0_t (KeyArray_outS03ser[4]), .B0_f (new_AGEMA_signal_4545), .B1_t (new_AGEMA_signal_4546), .B1_f (new_AGEMA_signal_4547), .Z0_t (KeyArray_MUX_inS02ser_mux_inst_4_X), .Z0_f (new_AGEMA_signal_4548), .Z1_t (new_AGEMA_signal_4549), .Z1_f (new_AGEMA_signal_4550) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS02ser_mux_inst_4_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS02ser_mux_inst_4_X), .B0_f (new_AGEMA_signal_4548), .B1_t (new_AGEMA_signal_4549), .B1_f (new_AGEMA_signal_4550), .Z0_t (KeyArray_MUX_inS02ser_mux_inst_4_Y), .Z0_f (new_AGEMA_signal_6172), .Z1_t (new_AGEMA_signal_6173), .Z1_f (new_AGEMA_signal_6174) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS02ser_mux_inst_4_XOR2_U1 ( .A0_t (KeyArray_MUX_inS02ser_mux_inst_4_Y), .A0_f (new_AGEMA_signal_6172), .A1_t (new_AGEMA_signal_6173), .A1_f (new_AGEMA_signal_6174), .B0_t (key_s0_t[60]), .B0_f (key_s0_f[60]), .B1_t (key_s1_t[60]), .B1_f (key_s1_f[60]), .Z0_t (KeyArray_inS02ser[4]), .Z0_f (new_AGEMA_signal_6946), .Z1_t (new_AGEMA_signal_6947), .Z1_f (new_AGEMA_signal_6948) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS02ser_mux_inst_5_XOR1_U1 ( .A0_t (key_s0_t[61]), .A0_f (key_s0_f[61]), .A1_t (key_s1_t[61]), .A1_f (key_s1_f[61]), .B0_t (KeyArray_outS03ser[5]), .B0_f (new_AGEMA_signal_4554), .B1_t (new_AGEMA_signal_4555), .B1_f (new_AGEMA_signal_4556), .Z0_t (KeyArray_MUX_inS02ser_mux_inst_5_X), .Z0_f (new_AGEMA_signal_4557), .Z1_t (new_AGEMA_signal_4558), .Z1_f (new_AGEMA_signal_4559) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS02ser_mux_inst_5_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS02ser_mux_inst_5_X), .B0_f (new_AGEMA_signal_4557), .B1_t (new_AGEMA_signal_4558), .B1_f (new_AGEMA_signal_4559), .Z0_t (KeyArray_MUX_inS02ser_mux_inst_5_Y), .Z0_f (new_AGEMA_signal_6175), .Z1_t (new_AGEMA_signal_6176), .Z1_f (new_AGEMA_signal_6177) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS02ser_mux_inst_5_XOR2_U1 ( .A0_t (KeyArray_MUX_inS02ser_mux_inst_5_Y), .A0_f (new_AGEMA_signal_6175), .A1_t (new_AGEMA_signal_6176), .A1_f (new_AGEMA_signal_6177), .B0_t (key_s0_t[61]), .B0_f (key_s0_f[61]), .B1_t (key_s1_t[61]), .B1_f (key_s1_f[61]), .Z0_t (KeyArray_inS02ser[5]), .Z0_f (new_AGEMA_signal_6949), .Z1_t (new_AGEMA_signal_6950), .Z1_f (new_AGEMA_signal_6951) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS02ser_mux_inst_6_XOR1_U1 ( .A0_t (key_s0_t[62]), .A0_f (key_s0_f[62]), .A1_t (key_s1_t[62]), .A1_f (key_s1_f[62]), .B0_t (KeyArray_outS03ser[6]), .B0_f (new_AGEMA_signal_4563), .B1_t (new_AGEMA_signal_4564), .B1_f (new_AGEMA_signal_4565), .Z0_t (KeyArray_MUX_inS02ser_mux_inst_6_X), .Z0_f (new_AGEMA_signal_4566), .Z1_t (new_AGEMA_signal_4567), .Z1_f (new_AGEMA_signal_4568) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS02ser_mux_inst_6_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS02ser_mux_inst_6_X), .B0_f (new_AGEMA_signal_4566), .B1_t (new_AGEMA_signal_4567), .B1_f (new_AGEMA_signal_4568), .Z0_t (KeyArray_MUX_inS02ser_mux_inst_6_Y), .Z0_f (new_AGEMA_signal_6178), .Z1_t (new_AGEMA_signal_6179), .Z1_f (new_AGEMA_signal_6180) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS02ser_mux_inst_6_XOR2_U1 ( .A0_t (KeyArray_MUX_inS02ser_mux_inst_6_Y), .A0_f (new_AGEMA_signal_6178), .A1_t (new_AGEMA_signal_6179), .A1_f (new_AGEMA_signal_6180), .B0_t (key_s0_t[62]), .B0_f (key_s0_f[62]), .B1_t (key_s1_t[62]), .B1_f (key_s1_f[62]), .Z0_t (KeyArray_inS02ser[6]), .Z0_f (new_AGEMA_signal_6952), .Z1_t (new_AGEMA_signal_6953), .Z1_f (new_AGEMA_signal_6954) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS02ser_mux_inst_7_XOR1_U1 ( .A0_t (key_s0_t[63]), .A0_f (key_s0_f[63]), .A1_t (key_s1_t[63]), .A1_f (key_s1_f[63]), .B0_t (KeyArray_outS03ser[7]), .B0_f (new_AGEMA_signal_4572), .B1_t (new_AGEMA_signal_4573), .B1_f (new_AGEMA_signal_4574), .Z0_t (KeyArray_MUX_inS02ser_mux_inst_7_X), .Z0_f (new_AGEMA_signal_4575), .Z1_t (new_AGEMA_signal_4576), .Z1_f (new_AGEMA_signal_4577) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS02ser_mux_inst_7_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS02ser_mux_inst_7_X), .B0_f (new_AGEMA_signal_4575), .B1_t (new_AGEMA_signal_4576), .B1_f (new_AGEMA_signal_4577), .Z0_t (KeyArray_MUX_inS02ser_mux_inst_7_Y), .Z0_f (new_AGEMA_signal_6181), .Z1_t (new_AGEMA_signal_6182), .Z1_f (new_AGEMA_signal_6183) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS02ser_mux_inst_7_XOR2_U1 ( .A0_t (KeyArray_MUX_inS02ser_mux_inst_7_Y), .A0_f (new_AGEMA_signal_6181), .A1_t (new_AGEMA_signal_6182), .A1_f (new_AGEMA_signal_6183), .B0_t (key_s0_t[63]), .B0_f (key_s0_f[63]), .B1_t (key_s1_t[63]), .B1_f (key_s1_f[63]), .Z0_t (KeyArray_inS02ser[7]), .Z0_f (new_AGEMA_signal_6955), .Z1_t (new_AGEMA_signal_6956), .Z1_f (new_AGEMA_signal_6957) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS03ser_mux_inst_0_XOR1_U1 ( .A0_t (key_s0_t[24]), .A0_f (key_s0_f[24]), .A1_t (key_s1_t[24]), .A1_f (key_s1_f[24]), .B0_t (KeyArray_outS10ser[0]), .B0_f (new_AGEMA_signal_4581), .B1_t (new_AGEMA_signal_4582), .B1_f (new_AGEMA_signal_4583), .Z0_t (KeyArray_MUX_inS03ser_mux_inst_0_X), .Z0_f (new_AGEMA_signal_4584), .Z1_t (new_AGEMA_signal_4585), .Z1_f (new_AGEMA_signal_4586) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS03ser_mux_inst_0_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS03ser_mux_inst_0_X), .B0_f (new_AGEMA_signal_4584), .B1_t (new_AGEMA_signal_4585), .B1_f (new_AGEMA_signal_4586), .Z0_t (KeyArray_MUX_inS03ser_mux_inst_0_Y), .Z0_f (new_AGEMA_signal_6184), .Z1_t (new_AGEMA_signal_6185), .Z1_f (new_AGEMA_signal_6186) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS03ser_mux_inst_0_XOR2_U1 ( .A0_t (KeyArray_MUX_inS03ser_mux_inst_0_Y), .A0_f (new_AGEMA_signal_6184), .A1_t (new_AGEMA_signal_6185), .A1_f (new_AGEMA_signal_6186), .B0_t (key_s0_t[24]), .B0_f (key_s0_f[24]), .B1_t (key_s1_t[24]), .B1_f (key_s1_f[24]), .Z0_t (KeyArray_inS03ser[0]), .Z0_f (new_AGEMA_signal_6958), .Z1_t (new_AGEMA_signal_6959), .Z1_f (new_AGEMA_signal_6960) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS03ser_mux_inst_1_XOR1_U1 ( .A0_t (key_s0_t[25]), .A0_f (key_s0_f[25]), .A1_t (key_s1_t[25]), .A1_f (key_s1_f[25]), .B0_t (KeyArray_outS10ser[1]), .B0_f (new_AGEMA_signal_4590), .B1_t (new_AGEMA_signal_4591), .B1_f (new_AGEMA_signal_4592), .Z0_t (KeyArray_MUX_inS03ser_mux_inst_1_X), .Z0_f (new_AGEMA_signal_4593), .Z1_t (new_AGEMA_signal_4594), .Z1_f (new_AGEMA_signal_4595) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS03ser_mux_inst_1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS03ser_mux_inst_1_X), .B0_f (new_AGEMA_signal_4593), .B1_t (new_AGEMA_signal_4594), .B1_f (new_AGEMA_signal_4595), .Z0_t (KeyArray_MUX_inS03ser_mux_inst_1_Y), .Z0_f (new_AGEMA_signal_6187), .Z1_t (new_AGEMA_signal_6188), .Z1_f (new_AGEMA_signal_6189) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS03ser_mux_inst_1_XOR2_U1 ( .A0_t (KeyArray_MUX_inS03ser_mux_inst_1_Y), .A0_f (new_AGEMA_signal_6187), .A1_t (new_AGEMA_signal_6188), .A1_f (new_AGEMA_signal_6189), .B0_t (key_s0_t[25]), .B0_f (key_s0_f[25]), .B1_t (key_s1_t[25]), .B1_f (key_s1_f[25]), .Z0_t (KeyArray_inS03ser[1]), .Z0_f (new_AGEMA_signal_6961), .Z1_t (new_AGEMA_signal_6962), .Z1_f (new_AGEMA_signal_6963) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS03ser_mux_inst_2_XOR1_U1 ( .A0_t (key_s0_t[26]), .A0_f (key_s0_f[26]), .A1_t (key_s1_t[26]), .A1_f (key_s1_f[26]), .B0_t (KeyArray_outS10ser[2]), .B0_f (new_AGEMA_signal_4599), .B1_t (new_AGEMA_signal_4600), .B1_f (new_AGEMA_signal_4601), .Z0_t (KeyArray_MUX_inS03ser_mux_inst_2_X), .Z0_f (new_AGEMA_signal_4602), .Z1_t (new_AGEMA_signal_4603), .Z1_f (new_AGEMA_signal_4604) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS03ser_mux_inst_2_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS03ser_mux_inst_2_X), .B0_f (new_AGEMA_signal_4602), .B1_t (new_AGEMA_signal_4603), .B1_f (new_AGEMA_signal_4604), .Z0_t (KeyArray_MUX_inS03ser_mux_inst_2_Y), .Z0_f (new_AGEMA_signal_6190), .Z1_t (new_AGEMA_signal_6191), .Z1_f (new_AGEMA_signal_6192) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS03ser_mux_inst_2_XOR2_U1 ( .A0_t (KeyArray_MUX_inS03ser_mux_inst_2_Y), .A0_f (new_AGEMA_signal_6190), .A1_t (new_AGEMA_signal_6191), .A1_f (new_AGEMA_signal_6192), .B0_t (key_s0_t[26]), .B0_f (key_s0_f[26]), .B1_t (key_s1_t[26]), .B1_f (key_s1_f[26]), .Z0_t (KeyArray_inS03ser[2]), .Z0_f (new_AGEMA_signal_6964), .Z1_t (new_AGEMA_signal_6965), .Z1_f (new_AGEMA_signal_6966) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS03ser_mux_inst_3_XOR1_U1 ( .A0_t (key_s0_t[27]), .A0_f (key_s0_f[27]), .A1_t (key_s1_t[27]), .A1_f (key_s1_f[27]), .B0_t (KeyArray_outS10ser[3]), .B0_f (new_AGEMA_signal_4608), .B1_t (new_AGEMA_signal_4609), .B1_f (new_AGEMA_signal_4610), .Z0_t (KeyArray_MUX_inS03ser_mux_inst_3_X), .Z0_f (new_AGEMA_signal_4611), .Z1_t (new_AGEMA_signal_4612), .Z1_f (new_AGEMA_signal_4613) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS03ser_mux_inst_3_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS03ser_mux_inst_3_X), .B0_f (new_AGEMA_signal_4611), .B1_t (new_AGEMA_signal_4612), .B1_f (new_AGEMA_signal_4613), .Z0_t (KeyArray_MUX_inS03ser_mux_inst_3_Y), .Z0_f (new_AGEMA_signal_6193), .Z1_t (new_AGEMA_signal_6194), .Z1_f (new_AGEMA_signal_6195) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS03ser_mux_inst_3_XOR2_U1 ( .A0_t (KeyArray_MUX_inS03ser_mux_inst_3_Y), .A0_f (new_AGEMA_signal_6193), .A1_t (new_AGEMA_signal_6194), .A1_f (new_AGEMA_signal_6195), .B0_t (key_s0_t[27]), .B0_f (key_s0_f[27]), .B1_t (key_s1_t[27]), .B1_f (key_s1_f[27]), .Z0_t (KeyArray_inS03ser[3]), .Z0_f (new_AGEMA_signal_6967), .Z1_t (new_AGEMA_signal_6968), .Z1_f (new_AGEMA_signal_6969) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS03ser_mux_inst_4_XOR1_U1 ( .A0_t (key_s0_t[28]), .A0_f (key_s0_f[28]), .A1_t (key_s1_t[28]), .A1_f (key_s1_f[28]), .B0_t (KeyArray_outS10ser[4]), .B0_f (new_AGEMA_signal_4617), .B1_t (new_AGEMA_signal_4618), .B1_f (new_AGEMA_signal_4619), .Z0_t (KeyArray_MUX_inS03ser_mux_inst_4_X), .Z0_f (new_AGEMA_signal_4620), .Z1_t (new_AGEMA_signal_4621), .Z1_f (new_AGEMA_signal_4622) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS03ser_mux_inst_4_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS03ser_mux_inst_4_X), .B0_f (new_AGEMA_signal_4620), .B1_t (new_AGEMA_signal_4621), .B1_f (new_AGEMA_signal_4622), .Z0_t (KeyArray_MUX_inS03ser_mux_inst_4_Y), .Z0_f (new_AGEMA_signal_6196), .Z1_t (new_AGEMA_signal_6197), .Z1_f (new_AGEMA_signal_6198) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS03ser_mux_inst_4_XOR2_U1 ( .A0_t (KeyArray_MUX_inS03ser_mux_inst_4_Y), .A0_f (new_AGEMA_signal_6196), .A1_t (new_AGEMA_signal_6197), .A1_f (new_AGEMA_signal_6198), .B0_t (key_s0_t[28]), .B0_f (key_s0_f[28]), .B1_t (key_s1_t[28]), .B1_f (key_s1_f[28]), .Z0_t (KeyArray_inS03ser[4]), .Z0_f (new_AGEMA_signal_6970), .Z1_t (new_AGEMA_signal_6971), .Z1_f (new_AGEMA_signal_6972) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS03ser_mux_inst_5_XOR1_U1 ( .A0_t (key_s0_t[29]), .A0_f (key_s0_f[29]), .A1_t (key_s1_t[29]), .A1_f (key_s1_f[29]), .B0_t (KeyArray_outS10ser[5]), .B0_f (new_AGEMA_signal_4626), .B1_t (new_AGEMA_signal_4627), .B1_f (new_AGEMA_signal_4628), .Z0_t (KeyArray_MUX_inS03ser_mux_inst_5_X), .Z0_f (new_AGEMA_signal_4629), .Z1_t (new_AGEMA_signal_4630), .Z1_f (new_AGEMA_signal_4631) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS03ser_mux_inst_5_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS03ser_mux_inst_5_X), .B0_f (new_AGEMA_signal_4629), .B1_t (new_AGEMA_signal_4630), .B1_f (new_AGEMA_signal_4631), .Z0_t (KeyArray_MUX_inS03ser_mux_inst_5_Y), .Z0_f (new_AGEMA_signal_6199), .Z1_t (new_AGEMA_signal_6200), .Z1_f (new_AGEMA_signal_6201) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS03ser_mux_inst_5_XOR2_U1 ( .A0_t (KeyArray_MUX_inS03ser_mux_inst_5_Y), .A0_f (new_AGEMA_signal_6199), .A1_t (new_AGEMA_signal_6200), .A1_f (new_AGEMA_signal_6201), .B0_t (key_s0_t[29]), .B0_f (key_s0_f[29]), .B1_t (key_s1_t[29]), .B1_f (key_s1_f[29]), .Z0_t (KeyArray_inS03ser[5]), .Z0_f (new_AGEMA_signal_6973), .Z1_t (new_AGEMA_signal_6974), .Z1_f (new_AGEMA_signal_6975) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS03ser_mux_inst_6_XOR1_U1 ( .A0_t (key_s0_t[30]), .A0_f (key_s0_f[30]), .A1_t (key_s1_t[30]), .A1_f (key_s1_f[30]), .B0_t (KeyArray_outS10ser[6]), .B0_f (new_AGEMA_signal_4635), .B1_t (new_AGEMA_signal_4636), .B1_f (new_AGEMA_signal_4637), .Z0_t (KeyArray_MUX_inS03ser_mux_inst_6_X), .Z0_f (new_AGEMA_signal_4638), .Z1_t (new_AGEMA_signal_4639), .Z1_f (new_AGEMA_signal_4640) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS03ser_mux_inst_6_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS03ser_mux_inst_6_X), .B0_f (new_AGEMA_signal_4638), .B1_t (new_AGEMA_signal_4639), .B1_f (new_AGEMA_signal_4640), .Z0_t (KeyArray_MUX_inS03ser_mux_inst_6_Y), .Z0_f (new_AGEMA_signal_6202), .Z1_t (new_AGEMA_signal_6203), .Z1_f (new_AGEMA_signal_6204) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS03ser_mux_inst_6_XOR2_U1 ( .A0_t (KeyArray_MUX_inS03ser_mux_inst_6_Y), .A0_f (new_AGEMA_signal_6202), .A1_t (new_AGEMA_signal_6203), .A1_f (new_AGEMA_signal_6204), .B0_t (key_s0_t[30]), .B0_f (key_s0_f[30]), .B1_t (key_s1_t[30]), .B1_f (key_s1_f[30]), .Z0_t (KeyArray_inS03ser[6]), .Z0_f (new_AGEMA_signal_6976), .Z1_t (new_AGEMA_signal_6977), .Z1_f (new_AGEMA_signal_6978) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS03ser_mux_inst_7_XOR1_U1 ( .A0_t (key_s0_t[31]), .A0_f (key_s0_f[31]), .A1_t (key_s1_t[31]), .A1_f (key_s1_f[31]), .B0_t (KeyArray_outS10ser[7]), .B0_f (new_AGEMA_signal_4644), .B1_t (new_AGEMA_signal_4645), .B1_f (new_AGEMA_signal_4646), .Z0_t (KeyArray_MUX_inS03ser_mux_inst_7_X), .Z0_f (new_AGEMA_signal_4647), .Z1_t (new_AGEMA_signal_4648), .Z1_f (new_AGEMA_signal_4649) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS03ser_mux_inst_7_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS03ser_mux_inst_7_X), .B0_f (new_AGEMA_signal_4647), .B1_t (new_AGEMA_signal_4648), .B1_f (new_AGEMA_signal_4649), .Z0_t (KeyArray_MUX_inS03ser_mux_inst_7_Y), .Z0_f (new_AGEMA_signal_6205), .Z1_t (new_AGEMA_signal_6206), .Z1_f (new_AGEMA_signal_6207) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS03ser_mux_inst_7_XOR2_U1 ( .A0_t (KeyArray_MUX_inS03ser_mux_inst_7_Y), .A0_f (new_AGEMA_signal_6205), .A1_t (new_AGEMA_signal_6206), .A1_f (new_AGEMA_signal_6207), .B0_t (key_s0_t[31]), .B0_f (key_s0_f[31]), .B1_t (key_s1_t[31]), .B1_f (key_s1_f[31]), .Z0_t (KeyArray_inS03ser[7]), .Z0_f (new_AGEMA_signal_6979), .Z1_t (new_AGEMA_signal_6980), .Z1_f (new_AGEMA_signal_6981) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS10ser_mux_inst_0_XOR1_U1 ( .A0_t (key_s0_t[112]), .A0_f (key_s0_f[112]), .A1_t (key_s1_t[112]), .A1_f (key_s1_f[112]), .B0_t (KeyArray_outS11ser[0]), .B0_f (new_AGEMA_signal_4653), .B1_t (new_AGEMA_signal_4654), .B1_f (new_AGEMA_signal_4655), .Z0_t (KeyArray_MUX_inS10ser_mux_inst_0_X), .Z0_f (new_AGEMA_signal_4656), .Z1_t (new_AGEMA_signal_4657), .Z1_f (new_AGEMA_signal_4658) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS10ser_mux_inst_0_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS10ser_mux_inst_0_X), .B0_f (new_AGEMA_signal_4656), .B1_t (new_AGEMA_signal_4657), .B1_f (new_AGEMA_signal_4658), .Z0_t (KeyArray_MUX_inS10ser_mux_inst_0_Y), .Z0_f (new_AGEMA_signal_6208), .Z1_t (new_AGEMA_signal_6209), .Z1_f (new_AGEMA_signal_6210) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS10ser_mux_inst_0_XOR2_U1 ( .A0_t (KeyArray_MUX_inS10ser_mux_inst_0_Y), .A0_f (new_AGEMA_signal_6208), .A1_t (new_AGEMA_signal_6209), .A1_f (new_AGEMA_signal_6210), .B0_t (key_s0_t[112]), .B0_f (key_s0_f[112]), .B1_t (key_s1_t[112]), .B1_f (key_s1_f[112]), .Z0_t (KeyArray_inS10ser[0]), .Z0_f (new_AGEMA_signal_6982), .Z1_t (new_AGEMA_signal_6983), .Z1_f (new_AGEMA_signal_6984) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS10ser_mux_inst_1_XOR1_U1 ( .A0_t (key_s0_t[113]), .A0_f (key_s0_f[113]), .A1_t (key_s1_t[113]), .A1_f (key_s1_f[113]), .B0_t (KeyArray_outS11ser[1]), .B0_f (new_AGEMA_signal_4662), .B1_t (new_AGEMA_signal_4663), .B1_f (new_AGEMA_signal_4664), .Z0_t (KeyArray_MUX_inS10ser_mux_inst_1_X), .Z0_f (new_AGEMA_signal_4665), .Z1_t (new_AGEMA_signal_4666), .Z1_f (new_AGEMA_signal_4667) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS10ser_mux_inst_1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS10ser_mux_inst_1_X), .B0_f (new_AGEMA_signal_4665), .B1_t (new_AGEMA_signal_4666), .B1_f (new_AGEMA_signal_4667), .Z0_t (KeyArray_MUX_inS10ser_mux_inst_1_Y), .Z0_f (new_AGEMA_signal_6211), .Z1_t (new_AGEMA_signal_6212), .Z1_f (new_AGEMA_signal_6213) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS10ser_mux_inst_1_XOR2_U1 ( .A0_t (KeyArray_MUX_inS10ser_mux_inst_1_Y), .A0_f (new_AGEMA_signal_6211), .A1_t (new_AGEMA_signal_6212), .A1_f (new_AGEMA_signal_6213), .B0_t (key_s0_t[113]), .B0_f (key_s0_f[113]), .B1_t (key_s1_t[113]), .B1_f (key_s1_f[113]), .Z0_t (KeyArray_inS10ser[1]), .Z0_f (new_AGEMA_signal_6985), .Z1_t (new_AGEMA_signal_6986), .Z1_f (new_AGEMA_signal_6987) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS10ser_mux_inst_2_XOR1_U1 ( .A0_t (key_s0_t[114]), .A0_f (key_s0_f[114]), .A1_t (key_s1_t[114]), .A1_f (key_s1_f[114]), .B0_t (KeyArray_outS11ser[2]), .B0_f (new_AGEMA_signal_4671), .B1_t (new_AGEMA_signal_4672), .B1_f (new_AGEMA_signal_4673), .Z0_t (KeyArray_MUX_inS10ser_mux_inst_2_X), .Z0_f (new_AGEMA_signal_4674), .Z1_t (new_AGEMA_signal_4675), .Z1_f (new_AGEMA_signal_4676) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS10ser_mux_inst_2_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS10ser_mux_inst_2_X), .B0_f (new_AGEMA_signal_4674), .B1_t (new_AGEMA_signal_4675), .B1_f (new_AGEMA_signal_4676), .Z0_t (KeyArray_MUX_inS10ser_mux_inst_2_Y), .Z0_f (new_AGEMA_signal_6214), .Z1_t (new_AGEMA_signal_6215), .Z1_f (new_AGEMA_signal_6216) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS10ser_mux_inst_2_XOR2_U1 ( .A0_t (KeyArray_MUX_inS10ser_mux_inst_2_Y), .A0_f (new_AGEMA_signal_6214), .A1_t (new_AGEMA_signal_6215), .A1_f (new_AGEMA_signal_6216), .B0_t (key_s0_t[114]), .B0_f (key_s0_f[114]), .B1_t (key_s1_t[114]), .B1_f (key_s1_f[114]), .Z0_t (KeyArray_inS10ser[2]), .Z0_f (new_AGEMA_signal_6988), .Z1_t (new_AGEMA_signal_6989), .Z1_f (new_AGEMA_signal_6990) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS10ser_mux_inst_3_XOR1_U1 ( .A0_t (key_s0_t[115]), .A0_f (key_s0_f[115]), .A1_t (key_s1_t[115]), .A1_f (key_s1_f[115]), .B0_t (KeyArray_outS11ser[3]), .B0_f (new_AGEMA_signal_4680), .B1_t (new_AGEMA_signal_4681), .B1_f (new_AGEMA_signal_4682), .Z0_t (KeyArray_MUX_inS10ser_mux_inst_3_X), .Z0_f (new_AGEMA_signal_4683), .Z1_t (new_AGEMA_signal_4684), .Z1_f (new_AGEMA_signal_4685) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS10ser_mux_inst_3_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS10ser_mux_inst_3_X), .B0_f (new_AGEMA_signal_4683), .B1_t (new_AGEMA_signal_4684), .B1_f (new_AGEMA_signal_4685), .Z0_t (KeyArray_MUX_inS10ser_mux_inst_3_Y), .Z0_f (new_AGEMA_signal_6217), .Z1_t (new_AGEMA_signal_6218), .Z1_f (new_AGEMA_signal_6219) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS10ser_mux_inst_3_XOR2_U1 ( .A0_t (KeyArray_MUX_inS10ser_mux_inst_3_Y), .A0_f (new_AGEMA_signal_6217), .A1_t (new_AGEMA_signal_6218), .A1_f (new_AGEMA_signal_6219), .B0_t (key_s0_t[115]), .B0_f (key_s0_f[115]), .B1_t (key_s1_t[115]), .B1_f (key_s1_f[115]), .Z0_t (KeyArray_inS10ser[3]), .Z0_f (new_AGEMA_signal_6991), .Z1_t (new_AGEMA_signal_6992), .Z1_f (new_AGEMA_signal_6993) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS10ser_mux_inst_4_XOR1_U1 ( .A0_t (key_s0_t[116]), .A0_f (key_s0_f[116]), .A1_t (key_s1_t[116]), .A1_f (key_s1_f[116]), .B0_t (KeyArray_outS11ser[4]), .B0_f (new_AGEMA_signal_4689), .B1_t (new_AGEMA_signal_4690), .B1_f (new_AGEMA_signal_4691), .Z0_t (KeyArray_MUX_inS10ser_mux_inst_4_X), .Z0_f (new_AGEMA_signal_4692), .Z1_t (new_AGEMA_signal_4693), .Z1_f (new_AGEMA_signal_4694) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS10ser_mux_inst_4_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS10ser_mux_inst_4_X), .B0_f (new_AGEMA_signal_4692), .B1_t (new_AGEMA_signal_4693), .B1_f (new_AGEMA_signal_4694), .Z0_t (KeyArray_MUX_inS10ser_mux_inst_4_Y), .Z0_f (new_AGEMA_signal_6220), .Z1_t (new_AGEMA_signal_6221), .Z1_f (new_AGEMA_signal_6222) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS10ser_mux_inst_4_XOR2_U1 ( .A0_t (KeyArray_MUX_inS10ser_mux_inst_4_Y), .A0_f (new_AGEMA_signal_6220), .A1_t (new_AGEMA_signal_6221), .A1_f (new_AGEMA_signal_6222), .B0_t (key_s0_t[116]), .B0_f (key_s0_f[116]), .B1_t (key_s1_t[116]), .B1_f (key_s1_f[116]), .Z0_t (KeyArray_inS10ser[4]), .Z0_f (new_AGEMA_signal_6994), .Z1_t (new_AGEMA_signal_6995), .Z1_f (new_AGEMA_signal_6996) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS10ser_mux_inst_5_XOR1_U1 ( .A0_t (key_s0_t[117]), .A0_f (key_s0_f[117]), .A1_t (key_s1_t[117]), .A1_f (key_s1_f[117]), .B0_t (KeyArray_outS11ser[5]), .B0_f (new_AGEMA_signal_4698), .B1_t (new_AGEMA_signal_4699), .B1_f (new_AGEMA_signal_4700), .Z0_t (KeyArray_MUX_inS10ser_mux_inst_5_X), .Z0_f (new_AGEMA_signal_4701), .Z1_t (new_AGEMA_signal_4702), .Z1_f (new_AGEMA_signal_4703) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS10ser_mux_inst_5_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS10ser_mux_inst_5_X), .B0_f (new_AGEMA_signal_4701), .B1_t (new_AGEMA_signal_4702), .B1_f (new_AGEMA_signal_4703), .Z0_t (KeyArray_MUX_inS10ser_mux_inst_5_Y), .Z0_f (new_AGEMA_signal_6223), .Z1_t (new_AGEMA_signal_6224), .Z1_f (new_AGEMA_signal_6225) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS10ser_mux_inst_5_XOR2_U1 ( .A0_t (KeyArray_MUX_inS10ser_mux_inst_5_Y), .A0_f (new_AGEMA_signal_6223), .A1_t (new_AGEMA_signal_6224), .A1_f (new_AGEMA_signal_6225), .B0_t (key_s0_t[117]), .B0_f (key_s0_f[117]), .B1_t (key_s1_t[117]), .B1_f (key_s1_f[117]), .Z0_t (KeyArray_inS10ser[5]), .Z0_f (new_AGEMA_signal_6997), .Z1_t (new_AGEMA_signal_6998), .Z1_f (new_AGEMA_signal_6999) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS10ser_mux_inst_6_XOR1_U1 ( .A0_t (key_s0_t[118]), .A0_f (key_s0_f[118]), .A1_t (key_s1_t[118]), .A1_f (key_s1_f[118]), .B0_t (KeyArray_outS11ser[6]), .B0_f (new_AGEMA_signal_4707), .B1_t (new_AGEMA_signal_4708), .B1_f (new_AGEMA_signal_4709), .Z0_t (KeyArray_MUX_inS10ser_mux_inst_6_X), .Z0_f (new_AGEMA_signal_4710), .Z1_t (new_AGEMA_signal_4711), .Z1_f (new_AGEMA_signal_4712) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS10ser_mux_inst_6_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS10ser_mux_inst_6_X), .B0_f (new_AGEMA_signal_4710), .B1_t (new_AGEMA_signal_4711), .B1_f (new_AGEMA_signal_4712), .Z0_t (KeyArray_MUX_inS10ser_mux_inst_6_Y), .Z0_f (new_AGEMA_signal_6226), .Z1_t (new_AGEMA_signal_6227), .Z1_f (new_AGEMA_signal_6228) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS10ser_mux_inst_6_XOR2_U1 ( .A0_t (KeyArray_MUX_inS10ser_mux_inst_6_Y), .A0_f (new_AGEMA_signal_6226), .A1_t (new_AGEMA_signal_6227), .A1_f (new_AGEMA_signal_6228), .B0_t (key_s0_t[118]), .B0_f (key_s0_f[118]), .B1_t (key_s1_t[118]), .B1_f (key_s1_f[118]), .Z0_t (KeyArray_inS10ser[6]), .Z0_f (new_AGEMA_signal_7000), .Z1_t (new_AGEMA_signal_7001), .Z1_f (new_AGEMA_signal_7002) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS10ser_mux_inst_7_XOR1_U1 ( .A0_t (key_s0_t[119]), .A0_f (key_s0_f[119]), .A1_t (key_s1_t[119]), .A1_f (key_s1_f[119]), .B0_t (KeyArray_outS11ser[7]), .B0_f (new_AGEMA_signal_4716), .B1_t (new_AGEMA_signal_4717), .B1_f (new_AGEMA_signal_4718), .Z0_t (KeyArray_MUX_inS10ser_mux_inst_7_X), .Z0_f (new_AGEMA_signal_4719), .Z1_t (new_AGEMA_signal_4720), .Z1_f (new_AGEMA_signal_4721) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS10ser_mux_inst_7_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS10ser_mux_inst_7_X), .B0_f (new_AGEMA_signal_4719), .B1_t (new_AGEMA_signal_4720), .B1_f (new_AGEMA_signal_4721), .Z0_t (KeyArray_MUX_inS10ser_mux_inst_7_Y), .Z0_f (new_AGEMA_signal_6229), .Z1_t (new_AGEMA_signal_6230), .Z1_f (new_AGEMA_signal_6231) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS10ser_mux_inst_7_XOR2_U1 ( .A0_t (KeyArray_MUX_inS10ser_mux_inst_7_Y), .A0_f (new_AGEMA_signal_6229), .A1_t (new_AGEMA_signal_6230), .A1_f (new_AGEMA_signal_6231), .B0_t (key_s0_t[119]), .B0_f (key_s0_f[119]), .B1_t (key_s1_t[119]), .B1_f (key_s1_f[119]), .Z0_t (KeyArray_inS10ser[7]), .Z0_f (new_AGEMA_signal_7003), .Z1_t (new_AGEMA_signal_7004), .Z1_f (new_AGEMA_signal_7005) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS11ser_mux_inst_0_XOR1_U1 ( .A0_t (key_s0_t[80]), .A0_f (key_s0_f[80]), .A1_t (key_s1_t[80]), .A1_f (key_s1_f[80]), .B0_t (KeyArray_outS12ser[0]), .B0_f (new_AGEMA_signal_4725), .B1_t (new_AGEMA_signal_4726), .B1_f (new_AGEMA_signal_4727), .Z0_t (KeyArray_MUX_inS11ser_mux_inst_0_X), .Z0_f (new_AGEMA_signal_4728), .Z1_t (new_AGEMA_signal_4729), .Z1_f (new_AGEMA_signal_4730) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS11ser_mux_inst_0_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS11ser_mux_inst_0_X), .B0_f (new_AGEMA_signal_4728), .B1_t (new_AGEMA_signal_4729), .B1_f (new_AGEMA_signal_4730), .Z0_t (KeyArray_MUX_inS11ser_mux_inst_0_Y), .Z0_f (new_AGEMA_signal_6232), .Z1_t (new_AGEMA_signal_6233), .Z1_f (new_AGEMA_signal_6234) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS11ser_mux_inst_0_XOR2_U1 ( .A0_t (KeyArray_MUX_inS11ser_mux_inst_0_Y), .A0_f (new_AGEMA_signal_6232), .A1_t (new_AGEMA_signal_6233), .A1_f (new_AGEMA_signal_6234), .B0_t (key_s0_t[80]), .B0_f (key_s0_f[80]), .B1_t (key_s1_t[80]), .B1_f (key_s1_f[80]), .Z0_t (KeyArray_inS11ser[0]), .Z0_f (new_AGEMA_signal_7006), .Z1_t (new_AGEMA_signal_7007), .Z1_f (new_AGEMA_signal_7008) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS11ser_mux_inst_1_XOR1_U1 ( .A0_t (key_s0_t[81]), .A0_f (key_s0_f[81]), .A1_t (key_s1_t[81]), .A1_f (key_s1_f[81]), .B0_t (KeyArray_outS12ser[1]), .B0_f (new_AGEMA_signal_4734), .B1_t (new_AGEMA_signal_4735), .B1_f (new_AGEMA_signal_4736), .Z0_t (KeyArray_MUX_inS11ser_mux_inst_1_X), .Z0_f (new_AGEMA_signal_4737), .Z1_t (new_AGEMA_signal_4738), .Z1_f (new_AGEMA_signal_4739) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS11ser_mux_inst_1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS11ser_mux_inst_1_X), .B0_f (new_AGEMA_signal_4737), .B1_t (new_AGEMA_signal_4738), .B1_f (new_AGEMA_signal_4739), .Z0_t (KeyArray_MUX_inS11ser_mux_inst_1_Y), .Z0_f (new_AGEMA_signal_6235), .Z1_t (new_AGEMA_signal_6236), .Z1_f (new_AGEMA_signal_6237) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS11ser_mux_inst_1_XOR2_U1 ( .A0_t (KeyArray_MUX_inS11ser_mux_inst_1_Y), .A0_f (new_AGEMA_signal_6235), .A1_t (new_AGEMA_signal_6236), .A1_f (new_AGEMA_signal_6237), .B0_t (key_s0_t[81]), .B0_f (key_s0_f[81]), .B1_t (key_s1_t[81]), .B1_f (key_s1_f[81]), .Z0_t (KeyArray_inS11ser[1]), .Z0_f (new_AGEMA_signal_7009), .Z1_t (new_AGEMA_signal_7010), .Z1_f (new_AGEMA_signal_7011) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS11ser_mux_inst_2_XOR1_U1 ( .A0_t (key_s0_t[82]), .A0_f (key_s0_f[82]), .A1_t (key_s1_t[82]), .A1_f (key_s1_f[82]), .B0_t (KeyArray_outS12ser[2]), .B0_f (new_AGEMA_signal_4743), .B1_t (new_AGEMA_signal_4744), .B1_f (new_AGEMA_signal_4745), .Z0_t (KeyArray_MUX_inS11ser_mux_inst_2_X), .Z0_f (new_AGEMA_signal_4746), .Z1_t (new_AGEMA_signal_4747), .Z1_f (new_AGEMA_signal_4748) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS11ser_mux_inst_2_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS11ser_mux_inst_2_X), .B0_f (new_AGEMA_signal_4746), .B1_t (new_AGEMA_signal_4747), .B1_f (new_AGEMA_signal_4748), .Z0_t (KeyArray_MUX_inS11ser_mux_inst_2_Y), .Z0_f (new_AGEMA_signal_6238), .Z1_t (new_AGEMA_signal_6239), .Z1_f (new_AGEMA_signal_6240) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS11ser_mux_inst_2_XOR2_U1 ( .A0_t (KeyArray_MUX_inS11ser_mux_inst_2_Y), .A0_f (new_AGEMA_signal_6238), .A1_t (new_AGEMA_signal_6239), .A1_f (new_AGEMA_signal_6240), .B0_t (key_s0_t[82]), .B0_f (key_s0_f[82]), .B1_t (key_s1_t[82]), .B1_f (key_s1_f[82]), .Z0_t (KeyArray_inS11ser[2]), .Z0_f (new_AGEMA_signal_7012), .Z1_t (new_AGEMA_signal_7013), .Z1_f (new_AGEMA_signal_7014) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS11ser_mux_inst_3_XOR1_U1 ( .A0_t (key_s0_t[83]), .A0_f (key_s0_f[83]), .A1_t (key_s1_t[83]), .A1_f (key_s1_f[83]), .B0_t (KeyArray_outS12ser[3]), .B0_f (new_AGEMA_signal_4752), .B1_t (new_AGEMA_signal_4753), .B1_f (new_AGEMA_signal_4754), .Z0_t (KeyArray_MUX_inS11ser_mux_inst_3_X), .Z0_f (new_AGEMA_signal_4755), .Z1_t (new_AGEMA_signal_4756), .Z1_f (new_AGEMA_signal_4757) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS11ser_mux_inst_3_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS11ser_mux_inst_3_X), .B0_f (new_AGEMA_signal_4755), .B1_t (new_AGEMA_signal_4756), .B1_f (new_AGEMA_signal_4757), .Z0_t (KeyArray_MUX_inS11ser_mux_inst_3_Y), .Z0_f (new_AGEMA_signal_6241), .Z1_t (new_AGEMA_signal_6242), .Z1_f (new_AGEMA_signal_6243) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS11ser_mux_inst_3_XOR2_U1 ( .A0_t (KeyArray_MUX_inS11ser_mux_inst_3_Y), .A0_f (new_AGEMA_signal_6241), .A1_t (new_AGEMA_signal_6242), .A1_f (new_AGEMA_signal_6243), .B0_t (key_s0_t[83]), .B0_f (key_s0_f[83]), .B1_t (key_s1_t[83]), .B1_f (key_s1_f[83]), .Z0_t (KeyArray_inS11ser[3]), .Z0_f (new_AGEMA_signal_7015), .Z1_t (new_AGEMA_signal_7016), .Z1_f (new_AGEMA_signal_7017) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS11ser_mux_inst_4_XOR1_U1 ( .A0_t (key_s0_t[84]), .A0_f (key_s0_f[84]), .A1_t (key_s1_t[84]), .A1_f (key_s1_f[84]), .B0_t (KeyArray_outS12ser[4]), .B0_f (new_AGEMA_signal_4761), .B1_t (new_AGEMA_signal_4762), .B1_f (new_AGEMA_signal_4763), .Z0_t (KeyArray_MUX_inS11ser_mux_inst_4_X), .Z0_f (new_AGEMA_signal_4764), .Z1_t (new_AGEMA_signal_4765), .Z1_f (new_AGEMA_signal_4766) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS11ser_mux_inst_4_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS11ser_mux_inst_4_X), .B0_f (new_AGEMA_signal_4764), .B1_t (new_AGEMA_signal_4765), .B1_f (new_AGEMA_signal_4766), .Z0_t (KeyArray_MUX_inS11ser_mux_inst_4_Y), .Z0_f (new_AGEMA_signal_6244), .Z1_t (new_AGEMA_signal_6245), .Z1_f (new_AGEMA_signal_6246) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS11ser_mux_inst_4_XOR2_U1 ( .A0_t (KeyArray_MUX_inS11ser_mux_inst_4_Y), .A0_f (new_AGEMA_signal_6244), .A1_t (new_AGEMA_signal_6245), .A1_f (new_AGEMA_signal_6246), .B0_t (key_s0_t[84]), .B0_f (key_s0_f[84]), .B1_t (key_s1_t[84]), .B1_f (key_s1_f[84]), .Z0_t (KeyArray_inS11ser[4]), .Z0_f (new_AGEMA_signal_7018), .Z1_t (new_AGEMA_signal_7019), .Z1_f (new_AGEMA_signal_7020) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS11ser_mux_inst_5_XOR1_U1 ( .A0_t (key_s0_t[85]), .A0_f (key_s0_f[85]), .A1_t (key_s1_t[85]), .A1_f (key_s1_f[85]), .B0_t (KeyArray_outS12ser[5]), .B0_f (new_AGEMA_signal_4770), .B1_t (new_AGEMA_signal_4771), .B1_f (new_AGEMA_signal_4772), .Z0_t (KeyArray_MUX_inS11ser_mux_inst_5_X), .Z0_f (new_AGEMA_signal_4773), .Z1_t (new_AGEMA_signal_4774), .Z1_f (new_AGEMA_signal_4775) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS11ser_mux_inst_5_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS11ser_mux_inst_5_X), .B0_f (new_AGEMA_signal_4773), .B1_t (new_AGEMA_signal_4774), .B1_f (new_AGEMA_signal_4775), .Z0_t (KeyArray_MUX_inS11ser_mux_inst_5_Y), .Z0_f (new_AGEMA_signal_6247), .Z1_t (new_AGEMA_signal_6248), .Z1_f (new_AGEMA_signal_6249) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS11ser_mux_inst_5_XOR2_U1 ( .A0_t (KeyArray_MUX_inS11ser_mux_inst_5_Y), .A0_f (new_AGEMA_signal_6247), .A1_t (new_AGEMA_signal_6248), .A1_f (new_AGEMA_signal_6249), .B0_t (key_s0_t[85]), .B0_f (key_s0_f[85]), .B1_t (key_s1_t[85]), .B1_f (key_s1_f[85]), .Z0_t (KeyArray_inS11ser[5]), .Z0_f (new_AGEMA_signal_7021), .Z1_t (new_AGEMA_signal_7022), .Z1_f (new_AGEMA_signal_7023) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS11ser_mux_inst_6_XOR1_U1 ( .A0_t (key_s0_t[86]), .A0_f (key_s0_f[86]), .A1_t (key_s1_t[86]), .A1_f (key_s1_f[86]), .B0_t (KeyArray_outS12ser[6]), .B0_f (new_AGEMA_signal_4779), .B1_t (new_AGEMA_signal_4780), .B1_f (new_AGEMA_signal_4781), .Z0_t (KeyArray_MUX_inS11ser_mux_inst_6_X), .Z0_f (new_AGEMA_signal_4782), .Z1_t (new_AGEMA_signal_4783), .Z1_f (new_AGEMA_signal_4784) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS11ser_mux_inst_6_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS11ser_mux_inst_6_X), .B0_f (new_AGEMA_signal_4782), .B1_t (new_AGEMA_signal_4783), .B1_f (new_AGEMA_signal_4784), .Z0_t (KeyArray_MUX_inS11ser_mux_inst_6_Y), .Z0_f (new_AGEMA_signal_6250), .Z1_t (new_AGEMA_signal_6251), .Z1_f (new_AGEMA_signal_6252) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS11ser_mux_inst_6_XOR2_U1 ( .A0_t (KeyArray_MUX_inS11ser_mux_inst_6_Y), .A0_f (new_AGEMA_signal_6250), .A1_t (new_AGEMA_signal_6251), .A1_f (new_AGEMA_signal_6252), .B0_t (key_s0_t[86]), .B0_f (key_s0_f[86]), .B1_t (key_s1_t[86]), .B1_f (key_s1_f[86]), .Z0_t (KeyArray_inS11ser[6]), .Z0_f (new_AGEMA_signal_7024), .Z1_t (new_AGEMA_signal_7025), .Z1_f (new_AGEMA_signal_7026) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS11ser_mux_inst_7_XOR1_U1 ( .A0_t (key_s0_t[87]), .A0_f (key_s0_f[87]), .A1_t (key_s1_t[87]), .A1_f (key_s1_f[87]), .B0_t (KeyArray_outS12ser[7]), .B0_f (new_AGEMA_signal_4788), .B1_t (new_AGEMA_signal_4789), .B1_f (new_AGEMA_signal_4790), .Z0_t (KeyArray_MUX_inS11ser_mux_inst_7_X), .Z0_f (new_AGEMA_signal_4791), .Z1_t (new_AGEMA_signal_4792), .Z1_f (new_AGEMA_signal_4793) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS11ser_mux_inst_7_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS11ser_mux_inst_7_X), .B0_f (new_AGEMA_signal_4791), .B1_t (new_AGEMA_signal_4792), .B1_f (new_AGEMA_signal_4793), .Z0_t (KeyArray_MUX_inS11ser_mux_inst_7_Y), .Z0_f (new_AGEMA_signal_6253), .Z1_t (new_AGEMA_signal_6254), .Z1_f (new_AGEMA_signal_6255) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS11ser_mux_inst_7_XOR2_U1 ( .A0_t (KeyArray_MUX_inS11ser_mux_inst_7_Y), .A0_f (new_AGEMA_signal_6253), .A1_t (new_AGEMA_signal_6254), .A1_f (new_AGEMA_signal_6255), .B0_t (key_s0_t[87]), .B0_f (key_s0_f[87]), .B1_t (key_s1_t[87]), .B1_f (key_s1_f[87]), .Z0_t (KeyArray_inS11ser[7]), .Z0_f (new_AGEMA_signal_7027), .Z1_t (new_AGEMA_signal_7028), .Z1_f (new_AGEMA_signal_7029) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS12ser_mux_inst_0_XOR1_U1 ( .A0_t (key_s0_t[48]), .A0_f (key_s0_f[48]), .A1_t (key_s1_t[48]), .A1_f (key_s1_f[48]), .B0_t (keySBIn[0]), .B0_f (new_AGEMA_signal_4797), .B1_t (new_AGEMA_signal_4798), .B1_f (new_AGEMA_signal_4799), .Z0_t (KeyArray_MUX_inS12ser_mux_inst_0_X), .Z0_f (new_AGEMA_signal_4800), .Z1_t (new_AGEMA_signal_4801), .Z1_f (new_AGEMA_signal_4802) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS12ser_mux_inst_0_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS12ser_mux_inst_0_X), .B0_f (new_AGEMA_signal_4800), .B1_t (new_AGEMA_signal_4801), .B1_f (new_AGEMA_signal_4802), .Z0_t (KeyArray_MUX_inS12ser_mux_inst_0_Y), .Z0_f (new_AGEMA_signal_6256), .Z1_t (new_AGEMA_signal_6257), .Z1_f (new_AGEMA_signal_6258) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS12ser_mux_inst_0_XOR2_U1 ( .A0_t (KeyArray_MUX_inS12ser_mux_inst_0_Y), .A0_f (new_AGEMA_signal_6256), .A1_t (new_AGEMA_signal_6257), .A1_f (new_AGEMA_signal_6258), .B0_t (key_s0_t[48]), .B0_f (key_s0_f[48]), .B1_t (key_s1_t[48]), .B1_f (key_s1_f[48]), .Z0_t (KeyArray_inS12ser[0]), .Z0_f (new_AGEMA_signal_7030), .Z1_t (new_AGEMA_signal_7031), .Z1_f (new_AGEMA_signal_7032) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS12ser_mux_inst_1_XOR1_U1 ( .A0_t (key_s0_t[49]), .A0_f (key_s0_f[49]), .A1_t (key_s1_t[49]), .A1_f (key_s1_f[49]), .B0_t (keySBIn[1]), .B0_f (new_AGEMA_signal_4806), .B1_t (new_AGEMA_signal_4807), .B1_f (new_AGEMA_signal_4808), .Z0_t (KeyArray_MUX_inS12ser_mux_inst_1_X), .Z0_f (new_AGEMA_signal_4809), .Z1_t (new_AGEMA_signal_4810), .Z1_f (new_AGEMA_signal_4811) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS12ser_mux_inst_1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS12ser_mux_inst_1_X), .B0_f (new_AGEMA_signal_4809), .B1_t (new_AGEMA_signal_4810), .B1_f (new_AGEMA_signal_4811), .Z0_t (KeyArray_MUX_inS12ser_mux_inst_1_Y), .Z0_f (new_AGEMA_signal_6259), .Z1_t (new_AGEMA_signal_6260), .Z1_f (new_AGEMA_signal_6261) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS12ser_mux_inst_1_XOR2_U1 ( .A0_t (KeyArray_MUX_inS12ser_mux_inst_1_Y), .A0_f (new_AGEMA_signal_6259), .A1_t (new_AGEMA_signal_6260), .A1_f (new_AGEMA_signal_6261), .B0_t (key_s0_t[49]), .B0_f (key_s0_f[49]), .B1_t (key_s1_t[49]), .B1_f (key_s1_f[49]), .Z0_t (KeyArray_inS12ser[1]), .Z0_f (new_AGEMA_signal_7033), .Z1_t (new_AGEMA_signal_7034), .Z1_f (new_AGEMA_signal_7035) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS12ser_mux_inst_2_XOR1_U1 ( .A0_t (key_s0_t[50]), .A0_f (key_s0_f[50]), .A1_t (key_s1_t[50]), .A1_f (key_s1_f[50]), .B0_t (keySBIn[2]), .B0_f (new_AGEMA_signal_4815), .B1_t (new_AGEMA_signal_4816), .B1_f (new_AGEMA_signal_4817), .Z0_t (KeyArray_MUX_inS12ser_mux_inst_2_X), .Z0_f (new_AGEMA_signal_4818), .Z1_t (new_AGEMA_signal_4819), .Z1_f (new_AGEMA_signal_4820) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS12ser_mux_inst_2_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS12ser_mux_inst_2_X), .B0_f (new_AGEMA_signal_4818), .B1_t (new_AGEMA_signal_4819), .B1_f (new_AGEMA_signal_4820), .Z0_t (KeyArray_MUX_inS12ser_mux_inst_2_Y), .Z0_f (new_AGEMA_signal_6262), .Z1_t (new_AGEMA_signal_6263), .Z1_f (new_AGEMA_signal_6264) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS12ser_mux_inst_2_XOR2_U1 ( .A0_t (KeyArray_MUX_inS12ser_mux_inst_2_Y), .A0_f (new_AGEMA_signal_6262), .A1_t (new_AGEMA_signal_6263), .A1_f (new_AGEMA_signal_6264), .B0_t (key_s0_t[50]), .B0_f (key_s0_f[50]), .B1_t (key_s1_t[50]), .B1_f (key_s1_f[50]), .Z0_t (KeyArray_inS12ser[2]), .Z0_f (new_AGEMA_signal_7036), .Z1_t (new_AGEMA_signal_7037), .Z1_f (new_AGEMA_signal_7038) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS12ser_mux_inst_3_XOR1_U1 ( .A0_t (key_s0_t[51]), .A0_f (key_s0_f[51]), .A1_t (key_s1_t[51]), .A1_f (key_s1_f[51]), .B0_t (keySBIn[3]), .B0_f (new_AGEMA_signal_4824), .B1_t (new_AGEMA_signal_4825), .B1_f (new_AGEMA_signal_4826), .Z0_t (KeyArray_MUX_inS12ser_mux_inst_3_X), .Z0_f (new_AGEMA_signal_4827), .Z1_t (new_AGEMA_signal_4828), .Z1_f (new_AGEMA_signal_4829) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS12ser_mux_inst_3_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS12ser_mux_inst_3_X), .B0_f (new_AGEMA_signal_4827), .B1_t (new_AGEMA_signal_4828), .B1_f (new_AGEMA_signal_4829), .Z0_t (KeyArray_MUX_inS12ser_mux_inst_3_Y), .Z0_f (new_AGEMA_signal_6265), .Z1_t (new_AGEMA_signal_6266), .Z1_f (new_AGEMA_signal_6267) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS12ser_mux_inst_3_XOR2_U1 ( .A0_t (KeyArray_MUX_inS12ser_mux_inst_3_Y), .A0_f (new_AGEMA_signal_6265), .A1_t (new_AGEMA_signal_6266), .A1_f (new_AGEMA_signal_6267), .B0_t (key_s0_t[51]), .B0_f (key_s0_f[51]), .B1_t (key_s1_t[51]), .B1_f (key_s1_f[51]), .Z0_t (KeyArray_inS12ser[3]), .Z0_f (new_AGEMA_signal_7039), .Z1_t (new_AGEMA_signal_7040), .Z1_f (new_AGEMA_signal_7041) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS12ser_mux_inst_4_XOR1_U1 ( .A0_t (key_s0_t[52]), .A0_f (key_s0_f[52]), .A1_t (key_s1_t[52]), .A1_f (key_s1_f[52]), .B0_t (keySBIn[4]), .B0_f (new_AGEMA_signal_4833), .B1_t (new_AGEMA_signal_4834), .B1_f (new_AGEMA_signal_4835), .Z0_t (KeyArray_MUX_inS12ser_mux_inst_4_X), .Z0_f (new_AGEMA_signal_4836), .Z1_t (new_AGEMA_signal_4837), .Z1_f (new_AGEMA_signal_4838) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS12ser_mux_inst_4_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS12ser_mux_inst_4_X), .B0_f (new_AGEMA_signal_4836), .B1_t (new_AGEMA_signal_4837), .B1_f (new_AGEMA_signal_4838), .Z0_t (KeyArray_MUX_inS12ser_mux_inst_4_Y), .Z0_f (new_AGEMA_signal_6268), .Z1_t (new_AGEMA_signal_6269), .Z1_f (new_AGEMA_signal_6270) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS12ser_mux_inst_4_XOR2_U1 ( .A0_t (KeyArray_MUX_inS12ser_mux_inst_4_Y), .A0_f (new_AGEMA_signal_6268), .A1_t (new_AGEMA_signal_6269), .A1_f (new_AGEMA_signal_6270), .B0_t (key_s0_t[52]), .B0_f (key_s0_f[52]), .B1_t (key_s1_t[52]), .B1_f (key_s1_f[52]), .Z0_t (KeyArray_inS12ser[4]), .Z0_f (new_AGEMA_signal_7042), .Z1_t (new_AGEMA_signal_7043), .Z1_f (new_AGEMA_signal_7044) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS12ser_mux_inst_5_XOR1_U1 ( .A0_t (key_s0_t[53]), .A0_f (key_s0_f[53]), .A1_t (key_s1_t[53]), .A1_f (key_s1_f[53]), .B0_t (keySBIn[5]), .B0_f (new_AGEMA_signal_4842), .B1_t (new_AGEMA_signal_4843), .B1_f (new_AGEMA_signal_4844), .Z0_t (KeyArray_MUX_inS12ser_mux_inst_5_X), .Z0_f (new_AGEMA_signal_4845), .Z1_t (new_AGEMA_signal_4846), .Z1_f (new_AGEMA_signal_4847) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS12ser_mux_inst_5_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS12ser_mux_inst_5_X), .B0_f (new_AGEMA_signal_4845), .B1_t (new_AGEMA_signal_4846), .B1_f (new_AGEMA_signal_4847), .Z0_t (KeyArray_MUX_inS12ser_mux_inst_5_Y), .Z0_f (new_AGEMA_signal_6271), .Z1_t (new_AGEMA_signal_6272), .Z1_f (new_AGEMA_signal_6273) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS12ser_mux_inst_5_XOR2_U1 ( .A0_t (KeyArray_MUX_inS12ser_mux_inst_5_Y), .A0_f (new_AGEMA_signal_6271), .A1_t (new_AGEMA_signal_6272), .A1_f (new_AGEMA_signal_6273), .B0_t (key_s0_t[53]), .B0_f (key_s0_f[53]), .B1_t (key_s1_t[53]), .B1_f (key_s1_f[53]), .Z0_t (KeyArray_inS12ser[5]), .Z0_f (new_AGEMA_signal_7045), .Z1_t (new_AGEMA_signal_7046), .Z1_f (new_AGEMA_signal_7047) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS12ser_mux_inst_6_XOR1_U1 ( .A0_t (key_s0_t[54]), .A0_f (key_s0_f[54]), .A1_t (key_s1_t[54]), .A1_f (key_s1_f[54]), .B0_t (keySBIn[6]), .B0_f (new_AGEMA_signal_4851), .B1_t (new_AGEMA_signal_4852), .B1_f (new_AGEMA_signal_4853), .Z0_t (KeyArray_MUX_inS12ser_mux_inst_6_X), .Z0_f (new_AGEMA_signal_4854), .Z1_t (new_AGEMA_signal_4855), .Z1_f (new_AGEMA_signal_4856) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS12ser_mux_inst_6_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS12ser_mux_inst_6_X), .B0_f (new_AGEMA_signal_4854), .B1_t (new_AGEMA_signal_4855), .B1_f (new_AGEMA_signal_4856), .Z0_t (KeyArray_MUX_inS12ser_mux_inst_6_Y), .Z0_f (new_AGEMA_signal_6274), .Z1_t (new_AGEMA_signal_6275), .Z1_f (new_AGEMA_signal_6276) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS12ser_mux_inst_6_XOR2_U1 ( .A0_t (KeyArray_MUX_inS12ser_mux_inst_6_Y), .A0_f (new_AGEMA_signal_6274), .A1_t (new_AGEMA_signal_6275), .A1_f (new_AGEMA_signal_6276), .B0_t (key_s0_t[54]), .B0_f (key_s0_f[54]), .B1_t (key_s1_t[54]), .B1_f (key_s1_f[54]), .Z0_t (KeyArray_inS12ser[6]), .Z0_f (new_AGEMA_signal_7048), .Z1_t (new_AGEMA_signal_7049), .Z1_f (new_AGEMA_signal_7050) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS12ser_mux_inst_7_XOR1_U1 ( .A0_t (key_s0_t[55]), .A0_f (key_s0_f[55]), .A1_t (key_s1_t[55]), .A1_f (key_s1_f[55]), .B0_t (keySBIn[7]), .B0_f (new_AGEMA_signal_4860), .B1_t (new_AGEMA_signal_4861), .B1_f (new_AGEMA_signal_4862), .Z0_t (KeyArray_MUX_inS12ser_mux_inst_7_X), .Z0_f (new_AGEMA_signal_4863), .Z1_t (new_AGEMA_signal_4864), .Z1_f (new_AGEMA_signal_4865) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS12ser_mux_inst_7_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS12ser_mux_inst_7_X), .B0_f (new_AGEMA_signal_4863), .B1_t (new_AGEMA_signal_4864), .B1_f (new_AGEMA_signal_4865), .Z0_t (KeyArray_MUX_inS12ser_mux_inst_7_Y), .Z0_f (new_AGEMA_signal_6277), .Z1_t (new_AGEMA_signal_6278), .Z1_f (new_AGEMA_signal_6279) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS12ser_mux_inst_7_XOR2_U1 ( .A0_t (KeyArray_MUX_inS12ser_mux_inst_7_Y), .A0_f (new_AGEMA_signal_6277), .A1_t (new_AGEMA_signal_6278), .A1_f (new_AGEMA_signal_6279), .B0_t (key_s0_t[55]), .B0_f (key_s0_f[55]), .B1_t (key_s1_t[55]), .B1_f (key_s1_f[55]), .Z0_t (KeyArray_inS12ser[7]), .Z0_f (new_AGEMA_signal_7051), .Z1_t (new_AGEMA_signal_7052), .Z1_f (new_AGEMA_signal_7053) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS13ser_mux_inst_0_XOR1_U1 ( .A0_t (key_s0_t[16]), .A0_f (key_s0_f[16]), .A1_t (key_s1_t[16]), .A1_f (key_s1_f[16]), .B0_t (KeyArray_outS20ser[0]), .B0_f (new_AGEMA_signal_4869), .B1_t (new_AGEMA_signal_4870), .B1_f (new_AGEMA_signal_4871), .Z0_t (KeyArray_MUX_inS13ser_mux_inst_0_X), .Z0_f (new_AGEMA_signal_4872), .Z1_t (new_AGEMA_signal_4873), .Z1_f (new_AGEMA_signal_4874) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS13ser_mux_inst_0_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS13ser_mux_inst_0_X), .B0_f (new_AGEMA_signal_4872), .B1_t (new_AGEMA_signal_4873), .B1_f (new_AGEMA_signal_4874), .Z0_t (KeyArray_MUX_inS13ser_mux_inst_0_Y), .Z0_f (new_AGEMA_signal_6280), .Z1_t (new_AGEMA_signal_6281), .Z1_f (new_AGEMA_signal_6282) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS13ser_mux_inst_0_XOR2_U1 ( .A0_t (KeyArray_MUX_inS13ser_mux_inst_0_Y), .A0_f (new_AGEMA_signal_6280), .A1_t (new_AGEMA_signal_6281), .A1_f (new_AGEMA_signal_6282), .B0_t (key_s0_t[16]), .B0_f (key_s0_f[16]), .B1_t (key_s1_t[16]), .B1_f (key_s1_f[16]), .Z0_t (KeyArray_inS13ser[0]), .Z0_f (new_AGEMA_signal_7054), .Z1_t (new_AGEMA_signal_7055), .Z1_f (new_AGEMA_signal_7056) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS13ser_mux_inst_1_XOR1_U1 ( .A0_t (key_s0_t[17]), .A0_f (key_s0_f[17]), .A1_t (key_s1_t[17]), .A1_f (key_s1_f[17]), .B0_t (KeyArray_outS20ser[1]), .B0_f (new_AGEMA_signal_4878), .B1_t (new_AGEMA_signal_4879), .B1_f (new_AGEMA_signal_4880), .Z0_t (KeyArray_MUX_inS13ser_mux_inst_1_X), .Z0_f (new_AGEMA_signal_4881), .Z1_t (new_AGEMA_signal_4882), .Z1_f (new_AGEMA_signal_4883) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS13ser_mux_inst_1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS13ser_mux_inst_1_X), .B0_f (new_AGEMA_signal_4881), .B1_t (new_AGEMA_signal_4882), .B1_f (new_AGEMA_signal_4883), .Z0_t (KeyArray_MUX_inS13ser_mux_inst_1_Y), .Z0_f (new_AGEMA_signal_6283), .Z1_t (new_AGEMA_signal_6284), .Z1_f (new_AGEMA_signal_6285) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS13ser_mux_inst_1_XOR2_U1 ( .A0_t (KeyArray_MUX_inS13ser_mux_inst_1_Y), .A0_f (new_AGEMA_signal_6283), .A1_t (new_AGEMA_signal_6284), .A1_f (new_AGEMA_signal_6285), .B0_t (key_s0_t[17]), .B0_f (key_s0_f[17]), .B1_t (key_s1_t[17]), .B1_f (key_s1_f[17]), .Z0_t (KeyArray_inS13ser[1]), .Z0_f (new_AGEMA_signal_7057), .Z1_t (new_AGEMA_signal_7058), .Z1_f (new_AGEMA_signal_7059) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS13ser_mux_inst_2_XOR1_U1 ( .A0_t (key_s0_t[18]), .A0_f (key_s0_f[18]), .A1_t (key_s1_t[18]), .A1_f (key_s1_f[18]), .B0_t (KeyArray_outS20ser[2]), .B0_f (new_AGEMA_signal_4887), .B1_t (new_AGEMA_signal_4888), .B1_f (new_AGEMA_signal_4889), .Z0_t (KeyArray_MUX_inS13ser_mux_inst_2_X), .Z0_f (new_AGEMA_signal_4890), .Z1_t (new_AGEMA_signal_4891), .Z1_f (new_AGEMA_signal_4892) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS13ser_mux_inst_2_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS13ser_mux_inst_2_X), .B0_f (new_AGEMA_signal_4890), .B1_t (new_AGEMA_signal_4891), .B1_f (new_AGEMA_signal_4892), .Z0_t (KeyArray_MUX_inS13ser_mux_inst_2_Y), .Z0_f (new_AGEMA_signal_6286), .Z1_t (new_AGEMA_signal_6287), .Z1_f (new_AGEMA_signal_6288) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS13ser_mux_inst_2_XOR2_U1 ( .A0_t (KeyArray_MUX_inS13ser_mux_inst_2_Y), .A0_f (new_AGEMA_signal_6286), .A1_t (new_AGEMA_signal_6287), .A1_f (new_AGEMA_signal_6288), .B0_t (key_s0_t[18]), .B0_f (key_s0_f[18]), .B1_t (key_s1_t[18]), .B1_f (key_s1_f[18]), .Z0_t (KeyArray_inS13ser[2]), .Z0_f (new_AGEMA_signal_7060), .Z1_t (new_AGEMA_signal_7061), .Z1_f (new_AGEMA_signal_7062) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS13ser_mux_inst_3_XOR1_U1 ( .A0_t (key_s0_t[19]), .A0_f (key_s0_f[19]), .A1_t (key_s1_t[19]), .A1_f (key_s1_f[19]), .B0_t (KeyArray_outS20ser[3]), .B0_f (new_AGEMA_signal_4896), .B1_t (new_AGEMA_signal_4897), .B1_f (new_AGEMA_signal_4898), .Z0_t (KeyArray_MUX_inS13ser_mux_inst_3_X), .Z0_f (new_AGEMA_signal_4899), .Z1_t (new_AGEMA_signal_4900), .Z1_f (new_AGEMA_signal_4901) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS13ser_mux_inst_3_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS13ser_mux_inst_3_X), .B0_f (new_AGEMA_signal_4899), .B1_t (new_AGEMA_signal_4900), .B1_f (new_AGEMA_signal_4901), .Z0_t (KeyArray_MUX_inS13ser_mux_inst_3_Y), .Z0_f (new_AGEMA_signal_6289), .Z1_t (new_AGEMA_signal_6290), .Z1_f (new_AGEMA_signal_6291) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS13ser_mux_inst_3_XOR2_U1 ( .A0_t (KeyArray_MUX_inS13ser_mux_inst_3_Y), .A0_f (new_AGEMA_signal_6289), .A1_t (new_AGEMA_signal_6290), .A1_f (new_AGEMA_signal_6291), .B0_t (key_s0_t[19]), .B0_f (key_s0_f[19]), .B1_t (key_s1_t[19]), .B1_f (key_s1_f[19]), .Z0_t (KeyArray_inS13ser[3]), .Z0_f (new_AGEMA_signal_7063), .Z1_t (new_AGEMA_signal_7064), .Z1_f (new_AGEMA_signal_7065) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS13ser_mux_inst_4_XOR1_U1 ( .A0_t (key_s0_t[20]), .A0_f (key_s0_f[20]), .A1_t (key_s1_t[20]), .A1_f (key_s1_f[20]), .B0_t (KeyArray_outS20ser[4]), .B0_f (new_AGEMA_signal_4905), .B1_t (new_AGEMA_signal_4906), .B1_f (new_AGEMA_signal_4907), .Z0_t (KeyArray_MUX_inS13ser_mux_inst_4_X), .Z0_f (new_AGEMA_signal_4908), .Z1_t (new_AGEMA_signal_4909), .Z1_f (new_AGEMA_signal_4910) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS13ser_mux_inst_4_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS13ser_mux_inst_4_X), .B0_f (new_AGEMA_signal_4908), .B1_t (new_AGEMA_signal_4909), .B1_f (new_AGEMA_signal_4910), .Z0_t (KeyArray_MUX_inS13ser_mux_inst_4_Y), .Z0_f (new_AGEMA_signal_6292), .Z1_t (new_AGEMA_signal_6293), .Z1_f (new_AGEMA_signal_6294) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS13ser_mux_inst_4_XOR2_U1 ( .A0_t (KeyArray_MUX_inS13ser_mux_inst_4_Y), .A0_f (new_AGEMA_signal_6292), .A1_t (new_AGEMA_signal_6293), .A1_f (new_AGEMA_signal_6294), .B0_t (key_s0_t[20]), .B0_f (key_s0_f[20]), .B1_t (key_s1_t[20]), .B1_f (key_s1_f[20]), .Z0_t (KeyArray_inS13ser[4]), .Z0_f (new_AGEMA_signal_7066), .Z1_t (new_AGEMA_signal_7067), .Z1_f (new_AGEMA_signal_7068) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS13ser_mux_inst_5_XOR1_U1 ( .A0_t (key_s0_t[21]), .A0_f (key_s0_f[21]), .A1_t (key_s1_t[21]), .A1_f (key_s1_f[21]), .B0_t (KeyArray_outS20ser[5]), .B0_f (new_AGEMA_signal_4914), .B1_t (new_AGEMA_signal_4915), .B1_f (new_AGEMA_signal_4916), .Z0_t (KeyArray_MUX_inS13ser_mux_inst_5_X), .Z0_f (new_AGEMA_signal_4917), .Z1_t (new_AGEMA_signal_4918), .Z1_f (new_AGEMA_signal_4919) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS13ser_mux_inst_5_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS13ser_mux_inst_5_X), .B0_f (new_AGEMA_signal_4917), .B1_t (new_AGEMA_signal_4918), .B1_f (new_AGEMA_signal_4919), .Z0_t (KeyArray_MUX_inS13ser_mux_inst_5_Y), .Z0_f (new_AGEMA_signal_6295), .Z1_t (new_AGEMA_signal_6296), .Z1_f (new_AGEMA_signal_6297) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS13ser_mux_inst_5_XOR2_U1 ( .A0_t (KeyArray_MUX_inS13ser_mux_inst_5_Y), .A0_f (new_AGEMA_signal_6295), .A1_t (new_AGEMA_signal_6296), .A1_f (new_AGEMA_signal_6297), .B0_t (key_s0_t[21]), .B0_f (key_s0_f[21]), .B1_t (key_s1_t[21]), .B1_f (key_s1_f[21]), .Z0_t (KeyArray_inS13ser[5]), .Z0_f (new_AGEMA_signal_7069), .Z1_t (new_AGEMA_signal_7070), .Z1_f (new_AGEMA_signal_7071) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS13ser_mux_inst_6_XOR1_U1 ( .A0_t (key_s0_t[22]), .A0_f (key_s0_f[22]), .A1_t (key_s1_t[22]), .A1_f (key_s1_f[22]), .B0_t (KeyArray_outS20ser[6]), .B0_f (new_AGEMA_signal_4923), .B1_t (new_AGEMA_signal_4924), .B1_f (new_AGEMA_signal_4925), .Z0_t (KeyArray_MUX_inS13ser_mux_inst_6_X), .Z0_f (new_AGEMA_signal_4926), .Z1_t (new_AGEMA_signal_4927), .Z1_f (new_AGEMA_signal_4928) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS13ser_mux_inst_6_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS13ser_mux_inst_6_X), .B0_f (new_AGEMA_signal_4926), .B1_t (new_AGEMA_signal_4927), .B1_f (new_AGEMA_signal_4928), .Z0_t (KeyArray_MUX_inS13ser_mux_inst_6_Y), .Z0_f (new_AGEMA_signal_6298), .Z1_t (new_AGEMA_signal_6299), .Z1_f (new_AGEMA_signal_6300) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS13ser_mux_inst_6_XOR2_U1 ( .A0_t (KeyArray_MUX_inS13ser_mux_inst_6_Y), .A0_f (new_AGEMA_signal_6298), .A1_t (new_AGEMA_signal_6299), .A1_f (new_AGEMA_signal_6300), .B0_t (key_s0_t[22]), .B0_f (key_s0_f[22]), .B1_t (key_s1_t[22]), .B1_f (key_s1_f[22]), .Z0_t (KeyArray_inS13ser[6]), .Z0_f (new_AGEMA_signal_7072), .Z1_t (new_AGEMA_signal_7073), .Z1_f (new_AGEMA_signal_7074) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS13ser_mux_inst_7_XOR1_U1 ( .A0_t (key_s0_t[23]), .A0_f (key_s0_f[23]), .A1_t (key_s1_t[23]), .A1_f (key_s1_f[23]), .B0_t (KeyArray_outS20ser[7]), .B0_f (new_AGEMA_signal_4932), .B1_t (new_AGEMA_signal_4933), .B1_f (new_AGEMA_signal_4934), .Z0_t (KeyArray_MUX_inS13ser_mux_inst_7_X), .Z0_f (new_AGEMA_signal_4935), .Z1_t (new_AGEMA_signal_4936), .Z1_f (new_AGEMA_signal_4937) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS13ser_mux_inst_7_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS13ser_mux_inst_7_X), .B0_f (new_AGEMA_signal_4935), .B1_t (new_AGEMA_signal_4936), .B1_f (new_AGEMA_signal_4937), .Z0_t (KeyArray_MUX_inS13ser_mux_inst_7_Y), .Z0_f (new_AGEMA_signal_6301), .Z1_t (new_AGEMA_signal_6302), .Z1_f (new_AGEMA_signal_6303) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS13ser_mux_inst_7_XOR2_U1 ( .A0_t (KeyArray_MUX_inS13ser_mux_inst_7_Y), .A0_f (new_AGEMA_signal_6301), .A1_t (new_AGEMA_signal_6302), .A1_f (new_AGEMA_signal_6303), .B0_t (key_s0_t[23]), .B0_f (key_s0_f[23]), .B1_t (key_s1_t[23]), .B1_f (key_s1_f[23]), .Z0_t (KeyArray_inS13ser[7]), .Z0_f (new_AGEMA_signal_7075), .Z1_t (new_AGEMA_signal_7076), .Z1_f (new_AGEMA_signal_7077) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS20ser_mux_inst_0_XOR1_U1 ( .A0_t (key_s0_t[104]), .A0_f (key_s0_f[104]), .A1_t (key_s1_t[104]), .A1_f (key_s1_f[104]), .B0_t (KeyArray_outS21ser[0]), .B0_f (new_AGEMA_signal_4941), .B1_t (new_AGEMA_signal_4942), .B1_f (new_AGEMA_signal_4943), .Z0_t (KeyArray_MUX_inS20ser_mux_inst_0_X), .Z0_f (new_AGEMA_signal_4944), .Z1_t (new_AGEMA_signal_4945), .Z1_f (new_AGEMA_signal_4946) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS20ser_mux_inst_0_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS20ser_mux_inst_0_X), .B0_f (new_AGEMA_signal_4944), .B1_t (new_AGEMA_signal_4945), .B1_f (new_AGEMA_signal_4946), .Z0_t (KeyArray_MUX_inS20ser_mux_inst_0_Y), .Z0_f (new_AGEMA_signal_6304), .Z1_t (new_AGEMA_signal_6305), .Z1_f (new_AGEMA_signal_6306) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS20ser_mux_inst_0_XOR2_U1 ( .A0_t (KeyArray_MUX_inS20ser_mux_inst_0_Y), .A0_f (new_AGEMA_signal_6304), .A1_t (new_AGEMA_signal_6305), .A1_f (new_AGEMA_signal_6306), .B0_t (key_s0_t[104]), .B0_f (key_s0_f[104]), .B1_t (key_s1_t[104]), .B1_f (key_s1_f[104]), .Z0_t (KeyArray_inS20ser[0]), .Z0_f (new_AGEMA_signal_7078), .Z1_t (new_AGEMA_signal_7079), .Z1_f (new_AGEMA_signal_7080) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS20ser_mux_inst_1_XOR1_U1 ( .A0_t (key_s0_t[105]), .A0_f (key_s0_f[105]), .A1_t (key_s1_t[105]), .A1_f (key_s1_f[105]), .B0_t (KeyArray_outS21ser[1]), .B0_f (new_AGEMA_signal_4950), .B1_t (new_AGEMA_signal_4951), .B1_f (new_AGEMA_signal_4952), .Z0_t (KeyArray_MUX_inS20ser_mux_inst_1_X), .Z0_f (new_AGEMA_signal_4953), .Z1_t (new_AGEMA_signal_4954), .Z1_f (new_AGEMA_signal_4955) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS20ser_mux_inst_1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS20ser_mux_inst_1_X), .B0_f (new_AGEMA_signal_4953), .B1_t (new_AGEMA_signal_4954), .B1_f (new_AGEMA_signal_4955), .Z0_t (KeyArray_MUX_inS20ser_mux_inst_1_Y), .Z0_f (new_AGEMA_signal_6307), .Z1_t (new_AGEMA_signal_6308), .Z1_f (new_AGEMA_signal_6309) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS20ser_mux_inst_1_XOR2_U1 ( .A0_t (KeyArray_MUX_inS20ser_mux_inst_1_Y), .A0_f (new_AGEMA_signal_6307), .A1_t (new_AGEMA_signal_6308), .A1_f (new_AGEMA_signal_6309), .B0_t (key_s0_t[105]), .B0_f (key_s0_f[105]), .B1_t (key_s1_t[105]), .B1_f (key_s1_f[105]), .Z0_t (KeyArray_inS20ser[1]), .Z0_f (new_AGEMA_signal_7081), .Z1_t (new_AGEMA_signal_7082), .Z1_f (new_AGEMA_signal_7083) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS20ser_mux_inst_2_XOR1_U1 ( .A0_t (key_s0_t[106]), .A0_f (key_s0_f[106]), .A1_t (key_s1_t[106]), .A1_f (key_s1_f[106]), .B0_t (KeyArray_outS21ser[2]), .B0_f (new_AGEMA_signal_4959), .B1_t (new_AGEMA_signal_4960), .B1_f (new_AGEMA_signal_4961), .Z0_t (KeyArray_MUX_inS20ser_mux_inst_2_X), .Z0_f (new_AGEMA_signal_4962), .Z1_t (new_AGEMA_signal_4963), .Z1_f (new_AGEMA_signal_4964) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS20ser_mux_inst_2_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS20ser_mux_inst_2_X), .B0_f (new_AGEMA_signal_4962), .B1_t (new_AGEMA_signal_4963), .B1_f (new_AGEMA_signal_4964), .Z0_t (KeyArray_MUX_inS20ser_mux_inst_2_Y), .Z0_f (new_AGEMA_signal_6310), .Z1_t (new_AGEMA_signal_6311), .Z1_f (new_AGEMA_signal_6312) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS20ser_mux_inst_2_XOR2_U1 ( .A0_t (KeyArray_MUX_inS20ser_mux_inst_2_Y), .A0_f (new_AGEMA_signal_6310), .A1_t (new_AGEMA_signal_6311), .A1_f (new_AGEMA_signal_6312), .B0_t (key_s0_t[106]), .B0_f (key_s0_f[106]), .B1_t (key_s1_t[106]), .B1_f (key_s1_f[106]), .Z0_t (KeyArray_inS20ser[2]), .Z0_f (new_AGEMA_signal_7084), .Z1_t (new_AGEMA_signal_7085), .Z1_f (new_AGEMA_signal_7086) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS20ser_mux_inst_3_XOR1_U1 ( .A0_t (key_s0_t[107]), .A0_f (key_s0_f[107]), .A1_t (key_s1_t[107]), .A1_f (key_s1_f[107]), .B0_t (KeyArray_outS21ser[3]), .B0_f (new_AGEMA_signal_4968), .B1_t (new_AGEMA_signal_4969), .B1_f (new_AGEMA_signal_4970), .Z0_t (KeyArray_MUX_inS20ser_mux_inst_3_X), .Z0_f (new_AGEMA_signal_4971), .Z1_t (new_AGEMA_signal_4972), .Z1_f (new_AGEMA_signal_4973) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS20ser_mux_inst_3_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS20ser_mux_inst_3_X), .B0_f (new_AGEMA_signal_4971), .B1_t (new_AGEMA_signal_4972), .B1_f (new_AGEMA_signal_4973), .Z0_t (KeyArray_MUX_inS20ser_mux_inst_3_Y), .Z0_f (new_AGEMA_signal_6313), .Z1_t (new_AGEMA_signal_6314), .Z1_f (new_AGEMA_signal_6315) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS20ser_mux_inst_3_XOR2_U1 ( .A0_t (KeyArray_MUX_inS20ser_mux_inst_3_Y), .A0_f (new_AGEMA_signal_6313), .A1_t (new_AGEMA_signal_6314), .A1_f (new_AGEMA_signal_6315), .B0_t (key_s0_t[107]), .B0_f (key_s0_f[107]), .B1_t (key_s1_t[107]), .B1_f (key_s1_f[107]), .Z0_t (KeyArray_inS20ser[3]), .Z0_f (new_AGEMA_signal_7087), .Z1_t (new_AGEMA_signal_7088), .Z1_f (new_AGEMA_signal_7089) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS20ser_mux_inst_4_XOR1_U1 ( .A0_t (key_s0_t[108]), .A0_f (key_s0_f[108]), .A1_t (key_s1_t[108]), .A1_f (key_s1_f[108]), .B0_t (KeyArray_outS21ser[4]), .B0_f (new_AGEMA_signal_4977), .B1_t (new_AGEMA_signal_4978), .B1_f (new_AGEMA_signal_4979), .Z0_t (KeyArray_MUX_inS20ser_mux_inst_4_X), .Z0_f (new_AGEMA_signal_4980), .Z1_t (new_AGEMA_signal_4981), .Z1_f (new_AGEMA_signal_4982) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS20ser_mux_inst_4_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS20ser_mux_inst_4_X), .B0_f (new_AGEMA_signal_4980), .B1_t (new_AGEMA_signal_4981), .B1_f (new_AGEMA_signal_4982), .Z0_t (KeyArray_MUX_inS20ser_mux_inst_4_Y), .Z0_f (new_AGEMA_signal_6316), .Z1_t (new_AGEMA_signal_6317), .Z1_f (new_AGEMA_signal_6318) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS20ser_mux_inst_4_XOR2_U1 ( .A0_t (KeyArray_MUX_inS20ser_mux_inst_4_Y), .A0_f (new_AGEMA_signal_6316), .A1_t (new_AGEMA_signal_6317), .A1_f (new_AGEMA_signal_6318), .B0_t (key_s0_t[108]), .B0_f (key_s0_f[108]), .B1_t (key_s1_t[108]), .B1_f (key_s1_f[108]), .Z0_t (KeyArray_inS20ser[4]), .Z0_f (new_AGEMA_signal_7090), .Z1_t (new_AGEMA_signal_7091), .Z1_f (new_AGEMA_signal_7092) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS20ser_mux_inst_5_XOR1_U1 ( .A0_t (key_s0_t[109]), .A0_f (key_s0_f[109]), .A1_t (key_s1_t[109]), .A1_f (key_s1_f[109]), .B0_t (KeyArray_outS21ser[5]), .B0_f (new_AGEMA_signal_4986), .B1_t (new_AGEMA_signal_4987), .B1_f (new_AGEMA_signal_4988), .Z0_t (KeyArray_MUX_inS20ser_mux_inst_5_X), .Z0_f (new_AGEMA_signal_4989), .Z1_t (new_AGEMA_signal_4990), .Z1_f (new_AGEMA_signal_4991) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS20ser_mux_inst_5_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS20ser_mux_inst_5_X), .B0_f (new_AGEMA_signal_4989), .B1_t (new_AGEMA_signal_4990), .B1_f (new_AGEMA_signal_4991), .Z0_t (KeyArray_MUX_inS20ser_mux_inst_5_Y), .Z0_f (new_AGEMA_signal_6319), .Z1_t (new_AGEMA_signal_6320), .Z1_f (new_AGEMA_signal_6321) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS20ser_mux_inst_5_XOR2_U1 ( .A0_t (KeyArray_MUX_inS20ser_mux_inst_5_Y), .A0_f (new_AGEMA_signal_6319), .A1_t (new_AGEMA_signal_6320), .A1_f (new_AGEMA_signal_6321), .B0_t (key_s0_t[109]), .B0_f (key_s0_f[109]), .B1_t (key_s1_t[109]), .B1_f (key_s1_f[109]), .Z0_t (KeyArray_inS20ser[5]), .Z0_f (new_AGEMA_signal_7093), .Z1_t (new_AGEMA_signal_7094), .Z1_f (new_AGEMA_signal_7095) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS20ser_mux_inst_6_XOR1_U1 ( .A0_t (key_s0_t[110]), .A0_f (key_s0_f[110]), .A1_t (key_s1_t[110]), .A1_f (key_s1_f[110]), .B0_t (KeyArray_outS21ser[6]), .B0_f (new_AGEMA_signal_4995), .B1_t (new_AGEMA_signal_4996), .B1_f (new_AGEMA_signal_4997), .Z0_t (KeyArray_MUX_inS20ser_mux_inst_6_X), .Z0_f (new_AGEMA_signal_4998), .Z1_t (new_AGEMA_signal_4999), .Z1_f (new_AGEMA_signal_5000) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS20ser_mux_inst_6_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS20ser_mux_inst_6_X), .B0_f (new_AGEMA_signal_4998), .B1_t (new_AGEMA_signal_4999), .B1_f (new_AGEMA_signal_5000), .Z0_t (KeyArray_MUX_inS20ser_mux_inst_6_Y), .Z0_f (new_AGEMA_signal_6322), .Z1_t (new_AGEMA_signal_6323), .Z1_f (new_AGEMA_signal_6324) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS20ser_mux_inst_6_XOR2_U1 ( .A0_t (KeyArray_MUX_inS20ser_mux_inst_6_Y), .A0_f (new_AGEMA_signal_6322), .A1_t (new_AGEMA_signal_6323), .A1_f (new_AGEMA_signal_6324), .B0_t (key_s0_t[110]), .B0_f (key_s0_f[110]), .B1_t (key_s1_t[110]), .B1_f (key_s1_f[110]), .Z0_t (KeyArray_inS20ser[6]), .Z0_f (new_AGEMA_signal_7096), .Z1_t (new_AGEMA_signal_7097), .Z1_f (new_AGEMA_signal_7098) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS20ser_mux_inst_7_XOR1_U1 ( .A0_t (key_s0_t[111]), .A0_f (key_s0_f[111]), .A1_t (key_s1_t[111]), .A1_f (key_s1_f[111]), .B0_t (KeyArray_outS21ser[7]), .B0_f (new_AGEMA_signal_5004), .B1_t (new_AGEMA_signal_5005), .B1_f (new_AGEMA_signal_5006), .Z0_t (KeyArray_MUX_inS20ser_mux_inst_7_X), .Z0_f (new_AGEMA_signal_5007), .Z1_t (new_AGEMA_signal_5008), .Z1_f (new_AGEMA_signal_5009) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS20ser_mux_inst_7_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS20ser_mux_inst_7_X), .B0_f (new_AGEMA_signal_5007), .B1_t (new_AGEMA_signal_5008), .B1_f (new_AGEMA_signal_5009), .Z0_t (KeyArray_MUX_inS20ser_mux_inst_7_Y), .Z0_f (new_AGEMA_signal_6325), .Z1_t (new_AGEMA_signal_6326), .Z1_f (new_AGEMA_signal_6327) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS20ser_mux_inst_7_XOR2_U1 ( .A0_t (KeyArray_MUX_inS20ser_mux_inst_7_Y), .A0_f (new_AGEMA_signal_6325), .A1_t (new_AGEMA_signal_6326), .A1_f (new_AGEMA_signal_6327), .B0_t (key_s0_t[111]), .B0_f (key_s0_f[111]), .B1_t (key_s1_t[111]), .B1_f (key_s1_f[111]), .Z0_t (KeyArray_inS20ser[7]), .Z0_f (new_AGEMA_signal_7099), .Z1_t (new_AGEMA_signal_7100), .Z1_f (new_AGEMA_signal_7101) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS21ser_mux_inst_0_XOR1_U1 ( .A0_t (key_s0_t[72]), .A0_f (key_s0_f[72]), .A1_t (key_s1_t[72]), .A1_f (key_s1_f[72]), .B0_t (KeyArray_outS22ser[0]), .B0_f (new_AGEMA_signal_5013), .B1_t (new_AGEMA_signal_5014), .B1_f (new_AGEMA_signal_5015), .Z0_t (KeyArray_MUX_inS21ser_mux_inst_0_X), .Z0_f (new_AGEMA_signal_5016), .Z1_t (new_AGEMA_signal_5017), .Z1_f (new_AGEMA_signal_5018) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS21ser_mux_inst_0_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS21ser_mux_inst_0_X), .B0_f (new_AGEMA_signal_5016), .B1_t (new_AGEMA_signal_5017), .B1_f (new_AGEMA_signal_5018), .Z0_t (KeyArray_MUX_inS21ser_mux_inst_0_Y), .Z0_f (new_AGEMA_signal_6328), .Z1_t (new_AGEMA_signal_6329), .Z1_f (new_AGEMA_signal_6330) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS21ser_mux_inst_0_XOR2_U1 ( .A0_t (KeyArray_MUX_inS21ser_mux_inst_0_Y), .A0_f (new_AGEMA_signal_6328), .A1_t (new_AGEMA_signal_6329), .A1_f (new_AGEMA_signal_6330), .B0_t (key_s0_t[72]), .B0_f (key_s0_f[72]), .B1_t (key_s1_t[72]), .B1_f (key_s1_f[72]), .Z0_t (KeyArray_inS21ser[0]), .Z0_f (new_AGEMA_signal_7102), .Z1_t (new_AGEMA_signal_7103), .Z1_f (new_AGEMA_signal_7104) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS21ser_mux_inst_1_XOR1_U1 ( .A0_t (key_s0_t[73]), .A0_f (key_s0_f[73]), .A1_t (key_s1_t[73]), .A1_f (key_s1_f[73]), .B0_t (KeyArray_outS22ser[1]), .B0_f (new_AGEMA_signal_5022), .B1_t (new_AGEMA_signal_5023), .B1_f (new_AGEMA_signal_5024), .Z0_t (KeyArray_MUX_inS21ser_mux_inst_1_X), .Z0_f (new_AGEMA_signal_5025), .Z1_t (new_AGEMA_signal_5026), .Z1_f (new_AGEMA_signal_5027) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS21ser_mux_inst_1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS21ser_mux_inst_1_X), .B0_f (new_AGEMA_signal_5025), .B1_t (new_AGEMA_signal_5026), .B1_f (new_AGEMA_signal_5027), .Z0_t (KeyArray_MUX_inS21ser_mux_inst_1_Y), .Z0_f (new_AGEMA_signal_6331), .Z1_t (new_AGEMA_signal_6332), .Z1_f (new_AGEMA_signal_6333) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS21ser_mux_inst_1_XOR2_U1 ( .A0_t (KeyArray_MUX_inS21ser_mux_inst_1_Y), .A0_f (new_AGEMA_signal_6331), .A1_t (new_AGEMA_signal_6332), .A1_f (new_AGEMA_signal_6333), .B0_t (key_s0_t[73]), .B0_f (key_s0_f[73]), .B1_t (key_s1_t[73]), .B1_f (key_s1_f[73]), .Z0_t (KeyArray_inS21ser[1]), .Z0_f (new_AGEMA_signal_7105), .Z1_t (new_AGEMA_signal_7106), .Z1_f (new_AGEMA_signal_7107) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS21ser_mux_inst_2_XOR1_U1 ( .A0_t (key_s0_t[74]), .A0_f (key_s0_f[74]), .A1_t (key_s1_t[74]), .A1_f (key_s1_f[74]), .B0_t (KeyArray_outS22ser[2]), .B0_f (new_AGEMA_signal_5031), .B1_t (new_AGEMA_signal_5032), .B1_f (new_AGEMA_signal_5033), .Z0_t (KeyArray_MUX_inS21ser_mux_inst_2_X), .Z0_f (new_AGEMA_signal_5034), .Z1_t (new_AGEMA_signal_5035), .Z1_f (new_AGEMA_signal_5036) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS21ser_mux_inst_2_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS21ser_mux_inst_2_X), .B0_f (new_AGEMA_signal_5034), .B1_t (new_AGEMA_signal_5035), .B1_f (new_AGEMA_signal_5036), .Z0_t (KeyArray_MUX_inS21ser_mux_inst_2_Y), .Z0_f (new_AGEMA_signal_6334), .Z1_t (new_AGEMA_signal_6335), .Z1_f (new_AGEMA_signal_6336) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS21ser_mux_inst_2_XOR2_U1 ( .A0_t (KeyArray_MUX_inS21ser_mux_inst_2_Y), .A0_f (new_AGEMA_signal_6334), .A1_t (new_AGEMA_signal_6335), .A1_f (new_AGEMA_signal_6336), .B0_t (key_s0_t[74]), .B0_f (key_s0_f[74]), .B1_t (key_s1_t[74]), .B1_f (key_s1_f[74]), .Z0_t (KeyArray_inS21ser[2]), .Z0_f (new_AGEMA_signal_7108), .Z1_t (new_AGEMA_signal_7109), .Z1_f (new_AGEMA_signal_7110) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS21ser_mux_inst_3_XOR1_U1 ( .A0_t (key_s0_t[75]), .A0_f (key_s0_f[75]), .A1_t (key_s1_t[75]), .A1_f (key_s1_f[75]), .B0_t (KeyArray_outS22ser[3]), .B0_f (new_AGEMA_signal_5040), .B1_t (new_AGEMA_signal_5041), .B1_f (new_AGEMA_signal_5042), .Z0_t (KeyArray_MUX_inS21ser_mux_inst_3_X), .Z0_f (new_AGEMA_signal_5043), .Z1_t (new_AGEMA_signal_5044), .Z1_f (new_AGEMA_signal_5045) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS21ser_mux_inst_3_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS21ser_mux_inst_3_X), .B0_f (new_AGEMA_signal_5043), .B1_t (new_AGEMA_signal_5044), .B1_f (new_AGEMA_signal_5045), .Z0_t (KeyArray_MUX_inS21ser_mux_inst_3_Y), .Z0_f (new_AGEMA_signal_6337), .Z1_t (new_AGEMA_signal_6338), .Z1_f (new_AGEMA_signal_6339) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS21ser_mux_inst_3_XOR2_U1 ( .A0_t (KeyArray_MUX_inS21ser_mux_inst_3_Y), .A0_f (new_AGEMA_signal_6337), .A1_t (new_AGEMA_signal_6338), .A1_f (new_AGEMA_signal_6339), .B0_t (key_s0_t[75]), .B0_f (key_s0_f[75]), .B1_t (key_s1_t[75]), .B1_f (key_s1_f[75]), .Z0_t (KeyArray_inS21ser[3]), .Z0_f (new_AGEMA_signal_7111), .Z1_t (new_AGEMA_signal_7112), .Z1_f (new_AGEMA_signal_7113) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS21ser_mux_inst_4_XOR1_U1 ( .A0_t (key_s0_t[76]), .A0_f (key_s0_f[76]), .A1_t (key_s1_t[76]), .A1_f (key_s1_f[76]), .B0_t (KeyArray_outS22ser[4]), .B0_f (new_AGEMA_signal_5049), .B1_t (new_AGEMA_signal_5050), .B1_f (new_AGEMA_signal_5051), .Z0_t (KeyArray_MUX_inS21ser_mux_inst_4_X), .Z0_f (new_AGEMA_signal_5052), .Z1_t (new_AGEMA_signal_5053), .Z1_f (new_AGEMA_signal_5054) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS21ser_mux_inst_4_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS21ser_mux_inst_4_X), .B0_f (new_AGEMA_signal_5052), .B1_t (new_AGEMA_signal_5053), .B1_f (new_AGEMA_signal_5054), .Z0_t (KeyArray_MUX_inS21ser_mux_inst_4_Y), .Z0_f (new_AGEMA_signal_6340), .Z1_t (new_AGEMA_signal_6341), .Z1_f (new_AGEMA_signal_6342) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS21ser_mux_inst_4_XOR2_U1 ( .A0_t (KeyArray_MUX_inS21ser_mux_inst_4_Y), .A0_f (new_AGEMA_signal_6340), .A1_t (new_AGEMA_signal_6341), .A1_f (new_AGEMA_signal_6342), .B0_t (key_s0_t[76]), .B0_f (key_s0_f[76]), .B1_t (key_s1_t[76]), .B1_f (key_s1_f[76]), .Z0_t (KeyArray_inS21ser[4]), .Z0_f (new_AGEMA_signal_7114), .Z1_t (new_AGEMA_signal_7115), .Z1_f (new_AGEMA_signal_7116) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS21ser_mux_inst_5_XOR1_U1 ( .A0_t (key_s0_t[77]), .A0_f (key_s0_f[77]), .A1_t (key_s1_t[77]), .A1_f (key_s1_f[77]), .B0_t (KeyArray_outS22ser[5]), .B0_f (new_AGEMA_signal_5058), .B1_t (new_AGEMA_signal_5059), .B1_f (new_AGEMA_signal_5060), .Z0_t (KeyArray_MUX_inS21ser_mux_inst_5_X), .Z0_f (new_AGEMA_signal_5061), .Z1_t (new_AGEMA_signal_5062), .Z1_f (new_AGEMA_signal_5063) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS21ser_mux_inst_5_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS21ser_mux_inst_5_X), .B0_f (new_AGEMA_signal_5061), .B1_t (new_AGEMA_signal_5062), .B1_f (new_AGEMA_signal_5063), .Z0_t (KeyArray_MUX_inS21ser_mux_inst_5_Y), .Z0_f (new_AGEMA_signal_6343), .Z1_t (new_AGEMA_signal_6344), .Z1_f (new_AGEMA_signal_6345) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS21ser_mux_inst_5_XOR2_U1 ( .A0_t (KeyArray_MUX_inS21ser_mux_inst_5_Y), .A0_f (new_AGEMA_signal_6343), .A1_t (new_AGEMA_signal_6344), .A1_f (new_AGEMA_signal_6345), .B0_t (key_s0_t[77]), .B0_f (key_s0_f[77]), .B1_t (key_s1_t[77]), .B1_f (key_s1_f[77]), .Z0_t (KeyArray_inS21ser[5]), .Z0_f (new_AGEMA_signal_7117), .Z1_t (new_AGEMA_signal_7118), .Z1_f (new_AGEMA_signal_7119) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS21ser_mux_inst_6_XOR1_U1 ( .A0_t (key_s0_t[78]), .A0_f (key_s0_f[78]), .A1_t (key_s1_t[78]), .A1_f (key_s1_f[78]), .B0_t (KeyArray_outS22ser[6]), .B0_f (new_AGEMA_signal_5067), .B1_t (new_AGEMA_signal_5068), .B1_f (new_AGEMA_signal_5069), .Z0_t (KeyArray_MUX_inS21ser_mux_inst_6_X), .Z0_f (new_AGEMA_signal_5070), .Z1_t (new_AGEMA_signal_5071), .Z1_f (new_AGEMA_signal_5072) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS21ser_mux_inst_6_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS21ser_mux_inst_6_X), .B0_f (new_AGEMA_signal_5070), .B1_t (new_AGEMA_signal_5071), .B1_f (new_AGEMA_signal_5072), .Z0_t (KeyArray_MUX_inS21ser_mux_inst_6_Y), .Z0_f (new_AGEMA_signal_6346), .Z1_t (new_AGEMA_signal_6347), .Z1_f (new_AGEMA_signal_6348) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS21ser_mux_inst_6_XOR2_U1 ( .A0_t (KeyArray_MUX_inS21ser_mux_inst_6_Y), .A0_f (new_AGEMA_signal_6346), .A1_t (new_AGEMA_signal_6347), .A1_f (new_AGEMA_signal_6348), .B0_t (key_s0_t[78]), .B0_f (key_s0_f[78]), .B1_t (key_s1_t[78]), .B1_f (key_s1_f[78]), .Z0_t (KeyArray_inS21ser[6]), .Z0_f (new_AGEMA_signal_7120), .Z1_t (new_AGEMA_signal_7121), .Z1_f (new_AGEMA_signal_7122) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS21ser_mux_inst_7_XOR1_U1 ( .A0_t (key_s0_t[79]), .A0_f (key_s0_f[79]), .A1_t (key_s1_t[79]), .A1_f (key_s1_f[79]), .B0_t (KeyArray_outS22ser[7]), .B0_f (new_AGEMA_signal_5076), .B1_t (new_AGEMA_signal_5077), .B1_f (new_AGEMA_signal_5078), .Z0_t (KeyArray_MUX_inS21ser_mux_inst_7_X), .Z0_f (new_AGEMA_signal_5079), .Z1_t (new_AGEMA_signal_5080), .Z1_f (new_AGEMA_signal_5081) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS21ser_mux_inst_7_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS21ser_mux_inst_7_X), .B0_f (new_AGEMA_signal_5079), .B1_t (new_AGEMA_signal_5080), .B1_f (new_AGEMA_signal_5081), .Z0_t (KeyArray_MUX_inS21ser_mux_inst_7_Y), .Z0_f (new_AGEMA_signal_6349), .Z1_t (new_AGEMA_signal_6350), .Z1_f (new_AGEMA_signal_6351) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS21ser_mux_inst_7_XOR2_U1 ( .A0_t (KeyArray_MUX_inS21ser_mux_inst_7_Y), .A0_f (new_AGEMA_signal_6349), .A1_t (new_AGEMA_signal_6350), .A1_f (new_AGEMA_signal_6351), .B0_t (key_s0_t[79]), .B0_f (key_s0_f[79]), .B1_t (key_s1_t[79]), .B1_f (key_s1_f[79]), .Z0_t (KeyArray_inS21ser[7]), .Z0_f (new_AGEMA_signal_7123), .Z1_t (new_AGEMA_signal_7124), .Z1_f (new_AGEMA_signal_7125) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS22ser_mux_inst_0_XOR1_U1 ( .A0_t (key_s0_t[40]), .A0_f (key_s0_f[40]), .A1_t (key_s1_t[40]), .A1_f (key_s1_f[40]), .B0_t (KeyArray_outS23ser[0]), .B0_f (new_AGEMA_signal_5085), .B1_t (new_AGEMA_signal_5086), .B1_f (new_AGEMA_signal_5087), .Z0_t (KeyArray_MUX_inS22ser_mux_inst_0_X), .Z0_f (new_AGEMA_signal_5088), .Z1_t (new_AGEMA_signal_5089), .Z1_f (new_AGEMA_signal_5090) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS22ser_mux_inst_0_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS22ser_mux_inst_0_X), .B0_f (new_AGEMA_signal_5088), .B1_t (new_AGEMA_signal_5089), .B1_f (new_AGEMA_signal_5090), .Z0_t (KeyArray_MUX_inS22ser_mux_inst_0_Y), .Z0_f (new_AGEMA_signal_6352), .Z1_t (new_AGEMA_signal_6353), .Z1_f (new_AGEMA_signal_6354) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS22ser_mux_inst_0_XOR2_U1 ( .A0_t (KeyArray_MUX_inS22ser_mux_inst_0_Y), .A0_f (new_AGEMA_signal_6352), .A1_t (new_AGEMA_signal_6353), .A1_f (new_AGEMA_signal_6354), .B0_t (key_s0_t[40]), .B0_f (key_s0_f[40]), .B1_t (key_s1_t[40]), .B1_f (key_s1_f[40]), .Z0_t (KeyArray_inS22ser[0]), .Z0_f (new_AGEMA_signal_7126), .Z1_t (new_AGEMA_signal_7127), .Z1_f (new_AGEMA_signal_7128) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS22ser_mux_inst_1_XOR1_U1 ( .A0_t (key_s0_t[41]), .A0_f (key_s0_f[41]), .A1_t (key_s1_t[41]), .A1_f (key_s1_f[41]), .B0_t (KeyArray_outS23ser[1]), .B0_f (new_AGEMA_signal_5094), .B1_t (new_AGEMA_signal_5095), .B1_f (new_AGEMA_signal_5096), .Z0_t (KeyArray_MUX_inS22ser_mux_inst_1_X), .Z0_f (new_AGEMA_signal_5097), .Z1_t (new_AGEMA_signal_5098), .Z1_f (new_AGEMA_signal_5099) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS22ser_mux_inst_1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS22ser_mux_inst_1_X), .B0_f (new_AGEMA_signal_5097), .B1_t (new_AGEMA_signal_5098), .B1_f (new_AGEMA_signal_5099), .Z0_t (KeyArray_MUX_inS22ser_mux_inst_1_Y), .Z0_f (new_AGEMA_signal_6355), .Z1_t (new_AGEMA_signal_6356), .Z1_f (new_AGEMA_signal_6357) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS22ser_mux_inst_1_XOR2_U1 ( .A0_t (KeyArray_MUX_inS22ser_mux_inst_1_Y), .A0_f (new_AGEMA_signal_6355), .A1_t (new_AGEMA_signal_6356), .A1_f (new_AGEMA_signal_6357), .B0_t (key_s0_t[41]), .B0_f (key_s0_f[41]), .B1_t (key_s1_t[41]), .B1_f (key_s1_f[41]), .Z0_t (KeyArray_inS22ser[1]), .Z0_f (new_AGEMA_signal_7129), .Z1_t (new_AGEMA_signal_7130), .Z1_f (new_AGEMA_signal_7131) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS22ser_mux_inst_2_XOR1_U1 ( .A0_t (key_s0_t[42]), .A0_f (key_s0_f[42]), .A1_t (key_s1_t[42]), .A1_f (key_s1_f[42]), .B0_t (KeyArray_outS23ser[2]), .B0_f (new_AGEMA_signal_5103), .B1_t (new_AGEMA_signal_5104), .B1_f (new_AGEMA_signal_5105), .Z0_t (KeyArray_MUX_inS22ser_mux_inst_2_X), .Z0_f (new_AGEMA_signal_5106), .Z1_t (new_AGEMA_signal_5107), .Z1_f (new_AGEMA_signal_5108) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS22ser_mux_inst_2_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS22ser_mux_inst_2_X), .B0_f (new_AGEMA_signal_5106), .B1_t (new_AGEMA_signal_5107), .B1_f (new_AGEMA_signal_5108), .Z0_t (KeyArray_MUX_inS22ser_mux_inst_2_Y), .Z0_f (new_AGEMA_signal_6358), .Z1_t (new_AGEMA_signal_6359), .Z1_f (new_AGEMA_signal_6360) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS22ser_mux_inst_2_XOR2_U1 ( .A0_t (KeyArray_MUX_inS22ser_mux_inst_2_Y), .A0_f (new_AGEMA_signal_6358), .A1_t (new_AGEMA_signal_6359), .A1_f (new_AGEMA_signal_6360), .B0_t (key_s0_t[42]), .B0_f (key_s0_f[42]), .B1_t (key_s1_t[42]), .B1_f (key_s1_f[42]), .Z0_t (KeyArray_inS22ser[2]), .Z0_f (new_AGEMA_signal_7132), .Z1_t (new_AGEMA_signal_7133), .Z1_f (new_AGEMA_signal_7134) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS22ser_mux_inst_3_XOR1_U1 ( .A0_t (key_s0_t[43]), .A0_f (key_s0_f[43]), .A1_t (key_s1_t[43]), .A1_f (key_s1_f[43]), .B0_t (KeyArray_outS23ser[3]), .B0_f (new_AGEMA_signal_5112), .B1_t (new_AGEMA_signal_5113), .B1_f (new_AGEMA_signal_5114), .Z0_t (KeyArray_MUX_inS22ser_mux_inst_3_X), .Z0_f (new_AGEMA_signal_5115), .Z1_t (new_AGEMA_signal_5116), .Z1_f (new_AGEMA_signal_5117) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS22ser_mux_inst_3_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS22ser_mux_inst_3_X), .B0_f (new_AGEMA_signal_5115), .B1_t (new_AGEMA_signal_5116), .B1_f (new_AGEMA_signal_5117), .Z0_t (KeyArray_MUX_inS22ser_mux_inst_3_Y), .Z0_f (new_AGEMA_signal_6361), .Z1_t (new_AGEMA_signal_6362), .Z1_f (new_AGEMA_signal_6363) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS22ser_mux_inst_3_XOR2_U1 ( .A0_t (KeyArray_MUX_inS22ser_mux_inst_3_Y), .A0_f (new_AGEMA_signal_6361), .A1_t (new_AGEMA_signal_6362), .A1_f (new_AGEMA_signal_6363), .B0_t (key_s0_t[43]), .B0_f (key_s0_f[43]), .B1_t (key_s1_t[43]), .B1_f (key_s1_f[43]), .Z0_t (KeyArray_inS22ser[3]), .Z0_f (new_AGEMA_signal_7135), .Z1_t (new_AGEMA_signal_7136), .Z1_f (new_AGEMA_signal_7137) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS22ser_mux_inst_4_XOR1_U1 ( .A0_t (key_s0_t[44]), .A0_f (key_s0_f[44]), .A1_t (key_s1_t[44]), .A1_f (key_s1_f[44]), .B0_t (KeyArray_outS23ser[4]), .B0_f (new_AGEMA_signal_5121), .B1_t (new_AGEMA_signal_5122), .B1_f (new_AGEMA_signal_5123), .Z0_t (KeyArray_MUX_inS22ser_mux_inst_4_X), .Z0_f (new_AGEMA_signal_5124), .Z1_t (new_AGEMA_signal_5125), .Z1_f (new_AGEMA_signal_5126) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS22ser_mux_inst_4_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS22ser_mux_inst_4_X), .B0_f (new_AGEMA_signal_5124), .B1_t (new_AGEMA_signal_5125), .B1_f (new_AGEMA_signal_5126), .Z0_t (KeyArray_MUX_inS22ser_mux_inst_4_Y), .Z0_f (new_AGEMA_signal_6364), .Z1_t (new_AGEMA_signal_6365), .Z1_f (new_AGEMA_signal_6366) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS22ser_mux_inst_4_XOR2_U1 ( .A0_t (KeyArray_MUX_inS22ser_mux_inst_4_Y), .A0_f (new_AGEMA_signal_6364), .A1_t (new_AGEMA_signal_6365), .A1_f (new_AGEMA_signal_6366), .B0_t (key_s0_t[44]), .B0_f (key_s0_f[44]), .B1_t (key_s1_t[44]), .B1_f (key_s1_f[44]), .Z0_t (KeyArray_inS22ser[4]), .Z0_f (new_AGEMA_signal_7138), .Z1_t (new_AGEMA_signal_7139), .Z1_f (new_AGEMA_signal_7140) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS22ser_mux_inst_5_XOR1_U1 ( .A0_t (key_s0_t[45]), .A0_f (key_s0_f[45]), .A1_t (key_s1_t[45]), .A1_f (key_s1_f[45]), .B0_t (KeyArray_outS23ser[5]), .B0_f (new_AGEMA_signal_5130), .B1_t (new_AGEMA_signal_5131), .B1_f (new_AGEMA_signal_5132), .Z0_t (KeyArray_MUX_inS22ser_mux_inst_5_X), .Z0_f (new_AGEMA_signal_5133), .Z1_t (new_AGEMA_signal_5134), .Z1_f (new_AGEMA_signal_5135) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS22ser_mux_inst_5_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS22ser_mux_inst_5_X), .B0_f (new_AGEMA_signal_5133), .B1_t (new_AGEMA_signal_5134), .B1_f (new_AGEMA_signal_5135), .Z0_t (KeyArray_MUX_inS22ser_mux_inst_5_Y), .Z0_f (new_AGEMA_signal_6367), .Z1_t (new_AGEMA_signal_6368), .Z1_f (new_AGEMA_signal_6369) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS22ser_mux_inst_5_XOR2_U1 ( .A0_t (KeyArray_MUX_inS22ser_mux_inst_5_Y), .A0_f (new_AGEMA_signal_6367), .A1_t (new_AGEMA_signal_6368), .A1_f (new_AGEMA_signal_6369), .B0_t (key_s0_t[45]), .B0_f (key_s0_f[45]), .B1_t (key_s1_t[45]), .B1_f (key_s1_f[45]), .Z0_t (KeyArray_inS22ser[5]), .Z0_f (new_AGEMA_signal_7141), .Z1_t (new_AGEMA_signal_7142), .Z1_f (new_AGEMA_signal_7143) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS22ser_mux_inst_6_XOR1_U1 ( .A0_t (key_s0_t[46]), .A0_f (key_s0_f[46]), .A1_t (key_s1_t[46]), .A1_f (key_s1_f[46]), .B0_t (KeyArray_outS23ser[6]), .B0_f (new_AGEMA_signal_5139), .B1_t (new_AGEMA_signal_5140), .B1_f (new_AGEMA_signal_5141), .Z0_t (KeyArray_MUX_inS22ser_mux_inst_6_X), .Z0_f (new_AGEMA_signal_5142), .Z1_t (new_AGEMA_signal_5143), .Z1_f (new_AGEMA_signal_5144) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS22ser_mux_inst_6_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS22ser_mux_inst_6_X), .B0_f (new_AGEMA_signal_5142), .B1_t (new_AGEMA_signal_5143), .B1_f (new_AGEMA_signal_5144), .Z0_t (KeyArray_MUX_inS22ser_mux_inst_6_Y), .Z0_f (new_AGEMA_signal_6370), .Z1_t (new_AGEMA_signal_6371), .Z1_f (new_AGEMA_signal_6372) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS22ser_mux_inst_6_XOR2_U1 ( .A0_t (KeyArray_MUX_inS22ser_mux_inst_6_Y), .A0_f (new_AGEMA_signal_6370), .A1_t (new_AGEMA_signal_6371), .A1_f (new_AGEMA_signal_6372), .B0_t (key_s0_t[46]), .B0_f (key_s0_f[46]), .B1_t (key_s1_t[46]), .B1_f (key_s1_f[46]), .Z0_t (KeyArray_inS22ser[6]), .Z0_f (new_AGEMA_signal_7144), .Z1_t (new_AGEMA_signal_7145), .Z1_f (new_AGEMA_signal_7146) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS22ser_mux_inst_7_XOR1_U1 ( .A0_t (key_s0_t[47]), .A0_f (key_s0_f[47]), .A1_t (key_s1_t[47]), .A1_f (key_s1_f[47]), .B0_t (KeyArray_outS23ser[7]), .B0_f (new_AGEMA_signal_5148), .B1_t (new_AGEMA_signal_5149), .B1_f (new_AGEMA_signal_5150), .Z0_t (KeyArray_MUX_inS22ser_mux_inst_7_X), .Z0_f (new_AGEMA_signal_5151), .Z1_t (new_AGEMA_signal_5152), .Z1_f (new_AGEMA_signal_5153) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS22ser_mux_inst_7_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS22ser_mux_inst_7_X), .B0_f (new_AGEMA_signal_5151), .B1_t (new_AGEMA_signal_5152), .B1_f (new_AGEMA_signal_5153), .Z0_t (KeyArray_MUX_inS22ser_mux_inst_7_Y), .Z0_f (new_AGEMA_signal_6373), .Z1_t (new_AGEMA_signal_6374), .Z1_f (new_AGEMA_signal_6375) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS22ser_mux_inst_7_XOR2_U1 ( .A0_t (KeyArray_MUX_inS22ser_mux_inst_7_Y), .A0_f (new_AGEMA_signal_6373), .A1_t (new_AGEMA_signal_6374), .A1_f (new_AGEMA_signal_6375), .B0_t (key_s0_t[47]), .B0_f (key_s0_f[47]), .B1_t (key_s1_t[47]), .B1_f (key_s1_f[47]), .Z0_t (KeyArray_inS22ser[7]), .Z0_f (new_AGEMA_signal_7147), .Z1_t (new_AGEMA_signal_7148), .Z1_f (new_AGEMA_signal_7149) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS23ser_mux_inst_0_XOR1_U1 ( .A0_t (key_s0_t[8]), .A0_f (key_s0_f[8]), .A1_t (key_s1_t[8]), .A1_f (key_s1_f[8]), .B0_t (KeyArray_outS30ser[0]), .B0_f (new_AGEMA_signal_5157), .B1_t (new_AGEMA_signal_5158), .B1_f (new_AGEMA_signal_5159), .Z0_t (KeyArray_MUX_inS23ser_mux_inst_0_X), .Z0_f (new_AGEMA_signal_5160), .Z1_t (new_AGEMA_signal_5161), .Z1_f (new_AGEMA_signal_5162) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS23ser_mux_inst_0_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS23ser_mux_inst_0_X), .B0_f (new_AGEMA_signal_5160), .B1_t (new_AGEMA_signal_5161), .B1_f (new_AGEMA_signal_5162), .Z0_t (KeyArray_MUX_inS23ser_mux_inst_0_Y), .Z0_f (new_AGEMA_signal_6376), .Z1_t (new_AGEMA_signal_6377), .Z1_f (new_AGEMA_signal_6378) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS23ser_mux_inst_0_XOR2_U1 ( .A0_t (KeyArray_MUX_inS23ser_mux_inst_0_Y), .A0_f (new_AGEMA_signal_6376), .A1_t (new_AGEMA_signal_6377), .A1_f (new_AGEMA_signal_6378), .B0_t (key_s0_t[8]), .B0_f (key_s0_f[8]), .B1_t (key_s1_t[8]), .B1_f (key_s1_f[8]), .Z0_t (KeyArray_inS23ser[0]), .Z0_f (new_AGEMA_signal_7150), .Z1_t (new_AGEMA_signal_7151), .Z1_f (new_AGEMA_signal_7152) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS23ser_mux_inst_1_XOR1_U1 ( .A0_t (key_s0_t[9]), .A0_f (key_s0_f[9]), .A1_t (key_s1_t[9]), .A1_f (key_s1_f[9]), .B0_t (KeyArray_outS30ser[1]), .B0_f (new_AGEMA_signal_5166), .B1_t (new_AGEMA_signal_5167), .B1_f (new_AGEMA_signal_5168), .Z0_t (KeyArray_MUX_inS23ser_mux_inst_1_X), .Z0_f (new_AGEMA_signal_5169), .Z1_t (new_AGEMA_signal_5170), .Z1_f (new_AGEMA_signal_5171) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS23ser_mux_inst_1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS23ser_mux_inst_1_X), .B0_f (new_AGEMA_signal_5169), .B1_t (new_AGEMA_signal_5170), .B1_f (new_AGEMA_signal_5171), .Z0_t (KeyArray_MUX_inS23ser_mux_inst_1_Y), .Z0_f (new_AGEMA_signal_6379), .Z1_t (new_AGEMA_signal_6380), .Z1_f (new_AGEMA_signal_6381) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS23ser_mux_inst_1_XOR2_U1 ( .A0_t (KeyArray_MUX_inS23ser_mux_inst_1_Y), .A0_f (new_AGEMA_signal_6379), .A1_t (new_AGEMA_signal_6380), .A1_f (new_AGEMA_signal_6381), .B0_t (key_s0_t[9]), .B0_f (key_s0_f[9]), .B1_t (key_s1_t[9]), .B1_f (key_s1_f[9]), .Z0_t (KeyArray_inS23ser[1]), .Z0_f (new_AGEMA_signal_7153), .Z1_t (new_AGEMA_signal_7154), .Z1_f (new_AGEMA_signal_7155) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS23ser_mux_inst_2_XOR1_U1 ( .A0_t (key_s0_t[10]), .A0_f (key_s0_f[10]), .A1_t (key_s1_t[10]), .A1_f (key_s1_f[10]), .B0_t (KeyArray_outS30ser[2]), .B0_f (new_AGEMA_signal_5175), .B1_t (new_AGEMA_signal_5176), .B1_f (new_AGEMA_signal_5177), .Z0_t (KeyArray_MUX_inS23ser_mux_inst_2_X), .Z0_f (new_AGEMA_signal_5178), .Z1_t (new_AGEMA_signal_5179), .Z1_f (new_AGEMA_signal_5180) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS23ser_mux_inst_2_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS23ser_mux_inst_2_X), .B0_f (new_AGEMA_signal_5178), .B1_t (new_AGEMA_signal_5179), .B1_f (new_AGEMA_signal_5180), .Z0_t (KeyArray_MUX_inS23ser_mux_inst_2_Y), .Z0_f (new_AGEMA_signal_6382), .Z1_t (new_AGEMA_signal_6383), .Z1_f (new_AGEMA_signal_6384) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS23ser_mux_inst_2_XOR2_U1 ( .A0_t (KeyArray_MUX_inS23ser_mux_inst_2_Y), .A0_f (new_AGEMA_signal_6382), .A1_t (new_AGEMA_signal_6383), .A1_f (new_AGEMA_signal_6384), .B0_t (key_s0_t[10]), .B0_f (key_s0_f[10]), .B1_t (key_s1_t[10]), .B1_f (key_s1_f[10]), .Z0_t (KeyArray_inS23ser[2]), .Z0_f (new_AGEMA_signal_7156), .Z1_t (new_AGEMA_signal_7157), .Z1_f (new_AGEMA_signal_7158) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS23ser_mux_inst_3_XOR1_U1 ( .A0_t (key_s0_t[11]), .A0_f (key_s0_f[11]), .A1_t (key_s1_t[11]), .A1_f (key_s1_f[11]), .B0_t (KeyArray_outS30ser[3]), .B0_f (new_AGEMA_signal_5184), .B1_t (new_AGEMA_signal_5185), .B1_f (new_AGEMA_signal_5186), .Z0_t (KeyArray_MUX_inS23ser_mux_inst_3_X), .Z0_f (new_AGEMA_signal_5187), .Z1_t (new_AGEMA_signal_5188), .Z1_f (new_AGEMA_signal_5189) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS23ser_mux_inst_3_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS23ser_mux_inst_3_X), .B0_f (new_AGEMA_signal_5187), .B1_t (new_AGEMA_signal_5188), .B1_f (new_AGEMA_signal_5189), .Z0_t (KeyArray_MUX_inS23ser_mux_inst_3_Y), .Z0_f (new_AGEMA_signal_6385), .Z1_t (new_AGEMA_signal_6386), .Z1_f (new_AGEMA_signal_6387) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS23ser_mux_inst_3_XOR2_U1 ( .A0_t (KeyArray_MUX_inS23ser_mux_inst_3_Y), .A0_f (new_AGEMA_signal_6385), .A1_t (new_AGEMA_signal_6386), .A1_f (new_AGEMA_signal_6387), .B0_t (key_s0_t[11]), .B0_f (key_s0_f[11]), .B1_t (key_s1_t[11]), .B1_f (key_s1_f[11]), .Z0_t (KeyArray_inS23ser[3]), .Z0_f (new_AGEMA_signal_7159), .Z1_t (new_AGEMA_signal_7160), .Z1_f (new_AGEMA_signal_7161) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS23ser_mux_inst_4_XOR1_U1 ( .A0_t (key_s0_t[12]), .A0_f (key_s0_f[12]), .A1_t (key_s1_t[12]), .A1_f (key_s1_f[12]), .B0_t (KeyArray_outS30ser[4]), .B0_f (new_AGEMA_signal_5193), .B1_t (new_AGEMA_signal_5194), .B1_f (new_AGEMA_signal_5195), .Z0_t (KeyArray_MUX_inS23ser_mux_inst_4_X), .Z0_f (new_AGEMA_signal_5196), .Z1_t (new_AGEMA_signal_5197), .Z1_f (new_AGEMA_signal_5198) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS23ser_mux_inst_4_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS23ser_mux_inst_4_X), .B0_f (new_AGEMA_signal_5196), .B1_t (new_AGEMA_signal_5197), .B1_f (new_AGEMA_signal_5198), .Z0_t (KeyArray_MUX_inS23ser_mux_inst_4_Y), .Z0_f (new_AGEMA_signal_6388), .Z1_t (new_AGEMA_signal_6389), .Z1_f (new_AGEMA_signal_6390) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS23ser_mux_inst_4_XOR2_U1 ( .A0_t (KeyArray_MUX_inS23ser_mux_inst_4_Y), .A0_f (new_AGEMA_signal_6388), .A1_t (new_AGEMA_signal_6389), .A1_f (new_AGEMA_signal_6390), .B0_t (key_s0_t[12]), .B0_f (key_s0_f[12]), .B1_t (key_s1_t[12]), .B1_f (key_s1_f[12]), .Z0_t (KeyArray_inS23ser[4]), .Z0_f (new_AGEMA_signal_7162), .Z1_t (new_AGEMA_signal_7163), .Z1_f (new_AGEMA_signal_7164) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS23ser_mux_inst_5_XOR1_U1 ( .A0_t (key_s0_t[13]), .A0_f (key_s0_f[13]), .A1_t (key_s1_t[13]), .A1_f (key_s1_f[13]), .B0_t (KeyArray_outS30ser[5]), .B0_f (new_AGEMA_signal_5202), .B1_t (new_AGEMA_signal_5203), .B1_f (new_AGEMA_signal_5204), .Z0_t (KeyArray_MUX_inS23ser_mux_inst_5_X), .Z0_f (new_AGEMA_signal_5205), .Z1_t (new_AGEMA_signal_5206), .Z1_f (new_AGEMA_signal_5207) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS23ser_mux_inst_5_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS23ser_mux_inst_5_X), .B0_f (new_AGEMA_signal_5205), .B1_t (new_AGEMA_signal_5206), .B1_f (new_AGEMA_signal_5207), .Z0_t (KeyArray_MUX_inS23ser_mux_inst_5_Y), .Z0_f (new_AGEMA_signal_6391), .Z1_t (new_AGEMA_signal_6392), .Z1_f (new_AGEMA_signal_6393) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS23ser_mux_inst_5_XOR2_U1 ( .A0_t (KeyArray_MUX_inS23ser_mux_inst_5_Y), .A0_f (new_AGEMA_signal_6391), .A1_t (new_AGEMA_signal_6392), .A1_f (new_AGEMA_signal_6393), .B0_t (key_s0_t[13]), .B0_f (key_s0_f[13]), .B1_t (key_s1_t[13]), .B1_f (key_s1_f[13]), .Z0_t (KeyArray_inS23ser[5]), .Z0_f (new_AGEMA_signal_7165), .Z1_t (new_AGEMA_signal_7166), .Z1_f (new_AGEMA_signal_7167) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS23ser_mux_inst_6_XOR1_U1 ( .A0_t (key_s0_t[14]), .A0_f (key_s0_f[14]), .A1_t (key_s1_t[14]), .A1_f (key_s1_f[14]), .B0_t (KeyArray_outS30ser[6]), .B0_f (new_AGEMA_signal_5211), .B1_t (new_AGEMA_signal_5212), .B1_f (new_AGEMA_signal_5213), .Z0_t (KeyArray_MUX_inS23ser_mux_inst_6_X), .Z0_f (new_AGEMA_signal_5214), .Z1_t (new_AGEMA_signal_5215), .Z1_f (new_AGEMA_signal_5216) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS23ser_mux_inst_6_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS23ser_mux_inst_6_X), .B0_f (new_AGEMA_signal_5214), .B1_t (new_AGEMA_signal_5215), .B1_f (new_AGEMA_signal_5216), .Z0_t (KeyArray_MUX_inS23ser_mux_inst_6_Y), .Z0_f (new_AGEMA_signal_6394), .Z1_t (new_AGEMA_signal_6395), .Z1_f (new_AGEMA_signal_6396) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS23ser_mux_inst_6_XOR2_U1 ( .A0_t (KeyArray_MUX_inS23ser_mux_inst_6_Y), .A0_f (new_AGEMA_signal_6394), .A1_t (new_AGEMA_signal_6395), .A1_f (new_AGEMA_signal_6396), .B0_t (key_s0_t[14]), .B0_f (key_s0_f[14]), .B1_t (key_s1_t[14]), .B1_f (key_s1_f[14]), .Z0_t (KeyArray_inS23ser[6]), .Z0_f (new_AGEMA_signal_7168), .Z1_t (new_AGEMA_signal_7169), .Z1_f (new_AGEMA_signal_7170) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS23ser_mux_inst_7_XOR1_U1 ( .A0_t (key_s0_t[15]), .A0_f (key_s0_f[15]), .A1_t (key_s1_t[15]), .A1_f (key_s1_f[15]), .B0_t (KeyArray_outS30ser[7]), .B0_f (new_AGEMA_signal_5220), .B1_t (new_AGEMA_signal_5221), .B1_f (new_AGEMA_signal_5222), .Z0_t (KeyArray_MUX_inS23ser_mux_inst_7_X), .Z0_f (new_AGEMA_signal_5223), .Z1_t (new_AGEMA_signal_5224), .Z1_f (new_AGEMA_signal_5225) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS23ser_mux_inst_7_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS23ser_mux_inst_7_X), .B0_f (new_AGEMA_signal_5223), .B1_t (new_AGEMA_signal_5224), .B1_f (new_AGEMA_signal_5225), .Z0_t (KeyArray_MUX_inS23ser_mux_inst_7_Y), .Z0_f (new_AGEMA_signal_6397), .Z1_t (new_AGEMA_signal_6398), .Z1_f (new_AGEMA_signal_6399) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS23ser_mux_inst_7_XOR2_U1 ( .A0_t (KeyArray_MUX_inS23ser_mux_inst_7_Y), .A0_f (new_AGEMA_signal_6397), .A1_t (new_AGEMA_signal_6398), .A1_f (new_AGEMA_signal_6399), .B0_t (key_s0_t[15]), .B0_f (key_s0_f[15]), .B1_t (key_s1_t[15]), .B1_f (key_s1_f[15]), .Z0_t (KeyArray_inS23ser[7]), .Z0_f (new_AGEMA_signal_7171), .Z1_t (new_AGEMA_signal_7172), .Z1_f (new_AGEMA_signal_7173) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS30ser_mux_inst_0_XOR1_U1 ( .A0_t (key_s0_t[96]), .A0_f (key_s0_f[96]), .A1_t (key_s1_t[96]), .A1_f (key_s1_f[96]), .B0_t (KeyArray_outS31ser[0]), .B0_f (new_AGEMA_signal_5229), .B1_t (new_AGEMA_signal_5230), .B1_f (new_AGEMA_signal_5231), .Z0_t (KeyArray_MUX_inS30ser_mux_inst_0_X), .Z0_f (new_AGEMA_signal_5232), .Z1_t (new_AGEMA_signal_5233), .Z1_f (new_AGEMA_signal_5234) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS30ser_mux_inst_0_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS30ser_mux_inst_0_X), .B0_f (new_AGEMA_signal_5232), .B1_t (new_AGEMA_signal_5233), .B1_f (new_AGEMA_signal_5234), .Z0_t (KeyArray_MUX_inS30ser_mux_inst_0_Y), .Z0_f (new_AGEMA_signal_6400), .Z1_t (new_AGEMA_signal_6401), .Z1_f (new_AGEMA_signal_6402) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS30ser_mux_inst_0_XOR2_U1 ( .A0_t (KeyArray_MUX_inS30ser_mux_inst_0_Y), .A0_f (new_AGEMA_signal_6400), .A1_t (new_AGEMA_signal_6401), .A1_f (new_AGEMA_signal_6402), .B0_t (key_s0_t[96]), .B0_f (key_s0_f[96]), .B1_t (key_s1_t[96]), .B1_f (key_s1_f[96]), .Z0_t (KeyArray_inS30ser[0]), .Z0_f (new_AGEMA_signal_7174), .Z1_t (new_AGEMA_signal_7175), .Z1_f (new_AGEMA_signal_7176) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS30ser_mux_inst_1_XOR1_U1 ( .A0_t (key_s0_t[97]), .A0_f (key_s0_f[97]), .A1_t (key_s1_t[97]), .A1_f (key_s1_f[97]), .B0_t (KeyArray_outS31ser[1]), .B0_f (new_AGEMA_signal_5238), .B1_t (new_AGEMA_signal_5239), .B1_f (new_AGEMA_signal_5240), .Z0_t (KeyArray_MUX_inS30ser_mux_inst_1_X), .Z0_f (new_AGEMA_signal_5241), .Z1_t (new_AGEMA_signal_5242), .Z1_f (new_AGEMA_signal_5243) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS30ser_mux_inst_1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS30ser_mux_inst_1_X), .B0_f (new_AGEMA_signal_5241), .B1_t (new_AGEMA_signal_5242), .B1_f (new_AGEMA_signal_5243), .Z0_t (KeyArray_MUX_inS30ser_mux_inst_1_Y), .Z0_f (new_AGEMA_signal_6403), .Z1_t (new_AGEMA_signal_6404), .Z1_f (new_AGEMA_signal_6405) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS30ser_mux_inst_1_XOR2_U1 ( .A0_t (KeyArray_MUX_inS30ser_mux_inst_1_Y), .A0_f (new_AGEMA_signal_6403), .A1_t (new_AGEMA_signal_6404), .A1_f (new_AGEMA_signal_6405), .B0_t (key_s0_t[97]), .B0_f (key_s0_f[97]), .B1_t (key_s1_t[97]), .B1_f (key_s1_f[97]), .Z0_t (KeyArray_inS30ser[1]), .Z0_f (new_AGEMA_signal_7177), .Z1_t (new_AGEMA_signal_7178), .Z1_f (new_AGEMA_signal_7179) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS30ser_mux_inst_2_XOR1_U1 ( .A0_t (key_s0_t[98]), .A0_f (key_s0_f[98]), .A1_t (key_s1_t[98]), .A1_f (key_s1_f[98]), .B0_t (KeyArray_outS31ser[2]), .B0_f (new_AGEMA_signal_5247), .B1_t (new_AGEMA_signal_5248), .B1_f (new_AGEMA_signal_5249), .Z0_t (KeyArray_MUX_inS30ser_mux_inst_2_X), .Z0_f (new_AGEMA_signal_5250), .Z1_t (new_AGEMA_signal_5251), .Z1_f (new_AGEMA_signal_5252) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS30ser_mux_inst_2_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS30ser_mux_inst_2_X), .B0_f (new_AGEMA_signal_5250), .B1_t (new_AGEMA_signal_5251), .B1_f (new_AGEMA_signal_5252), .Z0_t (KeyArray_MUX_inS30ser_mux_inst_2_Y), .Z0_f (new_AGEMA_signal_6406), .Z1_t (new_AGEMA_signal_6407), .Z1_f (new_AGEMA_signal_6408) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS30ser_mux_inst_2_XOR2_U1 ( .A0_t (KeyArray_MUX_inS30ser_mux_inst_2_Y), .A0_f (new_AGEMA_signal_6406), .A1_t (new_AGEMA_signal_6407), .A1_f (new_AGEMA_signal_6408), .B0_t (key_s0_t[98]), .B0_f (key_s0_f[98]), .B1_t (key_s1_t[98]), .B1_f (key_s1_f[98]), .Z0_t (KeyArray_inS30ser[2]), .Z0_f (new_AGEMA_signal_7180), .Z1_t (new_AGEMA_signal_7181), .Z1_f (new_AGEMA_signal_7182) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS30ser_mux_inst_3_XOR1_U1 ( .A0_t (key_s0_t[99]), .A0_f (key_s0_f[99]), .A1_t (key_s1_t[99]), .A1_f (key_s1_f[99]), .B0_t (KeyArray_outS31ser[3]), .B0_f (new_AGEMA_signal_5256), .B1_t (new_AGEMA_signal_5257), .B1_f (new_AGEMA_signal_5258), .Z0_t (KeyArray_MUX_inS30ser_mux_inst_3_X), .Z0_f (new_AGEMA_signal_5259), .Z1_t (new_AGEMA_signal_5260), .Z1_f (new_AGEMA_signal_5261) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS30ser_mux_inst_3_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS30ser_mux_inst_3_X), .B0_f (new_AGEMA_signal_5259), .B1_t (new_AGEMA_signal_5260), .B1_f (new_AGEMA_signal_5261), .Z0_t (KeyArray_MUX_inS30ser_mux_inst_3_Y), .Z0_f (new_AGEMA_signal_6409), .Z1_t (new_AGEMA_signal_6410), .Z1_f (new_AGEMA_signal_6411) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS30ser_mux_inst_3_XOR2_U1 ( .A0_t (KeyArray_MUX_inS30ser_mux_inst_3_Y), .A0_f (new_AGEMA_signal_6409), .A1_t (new_AGEMA_signal_6410), .A1_f (new_AGEMA_signal_6411), .B0_t (key_s0_t[99]), .B0_f (key_s0_f[99]), .B1_t (key_s1_t[99]), .B1_f (key_s1_f[99]), .Z0_t (KeyArray_inS30ser[3]), .Z0_f (new_AGEMA_signal_7183), .Z1_t (new_AGEMA_signal_7184), .Z1_f (new_AGEMA_signal_7185) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS30ser_mux_inst_4_XOR1_U1 ( .A0_t (key_s0_t[100]), .A0_f (key_s0_f[100]), .A1_t (key_s1_t[100]), .A1_f (key_s1_f[100]), .B0_t (KeyArray_outS31ser[4]), .B0_f (new_AGEMA_signal_5265), .B1_t (new_AGEMA_signal_5266), .B1_f (new_AGEMA_signal_5267), .Z0_t (KeyArray_MUX_inS30ser_mux_inst_4_X), .Z0_f (new_AGEMA_signal_5268), .Z1_t (new_AGEMA_signal_5269), .Z1_f (new_AGEMA_signal_5270) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS30ser_mux_inst_4_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS30ser_mux_inst_4_X), .B0_f (new_AGEMA_signal_5268), .B1_t (new_AGEMA_signal_5269), .B1_f (new_AGEMA_signal_5270), .Z0_t (KeyArray_MUX_inS30ser_mux_inst_4_Y), .Z0_f (new_AGEMA_signal_6412), .Z1_t (new_AGEMA_signal_6413), .Z1_f (new_AGEMA_signal_6414) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS30ser_mux_inst_4_XOR2_U1 ( .A0_t (KeyArray_MUX_inS30ser_mux_inst_4_Y), .A0_f (new_AGEMA_signal_6412), .A1_t (new_AGEMA_signal_6413), .A1_f (new_AGEMA_signal_6414), .B0_t (key_s0_t[100]), .B0_f (key_s0_f[100]), .B1_t (key_s1_t[100]), .B1_f (key_s1_f[100]), .Z0_t (KeyArray_inS30ser[4]), .Z0_f (new_AGEMA_signal_7186), .Z1_t (new_AGEMA_signal_7187), .Z1_f (new_AGEMA_signal_7188) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS30ser_mux_inst_5_XOR1_U1 ( .A0_t (key_s0_t[101]), .A0_f (key_s0_f[101]), .A1_t (key_s1_t[101]), .A1_f (key_s1_f[101]), .B0_t (KeyArray_outS31ser[5]), .B0_f (new_AGEMA_signal_5274), .B1_t (new_AGEMA_signal_5275), .B1_f (new_AGEMA_signal_5276), .Z0_t (KeyArray_MUX_inS30ser_mux_inst_5_X), .Z0_f (new_AGEMA_signal_5277), .Z1_t (new_AGEMA_signal_5278), .Z1_f (new_AGEMA_signal_5279) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS30ser_mux_inst_5_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS30ser_mux_inst_5_X), .B0_f (new_AGEMA_signal_5277), .B1_t (new_AGEMA_signal_5278), .B1_f (new_AGEMA_signal_5279), .Z0_t (KeyArray_MUX_inS30ser_mux_inst_5_Y), .Z0_f (new_AGEMA_signal_6415), .Z1_t (new_AGEMA_signal_6416), .Z1_f (new_AGEMA_signal_6417) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS30ser_mux_inst_5_XOR2_U1 ( .A0_t (KeyArray_MUX_inS30ser_mux_inst_5_Y), .A0_f (new_AGEMA_signal_6415), .A1_t (new_AGEMA_signal_6416), .A1_f (new_AGEMA_signal_6417), .B0_t (key_s0_t[101]), .B0_f (key_s0_f[101]), .B1_t (key_s1_t[101]), .B1_f (key_s1_f[101]), .Z0_t (KeyArray_inS30ser[5]), .Z0_f (new_AGEMA_signal_7189), .Z1_t (new_AGEMA_signal_7190), .Z1_f (new_AGEMA_signal_7191) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS30ser_mux_inst_6_XOR1_U1 ( .A0_t (key_s0_t[102]), .A0_f (key_s0_f[102]), .A1_t (key_s1_t[102]), .A1_f (key_s1_f[102]), .B0_t (KeyArray_outS31ser[6]), .B0_f (new_AGEMA_signal_5283), .B1_t (new_AGEMA_signal_5284), .B1_f (new_AGEMA_signal_5285), .Z0_t (KeyArray_MUX_inS30ser_mux_inst_6_X), .Z0_f (new_AGEMA_signal_5286), .Z1_t (new_AGEMA_signal_5287), .Z1_f (new_AGEMA_signal_5288) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS30ser_mux_inst_6_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS30ser_mux_inst_6_X), .B0_f (new_AGEMA_signal_5286), .B1_t (new_AGEMA_signal_5287), .B1_f (new_AGEMA_signal_5288), .Z0_t (KeyArray_MUX_inS30ser_mux_inst_6_Y), .Z0_f (new_AGEMA_signal_6418), .Z1_t (new_AGEMA_signal_6419), .Z1_f (new_AGEMA_signal_6420) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS30ser_mux_inst_6_XOR2_U1 ( .A0_t (KeyArray_MUX_inS30ser_mux_inst_6_Y), .A0_f (new_AGEMA_signal_6418), .A1_t (new_AGEMA_signal_6419), .A1_f (new_AGEMA_signal_6420), .B0_t (key_s0_t[102]), .B0_f (key_s0_f[102]), .B1_t (key_s1_t[102]), .B1_f (key_s1_f[102]), .Z0_t (KeyArray_inS30ser[6]), .Z0_f (new_AGEMA_signal_7192), .Z1_t (new_AGEMA_signal_7193), .Z1_f (new_AGEMA_signal_7194) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS30ser_mux_inst_7_XOR1_U1 ( .A0_t (key_s0_t[103]), .A0_f (key_s0_f[103]), .A1_t (key_s1_t[103]), .A1_f (key_s1_f[103]), .B0_t (KeyArray_outS31ser[7]), .B0_f (new_AGEMA_signal_5292), .B1_t (new_AGEMA_signal_5293), .B1_f (new_AGEMA_signal_5294), .Z0_t (KeyArray_MUX_inS30ser_mux_inst_7_X), .Z0_f (new_AGEMA_signal_5295), .Z1_t (new_AGEMA_signal_5296), .Z1_f (new_AGEMA_signal_5297) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS30ser_mux_inst_7_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS30ser_mux_inst_7_X), .B0_f (new_AGEMA_signal_5295), .B1_t (new_AGEMA_signal_5296), .B1_f (new_AGEMA_signal_5297), .Z0_t (KeyArray_MUX_inS30ser_mux_inst_7_Y), .Z0_f (new_AGEMA_signal_6421), .Z1_t (new_AGEMA_signal_6422), .Z1_f (new_AGEMA_signal_6423) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS30ser_mux_inst_7_XOR2_U1 ( .A0_t (KeyArray_MUX_inS30ser_mux_inst_7_Y), .A0_f (new_AGEMA_signal_6421), .A1_t (new_AGEMA_signal_6422), .A1_f (new_AGEMA_signal_6423), .B0_t (key_s0_t[103]), .B0_f (key_s0_f[103]), .B1_t (key_s1_t[103]), .B1_f (key_s1_f[103]), .Z0_t (KeyArray_inS30ser[7]), .Z0_f (new_AGEMA_signal_7195), .Z1_t (new_AGEMA_signal_7196), .Z1_f (new_AGEMA_signal_7197) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS31ser_mux_inst_0_XOR1_U1 ( .A0_t (key_s0_t[64]), .A0_f (key_s0_f[64]), .A1_t (key_s1_t[64]), .A1_f (key_s1_f[64]), .B0_t (KeyArray_outS32ser[0]), .B0_f (new_AGEMA_signal_5301), .B1_t (new_AGEMA_signal_5302), .B1_f (new_AGEMA_signal_5303), .Z0_t (KeyArray_MUX_inS31ser_mux_inst_0_X), .Z0_f (new_AGEMA_signal_5304), .Z1_t (new_AGEMA_signal_5305), .Z1_f (new_AGEMA_signal_5306) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS31ser_mux_inst_0_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS31ser_mux_inst_0_X), .B0_f (new_AGEMA_signal_5304), .B1_t (new_AGEMA_signal_5305), .B1_f (new_AGEMA_signal_5306), .Z0_t (KeyArray_MUX_inS31ser_mux_inst_0_Y), .Z0_f (new_AGEMA_signal_6424), .Z1_t (new_AGEMA_signal_6425), .Z1_f (new_AGEMA_signal_6426) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS31ser_mux_inst_0_XOR2_U1 ( .A0_t (KeyArray_MUX_inS31ser_mux_inst_0_Y), .A0_f (new_AGEMA_signal_6424), .A1_t (new_AGEMA_signal_6425), .A1_f (new_AGEMA_signal_6426), .B0_t (key_s0_t[64]), .B0_f (key_s0_f[64]), .B1_t (key_s1_t[64]), .B1_f (key_s1_f[64]), .Z0_t (KeyArray_inS31ser[0]), .Z0_f (new_AGEMA_signal_7198), .Z1_t (new_AGEMA_signal_7199), .Z1_f (new_AGEMA_signal_7200) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS31ser_mux_inst_1_XOR1_U1 ( .A0_t (key_s0_t[65]), .A0_f (key_s0_f[65]), .A1_t (key_s1_t[65]), .A1_f (key_s1_f[65]), .B0_t (KeyArray_outS32ser[1]), .B0_f (new_AGEMA_signal_5310), .B1_t (new_AGEMA_signal_5311), .B1_f (new_AGEMA_signal_5312), .Z0_t (KeyArray_MUX_inS31ser_mux_inst_1_X), .Z0_f (new_AGEMA_signal_5313), .Z1_t (new_AGEMA_signal_5314), .Z1_f (new_AGEMA_signal_5315) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS31ser_mux_inst_1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS31ser_mux_inst_1_X), .B0_f (new_AGEMA_signal_5313), .B1_t (new_AGEMA_signal_5314), .B1_f (new_AGEMA_signal_5315), .Z0_t (KeyArray_MUX_inS31ser_mux_inst_1_Y), .Z0_f (new_AGEMA_signal_6427), .Z1_t (new_AGEMA_signal_6428), .Z1_f (new_AGEMA_signal_6429) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS31ser_mux_inst_1_XOR2_U1 ( .A0_t (KeyArray_MUX_inS31ser_mux_inst_1_Y), .A0_f (new_AGEMA_signal_6427), .A1_t (new_AGEMA_signal_6428), .A1_f (new_AGEMA_signal_6429), .B0_t (key_s0_t[65]), .B0_f (key_s0_f[65]), .B1_t (key_s1_t[65]), .B1_f (key_s1_f[65]), .Z0_t (KeyArray_inS31ser[1]), .Z0_f (new_AGEMA_signal_7201), .Z1_t (new_AGEMA_signal_7202), .Z1_f (new_AGEMA_signal_7203) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS31ser_mux_inst_2_XOR1_U1 ( .A0_t (key_s0_t[66]), .A0_f (key_s0_f[66]), .A1_t (key_s1_t[66]), .A1_f (key_s1_f[66]), .B0_t (KeyArray_outS32ser[2]), .B0_f (new_AGEMA_signal_5319), .B1_t (new_AGEMA_signal_5320), .B1_f (new_AGEMA_signal_5321), .Z0_t (KeyArray_MUX_inS31ser_mux_inst_2_X), .Z0_f (new_AGEMA_signal_5322), .Z1_t (new_AGEMA_signal_5323), .Z1_f (new_AGEMA_signal_5324) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS31ser_mux_inst_2_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS31ser_mux_inst_2_X), .B0_f (new_AGEMA_signal_5322), .B1_t (new_AGEMA_signal_5323), .B1_f (new_AGEMA_signal_5324), .Z0_t (KeyArray_MUX_inS31ser_mux_inst_2_Y), .Z0_f (new_AGEMA_signal_6430), .Z1_t (new_AGEMA_signal_6431), .Z1_f (new_AGEMA_signal_6432) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS31ser_mux_inst_2_XOR2_U1 ( .A0_t (KeyArray_MUX_inS31ser_mux_inst_2_Y), .A0_f (new_AGEMA_signal_6430), .A1_t (new_AGEMA_signal_6431), .A1_f (new_AGEMA_signal_6432), .B0_t (key_s0_t[66]), .B0_f (key_s0_f[66]), .B1_t (key_s1_t[66]), .B1_f (key_s1_f[66]), .Z0_t (KeyArray_inS31ser[2]), .Z0_f (new_AGEMA_signal_7204), .Z1_t (new_AGEMA_signal_7205), .Z1_f (new_AGEMA_signal_7206) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS31ser_mux_inst_3_XOR1_U1 ( .A0_t (key_s0_t[67]), .A0_f (key_s0_f[67]), .A1_t (key_s1_t[67]), .A1_f (key_s1_f[67]), .B0_t (KeyArray_outS32ser[3]), .B0_f (new_AGEMA_signal_5328), .B1_t (new_AGEMA_signal_5329), .B1_f (new_AGEMA_signal_5330), .Z0_t (KeyArray_MUX_inS31ser_mux_inst_3_X), .Z0_f (new_AGEMA_signal_5331), .Z1_t (new_AGEMA_signal_5332), .Z1_f (new_AGEMA_signal_5333) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS31ser_mux_inst_3_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS31ser_mux_inst_3_X), .B0_f (new_AGEMA_signal_5331), .B1_t (new_AGEMA_signal_5332), .B1_f (new_AGEMA_signal_5333), .Z0_t (KeyArray_MUX_inS31ser_mux_inst_3_Y), .Z0_f (new_AGEMA_signal_6433), .Z1_t (new_AGEMA_signal_6434), .Z1_f (new_AGEMA_signal_6435) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS31ser_mux_inst_3_XOR2_U1 ( .A0_t (KeyArray_MUX_inS31ser_mux_inst_3_Y), .A0_f (new_AGEMA_signal_6433), .A1_t (new_AGEMA_signal_6434), .A1_f (new_AGEMA_signal_6435), .B0_t (key_s0_t[67]), .B0_f (key_s0_f[67]), .B1_t (key_s1_t[67]), .B1_f (key_s1_f[67]), .Z0_t (KeyArray_inS31ser[3]), .Z0_f (new_AGEMA_signal_7207), .Z1_t (new_AGEMA_signal_7208), .Z1_f (new_AGEMA_signal_7209) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS31ser_mux_inst_4_XOR1_U1 ( .A0_t (key_s0_t[68]), .A0_f (key_s0_f[68]), .A1_t (key_s1_t[68]), .A1_f (key_s1_f[68]), .B0_t (KeyArray_outS32ser[4]), .B0_f (new_AGEMA_signal_5337), .B1_t (new_AGEMA_signal_5338), .B1_f (new_AGEMA_signal_5339), .Z0_t (KeyArray_MUX_inS31ser_mux_inst_4_X), .Z0_f (new_AGEMA_signal_5340), .Z1_t (new_AGEMA_signal_5341), .Z1_f (new_AGEMA_signal_5342) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS31ser_mux_inst_4_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS31ser_mux_inst_4_X), .B0_f (new_AGEMA_signal_5340), .B1_t (new_AGEMA_signal_5341), .B1_f (new_AGEMA_signal_5342), .Z0_t (KeyArray_MUX_inS31ser_mux_inst_4_Y), .Z0_f (new_AGEMA_signal_6436), .Z1_t (new_AGEMA_signal_6437), .Z1_f (new_AGEMA_signal_6438) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS31ser_mux_inst_4_XOR2_U1 ( .A0_t (KeyArray_MUX_inS31ser_mux_inst_4_Y), .A0_f (new_AGEMA_signal_6436), .A1_t (new_AGEMA_signal_6437), .A1_f (new_AGEMA_signal_6438), .B0_t (key_s0_t[68]), .B0_f (key_s0_f[68]), .B1_t (key_s1_t[68]), .B1_f (key_s1_f[68]), .Z0_t (KeyArray_inS31ser[4]), .Z0_f (new_AGEMA_signal_7210), .Z1_t (new_AGEMA_signal_7211), .Z1_f (new_AGEMA_signal_7212) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS31ser_mux_inst_5_XOR1_U1 ( .A0_t (key_s0_t[69]), .A0_f (key_s0_f[69]), .A1_t (key_s1_t[69]), .A1_f (key_s1_f[69]), .B0_t (KeyArray_outS32ser[5]), .B0_f (new_AGEMA_signal_5346), .B1_t (new_AGEMA_signal_5347), .B1_f (new_AGEMA_signal_5348), .Z0_t (KeyArray_MUX_inS31ser_mux_inst_5_X), .Z0_f (new_AGEMA_signal_5349), .Z1_t (new_AGEMA_signal_5350), .Z1_f (new_AGEMA_signal_5351) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS31ser_mux_inst_5_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS31ser_mux_inst_5_X), .B0_f (new_AGEMA_signal_5349), .B1_t (new_AGEMA_signal_5350), .B1_f (new_AGEMA_signal_5351), .Z0_t (KeyArray_MUX_inS31ser_mux_inst_5_Y), .Z0_f (new_AGEMA_signal_6439), .Z1_t (new_AGEMA_signal_6440), .Z1_f (new_AGEMA_signal_6441) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS31ser_mux_inst_5_XOR2_U1 ( .A0_t (KeyArray_MUX_inS31ser_mux_inst_5_Y), .A0_f (new_AGEMA_signal_6439), .A1_t (new_AGEMA_signal_6440), .A1_f (new_AGEMA_signal_6441), .B0_t (key_s0_t[69]), .B0_f (key_s0_f[69]), .B1_t (key_s1_t[69]), .B1_f (key_s1_f[69]), .Z0_t (KeyArray_inS31ser[5]), .Z0_f (new_AGEMA_signal_7213), .Z1_t (new_AGEMA_signal_7214), .Z1_f (new_AGEMA_signal_7215) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS31ser_mux_inst_6_XOR1_U1 ( .A0_t (key_s0_t[70]), .A0_f (key_s0_f[70]), .A1_t (key_s1_t[70]), .A1_f (key_s1_f[70]), .B0_t (KeyArray_outS32ser[6]), .B0_f (new_AGEMA_signal_5355), .B1_t (new_AGEMA_signal_5356), .B1_f (new_AGEMA_signal_5357), .Z0_t (KeyArray_MUX_inS31ser_mux_inst_6_X), .Z0_f (new_AGEMA_signal_5358), .Z1_t (new_AGEMA_signal_5359), .Z1_f (new_AGEMA_signal_5360) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS31ser_mux_inst_6_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS31ser_mux_inst_6_X), .B0_f (new_AGEMA_signal_5358), .B1_t (new_AGEMA_signal_5359), .B1_f (new_AGEMA_signal_5360), .Z0_t (KeyArray_MUX_inS31ser_mux_inst_6_Y), .Z0_f (new_AGEMA_signal_6442), .Z1_t (new_AGEMA_signal_6443), .Z1_f (new_AGEMA_signal_6444) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS31ser_mux_inst_6_XOR2_U1 ( .A0_t (KeyArray_MUX_inS31ser_mux_inst_6_Y), .A0_f (new_AGEMA_signal_6442), .A1_t (new_AGEMA_signal_6443), .A1_f (new_AGEMA_signal_6444), .B0_t (key_s0_t[70]), .B0_f (key_s0_f[70]), .B1_t (key_s1_t[70]), .B1_f (key_s1_f[70]), .Z0_t (KeyArray_inS31ser[6]), .Z0_f (new_AGEMA_signal_7216), .Z1_t (new_AGEMA_signal_7217), .Z1_f (new_AGEMA_signal_7218) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS31ser_mux_inst_7_XOR1_U1 ( .A0_t (key_s0_t[71]), .A0_f (key_s0_f[71]), .A1_t (key_s1_t[71]), .A1_f (key_s1_f[71]), .B0_t (KeyArray_outS32ser[7]), .B0_f (new_AGEMA_signal_5364), .B1_t (new_AGEMA_signal_5365), .B1_f (new_AGEMA_signal_5366), .Z0_t (KeyArray_MUX_inS31ser_mux_inst_7_X), .Z0_f (new_AGEMA_signal_5367), .Z1_t (new_AGEMA_signal_5368), .Z1_f (new_AGEMA_signal_5369) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS31ser_mux_inst_7_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS31ser_mux_inst_7_X), .B0_f (new_AGEMA_signal_5367), .B1_t (new_AGEMA_signal_5368), .B1_f (new_AGEMA_signal_5369), .Z0_t (KeyArray_MUX_inS31ser_mux_inst_7_Y), .Z0_f (new_AGEMA_signal_6445), .Z1_t (new_AGEMA_signal_6446), .Z1_f (new_AGEMA_signal_6447) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS31ser_mux_inst_7_XOR2_U1 ( .A0_t (KeyArray_MUX_inS31ser_mux_inst_7_Y), .A0_f (new_AGEMA_signal_6445), .A1_t (new_AGEMA_signal_6446), .A1_f (new_AGEMA_signal_6447), .B0_t (key_s0_t[71]), .B0_f (key_s0_f[71]), .B1_t (key_s1_t[71]), .B1_f (key_s1_f[71]), .Z0_t (KeyArray_inS31ser[7]), .Z0_f (new_AGEMA_signal_7219), .Z1_t (new_AGEMA_signal_7220), .Z1_f (new_AGEMA_signal_7221) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS32ser_mux_inst_0_XOR1_U1 ( .A0_t (key_s0_t[32]), .A0_f (key_s0_f[32]), .A1_t (key_s1_t[32]), .A1_f (key_s1_f[32]), .B0_t (KeyArray_outS33ser[0]), .B0_f (new_AGEMA_signal_5373), .B1_t (new_AGEMA_signal_5374), .B1_f (new_AGEMA_signal_5375), .Z0_t (KeyArray_MUX_inS32ser_mux_inst_0_X), .Z0_f (new_AGEMA_signal_5376), .Z1_t (new_AGEMA_signal_5377), .Z1_f (new_AGEMA_signal_5378) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS32ser_mux_inst_0_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS32ser_mux_inst_0_X), .B0_f (new_AGEMA_signal_5376), .B1_t (new_AGEMA_signal_5377), .B1_f (new_AGEMA_signal_5378), .Z0_t (KeyArray_MUX_inS32ser_mux_inst_0_Y), .Z0_f (new_AGEMA_signal_6448), .Z1_t (new_AGEMA_signal_6449), .Z1_f (new_AGEMA_signal_6450) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS32ser_mux_inst_0_XOR2_U1 ( .A0_t (KeyArray_MUX_inS32ser_mux_inst_0_Y), .A0_f (new_AGEMA_signal_6448), .A1_t (new_AGEMA_signal_6449), .A1_f (new_AGEMA_signal_6450), .B0_t (key_s0_t[32]), .B0_f (key_s0_f[32]), .B1_t (key_s1_t[32]), .B1_f (key_s1_f[32]), .Z0_t (KeyArray_inS32ser[0]), .Z0_f (new_AGEMA_signal_7222), .Z1_t (new_AGEMA_signal_7223), .Z1_f (new_AGEMA_signal_7224) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS32ser_mux_inst_1_XOR1_U1 ( .A0_t (key_s0_t[33]), .A0_f (key_s0_f[33]), .A1_t (key_s1_t[33]), .A1_f (key_s1_f[33]), .B0_t (KeyArray_outS33ser[1]), .B0_f (new_AGEMA_signal_5382), .B1_t (new_AGEMA_signal_5383), .B1_f (new_AGEMA_signal_5384), .Z0_t (KeyArray_MUX_inS32ser_mux_inst_1_X), .Z0_f (new_AGEMA_signal_5385), .Z1_t (new_AGEMA_signal_5386), .Z1_f (new_AGEMA_signal_5387) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS32ser_mux_inst_1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS32ser_mux_inst_1_X), .B0_f (new_AGEMA_signal_5385), .B1_t (new_AGEMA_signal_5386), .B1_f (new_AGEMA_signal_5387), .Z0_t (KeyArray_MUX_inS32ser_mux_inst_1_Y), .Z0_f (new_AGEMA_signal_6451), .Z1_t (new_AGEMA_signal_6452), .Z1_f (new_AGEMA_signal_6453) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS32ser_mux_inst_1_XOR2_U1 ( .A0_t (KeyArray_MUX_inS32ser_mux_inst_1_Y), .A0_f (new_AGEMA_signal_6451), .A1_t (new_AGEMA_signal_6452), .A1_f (new_AGEMA_signal_6453), .B0_t (key_s0_t[33]), .B0_f (key_s0_f[33]), .B1_t (key_s1_t[33]), .B1_f (key_s1_f[33]), .Z0_t (KeyArray_inS32ser[1]), .Z0_f (new_AGEMA_signal_7225), .Z1_t (new_AGEMA_signal_7226), .Z1_f (new_AGEMA_signal_7227) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS32ser_mux_inst_2_XOR1_U1 ( .A0_t (key_s0_t[34]), .A0_f (key_s0_f[34]), .A1_t (key_s1_t[34]), .A1_f (key_s1_f[34]), .B0_t (KeyArray_outS33ser[2]), .B0_f (new_AGEMA_signal_5391), .B1_t (new_AGEMA_signal_5392), .B1_f (new_AGEMA_signal_5393), .Z0_t (KeyArray_MUX_inS32ser_mux_inst_2_X), .Z0_f (new_AGEMA_signal_5394), .Z1_t (new_AGEMA_signal_5395), .Z1_f (new_AGEMA_signal_5396) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS32ser_mux_inst_2_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS32ser_mux_inst_2_X), .B0_f (new_AGEMA_signal_5394), .B1_t (new_AGEMA_signal_5395), .B1_f (new_AGEMA_signal_5396), .Z0_t (KeyArray_MUX_inS32ser_mux_inst_2_Y), .Z0_f (new_AGEMA_signal_6454), .Z1_t (new_AGEMA_signal_6455), .Z1_f (new_AGEMA_signal_6456) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS32ser_mux_inst_2_XOR2_U1 ( .A0_t (KeyArray_MUX_inS32ser_mux_inst_2_Y), .A0_f (new_AGEMA_signal_6454), .A1_t (new_AGEMA_signal_6455), .A1_f (new_AGEMA_signal_6456), .B0_t (key_s0_t[34]), .B0_f (key_s0_f[34]), .B1_t (key_s1_t[34]), .B1_f (key_s1_f[34]), .Z0_t (KeyArray_inS32ser[2]), .Z0_f (new_AGEMA_signal_7228), .Z1_t (new_AGEMA_signal_7229), .Z1_f (new_AGEMA_signal_7230) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS32ser_mux_inst_3_XOR1_U1 ( .A0_t (key_s0_t[35]), .A0_f (key_s0_f[35]), .A1_t (key_s1_t[35]), .A1_f (key_s1_f[35]), .B0_t (KeyArray_outS33ser[3]), .B0_f (new_AGEMA_signal_5400), .B1_t (new_AGEMA_signal_5401), .B1_f (new_AGEMA_signal_5402), .Z0_t (KeyArray_MUX_inS32ser_mux_inst_3_X), .Z0_f (new_AGEMA_signal_5403), .Z1_t (new_AGEMA_signal_5404), .Z1_f (new_AGEMA_signal_5405) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS32ser_mux_inst_3_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS32ser_mux_inst_3_X), .B0_f (new_AGEMA_signal_5403), .B1_t (new_AGEMA_signal_5404), .B1_f (new_AGEMA_signal_5405), .Z0_t (KeyArray_MUX_inS32ser_mux_inst_3_Y), .Z0_f (new_AGEMA_signal_6457), .Z1_t (new_AGEMA_signal_6458), .Z1_f (new_AGEMA_signal_6459) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS32ser_mux_inst_3_XOR2_U1 ( .A0_t (KeyArray_MUX_inS32ser_mux_inst_3_Y), .A0_f (new_AGEMA_signal_6457), .A1_t (new_AGEMA_signal_6458), .A1_f (new_AGEMA_signal_6459), .B0_t (key_s0_t[35]), .B0_f (key_s0_f[35]), .B1_t (key_s1_t[35]), .B1_f (key_s1_f[35]), .Z0_t (KeyArray_inS32ser[3]), .Z0_f (new_AGEMA_signal_7231), .Z1_t (new_AGEMA_signal_7232), .Z1_f (new_AGEMA_signal_7233) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS32ser_mux_inst_4_XOR1_U1 ( .A0_t (key_s0_t[36]), .A0_f (key_s0_f[36]), .A1_t (key_s1_t[36]), .A1_f (key_s1_f[36]), .B0_t (KeyArray_outS33ser[4]), .B0_f (new_AGEMA_signal_5409), .B1_t (new_AGEMA_signal_5410), .B1_f (new_AGEMA_signal_5411), .Z0_t (KeyArray_MUX_inS32ser_mux_inst_4_X), .Z0_f (new_AGEMA_signal_5412), .Z1_t (new_AGEMA_signal_5413), .Z1_f (new_AGEMA_signal_5414) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS32ser_mux_inst_4_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS32ser_mux_inst_4_X), .B0_f (new_AGEMA_signal_5412), .B1_t (new_AGEMA_signal_5413), .B1_f (new_AGEMA_signal_5414), .Z0_t (KeyArray_MUX_inS32ser_mux_inst_4_Y), .Z0_f (new_AGEMA_signal_6460), .Z1_t (new_AGEMA_signal_6461), .Z1_f (new_AGEMA_signal_6462) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS32ser_mux_inst_4_XOR2_U1 ( .A0_t (KeyArray_MUX_inS32ser_mux_inst_4_Y), .A0_f (new_AGEMA_signal_6460), .A1_t (new_AGEMA_signal_6461), .A1_f (new_AGEMA_signal_6462), .B0_t (key_s0_t[36]), .B0_f (key_s0_f[36]), .B1_t (key_s1_t[36]), .B1_f (key_s1_f[36]), .Z0_t (KeyArray_inS32ser[4]), .Z0_f (new_AGEMA_signal_7234), .Z1_t (new_AGEMA_signal_7235), .Z1_f (new_AGEMA_signal_7236) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS32ser_mux_inst_5_XOR1_U1 ( .A0_t (key_s0_t[37]), .A0_f (key_s0_f[37]), .A1_t (key_s1_t[37]), .A1_f (key_s1_f[37]), .B0_t (KeyArray_outS33ser[5]), .B0_f (new_AGEMA_signal_5418), .B1_t (new_AGEMA_signal_5419), .B1_f (new_AGEMA_signal_5420), .Z0_t (KeyArray_MUX_inS32ser_mux_inst_5_X), .Z0_f (new_AGEMA_signal_5421), .Z1_t (new_AGEMA_signal_5422), .Z1_f (new_AGEMA_signal_5423) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS32ser_mux_inst_5_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS32ser_mux_inst_5_X), .B0_f (new_AGEMA_signal_5421), .B1_t (new_AGEMA_signal_5422), .B1_f (new_AGEMA_signal_5423), .Z0_t (KeyArray_MUX_inS32ser_mux_inst_5_Y), .Z0_f (new_AGEMA_signal_6463), .Z1_t (new_AGEMA_signal_6464), .Z1_f (new_AGEMA_signal_6465) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS32ser_mux_inst_5_XOR2_U1 ( .A0_t (KeyArray_MUX_inS32ser_mux_inst_5_Y), .A0_f (new_AGEMA_signal_6463), .A1_t (new_AGEMA_signal_6464), .A1_f (new_AGEMA_signal_6465), .B0_t (key_s0_t[37]), .B0_f (key_s0_f[37]), .B1_t (key_s1_t[37]), .B1_f (key_s1_f[37]), .Z0_t (KeyArray_inS32ser[5]), .Z0_f (new_AGEMA_signal_7237), .Z1_t (new_AGEMA_signal_7238), .Z1_f (new_AGEMA_signal_7239) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS32ser_mux_inst_6_XOR1_U1 ( .A0_t (key_s0_t[38]), .A0_f (key_s0_f[38]), .A1_t (key_s1_t[38]), .A1_f (key_s1_f[38]), .B0_t (KeyArray_outS33ser[6]), .B0_f (new_AGEMA_signal_5427), .B1_t (new_AGEMA_signal_5428), .B1_f (new_AGEMA_signal_5429), .Z0_t (KeyArray_MUX_inS32ser_mux_inst_6_X), .Z0_f (new_AGEMA_signal_5430), .Z1_t (new_AGEMA_signal_5431), .Z1_f (new_AGEMA_signal_5432) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS32ser_mux_inst_6_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS32ser_mux_inst_6_X), .B0_f (new_AGEMA_signal_5430), .B1_t (new_AGEMA_signal_5431), .B1_f (new_AGEMA_signal_5432), .Z0_t (KeyArray_MUX_inS32ser_mux_inst_6_Y), .Z0_f (new_AGEMA_signal_6466), .Z1_t (new_AGEMA_signal_6467), .Z1_f (new_AGEMA_signal_6468) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS32ser_mux_inst_6_XOR2_U1 ( .A0_t (KeyArray_MUX_inS32ser_mux_inst_6_Y), .A0_f (new_AGEMA_signal_6466), .A1_t (new_AGEMA_signal_6467), .A1_f (new_AGEMA_signal_6468), .B0_t (key_s0_t[38]), .B0_f (key_s0_f[38]), .B1_t (key_s1_t[38]), .B1_f (key_s1_f[38]), .Z0_t (KeyArray_inS32ser[6]), .Z0_f (new_AGEMA_signal_7240), .Z1_t (new_AGEMA_signal_7241), .Z1_f (new_AGEMA_signal_7242) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS32ser_mux_inst_7_XOR1_U1 ( .A0_t (key_s0_t[39]), .A0_f (key_s0_f[39]), .A1_t (key_s1_t[39]), .A1_f (key_s1_f[39]), .B0_t (KeyArray_outS33ser[7]), .B0_f (new_AGEMA_signal_5436), .B1_t (new_AGEMA_signal_5437), .B1_f (new_AGEMA_signal_5438), .Z0_t (KeyArray_MUX_inS32ser_mux_inst_7_X), .Z0_f (new_AGEMA_signal_5439), .Z1_t (new_AGEMA_signal_5440), .Z1_f (new_AGEMA_signal_5441) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS32ser_mux_inst_7_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS32ser_mux_inst_7_X), .B0_f (new_AGEMA_signal_5439), .B1_t (new_AGEMA_signal_5440), .B1_f (new_AGEMA_signal_5441), .Z0_t (KeyArray_MUX_inS32ser_mux_inst_7_Y), .Z0_f (new_AGEMA_signal_6469), .Z1_t (new_AGEMA_signal_6470), .Z1_f (new_AGEMA_signal_6471) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS32ser_mux_inst_7_XOR2_U1 ( .A0_t (KeyArray_MUX_inS32ser_mux_inst_7_Y), .A0_f (new_AGEMA_signal_6469), .A1_t (new_AGEMA_signal_6470), .A1_f (new_AGEMA_signal_6471), .B0_t (key_s0_t[39]), .B0_f (key_s0_f[39]), .B1_t (key_s1_t[39]), .B1_f (key_s1_f[39]), .Z0_t (KeyArray_inS32ser[7]), .Z0_f (new_AGEMA_signal_7243), .Z1_t (new_AGEMA_signal_7244), .Z1_f (new_AGEMA_signal_7245) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_0_XOR1_U1 ( .A0_t (key_s0_t[0]), .A0_f (key_s0_f[0]), .A1_t (key_s1_t[0]), .A1_f (key_s1_f[0]), .B0_t (keyStateIn[0]), .B0_f (new_AGEMA_signal_3432), .B1_t (new_AGEMA_signal_3433), .B1_f (new_AGEMA_signal_3434), .Z0_t (KeyArray_MUX_inS33ser_mux_inst_0_X), .Z0_f (new_AGEMA_signal_5445), .Z1_t (new_AGEMA_signal_5446), .Z1_f (new_AGEMA_signal_5447) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_0_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS33ser_mux_inst_0_X), .B0_f (new_AGEMA_signal_5445), .B1_t (new_AGEMA_signal_5446), .B1_f (new_AGEMA_signal_5447), .Z0_t (KeyArray_MUX_inS33ser_mux_inst_0_Y), .Z0_f (new_AGEMA_signal_6472), .Z1_t (new_AGEMA_signal_6473), .Z1_f (new_AGEMA_signal_6474) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_0_XOR2_U1 ( .A0_t (KeyArray_MUX_inS33ser_mux_inst_0_Y), .A0_f (new_AGEMA_signal_6472), .A1_t (new_AGEMA_signal_6473), .A1_f (new_AGEMA_signal_6474), .B0_t (key_s0_t[0]), .B0_f (key_s0_f[0]), .B1_t (key_s1_t[0]), .B1_f (key_s1_f[0]), .Z0_t (KeyArray_inS33ser[0]), .Z0_f (new_AGEMA_signal_7246), .Z1_t (new_AGEMA_signal_7247), .Z1_f (new_AGEMA_signal_7248) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_1_XOR1_U1 ( .A0_t (key_s0_t[1]), .A0_f (key_s0_f[1]), .A1_t (key_s1_t[1]), .A1_f (key_s1_f[1]), .B0_t (keyStateIn[1]), .B0_f (new_AGEMA_signal_3441), .B1_t (new_AGEMA_signal_3442), .B1_f (new_AGEMA_signal_3443), .Z0_t (KeyArray_MUX_inS33ser_mux_inst_1_X), .Z0_f (new_AGEMA_signal_5451), .Z1_t (new_AGEMA_signal_5452), .Z1_f (new_AGEMA_signal_5453) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS33ser_mux_inst_1_X), .B0_f (new_AGEMA_signal_5451), .B1_t (new_AGEMA_signal_5452), .B1_f (new_AGEMA_signal_5453), .Z0_t (KeyArray_MUX_inS33ser_mux_inst_1_Y), .Z0_f (new_AGEMA_signal_6475), .Z1_t (new_AGEMA_signal_6476), .Z1_f (new_AGEMA_signal_6477) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_1_XOR2_U1 ( .A0_t (KeyArray_MUX_inS33ser_mux_inst_1_Y), .A0_f (new_AGEMA_signal_6475), .A1_t (new_AGEMA_signal_6476), .A1_f (new_AGEMA_signal_6477), .B0_t (key_s0_t[1]), .B0_f (key_s0_f[1]), .B1_t (key_s1_t[1]), .B1_f (key_s1_f[1]), .Z0_t (KeyArray_inS33ser[1]), .Z0_f (new_AGEMA_signal_7249), .Z1_t (new_AGEMA_signal_7250), .Z1_f (new_AGEMA_signal_7251) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_2_XOR1_U1 ( .A0_t (key_s0_t[2]), .A0_f (key_s0_f[2]), .A1_t (key_s1_t[2]), .A1_f (key_s1_f[2]), .B0_t (keyStateIn[2]), .B0_f (new_AGEMA_signal_3450), .B1_t (new_AGEMA_signal_3451), .B1_f (new_AGEMA_signal_3452), .Z0_t (KeyArray_MUX_inS33ser_mux_inst_2_X), .Z0_f (new_AGEMA_signal_5457), .Z1_t (new_AGEMA_signal_5458), .Z1_f (new_AGEMA_signal_5459) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_2_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS33ser_mux_inst_2_X), .B0_f (new_AGEMA_signal_5457), .B1_t (new_AGEMA_signal_5458), .B1_f (new_AGEMA_signal_5459), .Z0_t (KeyArray_MUX_inS33ser_mux_inst_2_Y), .Z0_f (new_AGEMA_signal_6478), .Z1_t (new_AGEMA_signal_6479), .Z1_f (new_AGEMA_signal_6480) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_2_XOR2_U1 ( .A0_t (KeyArray_MUX_inS33ser_mux_inst_2_Y), .A0_f (new_AGEMA_signal_6478), .A1_t (new_AGEMA_signal_6479), .A1_f (new_AGEMA_signal_6480), .B0_t (key_s0_t[2]), .B0_f (key_s0_f[2]), .B1_t (key_s1_t[2]), .B1_f (key_s1_f[2]), .Z0_t (KeyArray_inS33ser[2]), .Z0_f (new_AGEMA_signal_7252), .Z1_t (new_AGEMA_signal_7253), .Z1_f (new_AGEMA_signal_7254) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_3_XOR1_U1 ( .A0_t (key_s0_t[3]), .A0_f (key_s0_f[3]), .A1_t (key_s1_t[3]), .A1_f (key_s1_f[3]), .B0_t (keyStateIn[3]), .B0_f (new_AGEMA_signal_3459), .B1_t (new_AGEMA_signal_3460), .B1_f (new_AGEMA_signal_3461), .Z0_t (KeyArray_MUX_inS33ser_mux_inst_3_X), .Z0_f (new_AGEMA_signal_5463), .Z1_t (new_AGEMA_signal_5464), .Z1_f (new_AGEMA_signal_5465) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_3_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS33ser_mux_inst_3_X), .B0_f (new_AGEMA_signal_5463), .B1_t (new_AGEMA_signal_5464), .B1_f (new_AGEMA_signal_5465), .Z0_t (KeyArray_MUX_inS33ser_mux_inst_3_Y), .Z0_f (new_AGEMA_signal_6481), .Z1_t (new_AGEMA_signal_6482), .Z1_f (new_AGEMA_signal_6483) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_3_XOR2_U1 ( .A0_t (KeyArray_MUX_inS33ser_mux_inst_3_Y), .A0_f (new_AGEMA_signal_6481), .A1_t (new_AGEMA_signal_6482), .A1_f (new_AGEMA_signal_6483), .B0_t (key_s0_t[3]), .B0_f (key_s0_f[3]), .B1_t (key_s1_t[3]), .B1_f (key_s1_f[3]), .Z0_t (KeyArray_inS33ser[3]), .Z0_f (new_AGEMA_signal_7255), .Z1_t (new_AGEMA_signal_7256), .Z1_f (new_AGEMA_signal_7257) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_4_XOR1_U1 ( .A0_t (key_s0_t[4]), .A0_f (key_s0_f[4]), .A1_t (key_s1_t[4]), .A1_f (key_s1_f[4]), .B0_t (keyStateIn[4]), .B0_f (new_AGEMA_signal_3468), .B1_t (new_AGEMA_signal_3469), .B1_f (new_AGEMA_signal_3470), .Z0_t (KeyArray_MUX_inS33ser_mux_inst_4_X), .Z0_f (new_AGEMA_signal_5469), .Z1_t (new_AGEMA_signal_5470), .Z1_f (new_AGEMA_signal_5471) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_4_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS33ser_mux_inst_4_X), .B0_f (new_AGEMA_signal_5469), .B1_t (new_AGEMA_signal_5470), .B1_f (new_AGEMA_signal_5471), .Z0_t (KeyArray_MUX_inS33ser_mux_inst_4_Y), .Z0_f (new_AGEMA_signal_6484), .Z1_t (new_AGEMA_signal_6485), .Z1_f (new_AGEMA_signal_6486) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_4_XOR2_U1 ( .A0_t (KeyArray_MUX_inS33ser_mux_inst_4_Y), .A0_f (new_AGEMA_signal_6484), .A1_t (new_AGEMA_signal_6485), .A1_f (new_AGEMA_signal_6486), .B0_t (key_s0_t[4]), .B0_f (key_s0_f[4]), .B1_t (key_s1_t[4]), .B1_f (key_s1_f[4]), .Z0_t (KeyArray_inS33ser[4]), .Z0_f (new_AGEMA_signal_7258), .Z1_t (new_AGEMA_signal_7259), .Z1_f (new_AGEMA_signal_7260) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_5_XOR1_U1 ( .A0_t (key_s0_t[5]), .A0_f (key_s0_f[5]), .A1_t (key_s1_t[5]), .A1_f (key_s1_f[5]), .B0_t (keyStateIn[5]), .B0_f (new_AGEMA_signal_3477), .B1_t (new_AGEMA_signal_3478), .B1_f (new_AGEMA_signal_3479), .Z0_t (KeyArray_MUX_inS33ser_mux_inst_5_X), .Z0_f (new_AGEMA_signal_5475), .Z1_t (new_AGEMA_signal_5476), .Z1_f (new_AGEMA_signal_5477) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_5_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS33ser_mux_inst_5_X), .B0_f (new_AGEMA_signal_5475), .B1_t (new_AGEMA_signal_5476), .B1_f (new_AGEMA_signal_5477), .Z0_t (KeyArray_MUX_inS33ser_mux_inst_5_Y), .Z0_f (new_AGEMA_signal_6487), .Z1_t (new_AGEMA_signal_6488), .Z1_f (new_AGEMA_signal_6489) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_5_XOR2_U1 ( .A0_t (KeyArray_MUX_inS33ser_mux_inst_5_Y), .A0_f (new_AGEMA_signal_6487), .A1_t (new_AGEMA_signal_6488), .A1_f (new_AGEMA_signal_6489), .B0_t (key_s0_t[5]), .B0_f (key_s0_f[5]), .B1_t (key_s1_t[5]), .B1_f (key_s1_f[5]), .Z0_t (KeyArray_inS33ser[5]), .Z0_f (new_AGEMA_signal_7261), .Z1_t (new_AGEMA_signal_7262), .Z1_f (new_AGEMA_signal_7263) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_6_XOR1_U1 ( .A0_t (key_s0_t[6]), .A0_f (key_s0_f[6]), .A1_t (key_s1_t[6]), .A1_f (key_s1_f[6]), .B0_t (keyStateIn[6]), .B0_f (new_AGEMA_signal_3486), .B1_t (new_AGEMA_signal_3487), .B1_f (new_AGEMA_signal_3488), .Z0_t (KeyArray_MUX_inS33ser_mux_inst_6_X), .Z0_f (new_AGEMA_signal_5481), .Z1_t (new_AGEMA_signal_5482), .Z1_f (new_AGEMA_signal_5483) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_6_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS33ser_mux_inst_6_X), .B0_f (new_AGEMA_signal_5481), .B1_t (new_AGEMA_signal_5482), .B1_f (new_AGEMA_signal_5483), .Z0_t (KeyArray_MUX_inS33ser_mux_inst_6_Y), .Z0_f (new_AGEMA_signal_6490), .Z1_t (new_AGEMA_signal_6491), .Z1_f (new_AGEMA_signal_6492) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_6_XOR2_U1 ( .A0_t (KeyArray_MUX_inS33ser_mux_inst_6_Y), .A0_f (new_AGEMA_signal_6490), .A1_t (new_AGEMA_signal_6491), .A1_f (new_AGEMA_signal_6492), .B0_t (key_s0_t[6]), .B0_f (key_s0_f[6]), .B1_t (key_s1_t[6]), .B1_f (key_s1_f[6]), .Z0_t (KeyArray_inS33ser[6]), .Z0_f (new_AGEMA_signal_7264), .Z1_t (new_AGEMA_signal_7265), .Z1_f (new_AGEMA_signal_7266) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_7_XOR1_U1 ( .A0_t (key_s0_t[7]), .A0_f (key_s0_f[7]), .A1_t (key_s1_t[7]), .A1_f (key_s1_f[7]), .B0_t (keyStateIn[7]), .B0_f (new_AGEMA_signal_3495), .B1_t (new_AGEMA_signal_3496), .B1_f (new_AGEMA_signal_3497), .Z0_t (KeyArray_MUX_inS33ser_mux_inst_7_X), .Z0_f (new_AGEMA_signal_5487), .Z1_t (new_AGEMA_signal_5488), .Z1_f (new_AGEMA_signal_5489) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_7_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (nReset), .A1_f (new_AGEMA_signal_3502), .B0_t (KeyArray_MUX_inS33ser_mux_inst_7_X), .B0_f (new_AGEMA_signal_5487), .B1_t (new_AGEMA_signal_5488), .B1_f (new_AGEMA_signal_5489), .Z0_t (KeyArray_MUX_inS33ser_mux_inst_7_Y), .Z0_f (new_AGEMA_signal_6493), .Z1_t (new_AGEMA_signal_6494), .Z1_f (new_AGEMA_signal_6495) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_7_XOR2_U1 ( .A0_t (KeyArray_MUX_inS33ser_mux_inst_7_Y), .A0_f (new_AGEMA_signal_6493), .A1_t (new_AGEMA_signal_6494), .A1_f (new_AGEMA_signal_6495), .B0_t (key_s0_t[7]), .B0_f (key_s0_f[7]), .B1_t (key_s1_t[7]), .B1_f (key_s1_f[7]), .Z0_t (KeyArray_inS33ser[7]), .Z0_f (new_AGEMA_signal_7267), .Z1_t (new_AGEMA_signal_7268), .Z1_f (new_AGEMA_signal_7269) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line0_U24 ( .A0_t (MixColumns_line0_n16), .A0_f (new_AGEMA_signal_6496), .A1_t (new_AGEMA_signal_6497), .A1_f (new_AGEMA_signal_6498), .B0_t (MixColumns_line0_n15), .B0_f (new_AGEMA_signal_5496), .B1_t (new_AGEMA_signal_5497), .B1_f (new_AGEMA_signal_5498), .Z0_t (MCout[31]), .Z0_f (new_AGEMA_signal_7270), .Z1_t (new_AGEMA_signal_7271), .Z1_f (new_AGEMA_signal_7272) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line0_U23 ( .A0_t (ciphertext_s0_t[111]), .A0_f (ciphertext_s0_f[111]), .A1_t (ciphertext_s1_t[111]), .A1_f (ciphertext_s1_f[111]), .B0_t (ciphertext_s0_t[103]), .B0_f (ciphertext_s0_f[103]), .B1_t (ciphertext_s1_t[103]), .B1_f (ciphertext_s1_f[103]), .Z0_t (MixColumns_line0_n15), .Z0_f (new_AGEMA_signal_5496), .Z1_t (new_AGEMA_signal_5497), .Z1_f (new_AGEMA_signal_5498) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_U22 ( .A0_t (ciphertext_s0_t[126]), .A0_f (ciphertext_s0_f[126]), .A1_t (ciphertext_s1_t[126]), .A1_f (ciphertext_s1_f[126]), .B0_t (MixColumns_line0_S13[7]), .B0_f (new_AGEMA_signal_5577), .B1_t (new_AGEMA_signal_5578), .B1_f (new_AGEMA_signal_5579), .Z0_t (MixColumns_line0_n16), .Z0_f (new_AGEMA_signal_6496), .Z1_t (new_AGEMA_signal_6497), .Z1_f (new_AGEMA_signal_6498) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line0_U21 ( .A0_t (MixColumns_line0_n14), .A0_f (new_AGEMA_signal_6499), .A1_t (new_AGEMA_signal_6500), .A1_f (new_AGEMA_signal_6501), .B0_t (MixColumns_line0_n13), .B0_f (new_AGEMA_signal_5505), .B1_t (new_AGEMA_signal_5506), .B1_f (new_AGEMA_signal_5507), .Z0_t (MCout[30]), .Z0_f (new_AGEMA_signal_7273), .Z1_t (new_AGEMA_signal_7274), .Z1_f (new_AGEMA_signal_7275) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line0_U20 ( .A0_t (ciphertext_s0_t[110]), .A0_f (ciphertext_s0_f[110]), .A1_t (ciphertext_s1_t[110]), .A1_f (ciphertext_s1_f[110]), .B0_t (ciphertext_s0_t[102]), .B0_f (ciphertext_s0_f[102]), .B1_t (ciphertext_s1_t[102]), .B1_f (ciphertext_s1_f[102]), .Z0_t (MixColumns_line0_n13), .Z0_f (new_AGEMA_signal_5505), .Z1_t (new_AGEMA_signal_5506), .Z1_f (new_AGEMA_signal_5507) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_U19 ( .A0_t (ciphertext_s0_t[125]), .A0_f (ciphertext_s0_f[125]), .A1_t (ciphertext_s1_t[125]), .A1_f (ciphertext_s1_f[125]), .B0_t (MixColumns_line0_S13[6]), .B0_f (new_AGEMA_signal_5583), .B1_t (new_AGEMA_signal_5584), .B1_f (new_AGEMA_signal_5585), .Z0_t (MixColumns_line0_n14), .Z0_f (new_AGEMA_signal_6499), .Z1_t (new_AGEMA_signal_6500), .Z1_f (new_AGEMA_signal_6501) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line0_U18 ( .A0_t (MixColumns_line0_n12), .A0_f (new_AGEMA_signal_6502), .A1_t (new_AGEMA_signal_6503), .A1_f (new_AGEMA_signal_6504), .B0_t (MixColumns_line0_n11), .B0_f (new_AGEMA_signal_5514), .B1_t (new_AGEMA_signal_5515), .B1_f (new_AGEMA_signal_5516), .Z0_t (MCout[29]), .Z0_f (new_AGEMA_signal_7276), .Z1_t (new_AGEMA_signal_7277), .Z1_f (new_AGEMA_signal_7278) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line0_U17 ( .A0_t (ciphertext_s0_t[109]), .A0_f (ciphertext_s0_f[109]), .A1_t (ciphertext_s1_t[109]), .A1_f (ciphertext_s1_f[109]), .B0_t (ciphertext_s0_t[101]), .B0_f (ciphertext_s0_f[101]), .B1_t (ciphertext_s1_t[101]), .B1_f (ciphertext_s1_f[101]), .Z0_t (MixColumns_line0_n11), .Z0_f (new_AGEMA_signal_5514), .Z1_t (new_AGEMA_signal_5515), .Z1_f (new_AGEMA_signal_5516) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_U16 ( .A0_t (ciphertext_s0_t[124]), .A0_f (ciphertext_s0_f[124]), .A1_t (ciphertext_s1_t[124]), .A1_f (ciphertext_s1_f[124]), .B0_t (MixColumns_line0_S13[5]), .B0_f (new_AGEMA_signal_5589), .B1_t (new_AGEMA_signal_5590), .B1_f (new_AGEMA_signal_5591), .Z0_t (MixColumns_line0_n12), .Z0_f (new_AGEMA_signal_6502), .Z1_t (new_AGEMA_signal_6503), .Z1_f (new_AGEMA_signal_6504) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line0_U15 ( .A0_t (MixColumns_line0_n10), .A0_f (new_AGEMA_signal_7279), .A1_t (new_AGEMA_signal_7280), .A1_f (new_AGEMA_signal_7281), .B0_t (MixColumns_line0_n9), .B0_f (new_AGEMA_signal_5523), .B1_t (new_AGEMA_signal_5524), .B1_f (new_AGEMA_signal_5525), .Z0_t (MCout[28]), .Z0_f (new_AGEMA_signal_8079), .Z1_t (new_AGEMA_signal_8080), .Z1_f (new_AGEMA_signal_8081) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line0_U14 ( .A0_t (ciphertext_s0_t[108]), .A0_f (ciphertext_s0_f[108]), .A1_t (ciphertext_s1_t[108]), .A1_f (ciphertext_s1_f[108]), .B0_t (ciphertext_s0_t[100]), .B0_f (ciphertext_s0_f[100]), .B1_t (ciphertext_s1_t[100]), .B1_f (ciphertext_s1_f[100]), .Z0_t (MixColumns_line0_n9), .Z0_f (new_AGEMA_signal_5523), .Z1_t (new_AGEMA_signal_5524), .Z1_f (new_AGEMA_signal_5525) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_U13 ( .A0_t (MixColumns_line0_S02[4]), .A0_f (new_AGEMA_signal_5562), .A1_t (new_AGEMA_signal_5563), .A1_f (new_AGEMA_signal_5564), .B0_t (MixColumns_line0_S13[4]), .B0_f (new_AGEMA_signal_6511), .B1_t (new_AGEMA_signal_6512), .B1_f (new_AGEMA_signal_6513), .Z0_t (MixColumns_line0_n10), .Z0_f (new_AGEMA_signal_7279), .Z1_t (new_AGEMA_signal_7280), .Z1_f (new_AGEMA_signal_7281) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line0_U12 ( .A0_t (MixColumns_line0_n8), .A0_f (new_AGEMA_signal_7282), .A1_t (new_AGEMA_signal_7283), .A1_f (new_AGEMA_signal_7284), .B0_t (MixColumns_line0_n7), .B0_f (new_AGEMA_signal_5532), .B1_t (new_AGEMA_signal_5533), .B1_f (new_AGEMA_signal_5534), .Z0_t (MCout[27]), .Z0_f (new_AGEMA_signal_8082), .Z1_t (new_AGEMA_signal_8083), .Z1_f (new_AGEMA_signal_8084) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line0_U11 ( .A0_t (ciphertext_s0_t[107]), .A0_f (ciphertext_s0_f[107]), .A1_t (ciphertext_s1_t[107]), .A1_f (ciphertext_s1_f[107]), .B0_t (ciphertext_s0_t[99]), .B0_f (ciphertext_s0_f[99]), .B1_t (ciphertext_s1_t[99]), .B1_f (ciphertext_s1_f[99]), .Z0_t (MixColumns_line0_n7), .Z0_f (new_AGEMA_signal_5532), .Z1_t (new_AGEMA_signal_5533), .Z1_f (new_AGEMA_signal_5534) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_U10 ( .A0_t (MixColumns_line0_S02[3]), .A0_f (new_AGEMA_signal_5565), .A1_t (new_AGEMA_signal_5566), .A1_f (new_AGEMA_signal_5567), .B0_t (MixColumns_line0_S13[3]), .B0_f (new_AGEMA_signal_6514), .B1_t (new_AGEMA_signal_6515), .B1_f (new_AGEMA_signal_6516), .Z0_t (MixColumns_line0_n8), .Z0_f (new_AGEMA_signal_7282), .Z1_t (new_AGEMA_signal_7283), .Z1_f (new_AGEMA_signal_7284) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line0_U9 ( .A0_t (MixColumns_line0_n6), .A0_f (new_AGEMA_signal_6505), .A1_t (new_AGEMA_signal_6506), .A1_f (new_AGEMA_signal_6507), .B0_t (MixColumns_line0_n5), .B0_f (new_AGEMA_signal_5541), .B1_t (new_AGEMA_signal_5542), .B1_f (new_AGEMA_signal_5543), .Z0_t (MCout[26]), .Z0_f (new_AGEMA_signal_7285), .Z1_t (new_AGEMA_signal_7286), .Z1_f (new_AGEMA_signal_7287) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line0_U8 ( .A0_t (ciphertext_s0_t[106]), .A0_f (ciphertext_s0_f[106]), .A1_t (ciphertext_s1_t[106]), .A1_f (ciphertext_s1_f[106]), .B0_t (ciphertext_s0_t[98]), .B0_f (ciphertext_s0_f[98]), .B1_t (ciphertext_s1_t[98]), .B1_f (ciphertext_s1_f[98]), .Z0_t (MixColumns_line0_n5), .Z0_f (new_AGEMA_signal_5541), .Z1_t (new_AGEMA_signal_5542), .Z1_f (new_AGEMA_signal_5543) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_U7 ( .A0_t (ciphertext_s0_t[121]), .A0_f (ciphertext_s0_f[121]), .A1_t (ciphertext_s1_t[121]), .A1_f (ciphertext_s1_f[121]), .B0_t (MixColumns_line0_S13[2]), .B0_f (new_AGEMA_signal_5598), .B1_t (new_AGEMA_signal_5599), .B1_f (new_AGEMA_signal_5600), .Z0_t (MixColumns_line0_n6), .Z0_f (new_AGEMA_signal_6505), .Z1_t (new_AGEMA_signal_6506), .Z1_f (new_AGEMA_signal_6507) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line0_U6 ( .A0_t (MixColumns_line0_n4), .A0_f (new_AGEMA_signal_7288), .A1_t (new_AGEMA_signal_7289), .A1_f (new_AGEMA_signal_7290), .B0_t (MixColumns_line0_n3), .B0_f (new_AGEMA_signal_5550), .B1_t (new_AGEMA_signal_5551), .B1_f (new_AGEMA_signal_5552), .Z0_t (MCout[25]), .Z0_f (new_AGEMA_signal_8085), .Z1_t (new_AGEMA_signal_8086), .Z1_f (new_AGEMA_signal_8087) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line0_U5 ( .A0_t (ciphertext_s0_t[97]), .A0_f (ciphertext_s0_f[97]), .A1_t (ciphertext_s1_t[97]), .A1_f (ciphertext_s1_f[97]), .B0_t (ciphertext_s0_t[105]), .B0_f (ciphertext_s0_f[105]), .B1_t (ciphertext_s1_t[105]), .B1_f (ciphertext_s1_f[105]), .Z0_t (MixColumns_line0_n3), .Z0_f (new_AGEMA_signal_5550), .Z1_t (new_AGEMA_signal_5551), .Z1_f (new_AGEMA_signal_5552) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_U4 ( .A0_t (MixColumns_line0_S02[1]), .A0_f (new_AGEMA_signal_5568), .A1_t (new_AGEMA_signal_5569), .A1_f (new_AGEMA_signal_5570), .B0_t (MixColumns_line0_S13[1]), .B0_f (new_AGEMA_signal_6517), .B1_t (new_AGEMA_signal_6518), .B1_f (new_AGEMA_signal_6519), .Z0_t (MixColumns_line0_n4), .Z0_f (new_AGEMA_signal_7288), .Z1_t (new_AGEMA_signal_7289), .Z1_f (new_AGEMA_signal_7290) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line0_U3 ( .A0_t (MixColumns_line0_n2), .A0_f (new_AGEMA_signal_6508), .A1_t (new_AGEMA_signal_6509), .A1_f (new_AGEMA_signal_6510), .B0_t (MixColumns_line0_n1), .B0_f (new_AGEMA_signal_5559), .B1_t (new_AGEMA_signal_5560), .B1_f (new_AGEMA_signal_5561), .Z0_t (MCout[24]), .Z0_f (new_AGEMA_signal_7291), .Z1_t (new_AGEMA_signal_7292), .Z1_f (new_AGEMA_signal_7293) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line0_U2 ( .A0_t (ciphertext_s0_t[96]), .A0_f (ciphertext_s0_f[96]), .A1_t (ciphertext_s1_t[96]), .A1_f (ciphertext_s1_f[96]), .B0_t (ciphertext_s0_t[104]), .B0_f (ciphertext_s0_f[104]), .B1_t (ciphertext_s1_t[104]), .B1_f (ciphertext_s1_f[104]), .Z0_t (MixColumns_line0_n1), .Z0_f (new_AGEMA_signal_5559), .Z1_t (new_AGEMA_signal_5560), .Z1_f (new_AGEMA_signal_5561) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_U1 ( .A0_t (ciphertext_s0_t[127]), .A0_f (ciphertext_s0_f[127]), .A1_t (ciphertext_s1_t[127]), .A1_f (ciphertext_s1_f[127]), .B0_t (MixColumns_line0_S13[0]), .B0_f (new_AGEMA_signal_5604), .B1_t (new_AGEMA_signal_5605), .B1_f (new_AGEMA_signal_5606), .Z0_t (MixColumns_line0_n2), .Z0_f (new_AGEMA_signal_6508), .Z1_t (new_AGEMA_signal_6509), .Z1_f (new_AGEMA_signal_6510) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_timesTWO_U3 ( .A0_t (ciphertext_s0_t[127]), .A0_f (ciphertext_s0_f[127]), .A1_t (ciphertext_s1_t[127]), .A1_f (ciphertext_s1_f[127]), .B0_t (ciphertext_s0_t[123]), .B0_f (ciphertext_s0_f[123]), .B1_t (ciphertext_s1_t[123]), .B1_f (ciphertext_s1_f[123]), .Z0_t (MixColumns_line0_S02[4]), .Z0_f (new_AGEMA_signal_5562), .Z1_t (new_AGEMA_signal_5563), .Z1_f (new_AGEMA_signal_5564) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_timesTWO_U2 ( .A0_t (ciphertext_s0_t[127]), .A0_f (ciphertext_s0_f[127]), .A1_t (ciphertext_s1_t[127]), .A1_f (ciphertext_s1_f[127]), .B0_t (ciphertext_s0_t[122]), .B0_f (ciphertext_s0_f[122]), .B1_t (ciphertext_s1_t[122]), .B1_f (ciphertext_s1_f[122]), .Z0_t (MixColumns_line0_S02[3]), .Z0_f (new_AGEMA_signal_5565), .Z1_t (new_AGEMA_signal_5566), .Z1_f (new_AGEMA_signal_5567) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_timesTWO_U1 ( .A0_t (ciphertext_s0_t[127]), .A0_f (ciphertext_s0_f[127]), .A1_t (ciphertext_s1_t[127]), .A1_f (ciphertext_s1_f[127]), .B0_t (ciphertext_s0_t[120]), .B0_f (ciphertext_s0_f[120]), .B1_t (ciphertext_s1_t[120]), .B1_f (ciphertext_s1_f[120]), .Z0_t (MixColumns_line0_S02[1]), .Z0_f (new_AGEMA_signal_5568), .Z1_t (new_AGEMA_signal_5569), .Z1_f (new_AGEMA_signal_5570) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_timesTHREE_U8 ( .A0_t (ciphertext_s0_t[119]), .A0_f (ciphertext_s0_f[119]), .A1_t (ciphertext_s1_t[119]), .A1_f (ciphertext_s1_f[119]), .B0_t (ciphertext_s0_t[118]), .B0_f (ciphertext_s0_f[118]), .B1_t (ciphertext_s1_t[118]), .B1_f (ciphertext_s1_f[118]), .Z0_t (MixColumns_line0_S13[7]), .Z0_f (new_AGEMA_signal_5577), .Z1_t (new_AGEMA_signal_5578), .Z1_f (new_AGEMA_signal_5579) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_timesTHREE_U7 ( .A0_t (ciphertext_s0_t[118]), .A0_f (ciphertext_s0_f[118]), .A1_t (ciphertext_s1_t[118]), .A1_f (ciphertext_s1_f[118]), .B0_t (ciphertext_s0_t[117]), .B0_f (ciphertext_s0_f[117]), .B1_t (ciphertext_s1_t[117]), .B1_f (ciphertext_s1_f[117]), .Z0_t (MixColumns_line0_S13[6]), .Z0_f (new_AGEMA_signal_5583), .Z1_t (new_AGEMA_signal_5584), .Z1_f (new_AGEMA_signal_5585) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_timesTHREE_U6 ( .A0_t (ciphertext_s0_t[117]), .A0_f (ciphertext_s0_f[117]), .A1_t (ciphertext_s1_t[117]), .A1_f (ciphertext_s1_f[117]), .B0_t (ciphertext_s0_t[116]), .B0_f (ciphertext_s0_f[116]), .B1_t (ciphertext_s1_t[116]), .B1_f (ciphertext_s1_f[116]), .Z0_t (MixColumns_line0_S13[5]), .Z0_f (new_AGEMA_signal_5589), .Z1_t (new_AGEMA_signal_5590), .Z1_f (new_AGEMA_signal_5591) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_timesTHREE_U5 ( .A0_t (ciphertext_s0_t[116]), .A0_f (ciphertext_s0_f[116]), .A1_t (ciphertext_s1_t[116]), .A1_f (ciphertext_s1_f[116]), .B0_t (MixColumns_line0_timesTHREE_input2[4]), .B0_f (new_AGEMA_signal_5610), .B1_t (new_AGEMA_signal_5611), .B1_f (new_AGEMA_signal_5612), .Z0_t (MixColumns_line0_S13[4]), .Z0_f (new_AGEMA_signal_6511), .Z1_t (new_AGEMA_signal_6512), .Z1_f (new_AGEMA_signal_6513) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_timesTHREE_U4 ( .A0_t (ciphertext_s0_t[115]), .A0_f (ciphertext_s0_f[115]), .A1_t (ciphertext_s1_t[115]), .A1_f (ciphertext_s1_f[115]), .B0_t (MixColumns_line0_timesTHREE_input2[3]), .B0_f (new_AGEMA_signal_5613), .B1_t (new_AGEMA_signal_5614), .B1_f (new_AGEMA_signal_5615), .Z0_t (MixColumns_line0_S13[3]), .Z0_f (new_AGEMA_signal_6514), .Z1_t (new_AGEMA_signal_6515), .Z1_f (new_AGEMA_signal_6516) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_timesTHREE_U3 ( .A0_t (ciphertext_s0_t[114]), .A0_f (ciphertext_s0_f[114]), .A1_t (ciphertext_s1_t[114]), .A1_f (ciphertext_s1_f[114]), .B0_t (ciphertext_s0_t[113]), .B0_f (ciphertext_s0_f[113]), .B1_t (ciphertext_s1_t[113]), .B1_f (ciphertext_s1_f[113]), .Z0_t (MixColumns_line0_S13[2]), .Z0_f (new_AGEMA_signal_5598), .Z1_t (new_AGEMA_signal_5599), .Z1_f (new_AGEMA_signal_5600) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_timesTHREE_U2 ( .A0_t (ciphertext_s0_t[113]), .A0_f (ciphertext_s0_f[113]), .A1_t (ciphertext_s1_t[113]), .A1_f (ciphertext_s1_f[113]), .B0_t (MixColumns_line0_timesTHREE_input2[1]), .B0_f (new_AGEMA_signal_5616), .B1_t (new_AGEMA_signal_5617), .B1_f (new_AGEMA_signal_5618), .Z0_t (MixColumns_line0_S13[1]), .Z0_f (new_AGEMA_signal_6517), .Z1_t (new_AGEMA_signal_6518), .Z1_f (new_AGEMA_signal_6519) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_timesTHREE_U1 ( .A0_t (ciphertext_s0_t[112]), .A0_f (ciphertext_s0_f[112]), .A1_t (ciphertext_s1_t[112]), .A1_f (ciphertext_s1_f[112]), .B0_t (ciphertext_s0_t[119]), .B0_f (ciphertext_s0_f[119]), .B1_t (ciphertext_s1_t[119]), .B1_f (ciphertext_s1_f[119]), .Z0_t (MixColumns_line0_S13[0]), .Z0_f (new_AGEMA_signal_5604), .Z1_t (new_AGEMA_signal_5605), .Z1_f (new_AGEMA_signal_5606) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_timesTHREE_timesTWO_U3 ( .A0_t (ciphertext_s0_t[119]), .A0_f (ciphertext_s0_f[119]), .A1_t (ciphertext_s1_t[119]), .A1_f (ciphertext_s1_f[119]), .B0_t (ciphertext_s0_t[115]), .B0_f (ciphertext_s0_f[115]), .B1_t (ciphertext_s1_t[115]), .B1_f (ciphertext_s1_f[115]), .Z0_t (MixColumns_line0_timesTHREE_input2[4]), .Z0_f (new_AGEMA_signal_5610), .Z1_t (new_AGEMA_signal_5611), .Z1_f (new_AGEMA_signal_5612) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_timesTHREE_timesTWO_U2 ( .A0_t (ciphertext_s0_t[119]), .A0_f (ciphertext_s0_f[119]), .A1_t (ciphertext_s1_t[119]), .A1_f (ciphertext_s1_f[119]), .B0_t (ciphertext_s0_t[114]), .B0_f (ciphertext_s0_f[114]), .B1_t (ciphertext_s1_t[114]), .B1_f (ciphertext_s1_f[114]), .Z0_t (MixColumns_line0_timesTHREE_input2[3]), .Z0_f (new_AGEMA_signal_5613), .Z1_t (new_AGEMA_signal_5614), .Z1_f (new_AGEMA_signal_5615) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_timesTHREE_timesTWO_U1 ( .A0_t (ciphertext_s0_t[119]), .A0_f (ciphertext_s0_f[119]), .A1_t (ciphertext_s1_t[119]), .A1_f (ciphertext_s1_f[119]), .B0_t (ciphertext_s0_t[112]), .B0_f (ciphertext_s0_f[112]), .B1_t (ciphertext_s1_t[112]), .B1_f (ciphertext_s1_f[112]), .Z0_t (MixColumns_line0_timesTHREE_input2[1]), .Z0_f (new_AGEMA_signal_5616), .Z1_t (new_AGEMA_signal_5617), .Z1_f (new_AGEMA_signal_5618) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line1_U24 ( .A0_t (MixColumns_line1_n16), .A0_f (new_AGEMA_signal_6520), .A1_t (new_AGEMA_signal_6521), .A1_f (new_AGEMA_signal_6522), .B0_t (MixColumns_line1_n15), .B0_f (new_AGEMA_signal_5619), .B1_t (new_AGEMA_signal_5620), .B1_f (new_AGEMA_signal_5621), .Z0_t (MCout[23]), .Z0_f (new_AGEMA_signal_7294), .Z1_t (new_AGEMA_signal_7295), .Z1_f (new_AGEMA_signal_7296) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line1_U23 ( .A0_t (ciphertext_s0_t[103]), .A0_f (ciphertext_s0_f[103]), .A1_t (ciphertext_s1_t[103]), .A1_f (ciphertext_s1_f[103]), .B0_t (ciphertext_s0_t[127]), .B0_f (ciphertext_s0_f[127]), .B1_t (ciphertext_s1_t[127]), .B1_f (ciphertext_s1_f[127]), .Z0_t (MixColumns_line1_n15), .Z0_f (new_AGEMA_signal_5619), .Z1_t (new_AGEMA_signal_5620), .Z1_f (new_AGEMA_signal_5621) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_U22 ( .A0_t (ciphertext_s0_t[118]), .A0_f (ciphertext_s0_f[118]), .A1_t (ciphertext_s1_t[118]), .A1_f (ciphertext_s1_f[118]), .B0_t (MixColumns_line1_S13[7]), .B0_f (new_AGEMA_signal_5652), .B1_t (new_AGEMA_signal_5653), .B1_f (new_AGEMA_signal_5654), .Z0_t (MixColumns_line1_n16), .Z0_f (new_AGEMA_signal_6520), .Z1_t (new_AGEMA_signal_6521), .Z1_f (new_AGEMA_signal_6522) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line1_U21 ( .A0_t (MixColumns_line1_n14), .A0_f (new_AGEMA_signal_6523), .A1_t (new_AGEMA_signal_6524), .A1_f (new_AGEMA_signal_6525), .B0_t (MixColumns_line1_n13), .B0_f (new_AGEMA_signal_5622), .B1_t (new_AGEMA_signal_5623), .B1_f (new_AGEMA_signal_5624), .Z0_t (MCout[22]), .Z0_f (new_AGEMA_signal_7297), .Z1_t (new_AGEMA_signal_7298), .Z1_f (new_AGEMA_signal_7299) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line1_U20 ( .A0_t (ciphertext_s0_t[102]), .A0_f (ciphertext_s0_f[102]), .A1_t (ciphertext_s1_t[102]), .A1_f (ciphertext_s1_f[102]), .B0_t (ciphertext_s0_t[126]), .B0_f (ciphertext_s0_f[126]), .B1_t (ciphertext_s1_t[126]), .B1_f (ciphertext_s1_f[126]), .Z0_t (MixColumns_line1_n13), .Z0_f (new_AGEMA_signal_5622), .Z1_t (new_AGEMA_signal_5623), .Z1_f (new_AGEMA_signal_5624) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_U19 ( .A0_t (ciphertext_s0_t[117]), .A0_f (ciphertext_s0_f[117]), .A1_t (ciphertext_s1_t[117]), .A1_f (ciphertext_s1_f[117]), .B0_t (MixColumns_line1_S13[6]), .B0_f (new_AGEMA_signal_5655), .B1_t (new_AGEMA_signal_5656), .B1_f (new_AGEMA_signal_5657), .Z0_t (MixColumns_line1_n14), .Z0_f (new_AGEMA_signal_6523), .Z1_t (new_AGEMA_signal_6524), .Z1_f (new_AGEMA_signal_6525) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line1_U18 ( .A0_t (MixColumns_line1_n12), .A0_f (new_AGEMA_signal_6526), .A1_t (new_AGEMA_signal_6527), .A1_f (new_AGEMA_signal_6528), .B0_t (MixColumns_line1_n11), .B0_f (new_AGEMA_signal_5625), .B1_t (new_AGEMA_signal_5626), .B1_f (new_AGEMA_signal_5627), .Z0_t (MCout[21]), .Z0_f (new_AGEMA_signal_7300), .Z1_t (new_AGEMA_signal_7301), .Z1_f (new_AGEMA_signal_7302) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line1_U17 ( .A0_t (ciphertext_s0_t[101]), .A0_f (ciphertext_s0_f[101]), .A1_t (ciphertext_s1_t[101]), .A1_f (ciphertext_s1_f[101]), .B0_t (ciphertext_s0_t[125]), .B0_f (ciphertext_s0_f[125]), .B1_t (ciphertext_s1_t[125]), .B1_f (ciphertext_s1_f[125]), .Z0_t (MixColumns_line1_n11), .Z0_f (new_AGEMA_signal_5625), .Z1_t (new_AGEMA_signal_5626), .Z1_f (new_AGEMA_signal_5627) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_U16 ( .A0_t (ciphertext_s0_t[116]), .A0_f (ciphertext_s0_f[116]), .A1_t (ciphertext_s1_t[116]), .A1_f (ciphertext_s1_f[116]), .B0_t (MixColumns_line1_S13[5]), .B0_f (new_AGEMA_signal_5658), .B1_t (new_AGEMA_signal_5659), .B1_f (new_AGEMA_signal_5660), .Z0_t (MixColumns_line1_n12), .Z0_f (new_AGEMA_signal_6526), .Z1_t (new_AGEMA_signal_6527), .Z1_f (new_AGEMA_signal_6528) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line1_U15 ( .A0_t (MixColumns_line1_n10), .A0_f (new_AGEMA_signal_7303), .A1_t (new_AGEMA_signal_7304), .A1_f (new_AGEMA_signal_7305), .B0_t (MixColumns_line1_n9), .B0_f (new_AGEMA_signal_5628), .B1_t (new_AGEMA_signal_5629), .B1_f (new_AGEMA_signal_5630), .Z0_t (MCout[20]), .Z0_f (new_AGEMA_signal_8088), .Z1_t (new_AGEMA_signal_8089), .Z1_f (new_AGEMA_signal_8090) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line1_U14 ( .A0_t (ciphertext_s0_t[100]), .A0_f (ciphertext_s0_f[100]), .A1_t (ciphertext_s1_t[100]), .A1_f (ciphertext_s1_f[100]), .B0_t (ciphertext_s0_t[124]), .B0_f (ciphertext_s0_f[124]), .B1_t (ciphertext_s1_t[124]), .B1_f (ciphertext_s1_f[124]), .Z0_t (MixColumns_line1_n9), .Z0_f (new_AGEMA_signal_5628), .Z1_t (new_AGEMA_signal_5629), .Z1_f (new_AGEMA_signal_5630) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_U13 ( .A0_t (MixColumns_line1_S02_4_), .A0_f (new_AGEMA_signal_5643), .A1_t (new_AGEMA_signal_5644), .A1_f (new_AGEMA_signal_5645), .B0_t (MixColumns_line1_S13[4]), .B0_f (new_AGEMA_signal_6535), .B1_t (new_AGEMA_signal_6536), .B1_f (new_AGEMA_signal_6537), .Z0_t (MixColumns_line1_n10), .Z0_f (new_AGEMA_signal_7303), .Z1_t (new_AGEMA_signal_7304), .Z1_f (new_AGEMA_signal_7305) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line1_U12 ( .A0_t (MixColumns_line1_n8), .A0_f (new_AGEMA_signal_7306), .A1_t (new_AGEMA_signal_7307), .A1_f (new_AGEMA_signal_7308), .B0_t (MixColumns_line1_n7), .B0_f (new_AGEMA_signal_5631), .B1_t (new_AGEMA_signal_5632), .B1_f (new_AGEMA_signal_5633), .Z0_t (MCout[19]), .Z0_f (new_AGEMA_signal_8091), .Z1_t (new_AGEMA_signal_8092), .Z1_f (new_AGEMA_signal_8093) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line1_U11 ( .A0_t (ciphertext_s0_t[99]), .A0_f (ciphertext_s0_f[99]), .A1_t (ciphertext_s1_t[99]), .A1_f (ciphertext_s1_f[99]), .B0_t (ciphertext_s0_t[123]), .B0_f (ciphertext_s0_f[123]), .B1_t (ciphertext_s1_t[123]), .B1_f (ciphertext_s1_f[123]), .Z0_t (MixColumns_line1_n7), .Z0_f (new_AGEMA_signal_5631), .Z1_t (new_AGEMA_signal_5632), .Z1_f (new_AGEMA_signal_5633) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_U10 ( .A0_t (MixColumns_line1_S02_3_), .A0_f (new_AGEMA_signal_5646), .A1_t (new_AGEMA_signal_5647), .A1_f (new_AGEMA_signal_5648), .B0_t (MixColumns_line1_S13[3]), .B0_f (new_AGEMA_signal_6538), .B1_t (new_AGEMA_signal_6539), .B1_f (new_AGEMA_signal_6540), .Z0_t (MixColumns_line1_n8), .Z0_f (new_AGEMA_signal_7306), .Z1_t (new_AGEMA_signal_7307), .Z1_f (new_AGEMA_signal_7308) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line1_U9 ( .A0_t (MixColumns_line1_n6), .A0_f (new_AGEMA_signal_6529), .A1_t (new_AGEMA_signal_6530), .A1_f (new_AGEMA_signal_6531), .B0_t (MixColumns_line1_n5), .B0_f (new_AGEMA_signal_5634), .B1_t (new_AGEMA_signal_5635), .B1_f (new_AGEMA_signal_5636), .Z0_t (MCout[18]), .Z0_f (new_AGEMA_signal_7309), .Z1_t (new_AGEMA_signal_7310), .Z1_f (new_AGEMA_signal_7311) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line1_U8 ( .A0_t (ciphertext_s0_t[98]), .A0_f (ciphertext_s0_f[98]), .A1_t (ciphertext_s1_t[98]), .A1_f (ciphertext_s1_f[98]), .B0_t (ciphertext_s0_t[122]), .B0_f (ciphertext_s0_f[122]), .B1_t (ciphertext_s1_t[122]), .B1_f (ciphertext_s1_f[122]), .Z0_t (MixColumns_line1_n5), .Z0_f (new_AGEMA_signal_5634), .Z1_t (new_AGEMA_signal_5635), .Z1_f (new_AGEMA_signal_5636) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_U7 ( .A0_t (ciphertext_s0_t[113]), .A0_f (ciphertext_s0_f[113]), .A1_t (ciphertext_s1_t[113]), .A1_f (ciphertext_s1_f[113]), .B0_t (MixColumns_line1_S13[2]), .B0_f (new_AGEMA_signal_5661), .B1_t (new_AGEMA_signal_5662), .B1_f (new_AGEMA_signal_5663), .Z0_t (MixColumns_line1_n6), .Z0_f (new_AGEMA_signal_6529), .Z1_t (new_AGEMA_signal_6530), .Z1_f (new_AGEMA_signal_6531) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line1_U6 ( .A0_t (MixColumns_line1_n4), .A0_f (new_AGEMA_signal_7312), .A1_t (new_AGEMA_signal_7313), .A1_f (new_AGEMA_signal_7314), .B0_t (MixColumns_line1_n3), .B0_f (new_AGEMA_signal_5637), .B1_t (new_AGEMA_signal_5638), .B1_f (new_AGEMA_signal_5639), .Z0_t (MCout[17]), .Z0_f (new_AGEMA_signal_8094), .Z1_t (new_AGEMA_signal_8095), .Z1_f (new_AGEMA_signal_8096) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line1_U5 ( .A0_t (ciphertext_s0_t[121]), .A0_f (ciphertext_s0_f[121]), .A1_t (ciphertext_s1_t[121]), .A1_f (ciphertext_s1_f[121]), .B0_t (ciphertext_s0_t[97]), .B0_f (ciphertext_s0_f[97]), .B1_t (ciphertext_s1_t[97]), .B1_f (ciphertext_s1_f[97]), .Z0_t (MixColumns_line1_n3), .Z0_f (new_AGEMA_signal_5637), .Z1_t (new_AGEMA_signal_5638), .Z1_f (new_AGEMA_signal_5639) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_U4 ( .A0_t (MixColumns_line1_S02_1_), .A0_f (new_AGEMA_signal_5649), .A1_t (new_AGEMA_signal_5650), .A1_f (new_AGEMA_signal_5651), .B0_t (MixColumns_line1_S13[1]), .B0_f (new_AGEMA_signal_6541), .B1_t (new_AGEMA_signal_6542), .B1_f (new_AGEMA_signal_6543), .Z0_t (MixColumns_line1_n4), .Z0_f (new_AGEMA_signal_7312), .Z1_t (new_AGEMA_signal_7313), .Z1_f (new_AGEMA_signal_7314) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line1_U3 ( .A0_t (MixColumns_line1_n2), .A0_f (new_AGEMA_signal_6532), .A1_t (new_AGEMA_signal_6533), .A1_f (new_AGEMA_signal_6534), .B0_t (MixColumns_line1_n1), .B0_f (new_AGEMA_signal_5640), .B1_t (new_AGEMA_signal_5641), .B1_f (new_AGEMA_signal_5642), .Z0_t (MCout[16]), .Z0_f (new_AGEMA_signal_7315), .Z1_t (new_AGEMA_signal_7316), .Z1_f (new_AGEMA_signal_7317) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line1_U2 ( .A0_t (ciphertext_s0_t[120]), .A0_f (ciphertext_s0_f[120]), .A1_t (ciphertext_s1_t[120]), .A1_f (ciphertext_s1_f[120]), .B0_t (ciphertext_s0_t[96]), .B0_f (ciphertext_s0_f[96]), .B1_t (ciphertext_s1_t[96]), .B1_f (ciphertext_s1_f[96]), .Z0_t (MixColumns_line1_n1), .Z0_f (new_AGEMA_signal_5640), .Z1_t (new_AGEMA_signal_5641), .Z1_f (new_AGEMA_signal_5642) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_U1 ( .A0_t (ciphertext_s0_t[119]), .A0_f (ciphertext_s0_f[119]), .A1_t (ciphertext_s1_t[119]), .A1_f (ciphertext_s1_f[119]), .B0_t (MixColumns_line1_S13[0]), .B0_f (new_AGEMA_signal_5664), .B1_t (new_AGEMA_signal_5665), .B1_f (new_AGEMA_signal_5666), .Z0_t (MixColumns_line1_n2), .Z0_f (new_AGEMA_signal_6532), .Z1_t (new_AGEMA_signal_6533), .Z1_f (new_AGEMA_signal_6534) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_timesTWO_U3 ( .A0_t (ciphertext_s0_t[119]), .A0_f (ciphertext_s0_f[119]), .A1_t (ciphertext_s1_t[119]), .A1_f (ciphertext_s1_f[119]), .B0_t (ciphertext_s0_t[115]), .B0_f (ciphertext_s0_f[115]), .B1_t (ciphertext_s1_t[115]), .B1_f (ciphertext_s1_f[115]), .Z0_t (MixColumns_line1_S02_4_), .Z0_f (new_AGEMA_signal_5643), .Z1_t (new_AGEMA_signal_5644), .Z1_f (new_AGEMA_signal_5645) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_timesTWO_U2 ( .A0_t (ciphertext_s0_t[119]), .A0_f (ciphertext_s0_f[119]), .A1_t (ciphertext_s1_t[119]), .A1_f (ciphertext_s1_f[119]), .B0_t (ciphertext_s0_t[114]), .B0_f (ciphertext_s0_f[114]), .B1_t (ciphertext_s1_t[114]), .B1_f (ciphertext_s1_f[114]), .Z0_t (MixColumns_line1_S02_3_), .Z0_f (new_AGEMA_signal_5646), .Z1_t (new_AGEMA_signal_5647), .Z1_f (new_AGEMA_signal_5648) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_timesTWO_U1 ( .A0_t (ciphertext_s0_t[119]), .A0_f (ciphertext_s0_f[119]), .A1_t (ciphertext_s1_t[119]), .A1_f (ciphertext_s1_f[119]), .B0_t (ciphertext_s0_t[112]), .B0_f (ciphertext_s0_f[112]), .B1_t (ciphertext_s1_t[112]), .B1_f (ciphertext_s1_f[112]), .Z0_t (MixColumns_line1_S02_1_), .Z0_f (new_AGEMA_signal_5649), .Z1_t (new_AGEMA_signal_5650), .Z1_f (new_AGEMA_signal_5651) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_timesTHREE_U8 ( .A0_t (ciphertext_s0_t[111]), .A0_f (ciphertext_s0_f[111]), .A1_t (ciphertext_s1_t[111]), .A1_f (ciphertext_s1_f[111]), .B0_t (ciphertext_s0_t[110]), .B0_f (ciphertext_s0_f[110]), .B1_t (ciphertext_s1_t[110]), .B1_f (ciphertext_s1_f[110]), .Z0_t (MixColumns_line1_S13[7]), .Z0_f (new_AGEMA_signal_5652), .Z1_t (new_AGEMA_signal_5653), .Z1_f (new_AGEMA_signal_5654) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_timesTHREE_U7 ( .A0_t (ciphertext_s0_t[110]), .A0_f (ciphertext_s0_f[110]), .A1_t (ciphertext_s1_t[110]), .A1_f (ciphertext_s1_f[110]), .B0_t (ciphertext_s0_t[109]), .B0_f (ciphertext_s0_f[109]), .B1_t (ciphertext_s1_t[109]), .B1_f (ciphertext_s1_f[109]), .Z0_t (MixColumns_line1_S13[6]), .Z0_f (new_AGEMA_signal_5655), .Z1_t (new_AGEMA_signal_5656), .Z1_f (new_AGEMA_signal_5657) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_timesTHREE_U6 ( .A0_t (ciphertext_s0_t[109]), .A0_f (ciphertext_s0_f[109]), .A1_t (ciphertext_s1_t[109]), .A1_f (ciphertext_s1_f[109]), .B0_t (ciphertext_s0_t[108]), .B0_f (ciphertext_s0_f[108]), .B1_t (ciphertext_s1_t[108]), .B1_f (ciphertext_s1_f[108]), .Z0_t (MixColumns_line1_S13[5]), .Z0_f (new_AGEMA_signal_5658), .Z1_t (new_AGEMA_signal_5659), .Z1_f (new_AGEMA_signal_5660) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_timesTHREE_U5 ( .A0_t (ciphertext_s0_t[108]), .A0_f (ciphertext_s0_f[108]), .A1_t (ciphertext_s1_t[108]), .A1_f (ciphertext_s1_f[108]), .B0_t (MixColumns_line1_timesTHREE_input2[4]), .B0_f (new_AGEMA_signal_5667), .B1_t (new_AGEMA_signal_5668), .B1_f (new_AGEMA_signal_5669), .Z0_t (MixColumns_line1_S13[4]), .Z0_f (new_AGEMA_signal_6535), .Z1_t (new_AGEMA_signal_6536), .Z1_f (new_AGEMA_signal_6537) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_timesTHREE_U4 ( .A0_t (ciphertext_s0_t[107]), .A0_f (ciphertext_s0_f[107]), .A1_t (ciphertext_s1_t[107]), .A1_f (ciphertext_s1_f[107]), .B0_t (MixColumns_line1_timesTHREE_input2[3]), .B0_f (new_AGEMA_signal_5670), .B1_t (new_AGEMA_signal_5671), .B1_f (new_AGEMA_signal_5672), .Z0_t (MixColumns_line1_S13[3]), .Z0_f (new_AGEMA_signal_6538), .Z1_t (new_AGEMA_signal_6539), .Z1_f (new_AGEMA_signal_6540) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_timesTHREE_U3 ( .A0_t (ciphertext_s0_t[106]), .A0_f (ciphertext_s0_f[106]), .A1_t (ciphertext_s1_t[106]), .A1_f (ciphertext_s1_f[106]), .B0_t (ciphertext_s0_t[105]), .B0_f (ciphertext_s0_f[105]), .B1_t (ciphertext_s1_t[105]), .B1_f (ciphertext_s1_f[105]), .Z0_t (MixColumns_line1_S13[2]), .Z0_f (new_AGEMA_signal_5661), .Z1_t (new_AGEMA_signal_5662), .Z1_f (new_AGEMA_signal_5663) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_timesTHREE_U2 ( .A0_t (ciphertext_s0_t[105]), .A0_f (ciphertext_s0_f[105]), .A1_t (ciphertext_s1_t[105]), .A1_f (ciphertext_s1_f[105]), .B0_t (MixColumns_line1_timesTHREE_input2[1]), .B0_f (new_AGEMA_signal_5673), .B1_t (new_AGEMA_signal_5674), .B1_f (new_AGEMA_signal_5675), .Z0_t (MixColumns_line1_S13[1]), .Z0_f (new_AGEMA_signal_6541), .Z1_t (new_AGEMA_signal_6542), .Z1_f (new_AGEMA_signal_6543) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_timesTHREE_U1 ( .A0_t (ciphertext_s0_t[104]), .A0_f (ciphertext_s0_f[104]), .A1_t (ciphertext_s1_t[104]), .A1_f (ciphertext_s1_f[104]), .B0_t (ciphertext_s0_t[111]), .B0_f (ciphertext_s0_f[111]), .B1_t (ciphertext_s1_t[111]), .B1_f (ciphertext_s1_f[111]), .Z0_t (MixColumns_line1_S13[0]), .Z0_f (new_AGEMA_signal_5664), .Z1_t (new_AGEMA_signal_5665), .Z1_f (new_AGEMA_signal_5666) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_timesTHREE_timesTWO_U3 ( .A0_t (ciphertext_s0_t[111]), .A0_f (ciphertext_s0_f[111]), .A1_t (ciphertext_s1_t[111]), .A1_f (ciphertext_s1_f[111]), .B0_t (ciphertext_s0_t[107]), .B0_f (ciphertext_s0_f[107]), .B1_t (ciphertext_s1_t[107]), .B1_f (ciphertext_s1_f[107]), .Z0_t (MixColumns_line1_timesTHREE_input2[4]), .Z0_f (new_AGEMA_signal_5667), .Z1_t (new_AGEMA_signal_5668), .Z1_f (new_AGEMA_signal_5669) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_timesTHREE_timesTWO_U2 ( .A0_t (ciphertext_s0_t[111]), .A0_f (ciphertext_s0_f[111]), .A1_t (ciphertext_s1_t[111]), .A1_f (ciphertext_s1_f[111]), .B0_t (ciphertext_s0_t[106]), .B0_f (ciphertext_s0_f[106]), .B1_t (ciphertext_s1_t[106]), .B1_f (ciphertext_s1_f[106]), .Z0_t (MixColumns_line1_timesTHREE_input2[3]), .Z0_f (new_AGEMA_signal_5670), .Z1_t (new_AGEMA_signal_5671), .Z1_f (new_AGEMA_signal_5672) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_timesTHREE_timesTWO_U1 ( .A0_t (ciphertext_s0_t[111]), .A0_f (ciphertext_s0_f[111]), .A1_t (ciphertext_s1_t[111]), .A1_f (ciphertext_s1_f[111]), .B0_t (ciphertext_s0_t[104]), .B0_f (ciphertext_s0_f[104]), .B1_t (ciphertext_s1_t[104]), .B1_f (ciphertext_s1_f[104]), .Z0_t (MixColumns_line1_timesTHREE_input2[1]), .Z0_f (new_AGEMA_signal_5673), .Z1_t (new_AGEMA_signal_5674), .Z1_f (new_AGEMA_signal_5675) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line2_U24 ( .A0_t (MixColumns_line2_n16), .A0_f (new_AGEMA_signal_6544), .A1_t (new_AGEMA_signal_6545), .A1_f (new_AGEMA_signal_6546), .B0_t (MixColumns_line2_n15), .B0_f (new_AGEMA_signal_5676), .B1_t (new_AGEMA_signal_5677), .B1_f (new_AGEMA_signal_5678), .Z0_t (MCout[15]), .Z0_f (new_AGEMA_signal_7318), .Z1_t (new_AGEMA_signal_7319), .Z1_f (new_AGEMA_signal_7320) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line2_U23 ( .A0_t (ciphertext_s0_t[127]), .A0_f (ciphertext_s0_f[127]), .A1_t (ciphertext_s1_t[127]), .A1_f (ciphertext_s1_f[127]), .B0_t (ciphertext_s0_t[119]), .B0_f (ciphertext_s0_f[119]), .B1_t (ciphertext_s1_t[119]), .B1_f (ciphertext_s1_f[119]), .Z0_t (MixColumns_line2_n15), .Z0_f (new_AGEMA_signal_5676), .Z1_t (new_AGEMA_signal_5677), .Z1_f (new_AGEMA_signal_5678) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_U22 ( .A0_t (ciphertext_s0_t[110]), .A0_f (ciphertext_s0_f[110]), .A1_t (ciphertext_s1_t[110]), .A1_f (ciphertext_s1_f[110]), .B0_t (MixColumns_line2_S13[7]), .B0_f (new_AGEMA_signal_5709), .B1_t (new_AGEMA_signal_5710), .B1_f (new_AGEMA_signal_5711), .Z0_t (MixColumns_line2_n16), .Z0_f (new_AGEMA_signal_6544), .Z1_t (new_AGEMA_signal_6545), .Z1_f (new_AGEMA_signal_6546) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line2_U21 ( .A0_t (MixColumns_line2_n14), .A0_f (new_AGEMA_signal_6547), .A1_t (new_AGEMA_signal_6548), .A1_f (new_AGEMA_signal_6549), .B0_t (MixColumns_line2_n13), .B0_f (new_AGEMA_signal_5679), .B1_t (new_AGEMA_signal_5680), .B1_f (new_AGEMA_signal_5681), .Z0_t (MCout[14]), .Z0_f (new_AGEMA_signal_7321), .Z1_t (new_AGEMA_signal_7322), .Z1_f (new_AGEMA_signal_7323) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line2_U20 ( .A0_t (ciphertext_s0_t[126]), .A0_f (ciphertext_s0_f[126]), .A1_t (ciphertext_s1_t[126]), .A1_f (ciphertext_s1_f[126]), .B0_t (ciphertext_s0_t[118]), .B0_f (ciphertext_s0_f[118]), .B1_t (ciphertext_s1_t[118]), .B1_f (ciphertext_s1_f[118]), .Z0_t (MixColumns_line2_n13), .Z0_f (new_AGEMA_signal_5679), .Z1_t (new_AGEMA_signal_5680), .Z1_f (new_AGEMA_signal_5681) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_U19 ( .A0_t (ciphertext_s0_t[109]), .A0_f (ciphertext_s0_f[109]), .A1_t (ciphertext_s1_t[109]), .A1_f (ciphertext_s1_f[109]), .B0_t (MixColumns_line2_S13[6]), .B0_f (new_AGEMA_signal_5712), .B1_t (new_AGEMA_signal_5713), .B1_f (new_AGEMA_signal_5714), .Z0_t (MixColumns_line2_n14), .Z0_f (new_AGEMA_signal_6547), .Z1_t (new_AGEMA_signal_6548), .Z1_f (new_AGEMA_signal_6549) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line2_U18 ( .A0_t (MixColumns_line2_n12), .A0_f (new_AGEMA_signal_6550), .A1_t (new_AGEMA_signal_6551), .A1_f (new_AGEMA_signal_6552), .B0_t (MixColumns_line2_n11), .B0_f (new_AGEMA_signal_5682), .B1_t (new_AGEMA_signal_5683), .B1_f (new_AGEMA_signal_5684), .Z0_t (MCout[13]), .Z0_f (new_AGEMA_signal_7324), .Z1_t (new_AGEMA_signal_7325), .Z1_f (new_AGEMA_signal_7326) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line2_U17 ( .A0_t (ciphertext_s0_t[125]), .A0_f (ciphertext_s0_f[125]), .A1_t (ciphertext_s1_t[125]), .A1_f (ciphertext_s1_f[125]), .B0_t (ciphertext_s0_t[117]), .B0_f (ciphertext_s0_f[117]), .B1_t (ciphertext_s1_t[117]), .B1_f (ciphertext_s1_f[117]), .Z0_t (MixColumns_line2_n11), .Z0_f (new_AGEMA_signal_5682), .Z1_t (new_AGEMA_signal_5683), .Z1_f (new_AGEMA_signal_5684) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_U16 ( .A0_t (ciphertext_s0_t[108]), .A0_f (ciphertext_s0_f[108]), .A1_t (ciphertext_s1_t[108]), .A1_f (ciphertext_s1_f[108]), .B0_t (MixColumns_line2_S13[5]), .B0_f (new_AGEMA_signal_5715), .B1_t (new_AGEMA_signal_5716), .B1_f (new_AGEMA_signal_5717), .Z0_t (MixColumns_line2_n12), .Z0_f (new_AGEMA_signal_6550), .Z1_t (new_AGEMA_signal_6551), .Z1_f (new_AGEMA_signal_6552) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line2_U15 ( .A0_t (MixColumns_line2_n10), .A0_f (new_AGEMA_signal_7327), .A1_t (new_AGEMA_signal_7328), .A1_f (new_AGEMA_signal_7329), .B0_t (MixColumns_line2_n9), .B0_f (new_AGEMA_signal_5685), .B1_t (new_AGEMA_signal_5686), .B1_f (new_AGEMA_signal_5687), .Z0_t (MCout[12]), .Z0_f (new_AGEMA_signal_8097), .Z1_t (new_AGEMA_signal_8098), .Z1_f (new_AGEMA_signal_8099) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line2_U14 ( .A0_t (ciphertext_s0_t[124]), .A0_f (ciphertext_s0_f[124]), .A1_t (ciphertext_s1_t[124]), .A1_f (ciphertext_s1_f[124]), .B0_t (ciphertext_s0_t[116]), .B0_f (ciphertext_s0_f[116]), .B1_t (ciphertext_s1_t[116]), .B1_f (ciphertext_s1_f[116]), .Z0_t (MixColumns_line2_n9), .Z0_f (new_AGEMA_signal_5685), .Z1_t (new_AGEMA_signal_5686), .Z1_f (new_AGEMA_signal_5687) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_U13 ( .A0_t (MixColumns_line2_S02_4_), .A0_f (new_AGEMA_signal_5700), .A1_t (new_AGEMA_signal_5701), .A1_f (new_AGEMA_signal_5702), .B0_t (MixColumns_line2_S13[4]), .B0_f (new_AGEMA_signal_6559), .B1_t (new_AGEMA_signal_6560), .B1_f (new_AGEMA_signal_6561), .Z0_t (MixColumns_line2_n10), .Z0_f (new_AGEMA_signal_7327), .Z1_t (new_AGEMA_signal_7328), .Z1_f (new_AGEMA_signal_7329) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line2_U12 ( .A0_t (MixColumns_line2_n8), .A0_f (new_AGEMA_signal_7330), .A1_t (new_AGEMA_signal_7331), .A1_f (new_AGEMA_signal_7332), .B0_t (MixColumns_line2_n7), .B0_f (new_AGEMA_signal_5688), .B1_t (new_AGEMA_signal_5689), .B1_f (new_AGEMA_signal_5690), .Z0_t (MCout[11]), .Z0_f (new_AGEMA_signal_8100), .Z1_t (new_AGEMA_signal_8101), .Z1_f (new_AGEMA_signal_8102) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line2_U11 ( .A0_t (ciphertext_s0_t[123]), .A0_f (ciphertext_s0_f[123]), .A1_t (ciphertext_s1_t[123]), .A1_f (ciphertext_s1_f[123]), .B0_t (ciphertext_s0_t[115]), .B0_f (ciphertext_s0_f[115]), .B1_t (ciphertext_s1_t[115]), .B1_f (ciphertext_s1_f[115]), .Z0_t (MixColumns_line2_n7), .Z0_f (new_AGEMA_signal_5688), .Z1_t (new_AGEMA_signal_5689), .Z1_f (new_AGEMA_signal_5690) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_U10 ( .A0_t (MixColumns_line2_S02_3_), .A0_f (new_AGEMA_signal_5703), .A1_t (new_AGEMA_signal_5704), .A1_f (new_AGEMA_signal_5705), .B0_t (MixColumns_line2_S13[3]), .B0_f (new_AGEMA_signal_6562), .B1_t (new_AGEMA_signal_6563), .B1_f (new_AGEMA_signal_6564), .Z0_t (MixColumns_line2_n8), .Z0_f (new_AGEMA_signal_7330), .Z1_t (new_AGEMA_signal_7331), .Z1_f (new_AGEMA_signal_7332) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line2_U9 ( .A0_t (MixColumns_line2_n6), .A0_f (new_AGEMA_signal_6553), .A1_t (new_AGEMA_signal_6554), .A1_f (new_AGEMA_signal_6555), .B0_t (MixColumns_line2_n5), .B0_f (new_AGEMA_signal_5691), .B1_t (new_AGEMA_signal_5692), .B1_f (new_AGEMA_signal_5693), .Z0_t (MCout[10]), .Z0_f (new_AGEMA_signal_7333), .Z1_t (new_AGEMA_signal_7334), .Z1_f (new_AGEMA_signal_7335) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line2_U8 ( .A0_t (ciphertext_s0_t[122]), .A0_f (ciphertext_s0_f[122]), .A1_t (ciphertext_s1_t[122]), .A1_f (ciphertext_s1_f[122]), .B0_t (ciphertext_s0_t[114]), .B0_f (ciphertext_s0_f[114]), .B1_t (ciphertext_s1_t[114]), .B1_f (ciphertext_s1_f[114]), .Z0_t (MixColumns_line2_n5), .Z0_f (new_AGEMA_signal_5691), .Z1_t (new_AGEMA_signal_5692), .Z1_f (new_AGEMA_signal_5693) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_U7 ( .A0_t (ciphertext_s0_t[105]), .A0_f (ciphertext_s0_f[105]), .A1_t (ciphertext_s1_t[105]), .A1_f (ciphertext_s1_f[105]), .B0_t (MixColumns_line2_S13[2]), .B0_f (new_AGEMA_signal_5718), .B1_t (new_AGEMA_signal_5719), .B1_f (new_AGEMA_signal_5720), .Z0_t (MixColumns_line2_n6), .Z0_f (new_AGEMA_signal_6553), .Z1_t (new_AGEMA_signal_6554), .Z1_f (new_AGEMA_signal_6555) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line2_U6 ( .A0_t (MixColumns_line2_n4), .A0_f (new_AGEMA_signal_7336), .A1_t (new_AGEMA_signal_7337), .A1_f (new_AGEMA_signal_7338), .B0_t (MixColumns_line2_n3), .B0_f (new_AGEMA_signal_5694), .B1_t (new_AGEMA_signal_5695), .B1_f (new_AGEMA_signal_5696), .Z0_t (MCout[9]), .Z0_f (new_AGEMA_signal_8103), .Z1_t (new_AGEMA_signal_8104), .Z1_f (new_AGEMA_signal_8105) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line2_U5 ( .A0_t (ciphertext_s0_t[113]), .A0_f (ciphertext_s0_f[113]), .A1_t (ciphertext_s1_t[113]), .A1_f (ciphertext_s1_f[113]), .B0_t (ciphertext_s0_t[121]), .B0_f (ciphertext_s0_f[121]), .B1_t (ciphertext_s1_t[121]), .B1_f (ciphertext_s1_f[121]), .Z0_t (MixColumns_line2_n3), .Z0_f (new_AGEMA_signal_5694), .Z1_t (new_AGEMA_signal_5695), .Z1_f (new_AGEMA_signal_5696) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_U4 ( .A0_t (MixColumns_line2_S02_1_), .A0_f (new_AGEMA_signal_5706), .A1_t (new_AGEMA_signal_5707), .A1_f (new_AGEMA_signal_5708), .B0_t (MixColumns_line2_S13[1]), .B0_f (new_AGEMA_signal_6565), .B1_t (new_AGEMA_signal_6566), .B1_f (new_AGEMA_signal_6567), .Z0_t (MixColumns_line2_n4), .Z0_f (new_AGEMA_signal_7336), .Z1_t (new_AGEMA_signal_7337), .Z1_f (new_AGEMA_signal_7338) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line2_U3 ( .A0_t (MixColumns_line2_n2), .A0_f (new_AGEMA_signal_6556), .A1_t (new_AGEMA_signal_6557), .A1_f (new_AGEMA_signal_6558), .B0_t (MixColumns_line2_n1), .B0_f (new_AGEMA_signal_5697), .B1_t (new_AGEMA_signal_5698), .B1_f (new_AGEMA_signal_5699), .Z0_t (MCout[8]), .Z0_f (new_AGEMA_signal_7339), .Z1_t (new_AGEMA_signal_7340), .Z1_f (new_AGEMA_signal_7341) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line2_U2 ( .A0_t (ciphertext_s0_t[112]), .A0_f (ciphertext_s0_f[112]), .A1_t (ciphertext_s1_t[112]), .A1_f (ciphertext_s1_f[112]), .B0_t (ciphertext_s0_t[120]), .B0_f (ciphertext_s0_f[120]), .B1_t (ciphertext_s1_t[120]), .B1_f (ciphertext_s1_f[120]), .Z0_t (MixColumns_line2_n1), .Z0_f (new_AGEMA_signal_5697), .Z1_t (new_AGEMA_signal_5698), .Z1_f (new_AGEMA_signal_5699) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_U1 ( .A0_t (ciphertext_s0_t[111]), .A0_f (ciphertext_s0_f[111]), .A1_t (ciphertext_s1_t[111]), .A1_f (ciphertext_s1_f[111]), .B0_t (MixColumns_line2_S13[0]), .B0_f (new_AGEMA_signal_5721), .B1_t (new_AGEMA_signal_5722), .B1_f (new_AGEMA_signal_5723), .Z0_t (MixColumns_line2_n2), .Z0_f (new_AGEMA_signal_6556), .Z1_t (new_AGEMA_signal_6557), .Z1_f (new_AGEMA_signal_6558) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_timesTWO_U3 ( .A0_t (ciphertext_s0_t[111]), .A0_f (ciphertext_s0_f[111]), .A1_t (ciphertext_s1_t[111]), .A1_f (ciphertext_s1_f[111]), .B0_t (ciphertext_s0_t[107]), .B0_f (ciphertext_s0_f[107]), .B1_t (ciphertext_s1_t[107]), .B1_f (ciphertext_s1_f[107]), .Z0_t (MixColumns_line2_S02_4_), .Z0_f (new_AGEMA_signal_5700), .Z1_t (new_AGEMA_signal_5701), .Z1_f (new_AGEMA_signal_5702) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_timesTWO_U2 ( .A0_t (ciphertext_s0_t[111]), .A0_f (ciphertext_s0_f[111]), .A1_t (ciphertext_s1_t[111]), .A1_f (ciphertext_s1_f[111]), .B0_t (ciphertext_s0_t[106]), .B0_f (ciphertext_s0_f[106]), .B1_t (ciphertext_s1_t[106]), .B1_f (ciphertext_s1_f[106]), .Z0_t (MixColumns_line2_S02_3_), .Z0_f (new_AGEMA_signal_5703), .Z1_t (new_AGEMA_signal_5704), .Z1_f (new_AGEMA_signal_5705) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_timesTWO_U1 ( .A0_t (ciphertext_s0_t[111]), .A0_f (ciphertext_s0_f[111]), .A1_t (ciphertext_s1_t[111]), .A1_f (ciphertext_s1_f[111]), .B0_t (ciphertext_s0_t[104]), .B0_f (ciphertext_s0_f[104]), .B1_t (ciphertext_s1_t[104]), .B1_f (ciphertext_s1_f[104]), .Z0_t (MixColumns_line2_S02_1_), .Z0_f (new_AGEMA_signal_5706), .Z1_t (new_AGEMA_signal_5707), .Z1_f (new_AGEMA_signal_5708) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_timesTHREE_U8 ( .A0_t (ciphertext_s0_t[103]), .A0_f (ciphertext_s0_f[103]), .A1_t (ciphertext_s1_t[103]), .A1_f (ciphertext_s1_f[103]), .B0_t (ciphertext_s0_t[102]), .B0_f (ciphertext_s0_f[102]), .B1_t (ciphertext_s1_t[102]), .B1_f (ciphertext_s1_f[102]), .Z0_t (MixColumns_line2_S13[7]), .Z0_f (new_AGEMA_signal_5709), .Z1_t (new_AGEMA_signal_5710), .Z1_f (new_AGEMA_signal_5711) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_timesTHREE_U7 ( .A0_t (ciphertext_s0_t[102]), .A0_f (ciphertext_s0_f[102]), .A1_t (ciphertext_s1_t[102]), .A1_f (ciphertext_s1_f[102]), .B0_t (ciphertext_s0_t[101]), .B0_f (ciphertext_s0_f[101]), .B1_t (ciphertext_s1_t[101]), .B1_f (ciphertext_s1_f[101]), .Z0_t (MixColumns_line2_S13[6]), .Z0_f (new_AGEMA_signal_5712), .Z1_t (new_AGEMA_signal_5713), .Z1_f (new_AGEMA_signal_5714) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_timesTHREE_U6 ( .A0_t (ciphertext_s0_t[101]), .A0_f (ciphertext_s0_f[101]), .A1_t (ciphertext_s1_t[101]), .A1_f (ciphertext_s1_f[101]), .B0_t (ciphertext_s0_t[100]), .B0_f (ciphertext_s0_f[100]), .B1_t (ciphertext_s1_t[100]), .B1_f (ciphertext_s1_f[100]), .Z0_t (MixColumns_line2_S13[5]), .Z0_f (new_AGEMA_signal_5715), .Z1_t (new_AGEMA_signal_5716), .Z1_f (new_AGEMA_signal_5717) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_timesTHREE_U5 ( .A0_t (ciphertext_s0_t[100]), .A0_f (ciphertext_s0_f[100]), .A1_t (ciphertext_s1_t[100]), .A1_f (ciphertext_s1_f[100]), .B0_t (MixColumns_line2_timesTHREE_input2[4]), .B0_f (new_AGEMA_signal_5724), .B1_t (new_AGEMA_signal_5725), .B1_f (new_AGEMA_signal_5726), .Z0_t (MixColumns_line2_S13[4]), .Z0_f (new_AGEMA_signal_6559), .Z1_t (new_AGEMA_signal_6560), .Z1_f (new_AGEMA_signal_6561) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_timesTHREE_U4 ( .A0_t (ciphertext_s0_t[99]), .A0_f (ciphertext_s0_f[99]), .A1_t (ciphertext_s1_t[99]), .A1_f (ciphertext_s1_f[99]), .B0_t (MixColumns_line2_timesTHREE_input2[3]), .B0_f (new_AGEMA_signal_5727), .B1_t (new_AGEMA_signal_5728), .B1_f (new_AGEMA_signal_5729), .Z0_t (MixColumns_line2_S13[3]), .Z0_f (new_AGEMA_signal_6562), .Z1_t (new_AGEMA_signal_6563), .Z1_f (new_AGEMA_signal_6564) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_timesTHREE_U3 ( .A0_t (ciphertext_s0_t[98]), .A0_f (ciphertext_s0_f[98]), .A1_t (ciphertext_s1_t[98]), .A1_f (ciphertext_s1_f[98]), .B0_t (ciphertext_s0_t[97]), .B0_f (ciphertext_s0_f[97]), .B1_t (ciphertext_s1_t[97]), .B1_f (ciphertext_s1_f[97]), .Z0_t (MixColumns_line2_S13[2]), .Z0_f (new_AGEMA_signal_5718), .Z1_t (new_AGEMA_signal_5719), .Z1_f (new_AGEMA_signal_5720) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_timesTHREE_U2 ( .A0_t (ciphertext_s0_t[97]), .A0_f (ciphertext_s0_f[97]), .A1_t (ciphertext_s1_t[97]), .A1_f (ciphertext_s1_f[97]), .B0_t (MixColumns_line2_timesTHREE_input2[1]), .B0_f (new_AGEMA_signal_5730), .B1_t (new_AGEMA_signal_5731), .B1_f (new_AGEMA_signal_5732), .Z0_t (MixColumns_line2_S13[1]), .Z0_f (new_AGEMA_signal_6565), .Z1_t (new_AGEMA_signal_6566), .Z1_f (new_AGEMA_signal_6567) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_timesTHREE_U1 ( .A0_t (ciphertext_s0_t[96]), .A0_f (ciphertext_s0_f[96]), .A1_t (ciphertext_s1_t[96]), .A1_f (ciphertext_s1_f[96]), .B0_t (ciphertext_s0_t[103]), .B0_f (ciphertext_s0_f[103]), .B1_t (ciphertext_s1_t[103]), .B1_f (ciphertext_s1_f[103]), .Z0_t (MixColumns_line2_S13[0]), .Z0_f (new_AGEMA_signal_5721), .Z1_t (new_AGEMA_signal_5722), .Z1_f (new_AGEMA_signal_5723) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_timesTHREE_timesTWO_U3 ( .A0_t (ciphertext_s0_t[103]), .A0_f (ciphertext_s0_f[103]), .A1_t (ciphertext_s1_t[103]), .A1_f (ciphertext_s1_f[103]), .B0_t (ciphertext_s0_t[99]), .B0_f (ciphertext_s0_f[99]), .B1_t (ciphertext_s1_t[99]), .B1_f (ciphertext_s1_f[99]), .Z0_t (MixColumns_line2_timesTHREE_input2[4]), .Z0_f (new_AGEMA_signal_5724), .Z1_t (new_AGEMA_signal_5725), .Z1_f (new_AGEMA_signal_5726) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_timesTHREE_timesTWO_U2 ( .A0_t (ciphertext_s0_t[103]), .A0_f (ciphertext_s0_f[103]), .A1_t (ciphertext_s1_t[103]), .A1_f (ciphertext_s1_f[103]), .B0_t (ciphertext_s0_t[98]), .B0_f (ciphertext_s0_f[98]), .B1_t (ciphertext_s1_t[98]), .B1_f (ciphertext_s1_f[98]), .Z0_t (MixColumns_line2_timesTHREE_input2[3]), .Z0_f (new_AGEMA_signal_5727), .Z1_t (new_AGEMA_signal_5728), .Z1_f (new_AGEMA_signal_5729) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_timesTHREE_timesTWO_U1 ( .A0_t (ciphertext_s0_t[103]), .A0_f (ciphertext_s0_f[103]), .A1_t (ciphertext_s1_t[103]), .A1_f (ciphertext_s1_f[103]), .B0_t (ciphertext_s0_t[96]), .B0_f (ciphertext_s0_f[96]), .B1_t (ciphertext_s1_t[96]), .B1_f (ciphertext_s1_f[96]), .Z0_t (MixColumns_line2_timesTHREE_input2[1]), .Z0_f (new_AGEMA_signal_5730), .Z1_t (new_AGEMA_signal_5731), .Z1_f (new_AGEMA_signal_5732) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line3_U24 ( .A0_t (MixColumns_line3_n16), .A0_f (new_AGEMA_signal_6568), .A1_t (new_AGEMA_signal_6569), .A1_f (new_AGEMA_signal_6570), .B0_t (MixColumns_line3_n15), .B0_f (new_AGEMA_signal_5733), .B1_t (new_AGEMA_signal_5734), .B1_f (new_AGEMA_signal_5735), .Z0_t (MCout[7]), .Z0_f (new_AGEMA_signal_7342), .Z1_t (new_AGEMA_signal_7343), .Z1_f (new_AGEMA_signal_7344) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line3_U23 ( .A0_t (ciphertext_s0_t[119]), .A0_f (ciphertext_s0_f[119]), .A1_t (ciphertext_s1_t[119]), .A1_f (ciphertext_s1_f[119]), .B0_t (ciphertext_s0_t[111]), .B0_f (ciphertext_s0_f[111]), .B1_t (ciphertext_s1_t[111]), .B1_f (ciphertext_s1_f[111]), .Z0_t (MixColumns_line3_n15), .Z0_f (new_AGEMA_signal_5733), .Z1_t (new_AGEMA_signal_5734), .Z1_f (new_AGEMA_signal_5735) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_U22 ( .A0_t (ciphertext_s0_t[102]), .A0_f (ciphertext_s0_f[102]), .A1_t (ciphertext_s1_t[102]), .A1_f (ciphertext_s1_f[102]), .B0_t (MixColumns_line3_S13[7]), .B0_f (new_AGEMA_signal_5766), .B1_t (new_AGEMA_signal_5767), .B1_f (new_AGEMA_signal_5768), .Z0_t (MixColumns_line3_n16), .Z0_f (new_AGEMA_signal_6568), .Z1_t (new_AGEMA_signal_6569), .Z1_f (new_AGEMA_signal_6570) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line3_U21 ( .A0_t (MixColumns_line3_n14), .A0_f (new_AGEMA_signal_6571), .A1_t (new_AGEMA_signal_6572), .A1_f (new_AGEMA_signal_6573), .B0_t (MixColumns_line3_n13), .B0_f (new_AGEMA_signal_5736), .B1_t (new_AGEMA_signal_5737), .B1_f (new_AGEMA_signal_5738), .Z0_t (MCout[6]), .Z0_f (new_AGEMA_signal_7345), .Z1_t (new_AGEMA_signal_7346), .Z1_f (new_AGEMA_signal_7347) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line3_U20 ( .A0_t (ciphertext_s0_t[118]), .A0_f (ciphertext_s0_f[118]), .A1_t (ciphertext_s1_t[118]), .A1_f (ciphertext_s1_f[118]), .B0_t (ciphertext_s0_t[110]), .B0_f (ciphertext_s0_f[110]), .B1_t (ciphertext_s1_t[110]), .B1_f (ciphertext_s1_f[110]), .Z0_t (MixColumns_line3_n13), .Z0_f (new_AGEMA_signal_5736), .Z1_t (new_AGEMA_signal_5737), .Z1_f (new_AGEMA_signal_5738) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_U19 ( .A0_t (ciphertext_s0_t[101]), .A0_f (ciphertext_s0_f[101]), .A1_t (ciphertext_s1_t[101]), .A1_f (ciphertext_s1_f[101]), .B0_t (MixColumns_line3_S13[6]), .B0_f (new_AGEMA_signal_5769), .B1_t (new_AGEMA_signal_5770), .B1_f (new_AGEMA_signal_5771), .Z0_t (MixColumns_line3_n14), .Z0_f (new_AGEMA_signal_6571), .Z1_t (new_AGEMA_signal_6572), .Z1_f (new_AGEMA_signal_6573) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line3_U18 ( .A0_t (MixColumns_line3_n12), .A0_f (new_AGEMA_signal_6574), .A1_t (new_AGEMA_signal_6575), .A1_f (new_AGEMA_signal_6576), .B0_t (MixColumns_line3_n11), .B0_f (new_AGEMA_signal_5739), .B1_t (new_AGEMA_signal_5740), .B1_f (new_AGEMA_signal_5741), .Z0_t (MCout[5]), .Z0_f (new_AGEMA_signal_7348), .Z1_t (new_AGEMA_signal_7349), .Z1_f (new_AGEMA_signal_7350) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line3_U17 ( .A0_t (ciphertext_s0_t[117]), .A0_f (ciphertext_s0_f[117]), .A1_t (ciphertext_s1_t[117]), .A1_f (ciphertext_s1_f[117]), .B0_t (ciphertext_s0_t[109]), .B0_f (ciphertext_s0_f[109]), .B1_t (ciphertext_s1_t[109]), .B1_f (ciphertext_s1_f[109]), .Z0_t (MixColumns_line3_n11), .Z0_f (new_AGEMA_signal_5739), .Z1_t (new_AGEMA_signal_5740), .Z1_f (new_AGEMA_signal_5741) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_U16 ( .A0_t (ciphertext_s0_t[100]), .A0_f (ciphertext_s0_f[100]), .A1_t (ciphertext_s1_t[100]), .A1_f (ciphertext_s1_f[100]), .B0_t (MixColumns_line3_S13[5]), .B0_f (new_AGEMA_signal_5772), .B1_t (new_AGEMA_signal_5773), .B1_f (new_AGEMA_signal_5774), .Z0_t (MixColumns_line3_n12), .Z0_f (new_AGEMA_signal_6574), .Z1_t (new_AGEMA_signal_6575), .Z1_f (new_AGEMA_signal_6576) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line3_U15 ( .A0_t (MixColumns_line3_n10), .A0_f (new_AGEMA_signal_7351), .A1_t (new_AGEMA_signal_7352), .A1_f (new_AGEMA_signal_7353), .B0_t (MixColumns_line3_n9), .B0_f (new_AGEMA_signal_5742), .B1_t (new_AGEMA_signal_5743), .B1_f (new_AGEMA_signal_5744), .Z0_t (MCout[4]), .Z0_f (new_AGEMA_signal_8106), .Z1_t (new_AGEMA_signal_8107), .Z1_f (new_AGEMA_signal_8108) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line3_U14 ( .A0_t (ciphertext_s0_t[116]), .A0_f (ciphertext_s0_f[116]), .A1_t (ciphertext_s1_t[116]), .A1_f (ciphertext_s1_f[116]), .B0_t (ciphertext_s0_t[108]), .B0_f (ciphertext_s0_f[108]), .B1_t (ciphertext_s1_t[108]), .B1_f (ciphertext_s1_f[108]), .Z0_t (MixColumns_line3_n9), .Z0_f (new_AGEMA_signal_5742), .Z1_t (new_AGEMA_signal_5743), .Z1_f (new_AGEMA_signal_5744) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_U13 ( .A0_t (MixColumns_line3_S02_4_), .A0_f (new_AGEMA_signal_5757), .A1_t (new_AGEMA_signal_5758), .A1_f (new_AGEMA_signal_5759), .B0_t (MixColumns_line3_S13[4]), .B0_f (new_AGEMA_signal_6583), .B1_t (new_AGEMA_signal_6584), .B1_f (new_AGEMA_signal_6585), .Z0_t (MixColumns_line3_n10), .Z0_f (new_AGEMA_signal_7351), .Z1_t (new_AGEMA_signal_7352), .Z1_f (new_AGEMA_signal_7353) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line3_U12 ( .A0_t (MixColumns_line3_n8), .A0_f (new_AGEMA_signal_7354), .A1_t (new_AGEMA_signal_7355), .A1_f (new_AGEMA_signal_7356), .B0_t (MixColumns_line3_n7), .B0_f (new_AGEMA_signal_5745), .B1_t (new_AGEMA_signal_5746), .B1_f (new_AGEMA_signal_5747), .Z0_t (MCout[3]), .Z0_f (new_AGEMA_signal_8109), .Z1_t (new_AGEMA_signal_8110), .Z1_f (new_AGEMA_signal_8111) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line3_U11 ( .A0_t (ciphertext_s0_t[115]), .A0_f (ciphertext_s0_f[115]), .A1_t (ciphertext_s1_t[115]), .A1_f (ciphertext_s1_f[115]), .B0_t (ciphertext_s0_t[107]), .B0_f (ciphertext_s0_f[107]), .B1_t (ciphertext_s1_t[107]), .B1_f (ciphertext_s1_f[107]), .Z0_t (MixColumns_line3_n7), .Z0_f (new_AGEMA_signal_5745), .Z1_t (new_AGEMA_signal_5746), .Z1_f (new_AGEMA_signal_5747) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_U10 ( .A0_t (MixColumns_line3_S02_3_), .A0_f (new_AGEMA_signal_5760), .A1_t (new_AGEMA_signal_5761), .A1_f (new_AGEMA_signal_5762), .B0_t (MixColumns_line3_S13[3]), .B0_f (new_AGEMA_signal_6586), .B1_t (new_AGEMA_signal_6587), .B1_f (new_AGEMA_signal_6588), .Z0_t (MixColumns_line3_n8), .Z0_f (new_AGEMA_signal_7354), .Z1_t (new_AGEMA_signal_7355), .Z1_f (new_AGEMA_signal_7356) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line3_U9 ( .A0_t (MixColumns_line3_n6), .A0_f (new_AGEMA_signal_6577), .A1_t (new_AGEMA_signal_6578), .A1_f (new_AGEMA_signal_6579), .B0_t (MixColumns_line3_n5), .B0_f (new_AGEMA_signal_5748), .B1_t (new_AGEMA_signal_5749), .B1_f (new_AGEMA_signal_5750), .Z0_t (MCout[2]), .Z0_f (new_AGEMA_signal_7357), .Z1_t (new_AGEMA_signal_7358), .Z1_f (new_AGEMA_signal_7359) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line3_U8 ( .A0_t (ciphertext_s0_t[114]), .A0_f (ciphertext_s0_f[114]), .A1_t (ciphertext_s1_t[114]), .A1_f (ciphertext_s1_f[114]), .B0_t (ciphertext_s0_t[106]), .B0_f (ciphertext_s0_f[106]), .B1_t (ciphertext_s1_t[106]), .B1_f (ciphertext_s1_f[106]), .Z0_t (MixColumns_line3_n5), .Z0_f (new_AGEMA_signal_5748), .Z1_t (new_AGEMA_signal_5749), .Z1_f (new_AGEMA_signal_5750) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_U7 ( .A0_t (ciphertext_s0_t[97]), .A0_f (ciphertext_s0_f[97]), .A1_t (ciphertext_s1_t[97]), .A1_f (ciphertext_s1_f[97]), .B0_t (MixColumns_line3_S13[2]), .B0_f (new_AGEMA_signal_5775), .B1_t (new_AGEMA_signal_5776), .B1_f (new_AGEMA_signal_5777), .Z0_t (MixColumns_line3_n6), .Z0_f (new_AGEMA_signal_6577), .Z1_t (new_AGEMA_signal_6578), .Z1_f (new_AGEMA_signal_6579) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line3_U6 ( .A0_t (MixColumns_line3_n4), .A0_f (new_AGEMA_signal_7360), .A1_t (new_AGEMA_signal_7361), .A1_f (new_AGEMA_signal_7362), .B0_t (MixColumns_line3_n3), .B0_f (new_AGEMA_signal_5751), .B1_t (new_AGEMA_signal_5752), .B1_f (new_AGEMA_signal_5753), .Z0_t (MCout[1]), .Z0_f (new_AGEMA_signal_8112), .Z1_t (new_AGEMA_signal_8113), .Z1_f (new_AGEMA_signal_8114) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line3_U5 ( .A0_t (ciphertext_s0_t[105]), .A0_f (ciphertext_s0_f[105]), .A1_t (ciphertext_s1_t[105]), .A1_f (ciphertext_s1_f[105]), .B0_t (ciphertext_s0_t[113]), .B0_f (ciphertext_s0_f[113]), .B1_t (ciphertext_s1_t[113]), .B1_f (ciphertext_s1_f[113]), .Z0_t (MixColumns_line3_n3), .Z0_f (new_AGEMA_signal_5751), .Z1_t (new_AGEMA_signal_5752), .Z1_f (new_AGEMA_signal_5753) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_U4 ( .A0_t (MixColumns_line3_S02_1_), .A0_f (new_AGEMA_signal_5763), .A1_t (new_AGEMA_signal_5764), .A1_f (new_AGEMA_signal_5765), .B0_t (MixColumns_line3_S13[1]), .B0_f (new_AGEMA_signal_6589), .B1_t (new_AGEMA_signal_6590), .B1_f (new_AGEMA_signal_6591), .Z0_t (MixColumns_line3_n4), .Z0_f (new_AGEMA_signal_7360), .Z1_t (new_AGEMA_signal_7361), .Z1_f (new_AGEMA_signal_7362) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line3_U3 ( .A0_t (MixColumns_line3_n2), .A0_f (new_AGEMA_signal_6580), .A1_t (new_AGEMA_signal_6581), .A1_f (new_AGEMA_signal_6582), .B0_t (MixColumns_line3_n1), .B0_f (new_AGEMA_signal_5754), .B1_t (new_AGEMA_signal_5755), .B1_f (new_AGEMA_signal_5756), .Z0_t (MCout[0]), .Z0_f (new_AGEMA_signal_7363), .Z1_t (new_AGEMA_signal_7364), .Z1_f (new_AGEMA_signal_7365) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line3_U2 ( .A0_t (ciphertext_s0_t[104]), .A0_f (ciphertext_s0_f[104]), .A1_t (ciphertext_s1_t[104]), .A1_f (ciphertext_s1_f[104]), .B0_t (ciphertext_s0_t[112]), .B0_f (ciphertext_s0_f[112]), .B1_t (ciphertext_s1_t[112]), .B1_f (ciphertext_s1_f[112]), .Z0_t (MixColumns_line3_n1), .Z0_f (new_AGEMA_signal_5754), .Z1_t (new_AGEMA_signal_5755), .Z1_f (new_AGEMA_signal_5756) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_U1 ( .A0_t (ciphertext_s0_t[103]), .A0_f (ciphertext_s0_f[103]), .A1_t (ciphertext_s1_t[103]), .A1_f (ciphertext_s1_f[103]), .B0_t (MixColumns_line3_S13[0]), .B0_f (new_AGEMA_signal_5778), .B1_t (new_AGEMA_signal_5779), .B1_f (new_AGEMA_signal_5780), .Z0_t (MixColumns_line3_n2), .Z0_f (new_AGEMA_signal_6580), .Z1_t (new_AGEMA_signal_6581), .Z1_f (new_AGEMA_signal_6582) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_timesTWO_U3 ( .A0_t (ciphertext_s0_t[103]), .A0_f (ciphertext_s0_f[103]), .A1_t (ciphertext_s1_t[103]), .A1_f (ciphertext_s1_f[103]), .B0_t (ciphertext_s0_t[99]), .B0_f (ciphertext_s0_f[99]), .B1_t (ciphertext_s1_t[99]), .B1_f (ciphertext_s1_f[99]), .Z0_t (MixColumns_line3_S02_4_), .Z0_f (new_AGEMA_signal_5757), .Z1_t (new_AGEMA_signal_5758), .Z1_f (new_AGEMA_signal_5759) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_timesTWO_U2 ( .A0_t (ciphertext_s0_t[103]), .A0_f (ciphertext_s0_f[103]), .A1_t (ciphertext_s1_t[103]), .A1_f (ciphertext_s1_f[103]), .B0_t (ciphertext_s0_t[98]), .B0_f (ciphertext_s0_f[98]), .B1_t (ciphertext_s1_t[98]), .B1_f (ciphertext_s1_f[98]), .Z0_t (MixColumns_line3_S02_3_), .Z0_f (new_AGEMA_signal_5760), .Z1_t (new_AGEMA_signal_5761), .Z1_f (new_AGEMA_signal_5762) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_timesTWO_U1 ( .A0_t (ciphertext_s0_t[103]), .A0_f (ciphertext_s0_f[103]), .A1_t (ciphertext_s1_t[103]), .A1_f (ciphertext_s1_f[103]), .B0_t (ciphertext_s0_t[96]), .B0_f (ciphertext_s0_f[96]), .B1_t (ciphertext_s1_t[96]), .B1_f (ciphertext_s1_f[96]), .Z0_t (MixColumns_line3_S02_1_), .Z0_f (new_AGEMA_signal_5763), .Z1_t (new_AGEMA_signal_5764), .Z1_f (new_AGEMA_signal_5765) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_timesTHREE_U8 ( .A0_t (ciphertext_s0_t[127]), .A0_f (ciphertext_s0_f[127]), .A1_t (ciphertext_s1_t[127]), .A1_f (ciphertext_s1_f[127]), .B0_t (ciphertext_s0_t[126]), .B0_f (ciphertext_s0_f[126]), .B1_t (ciphertext_s1_t[126]), .B1_f (ciphertext_s1_f[126]), .Z0_t (MixColumns_line3_S13[7]), .Z0_f (new_AGEMA_signal_5766), .Z1_t (new_AGEMA_signal_5767), .Z1_f (new_AGEMA_signal_5768) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_timesTHREE_U7 ( .A0_t (ciphertext_s0_t[126]), .A0_f (ciphertext_s0_f[126]), .A1_t (ciphertext_s1_t[126]), .A1_f (ciphertext_s1_f[126]), .B0_t (ciphertext_s0_t[125]), .B0_f (ciphertext_s0_f[125]), .B1_t (ciphertext_s1_t[125]), .B1_f (ciphertext_s1_f[125]), .Z0_t (MixColumns_line3_S13[6]), .Z0_f (new_AGEMA_signal_5769), .Z1_t (new_AGEMA_signal_5770), .Z1_f (new_AGEMA_signal_5771) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_timesTHREE_U6 ( .A0_t (ciphertext_s0_t[125]), .A0_f (ciphertext_s0_f[125]), .A1_t (ciphertext_s1_t[125]), .A1_f (ciphertext_s1_f[125]), .B0_t (ciphertext_s0_t[124]), .B0_f (ciphertext_s0_f[124]), .B1_t (ciphertext_s1_t[124]), .B1_f (ciphertext_s1_f[124]), .Z0_t (MixColumns_line3_S13[5]), .Z0_f (new_AGEMA_signal_5772), .Z1_t (new_AGEMA_signal_5773), .Z1_f (new_AGEMA_signal_5774) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_timesTHREE_U5 ( .A0_t (ciphertext_s0_t[124]), .A0_f (ciphertext_s0_f[124]), .A1_t (ciphertext_s1_t[124]), .A1_f (ciphertext_s1_f[124]), .B0_t (MixColumns_line3_timesTHREE_input2_4_), .B0_f (new_AGEMA_signal_5781), .B1_t (new_AGEMA_signal_5782), .B1_f (new_AGEMA_signal_5783), .Z0_t (MixColumns_line3_S13[4]), .Z0_f (new_AGEMA_signal_6583), .Z1_t (new_AGEMA_signal_6584), .Z1_f (new_AGEMA_signal_6585) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_timesTHREE_U4 ( .A0_t (ciphertext_s0_t[123]), .A0_f (ciphertext_s0_f[123]), .A1_t (ciphertext_s1_t[123]), .A1_f (ciphertext_s1_f[123]), .B0_t (MixColumns_line3_timesTHREE_input2_3_), .B0_f (new_AGEMA_signal_5784), .B1_t (new_AGEMA_signal_5785), .B1_f (new_AGEMA_signal_5786), .Z0_t (MixColumns_line3_S13[3]), .Z0_f (new_AGEMA_signal_6586), .Z1_t (new_AGEMA_signal_6587), .Z1_f (new_AGEMA_signal_6588) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_timesTHREE_U3 ( .A0_t (ciphertext_s0_t[122]), .A0_f (ciphertext_s0_f[122]), .A1_t (ciphertext_s1_t[122]), .A1_f (ciphertext_s1_f[122]), .B0_t (ciphertext_s0_t[121]), .B0_f (ciphertext_s0_f[121]), .B1_t (ciphertext_s1_t[121]), .B1_f (ciphertext_s1_f[121]), .Z0_t (MixColumns_line3_S13[2]), .Z0_f (new_AGEMA_signal_5775), .Z1_t (new_AGEMA_signal_5776), .Z1_f (new_AGEMA_signal_5777) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_timesTHREE_U2 ( .A0_t (ciphertext_s0_t[121]), .A0_f (ciphertext_s0_f[121]), .A1_t (ciphertext_s1_t[121]), .A1_f (ciphertext_s1_f[121]), .B0_t (MixColumns_line3_timesTHREE_input2_1_), .B0_f (new_AGEMA_signal_5787), .B1_t (new_AGEMA_signal_5788), .B1_f (new_AGEMA_signal_5789), .Z0_t (MixColumns_line3_S13[1]), .Z0_f (new_AGEMA_signal_6589), .Z1_t (new_AGEMA_signal_6590), .Z1_f (new_AGEMA_signal_6591) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_timesTHREE_U1 ( .A0_t (ciphertext_s0_t[120]), .A0_f (ciphertext_s0_f[120]), .A1_t (ciphertext_s1_t[120]), .A1_f (ciphertext_s1_f[120]), .B0_t (ciphertext_s0_t[127]), .B0_f (ciphertext_s0_f[127]), .B1_t (ciphertext_s1_t[127]), .B1_f (ciphertext_s1_f[127]), .Z0_t (MixColumns_line3_S13[0]), .Z0_f (new_AGEMA_signal_5778), .Z1_t (new_AGEMA_signal_5779), .Z1_f (new_AGEMA_signal_5780) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_timesTHREE_timesTWO_U3 ( .A0_t (ciphertext_s0_t[127]), .A0_f (ciphertext_s0_f[127]), .A1_t (ciphertext_s1_t[127]), .A1_f (ciphertext_s1_f[127]), .B0_t (ciphertext_s0_t[123]), .B0_f (ciphertext_s0_f[123]), .B1_t (ciphertext_s1_t[123]), .B1_f (ciphertext_s1_f[123]), .Z0_t (MixColumns_line3_timesTHREE_input2_4_), .Z0_f (new_AGEMA_signal_5781), .Z1_t (new_AGEMA_signal_5782), .Z1_f (new_AGEMA_signal_5783) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_timesTHREE_timesTWO_U2 ( .A0_t (ciphertext_s0_t[127]), .A0_f (ciphertext_s0_f[127]), .A1_t (ciphertext_s1_t[127]), .A1_f (ciphertext_s1_f[127]), .B0_t (ciphertext_s0_t[122]), .B0_f (ciphertext_s0_f[122]), .B1_t (ciphertext_s1_t[122]), .B1_f (ciphertext_s1_f[122]), .Z0_t (MixColumns_line3_timesTHREE_input2_3_), .Z0_f (new_AGEMA_signal_5784), .Z1_t (new_AGEMA_signal_5785), .Z1_f (new_AGEMA_signal_5786) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_timesTHREE_timesTWO_U1 ( .A0_t (ciphertext_s0_t[127]), .A0_f (ciphertext_s0_f[127]), .A1_t (ciphertext_s1_t[127]), .A1_f (ciphertext_s1_f[127]), .B0_t (ciphertext_s0_t[120]), .B0_f (ciphertext_s0_f[120]), .B1_t (ciphertext_s1_t[120]), .B1_f (ciphertext_s1_f[120]), .Z0_t (MixColumns_line3_timesTHREE_input2_1_), .Z0_f (new_AGEMA_signal_5787), .Z1_t (new_AGEMA_signal_5788), .Z1_f (new_AGEMA_signal_5789) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U53 ( .A0_t (calcRCon_s_current_state_7_), .A0_f (new_AGEMA_signal_5790), .B0_t (enRCon), .B0_f (new_AGEMA_signal_5791), .Z0_t (roundConstant[7]), .Z0_f (new_AGEMA_signal_5792) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U52 ( .A0_t (calcRCon_s_current_state_6_), .A0_f (new_AGEMA_signal_5793), .B0_t (enRCon), .B0_f (new_AGEMA_signal_5791), .Z0_t (roundConstant[6]), .Z0_f (new_AGEMA_signal_5794) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U51 ( .A0_t (calcRCon_s_current_state_5_), .A0_f (new_AGEMA_signal_5795), .B0_t (enRCon), .B0_f (new_AGEMA_signal_5791), .Z0_t (roundConstant[5]), .Z0_f (new_AGEMA_signal_5796) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U50 ( .A0_t (calcRCon_s_current_state_4_), .A0_f (new_AGEMA_signal_5797), .B0_t (enRCon), .B0_f (new_AGEMA_signal_5791), .Z0_t (roundConstant[4]), .Z0_f (new_AGEMA_signal_5798) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U49 ( .A0_t (calcRCon_s_current_state_3_), .A0_f (new_AGEMA_signal_5799), .B0_t (enRCon), .B0_f (new_AGEMA_signal_5791), .Z0_t (roundConstant[3]), .Z0_f (new_AGEMA_signal_5800) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U48 ( .A0_t (calcRCon_s_current_state_2_), .A0_f (new_AGEMA_signal_5801), .B0_t (enRCon), .B0_f (new_AGEMA_signal_5791), .Z0_t (roundConstant[2]), .Z0_f (new_AGEMA_signal_5802) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U47 ( .A0_t (calcRCon_s_current_state_1_), .A0_f (new_AGEMA_signal_5803), .B0_t (enRCon), .B0_f (new_AGEMA_signal_5791), .Z0_t (roundConstant[1]), .Z0_f (new_AGEMA_signal_5804) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U46 ( .A0_t (calcRCon_s_current_state_0_), .A0_f (new_AGEMA_signal_5805), .B0_t (enRCon), .B0_f (new_AGEMA_signal_5791), .Z0_t (roundConstant[0]), .Z0_f (new_AGEMA_signal_5806) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) calcRCon_U44 ( .A0_t (calcRCon_n42), .A0_f (new_AGEMA_signal_6593), .B0_t (calcRCon_n41), .B0_f (new_AGEMA_signal_6592), .Z0_t (notFirst), .Z0_f (new_AGEMA_signal_7366) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U43 ( .A0_t (calcRCon_n40), .A0_f (new_AGEMA_signal_5808), .B0_t (calcRCon_n39), .B0_f (new_AGEMA_signal_5807), .Z0_t (calcRCon_n41), .Z0_f (new_AGEMA_signal_6592) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) calcRCon_U42 ( .A0_t (calcRCon_s_current_state_6_), .A0_f (new_AGEMA_signal_5793), .B0_t (calcRCon_s_current_state_5_), .B0_f (new_AGEMA_signal_5795), .Z0_t (calcRCon_n39), .Z0_f (new_AGEMA_signal_5807) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) calcRCon_U41 ( .A0_t (calcRCon_s_current_state_3_), .A0_f (new_AGEMA_signal_5799), .B0_t (calcRCon_s_current_state_7_), .B0_f (new_AGEMA_signal_5790), .Z0_t (calcRCon_n40), .Z0_f (new_AGEMA_signal_5808) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U40 ( .A0_t (calcRCon_n38), .A0_f (new_AGEMA_signal_5810), .B0_t (calcRCon_n37), .B0_f (new_AGEMA_signal_5809), .Z0_t (calcRCon_n42), .Z0_f (new_AGEMA_signal_6593) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) calcRCon_U39 ( .A0_t (calcRCon_s_current_state_2_), .A0_f (new_AGEMA_signal_5801), .B0_t (calcRCon_s_current_state_0_), .B0_f (new_AGEMA_signal_5805), .Z0_t (calcRCon_n37), .Z0_f (new_AGEMA_signal_5809) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) calcRCon_U38 ( .A0_t (calcRCon_s_current_state_1_), .A0_f (new_AGEMA_signal_5803), .B0_t (calcRCon_s_current_state_4_), .B0_f (new_AGEMA_signal_5797), .Z0_t (calcRCon_n38), .Z0_f (new_AGEMA_signal_5810) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1), .NL(1'b1)) calcRCon_U37 ( .A0_t (calcRCon_n36), .A0_f (new_AGEMA_signal_10260), .B0_t (calcRCon_n35), .B0_f (new_AGEMA_signal_9760), .Z0_t (calcRCon_s_current_state_0_), .Z0_f (new_AGEMA_signal_5805) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) calcRCon_U36 ( .A0_t (calcRCon_n34), .A0_f (new_AGEMA_signal_9272), .B0_t (calcRCon_s_current_state_0_), .B0_f (new_AGEMA_signal_5805), .Z0_t (calcRCon_n35), .Z0_f (new_AGEMA_signal_9760) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U35 ( .A0_t (nReset), .A0_f (new_AGEMA_signal_3502), .B0_t (calcRCon_n33), .B0_f (new_AGEMA_signal_9761), .Z0_t (calcRCon_n36), .Z0_f (new_AGEMA_signal_10260) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U34 ( .A0_t (calcRCon_n34), .A0_f (new_AGEMA_signal_9272), .B0_t (calcRCon_s_current_state_7_), .B0_f (new_AGEMA_signal_5790), .Z0_t (calcRCon_n33), .Z0_f (new_AGEMA_signal_9761) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1), .NL(1'b1)) calcRCon_U33 ( .A0_t (calcRCon_n32), .A0_f (new_AGEMA_signal_10261), .B0_t (calcRCon_n31), .B0_f (new_AGEMA_signal_9762), .Z0_t (calcRCon_s_current_state_1_), .Z0_f (new_AGEMA_signal_5803) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) calcRCon_U32 ( .A0_t (calcRCon_n34), .A0_f (new_AGEMA_signal_9272), .B0_t (calcRCon_s_current_state_1_), .B0_f (new_AGEMA_signal_5803), .Z0_t (calcRCon_n31), .Z0_f (new_AGEMA_signal_9762) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) calcRCon_U31 ( .A0_t (calcRCon_n30), .A0_f (new_AGEMA_signal_5811), .B0_t (calcRCon_n29), .B0_f (new_AGEMA_signal_9769), .Z0_t (calcRCon_n32), .Z0_f (new_AGEMA_signal_10261) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) calcRCon_U30 ( .A0_t (calcRCon_s_current_state_0_), .A0_f (new_AGEMA_signal_5805), .B0_t (calcRCon_s_current_state_7_), .B0_f (new_AGEMA_signal_5790), .Z0_t (calcRCon_n30), .Z0_f (new_AGEMA_signal_5811) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1), .NL(1'b1)) calcRCon_U29 ( .A0_t (nReset), .A0_f (new_AGEMA_signal_3502), .B0_t (calcRCon_n28), .B0_f (new_AGEMA_signal_10262), .Z0_t (calcRCon_s_current_state_2_), .Z0_f (new_AGEMA_signal_5801) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U28 ( .A0_t (calcRCon_n27), .A0_f (new_AGEMA_signal_9763), .B0_t (calcRCon_n26), .B0_f (new_AGEMA_signal_9270), .Z0_t (calcRCon_n28), .Z0_f (new_AGEMA_signal_10262) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U27 ( .A0_t (ctrl_n9), .A0_f (new_AGEMA_signal_7394), .B0_t (calcRCon_s_current_state_2_), .B0_f (new_AGEMA_signal_5801), .Z0_t (calcRCon_n26), .Z0_f (new_AGEMA_signal_9270) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U26 ( .A0_t (calcRCon_n34), .A0_f (new_AGEMA_signal_9272), .B0_t (calcRCon_s_current_state_1_), .B0_f (new_AGEMA_signal_5803), .Z0_t (calcRCon_n27), .Z0_f (new_AGEMA_signal_9763) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1), .NL(1'b1)) calcRCon_U25 ( .A0_t (calcRCon_n25), .A0_f (new_AGEMA_signal_10263), .B0_t (calcRCon_n24), .B0_f (new_AGEMA_signal_9764), .Z0_t (calcRCon_s_current_state_3_), .Z0_f (new_AGEMA_signal_5799) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) calcRCon_U24 ( .A0_t (calcRCon_n34), .A0_f (new_AGEMA_signal_9272), .B0_t (calcRCon_s_current_state_3_), .B0_f (new_AGEMA_signal_5799), .Z0_t (calcRCon_n24), .Z0_f (new_AGEMA_signal_9764) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U23 ( .A0_t (calcRCon_n23), .A0_f (new_AGEMA_signal_9765), .B0_t (nReset), .B0_f (new_AGEMA_signal_3502), .Z0_t (calcRCon_n25), .Z0_f (new_AGEMA_signal_10263) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U22 ( .A0_t (calcRCon_n34), .A0_f (new_AGEMA_signal_9272), .B0_t (calcRCon_n22), .B0_f (new_AGEMA_signal_5812), .Z0_t (calcRCon_n23), .Z0_f (new_AGEMA_signal_9765) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) calcRCon_U21 ( .A0_t (calcRCon_s_current_state_2_), .A0_f (new_AGEMA_signal_5801), .B0_t (calcRCon_s_current_state_7_), .B0_f (new_AGEMA_signal_5790), .Z0_t (calcRCon_n22), .Z0_f (new_AGEMA_signal_5812) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1), .NL(1'b1)) calcRCon_U20 ( .A0_t (calcRCon_n21), .A0_f (new_AGEMA_signal_10264), .B0_t (calcRCon_n20), .B0_f (new_AGEMA_signal_9766), .Z0_t (calcRCon_s_current_state_4_), .Z0_f (new_AGEMA_signal_5797) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) calcRCon_U19 ( .A0_t (calcRCon_n34), .A0_f (new_AGEMA_signal_9272), .B0_t (calcRCon_s_current_state_4_), .B0_f (new_AGEMA_signal_5797), .Z0_t (calcRCon_n20), .Z0_f (new_AGEMA_signal_9766) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) calcRCon_U18 ( .A0_t (calcRCon_n19), .A0_f (new_AGEMA_signal_5813), .B0_t (calcRCon_n29), .B0_f (new_AGEMA_signal_9769), .Z0_t (calcRCon_n21), .Z0_f (new_AGEMA_signal_10264) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) calcRCon_U17 ( .A0_t (calcRCon_s_current_state_3_), .A0_f (new_AGEMA_signal_5799), .B0_t (calcRCon_s_current_state_7_), .B0_f (new_AGEMA_signal_5790), .Z0_t (calcRCon_n19), .Z0_f (new_AGEMA_signal_5813) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1), .NL(1'b1)) calcRCon_U16 ( .A0_t (calcRCon_n18), .A0_f (new_AGEMA_signal_10265), .B0_t (calcRCon_n17), .B0_f (new_AGEMA_signal_9767), .Z0_t (calcRCon_s_current_state_5_), .Z0_f (new_AGEMA_signal_5795) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) calcRCon_U15 ( .A0_t (calcRCon_s_current_state_5_), .A0_f (new_AGEMA_signal_5795), .B0_t (calcRCon_n34), .B0_f (new_AGEMA_signal_9272), .Z0_t (calcRCon_n17), .Z0_f (new_AGEMA_signal_9767) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) calcRCon_U14 ( .A0_t (calcRCon_s_current_state_4_), .A0_f (new_AGEMA_signal_5797), .B0_t (calcRCon_n29), .B0_f (new_AGEMA_signal_9769), .Z0_t (calcRCon_n18), .Z0_f (new_AGEMA_signal_10265) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1), .NL(1'b1)) calcRCon_U13 ( .A0_t (calcRCon_n16), .A0_f (new_AGEMA_signal_10266), .B0_t (calcRCon_n15), .B0_f (new_AGEMA_signal_9768), .Z0_t (calcRCon_s_current_state_6_), .Z0_f (new_AGEMA_signal_5793) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) calcRCon_U12 ( .A0_t (calcRCon_s_current_state_6_), .A0_f (new_AGEMA_signal_5793), .B0_t (calcRCon_n34), .B0_f (new_AGEMA_signal_9272), .Z0_t (calcRCon_n15), .Z0_f (new_AGEMA_signal_9768) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) calcRCon_U11 ( .A0_t (calcRCon_s_current_state_5_), .A0_f (new_AGEMA_signal_5795), .B0_t (calcRCon_n29), .B0_f (new_AGEMA_signal_9769), .Z0_t (calcRCon_n16), .Z0_f (new_AGEMA_signal_10266) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U10 ( .A0_t (calcRCon_n34), .A0_f (new_AGEMA_signal_9272), .B0_t (nReset), .B0_f (new_AGEMA_signal_3502), .Z0_t (calcRCon_n29), .Z0_f (new_AGEMA_signal_9769) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1), .NL(1'b1)) calcRCon_U9 ( .A0_t (nReset), .A0_f (new_AGEMA_signal_3502), .B0_t (calcRCon_n14), .B0_f (new_AGEMA_signal_10267), .Z0_t (calcRCon_s_current_state_7_), .Z0_f (new_AGEMA_signal_5790) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U8 ( .A0_t (calcRCon_n13), .A0_f (new_AGEMA_signal_9770), .B0_t (calcRCon_n9), .B0_f (new_AGEMA_signal_9271), .Z0_t (calcRCon_n14), .Z0_f (new_AGEMA_signal_10267) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U7 ( .A0_t (ctrl_n9), .A0_f (new_AGEMA_signal_7394), .B0_t (calcRCon_s_current_state_7_), .B0_f (new_AGEMA_signal_5790), .Z0_t (calcRCon_n9), .Z0_f (new_AGEMA_signal_9271) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U6 ( .A0_t (calcRCon_n34), .A0_f (new_AGEMA_signal_9272), .B0_t (calcRCon_s_current_state_6_), .B0_f (new_AGEMA_signal_5793), .Z0_t (calcRCon_n13), .Z0_f (new_AGEMA_signal_9770) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U5 ( .A0_t (calcRCon_n8), .A0_f (new_AGEMA_signal_5815), .B0_t (calcRCon_n7), .B0_f (new_AGEMA_signal_5814), .Z0_t (intFinal), .Z0_f (new_AGEMA_signal_6594) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) calcRCon_U4 ( .A0_t (calcRCon_s_current_state_5_), .A0_f (new_AGEMA_signal_5795), .B0_t (calcRCon_s_current_state_4_), .B0_f (new_AGEMA_signal_5797), .Z0_t (calcRCon_n7), .Z0_f (new_AGEMA_signal_5814) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) calcRCon_U3 ( .A0_t (calcRCon_s_current_state_1_), .A0_f (new_AGEMA_signal_5803), .B0_t (calcRCon_s_current_state_2_), .B0_f (new_AGEMA_signal_5801), .Z0_t (calcRCon_n8), .Z0_f (new_AGEMA_signal_5815) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U1 ( .A0_t (ctrl_n9), .A0_f (new_AGEMA_signal_7394), .B0_t (nReset), .B0_f (new_AGEMA_signal_3502), .Z0_t (calcRCon_n34), .Z0_f (new_AGEMA_signal_9272) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_0_XOR1_U1 ( .A0_t (StateOutXORroundKey[0]), .A0_f (new_AGEMA_signal_3435), .A1_t (new_AGEMA_signal_3436), .A1_f (new_AGEMA_signal_3437), .B0_t (keySBIn[0]), .B0_f (new_AGEMA_signal_4797), .B1_t (new_AGEMA_signal_4798), .B1_f (new_AGEMA_signal_4799), .Z0_t (MUX_SboxIn_mux_inst_0_X), .Z0_f (new_AGEMA_signal_6595), .Z1_t (new_AGEMA_signal_6596), .Z1_f (new_AGEMA_signal_6597) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_0_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (MUX_SboxIn_mux_inst_0_X), .B0_f (new_AGEMA_signal_6595), .B1_t (new_AGEMA_signal_6596), .B1_f (new_AGEMA_signal_6597), .Z0_t (MUX_SboxIn_mux_inst_0_Y), .Z0_f (new_AGEMA_signal_7367), .Z1_t (new_AGEMA_signal_7368), .Z1_f (new_AGEMA_signal_7369) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_0_XOR2_U1 ( .A0_t (MUX_SboxIn_mux_inst_0_Y), .A0_f (new_AGEMA_signal_7367), .A1_t (new_AGEMA_signal_7368), .A1_f (new_AGEMA_signal_7369), .B0_t (StateOutXORroundKey[0]), .B0_f (new_AGEMA_signal_3435), .B1_t (new_AGEMA_signal_3436), .B1_f (new_AGEMA_signal_3437), .Z0_t (SboxIn[0]), .Z0_f (new_AGEMA_signal_8115), .Z1_t (new_AGEMA_signal_8116), .Z1_f (new_AGEMA_signal_8117) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_1_XOR1_U1 ( .A0_t (StateOutXORroundKey[1]), .A0_f (new_AGEMA_signal_3444), .A1_t (new_AGEMA_signal_3445), .A1_f (new_AGEMA_signal_3446), .B0_t (keySBIn[1]), .B0_f (new_AGEMA_signal_4806), .B1_t (new_AGEMA_signal_4807), .B1_f (new_AGEMA_signal_4808), .Z0_t (MUX_SboxIn_mux_inst_1_X), .Z0_f (new_AGEMA_signal_6598), .Z1_t (new_AGEMA_signal_6599), .Z1_f (new_AGEMA_signal_6600) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (MUX_SboxIn_mux_inst_1_X), .B0_f (new_AGEMA_signal_6598), .B1_t (new_AGEMA_signal_6599), .B1_f (new_AGEMA_signal_6600), .Z0_t (MUX_SboxIn_mux_inst_1_Y), .Z0_f (new_AGEMA_signal_7370), .Z1_t (new_AGEMA_signal_7371), .Z1_f (new_AGEMA_signal_7372) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_1_XOR2_U1 ( .A0_t (MUX_SboxIn_mux_inst_1_Y), .A0_f (new_AGEMA_signal_7370), .A1_t (new_AGEMA_signal_7371), .A1_f (new_AGEMA_signal_7372), .B0_t (StateOutXORroundKey[1]), .B0_f (new_AGEMA_signal_3444), .B1_t (new_AGEMA_signal_3445), .B1_f (new_AGEMA_signal_3446), .Z0_t (SboxIn[1]), .Z0_f (new_AGEMA_signal_8118), .Z1_t (new_AGEMA_signal_8119), .Z1_f (new_AGEMA_signal_8120) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_2_XOR1_U1 ( .A0_t (StateOutXORroundKey[2]), .A0_f (new_AGEMA_signal_3453), .A1_t (new_AGEMA_signal_3454), .A1_f (new_AGEMA_signal_3455), .B0_t (keySBIn[2]), .B0_f (new_AGEMA_signal_4815), .B1_t (new_AGEMA_signal_4816), .B1_f (new_AGEMA_signal_4817), .Z0_t (MUX_SboxIn_mux_inst_2_X), .Z0_f (new_AGEMA_signal_6601), .Z1_t (new_AGEMA_signal_6602), .Z1_f (new_AGEMA_signal_6603) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_2_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (MUX_SboxIn_mux_inst_2_X), .B0_f (new_AGEMA_signal_6601), .B1_t (new_AGEMA_signal_6602), .B1_f (new_AGEMA_signal_6603), .Z0_t (MUX_SboxIn_mux_inst_2_Y), .Z0_f (new_AGEMA_signal_7373), .Z1_t (new_AGEMA_signal_7374), .Z1_f (new_AGEMA_signal_7375) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_2_XOR2_U1 ( .A0_t (MUX_SboxIn_mux_inst_2_Y), .A0_f (new_AGEMA_signal_7373), .A1_t (new_AGEMA_signal_7374), .A1_f (new_AGEMA_signal_7375), .B0_t (StateOutXORroundKey[2]), .B0_f (new_AGEMA_signal_3453), .B1_t (new_AGEMA_signal_3454), .B1_f (new_AGEMA_signal_3455), .Z0_t (SboxIn[2]), .Z0_f (new_AGEMA_signal_8121), .Z1_t (new_AGEMA_signal_8122), .Z1_f (new_AGEMA_signal_8123) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_3_XOR1_U1 ( .A0_t (StateOutXORroundKey[3]), .A0_f (new_AGEMA_signal_3462), .A1_t (new_AGEMA_signal_3463), .A1_f (new_AGEMA_signal_3464), .B0_t (keySBIn[3]), .B0_f (new_AGEMA_signal_4824), .B1_t (new_AGEMA_signal_4825), .B1_f (new_AGEMA_signal_4826), .Z0_t (MUX_SboxIn_mux_inst_3_X), .Z0_f (new_AGEMA_signal_6604), .Z1_t (new_AGEMA_signal_6605), .Z1_f (new_AGEMA_signal_6606) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_3_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (MUX_SboxIn_mux_inst_3_X), .B0_f (new_AGEMA_signal_6604), .B1_t (new_AGEMA_signal_6605), .B1_f (new_AGEMA_signal_6606), .Z0_t (MUX_SboxIn_mux_inst_3_Y), .Z0_f (new_AGEMA_signal_7376), .Z1_t (new_AGEMA_signal_7377), .Z1_f (new_AGEMA_signal_7378) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_3_XOR2_U1 ( .A0_t (MUX_SboxIn_mux_inst_3_Y), .A0_f (new_AGEMA_signal_7376), .A1_t (new_AGEMA_signal_7377), .A1_f (new_AGEMA_signal_7378), .B0_t (StateOutXORroundKey[3]), .B0_f (new_AGEMA_signal_3462), .B1_t (new_AGEMA_signal_3463), .B1_f (new_AGEMA_signal_3464), .Z0_t (SboxIn[3]), .Z0_f (new_AGEMA_signal_8124), .Z1_t (new_AGEMA_signal_8125), .Z1_f (new_AGEMA_signal_8126) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_4_XOR1_U1 ( .A0_t (StateOutXORroundKey[4]), .A0_f (new_AGEMA_signal_3471), .A1_t (new_AGEMA_signal_3472), .A1_f (new_AGEMA_signal_3473), .B0_t (keySBIn[4]), .B0_f (new_AGEMA_signal_4833), .B1_t (new_AGEMA_signal_4834), .B1_f (new_AGEMA_signal_4835), .Z0_t (MUX_SboxIn_mux_inst_4_X), .Z0_f (new_AGEMA_signal_6607), .Z1_t (new_AGEMA_signal_6608), .Z1_f (new_AGEMA_signal_6609) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_4_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (MUX_SboxIn_mux_inst_4_X), .B0_f (new_AGEMA_signal_6607), .B1_t (new_AGEMA_signal_6608), .B1_f (new_AGEMA_signal_6609), .Z0_t (MUX_SboxIn_mux_inst_4_Y), .Z0_f (new_AGEMA_signal_7379), .Z1_t (new_AGEMA_signal_7380), .Z1_f (new_AGEMA_signal_7381) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_4_XOR2_U1 ( .A0_t (MUX_SboxIn_mux_inst_4_Y), .A0_f (new_AGEMA_signal_7379), .A1_t (new_AGEMA_signal_7380), .A1_f (new_AGEMA_signal_7381), .B0_t (StateOutXORroundKey[4]), .B0_f (new_AGEMA_signal_3471), .B1_t (new_AGEMA_signal_3472), .B1_f (new_AGEMA_signal_3473), .Z0_t (SboxIn[4]), .Z0_f (new_AGEMA_signal_8127), .Z1_t (new_AGEMA_signal_8128), .Z1_f (new_AGEMA_signal_8129) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_5_XOR1_U1 ( .A0_t (StateOutXORroundKey[5]), .A0_f (new_AGEMA_signal_3480), .A1_t (new_AGEMA_signal_3481), .A1_f (new_AGEMA_signal_3482), .B0_t (keySBIn[5]), .B0_f (new_AGEMA_signal_4842), .B1_t (new_AGEMA_signal_4843), .B1_f (new_AGEMA_signal_4844), .Z0_t (MUX_SboxIn_mux_inst_5_X), .Z0_f (new_AGEMA_signal_6610), .Z1_t (new_AGEMA_signal_6611), .Z1_f (new_AGEMA_signal_6612) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_5_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (MUX_SboxIn_mux_inst_5_X), .B0_f (new_AGEMA_signal_6610), .B1_t (new_AGEMA_signal_6611), .B1_f (new_AGEMA_signal_6612), .Z0_t (MUX_SboxIn_mux_inst_5_Y), .Z0_f (new_AGEMA_signal_7382), .Z1_t (new_AGEMA_signal_7383), .Z1_f (new_AGEMA_signal_7384) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_5_XOR2_U1 ( .A0_t (MUX_SboxIn_mux_inst_5_Y), .A0_f (new_AGEMA_signal_7382), .A1_t (new_AGEMA_signal_7383), .A1_f (new_AGEMA_signal_7384), .B0_t (StateOutXORroundKey[5]), .B0_f (new_AGEMA_signal_3480), .B1_t (new_AGEMA_signal_3481), .B1_f (new_AGEMA_signal_3482), .Z0_t (SboxIn[5]), .Z0_f (new_AGEMA_signal_8130), .Z1_t (new_AGEMA_signal_8131), .Z1_f (new_AGEMA_signal_8132) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_6_XOR1_U1 ( .A0_t (StateOutXORroundKey[6]), .A0_f (new_AGEMA_signal_3489), .A1_t (new_AGEMA_signal_3490), .A1_f (new_AGEMA_signal_3491), .B0_t (keySBIn[6]), .B0_f (new_AGEMA_signal_4851), .B1_t (new_AGEMA_signal_4852), .B1_f (new_AGEMA_signal_4853), .Z0_t (MUX_SboxIn_mux_inst_6_X), .Z0_f (new_AGEMA_signal_6613), .Z1_t (new_AGEMA_signal_6614), .Z1_f (new_AGEMA_signal_6615) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_6_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (MUX_SboxIn_mux_inst_6_X), .B0_f (new_AGEMA_signal_6613), .B1_t (new_AGEMA_signal_6614), .B1_f (new_AGEMA_signal_6615), .Z0_t (MUX_SboxIn_mux_inst_6_Y), .Z0_f (new_AGEMA_signal_7385), .Z1_t (new_AGEMA_signal_7386), .Z1_f (new_AGEMA_signal_7387) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_6_XOR2_U1 ( .A0_t (MUX_SboxIn_mux_inst_6_Y), .A0_f (new_AGEMA_signal_7385), .A1_t (new_AGEMA_signal_7386), .A1_f (new_AGEMA_signal_7387), .B0_t (StateOutXORroundKey[6]), .B0_f (new_AGEMA_signal_3489), .B1_t (new_AGEMA_signal_3490), .B1_f (new_AGEMA_signal_3491), .Z0_t (SboxIn[6]), .Z0_f (new_AGEMA_signal_8133), .Z1_t (new_AGEMA_signal_8134), .Z1_f (new_AGEMA_signal_8135) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_7_XOR1_U1 ( .A0_t (StateOutXORroundKey[7]), .A0_f (new_AGEMA_signal_3498), .A1_t (new_AGEMA_signal_3499), .A1_f (new_AGEMA_signal_3500), .B0_t (keySBIn[7]), .B0_f (new_AGEMA_signal_4860), .B1_t (new_AGEMA_signal_4861), .B1_f (new_AGEMA_signal_4862), .Z0_t (MUX_SboxIn_mux_inst_7_X), .Z0_f (new_AGEMA_signal_6616), .Z1_t (new_AGEMA_signal_6617), .Z1_f (new_AGEMA_signal_6618) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_7_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_3503), .B0_t (MUX_SboxIn_mux_inst_7_X), .B0_f (new_AGEMA_signal_6616), .B1_t (new_AGEMA_signal_6617), .B1_f (new_AGEMA_signal_6618), .Z0_t (MUX_SboxIn_mux_inst_7_Y), .Z0_f (new_AGEMA_signal_7388), .Z1_t (new_AGEMA_signal_7389), .Z1_f (new_AGEMA_signal_7390) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_7_XOR2_U1 ( .A0_t (MUX_SboxIn_mux_inst_7_Y), .A0_f (new_AGEMA_signal_7388), .A1_t (new_AGEMA_signal_7389), .A1_f (new_AGEMA_signal_7390), .B0_t (StateOutXORroundKey[7]), .B0_f (new_AGEMA_signal_3498), .B1_t (new_AGEMA_signal_3499), .B1_f (new_AGEMA_signal_3500), .Z0_t (SboxIn[7]), .Z0_f (new_AGEMA_signal_8136), .Z1_t (new_AGEMA_signal_8137), .Z1_f (new_AGEMA_signal_8138) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T1_U1 ( .A0_t (SboxIn[7]), .A0_f (new_AGEMA_signal_8136), .A1_t (new_AGEMA_signal_8137), .A1_f (new_AGEMA_signal_8138), .B0_t (SboxIn[4]), .B0_f (new_AGEMA_signal_8127), .B1_t (new_AGEMA_signal_8128), .B1_f (new_AGEMA_signal_8129), .Z0_t (Inst_bSbox_T1), .Z0_f (new_AGEMA_signal_9273), .Z1_t (new_AGEMA_signal_9274), .Z1_f (new_AGEMA_signal_9275) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T2_U1 ( .A0_t (SboxIn[7]), .A0_f (new_AGEMA_signal_8136), .A1_t (new_AGEMA_signal_8137), .A1_f (new_AGEMA_signal_8138), .B0_t (SboxIn[2]), .B0_f (new_AGEMA_signal_8121), .B1_t (new_AGEMA_signal_8122), .B1_f (new_AGEMA_signal_8123), .Z0_t (Inst_bSbox_T2), .Z0_f (new_AGEMA_signal_9276), .Z1_t (new_AGEMA_signal_9277), .Z1_f (new_AGEMA_signal_9278) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T3_U1 ( .A0_t (SboxIn[7]), .A0_f (new_AGEMA_signal_8136), .A1_t (new_AGEMA_signal_8137), .A1_f (new_AGEMA_signal_8138), .B0_t (SboxIn[1]), .B0_f (new_AGEMA_signal_8118), .B1_t (new_AGEMA_signal_8119), .B1_f (new_AGEMA_signal_8120), .Z0_t (Inst_bSbox_T3), .Z0_f (new_AGEMA_signal_9279), .Z1_t (new_AGEMA_signal_9280), .Z1_f (new_AGEMA_signal_9281) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T4_U1 ( .A0_t (SboxIn[4]), .A0_f (new_AGEMA_signal_8127), .A1_t (new_AGEMA_signal_8128), .A1_f (new_AGEMA_signal_8129), .B0_t (SboxIn[2]), .B0_f (new_AGEMA_signal_8121), .B1_t (new_AGEMA_signal_8122), .B1_f (new_AGEMA_signal_8123), .Z0_t (Inst_bSbox_T4), .Z0_f (new_AGEMA_signal_9282), .Z1_t (new_AGEMA_signal_9283), .Z1_f (new_AGEMA_signal_9284) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T5_U1 ( .A0_t (SboxIn[3]), .A0_f (new_AGEMA_signal_8124), .A1_t (new_AGEMA_signal_8125), .A1_f (new_AGEMA_signal_8126), .B0_t (SboxIn[1]), .B0_f (new_AGEMA_signal_8118), .B1_t (new_AGEMA_signal_8119), .B1_f (new_AGEMA_signal_8120), .Z0_t (Inst_bSbox_T5), .Z0_f (new_AGEMA_signal_9285), .Z1_t (new_AGEMA_signal_9286), .Z1_f (new_AGEMA_signal_9287) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T6_U1 ( .A0_t (Inst_bSbox_T1), .A0_f (new_AGEMA_signal_9273), .A1_t (new_AGEMA_signal_9274), .A1_f (new_AGEMA_signal_9275), .B0_t (Inst_bSbox_T5), .B0_f (new_AGEMA_signal_9285), .B1_t (new_AGEMA_signal_9286), .B1_f (new_AGEMA_signal_9287), .Z0_t (Inst_bSbox_T6), .Z0_f (new_AGEMA_signal_9771), .Z1_t (new_AGEMA_signal_9772), .Z1_f (new_AGEMA_signal_9773) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T7_U1 ( .A0_t (SboxIn[6]), .A0_f (new_AGEMA_signal_8133), .A1_t (new_AGEMA_signal_8134), .A1_f (new_AGEMA_signal_8135), .B0_t (SboxIn[5]), .B0_f (new_AGEMA_signal_8130), .B1_t (new_AGEMA_signal_8131), .B1_f (new_AGEMA_signal_8132), .Z0_t (Inst_bSbox_T7), .Z0_f (new_AGEMA_signal_9288), .Z1_t (new_AGEMA_signal_9289), .Z1_f (new_AGEMA_signal_9290) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T8_U1 ( .A0_t (SboxIn[0]), .A0_f (new_AGEMA_signal_8115), .A1_t (new_AGEMA_signal_8116), .A1_f (new_AGEMA_signal_8117), .B0_t (Inst_bSbox_T6), .B0_f (new_AGEMA_signal_9771), .B1_t (new_AGEMA_signal_9772), .B1_f (new_AGEMA_signal_9773), .Z0_t (Inst_bSbox_T8), .Z0_f (new_AGEMA_signal_10268), .Z1_t (new_AGEMA_signal_10269), .Z1_f (new_AGEMA_signal_10270) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T9_U1 ( .A0_t (SboxIn[0]), .A0_f (new_AGEMA_signal_8115), .A1_t (new_AGEMA_signal_8116), .A1_f (new_AGEMA_signal_8117), .B0_t (Inst_bSbox_T7), .B0_f (new_AGEMA_signal_9288), .B1_t (new_AGEMA_signal_9289), .B1_f (new_AGEMA_signal_9290), .Z0_t (Inst_bSbox_T9), .Z0_f (new_AGEMA_signal_9774), .Z1_t (new_AGEMA_signal_9775), .Z1_f (new_AGEMA_signal_9776) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T10_U1 ( .A0_t (Inst_bSbox_T6), .A0_f (new_AGEMA_signal_9771), .A1_t (new_AGEMA_signal_9772), .A1_f (new_AGEMA_signal_9773), .B0_t (Inst_bSbox_T7), .B0_f (new_AGEMA_signal_9288), .B1_t (new_AGEMA_signal_9289), .B1_f (new_AGEMA_signal_9290), .Z0_t (Inst_bSbox_T10), .Z0_f (new_AGEMA_signal_10271), .Z1_t (new_AGEMA_signal_10272), .Z1_f (new_AGEMA_signal_10273) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T11_U1 ( .A0_t (SboxIn[6]), .A0_f (new_AGEMA_signal_8133), .A1_t (new_AGEMA_signal_8134), .A1_f (new_AGEMA_signal_8135), .B0_t (SboxIn[2]), .B0_f (new_AGEMA_signal_8121), .B1_t (new_AGEMA_signal_8122), .B1_f (new_AGEMA_signal_8123), .Z0_t (Inst_bSbox_T11), .Z0_f (new_AGEMA_signal_9291), .Z1_t (new_AGEMA_signal_9292), .Z1_f (new_AGEMA_signal_9293) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T12_U1 ( .A0_t (SboxIn[5]), .A0_f (new_AGEMA_signal_8130), .A1_t (new_AGEMA_signal_8131), .A1_f (new_AGEMA_signal_8132), .B0_t (SboxIn[2]), .B0_f (new_AGEMA_signal_8121), .B1_t (new_AGEMA_signal_8122), .B1_f (new_AGEMA_signal_8123), .Z0_t (Inst_bSbox_T12), .Z0_f (new_AGEMA_signal_9294), .Z1_t (new_AGEMA_signal_9295), .Z1_f (new_AGEMA_signal_9296) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T13_U1 ( .A0_t (Inst_bSbox_T3), .A0_f (new_AGEMA_signal_9279), .A1_t (new_AGEMA_signal_9280), .A1_f (new_AGEMA_signal_9281), .B0_t (Inst_bSbox_T4), .B0_f (new_AGEMA_signal_9282), .B1_t (new_AGEMA_signal_9283), .B1_f (new_AGEMA_signal_9284), .Z0_t (Inst_bSbox_T13), .Z0_f (new_AGEMA_signal_9777), .Z1_t (new_AGEMA_signal_9778), .Z1_f (new_AGEMA_signal_9779) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T14_U1 ( .A0_t (Inst_bSbox_T6), .A0_f (new_AGEMA_signal_9771), .A1_t (new_AGEMA_signal_9772), .A1_f (new_AGEMA_signal_9773), .B0_t (Inst_bSbox_T11), .B0_f (new_AGEMA_signal_9291), .B1_t (new_AGEMA_signal_9292), .B1_f (new_AGEMA_signal_9293), .Z0_t (Inst_bSbox_T14), .Z0_f (new_AGEMA_signal_10274), .Z1_t (new_AGEMA_signal_10275), .Z1_f (new_AGEMA_signal_10276) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T15_U1 ( .A0_t (Inst_bSbox_T5), .A0_f (new_AGEMA_signal_9285), .A1_t (new_AGEMA_signal_9286), .A1_f (new_AGEMA_signal_9287), .B0_t (Inst_bSbox_T11), .B0_f (new_AGEMA_signal_9291), .B1_t (new_AGEMA_signal_9292), .B1_f (new_AGEMA_signal_9293), .Z0_t (Inst_bSbox_T15), .Z0_f (new_AGEMA_signal_9780), .Z1_t (new_AGEMA_signal_9781), .Z1_f (new_AGEMA_signal_9782) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T16_U1 ( .A0_t (Inst_bSbox_T5), .A0_f (new_AGEMA_signal_9285), .A1_t (new_AGEMA_signal_9286), .A1_f (new_AGEMA_signal_9287), .B0_t (Inst_bSbox_T12), .B0_f (new_AGEMA_signal_9294), .B1_t (new_AGEMA_signal_9295), .B1_f (new_AGEMA_signal_9296), .Z0_t (Inst_bSbox_T16), .Z0_f (new_AGEMA_signal_9783), .Z1_t (new_AGEMA_signal_9784), .Z1_f (new_AGEMA_signal_9785) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T17_U1 ( .A0_t (Inst_bSbox_T9), .A0_f (new_AGEMA_signal_9774), .A1_t (new_AGEMA_signal_9775), .A1_f (new_AGEMA_signal_9776), .B0_t (Inst_bSbox_T16), .B0_f (new_AGEMA_signal_9783), .B1_t (new_AGEMA_signal_9784), .B1_f (new_AGEMA_signal_9785), .Z0_t (Inst_bSbox_T17), .Z0_f (new_AGEMA_signal_10277), .Z1_t (new_AGEMA_signal_10278), .Z1_f (new_AGEMA_signal_10279) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T18_U1 ( .A0_t (SboxIn[4]), .A0_f (new_AGEMA_signal_8127), .A1_t (new_AGEMA_signal_8128), .A1_f (new_AGEMA_signal_8129), .B0_t (SboxIn[0]), .B0_f (new_AGEMA_signal_8115), .B1_t (new_AGEMA_signal_8116), .B1_f (new_AGEMA_signal_8117), .Z0_t (Inst_bSbox_T18), .Z0_f (new_AGEMA_signal_9297), .Z1_t (new_AGEMA_signal_9298), .Z1_f (new_AGEMA_signal_9299) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T19_U1 ( .A0_t (Inst_bSbox_T7), .A0_f (new_AGEMA_signal_9288), .A1_t (new_AGEMA_signal_9289), .A1_f (new_AGEMA_signal_9290), .B0_t (Inst_bSbox_T18), .B0_f (new_AGEMA_signal_9297), .B1_t (new_AGEMA_signal_9298), .B1_f (new_AGEMA_signal_9299), .Z0_t (Inst_bSbox_T19), .Z0_f (new_AGEMA_signal_9786), .Z1_t (new_AGEMA_signal_9787), .Z1_f (new_AGEMA_signal_9788) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T20_U1 ( .A0_t (Inst_bSbox_T1), .A0_f (new_AGEMA_signal_9273), .A1_t (new_AGEMA_signal_9274), .A1_f (new_AGEMA_signal_9275), .B0_t (Inst_bSbox_T19), .B0_f (new_AGEMA_signal_9786), .B1_t (new_AGEMA_signal_9787), .B1_f (new_AGEMA_signal_9788), .Z0_t (Inst_bSbox_T20), .Z0_f (new_AGEMA_signal_10280), .Z1_t (new_AGEMA_signal_10281), .Z1_f (new_AGEMA_signal_10282) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T21_U1 ( .A0_t (SboxIn[1]), .A0_f (new_AGEMA_signal_8118), .A1_t (new_AGEMA_signal_8119), .A1_f (new_AGEMA_signal_8120), .B0_t (SboxIn[0]), .B0_f (new_AGEMA_signal_8115), .B1_t (new_AGEMA_signal_8116), .B1_f (new_AGEMA_signal_8117), .Z0_t (Inst_bSbox_T21), .Z0_f (new_AGEMA_signal_9300), .Z1_t (new_AGEMA_signal_9301), .Z1_f (new_AGEMA_signal_9302) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T22_U1 ( .A0_t (Inst_bSbox_T7), .A0_f (new_AGEMA_signal_9288), .A1_t (new_AGEMA_signal_9289), .A1_f (new_AGEMA_signal_9290), .B0_t (Inst_bSbox_T21), .B0_f (new_AGEMA_signal_9300), .B1_t (new_AGEMA_signal_9301), .B1_f (new_AGEMA_signal_9302), .Z0_t (Inst_bSbox_T22), .Z0_f (new_AGEMA_signal_9789), .Z1_t (new_AGEMA_signal_9790), .Z1_f (new_AGEMA_signal_9791) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T23_U1 ( .A0_t (Inst_bSbox_T2), .A0_f (new_AGEMA_signal_9276), .A1_t (new_AGEMA_signal_9277), .A1_f (new_AGEMA_signal_9278), .B0_t (Inst_bSbox_T22), .B0_f (new_AGEMA_signal_9789), .B1_t (new_AGEMA_signal_9790), .B1_f (new_AGEMA_signal_9791), .Z0_t (Inst_bSbox_T23), .Z0_f (new_AGEMA_signal_10283), .Z1_t (new_AGEMA_signal_10284), .Z1_f (new_AGEMA_signal_10285) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T24_U1 ( .A0_t (Inst_bSbox_T2), .A0_f (new_AGEMA_signal_9276), .A1_t (new_AGEMA_signal_9277), .A1_f (new_AGEMA_signal_9278), .B0_t (Inst_bSbox_T10), .B0_f (new_AGEMA_signal_10271), .B1_t (new_AGEMA_signal_10272), .B1_f (new_AGEMA_signal_10273), .Z0_t (Inst_bSbox_T24), .Z0_f (new_AGEMA_signal_10403), .Z1_t (new_AGEMA_signal_10404), .Z1_f (new_AGEMA_signal_10405) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T25_U1 ( .A0_t (Inst_bSbox_T20), .A0_f (new_AGEMA_signal_10280), .A1_t (new_AGEMA_signal_10281), .A1_f (new_AGEMA_signal_10282), .B0_t (Inst_bSbox_T17), .B0_f (new_AGEMA_signal_10277), .B1_t (new_AGEMA_signal_10278), .B1_f (new_AGEMA_signal_10279), .Z0_t (Inst_bSbox_T25), .Z0_f (new_AGEMA_signal_10406), .Z1_t (new_AGEMA_signal_10407), .Z1_f (new_AGEMA_signal_10408) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T26_U1 ( .A0_t (Inst_bSbox_T3), .A0_f (new_AGEMA_signal_9279), .A1_t (new_AGEMA_signal_9280), .A1_f (new_AGEMA_signal_9281), .B0_t (Inst_bSbox_T16), .B0_f (new_AGEMA_signal_9783), .B1_t (new_AGEMA_signal_9784), .B1_f (new_AGEMA_signal_9785), .Z0_t (Inst_bSbox_T26), .Z0_f (new_AGEMA_signal_10286), .Z1_t (new_AGEMA_signal_10287), .Z1_f (new_AGEMA_signal_10288) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T27_U1 ( .A0_t (Inst_bSbox_T1), .A0_f (new_AGEMA_signal_9273), .A1_t (new_AGEMA_signal_9274), .A1_f (new_AGEMA_signal_9275), .B0_t (Inst_bSbox_T12), .B0_f (new_AGEMA_signal_9294), .B1_t (new_AGEMA_signal_9295), .B1_f (new_AGEMA_signal_9296), .Z0_t (Inst_bSbox_T27), .Z0_f (new_AGEMA_signal_9792), .Z1_t (new_AGEMA_signal_9793), .Z1_f (new_AGEMA_signal_9794) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M1_U1 ( .A0_t (Inst_bSbox_T13), .A0_f (new_AGEMA_signal_9777), .A1_t (new_AGEMA_signal_9778), .A1_f (new_AGEMA_signal_9779), .B0_t (Inst_bSbox_T6), .B0_f (new_AGEMA_signal_9771), .B1_t (new_AGEMA_signal_9772), .B1_f (new_AGEMA_signal_9773), .Z0_t (Inst_bSbox_M1), .Z0_f (new_AGEMA_signal_10289), .Z1_t (new_AGEMA_signal_10290), .Z1_f (new_AGEMA_signal_10291) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M2_U1 ( .A0_t (Inst_bSbox_T23), .A0_f (new_AGEMA_signal_10283), .A1_t (new_AGEMA_signal_10284), .A1_f (new_AGEMA_signal_10285), .B0_t (Inst_bSbox_T8), .B0_f (new_AGEMA_signal_10268), .B1_t (new_AGEMA_signal_10269), .B1_f (new_AGEMA_signal_10270), .Z0_t (Inst_bSbox_M2), .Z0_f (new_AGEMA_signal_10409), .Z1_t (new_AGEMA_signal_10410), .Z1_f (new_AGEMA_signal_10411) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M3_U1 ( .A0_t (Inst_bSbox_T14), .A0_f (new_AGEMA_signal_10274), .A1_t (new_AGEMA_signal_10275), .A1_f (new_AGEMA_signal_10276), .B0_t (Inst_bSbox_M1), .B0_f (new_AGEMA_signal_10289), .B1_t (new_AGEMA_signal_10290), .B1_f (new_AGEMA_signal_10291), .Z0_t (Inst_bSbox_M3), .Z0_f (new_AGEMA_signal_10412), .Z1_t (new_AGEMA_signal_10413), .Z1_f (new_AGEMA_signal_10414) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M4_U1 ( .A0_t (Inst_bSbox_T19), .A0_f (new_AGEMA_signal_9786), .A1_t (new_AGEMA_signal_9787), .A1_f (new_AGEMA_signal_9788), .B0_t (SboxIn[0]), .B0_f (new_AGEMA_signal_8115), .B1_t (new_AGEMA_signal_8116), .B1_f (new_AGEMA_signal_8117), .Z0_t (Inst_bSbox_M4), .Z0_f (new_AGEMA_signal_10292), .Z1_t (new_AGEMA_signal_10293), .Z1_f (new_AGEMA_signal_10294) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M5_U1 ( .A0_t (Inst_bSbox_M4), .A0_f (new_AGEMA_signal_10292), .A1_t (new_AGEMA_signal_10293), .A1_f (new_AGEMA_signal_10294), .B0_t (Inst_bSbox_M1), .B0_f (new_AGEMA_signal_10289), .B1_t (new_AGEMA_signal_10290), .B1_f (new_AGEMA_signal_10291), .Z0_t (Inst_bSbox_M5), .Z0_f (new_AGEMA_signal_10415), .Z1_t (new_AGEMA_signal_10416), .Z1_f (new_AGEMA_signal_10417) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M6_U1 ( .A0_t (Inst_bSbox_T3), .A0_f (new_AGEMA_signal_9279), .A1_t (new_AGEMA_signal_9280), .A1_f (new_AGEMA_signal_9281), .B0_t (Inst_bSbox_T16), .B0_f (new_AGEMA_signal_9783), .B1_t (new_AGEMA_signal_9784), .B1_f (new_AGEMA_signal_9785), .Z0_t (Inst_bSbox_M6), .Z0_f (new_AGEMA_signal_10295), .Z1_t (new_AGEMA_signal_10296), .Z1_f (new_AGEMA_signal_10297) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M7_U1 ( .A0_t (Inst_bSbox_T22), .A0_f (new_AGEMA_signal_9789), .A1_t (new_AGEMA_signal_9790), .A1_f (new_AGEMA_signal_9791), .B0_t (Inst_bSbox_T9), .B0_f (new_AGEMA_signal_9774), .B1_t (new_AGEMA_signal_9775), .B1_f (new_AGEMA_signal_9776), .Z0_t (Inst_bSbox_M7), .Z0_f (new_AGEMA_signal_10298), .Z1_t (new_AGEMA_signal_10299), .Z1_f (new_AGEMA_signal_10300) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M8_U1 ( .A0_t (Inst_bSbox_T26), .A0_f (new_AGEMA_signal_10286), .A1_t (new_AGEMA_signal_10287), .A1_f (new_AGEMA_signal_10288), .B0_t (Inst_bSbox_M6), .B0_f (new_AGEMA_signal_10295), .B1_t (new_AGEMA_signal_10296), .B1_f (new_AGEMA_signal_10297), .Z0_t (Inst_bSbox_M8), .Z0_f (new_AGEMA_signal_10418), .Z1_t (new_AGEMA_signal_10419), .Z1_f (new_AGEMA_signal_10420) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M9_U1 ( .A0_t (Inst_bSbox_T20), .A0_f (new_AGEMA_signal_10280), .A1_t (new_AGEMA_signal_10281), .A1_f (new_AGEMA_signal_10282), .B0_t (Inst_bSbox_T17), .B0_f (new_AGEMA_signal_10277), .B1_t (new_AGEMA_signal_10278), .B1_f (new_AGEMA_signal_10279), .Z0_t (Inst_bSbox_M9), .Z0_f (new_AGEMA_signal_10421), .Z1_t (new_AGEMA_signal_10422), .Z1_f (new_AGEMA_signal_10423) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M10_U1 ( .A0_t (Inst_bSbox_M9), .A0_f (new_AGEMA_signal_10421), .A1_t (new_AGEMA_signal_10422), .A1_f (new_AGEMA_signal_10423), .B0_t (Inst_bSbox_M6), .B0_f (new_AGEMA_signal_10295), .B1_t (new_AGEMA_signal_10296), .B1_f (new_AGEMA_signal_10297), .Z0_t (Inst_bSbox_M10), .Z0_f (new_AGEMA_signal_10526), .Z1_t (new_AGEMA_signal_10527), .Z1_f (new_AGEMA_signal_10528) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M11_U1 ( .A0_t (Inst_bSbox_T1), .A0_f (new_AGEMA_signal_9273), .A1_t (new_AGEMA_signal_9274), .A1_f (new_AGEMA_signal_9275), .B0_t (Inst_bSbox_T15), .B0_f (new_AGEMA_signal_9780), .B1_t (new_AGEMA_signal_9781), .B1_f (new_AGEMA_signal_9782), .Z0_t (Inst_bSbox_M11), .Z0_f (new_AGEMA_signal_10301), .Z1_t (new_AGEMA_signal_10302), .Z1_f (new_AGEMA_signal_10303) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M12_U1 ( .A0_t (Inst_bSbox_T4), .A0_f (new_AGEMA_signal_9282), .A1_t (new_AGEMA_signal_9283), .A1_f (new_AGEMA_signal_9284), .B0_t (Inst_bSbox_T27), .B0_f (new_AGEMA_signal_9792), .B1_t (new_AGEMA_signal_9793), .B1_f (new_AGEMA_signal_9794), .Z0_t (Inst_bSbox_M12), .Z0_f (new_AGEMA_signal_10304), .Z1_t (new_AGEMA_signal_10305), .Z1_f (new_AGEMA_signal_10306) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M13_U1 ( .A0_t (Inst_bSbox_M12), .A0_f (new_AGEMA_signal_10304), .A1_t (new_AGEMA_signal_10305), .A1_f (new_AGEMA_signal_10306), .B0_t (Inst_bSbox_M11), .B0_f (new_AGEMA_signal_10301), .B1_t (new_AGEMA_signal_10302), .B1_f (new_AGEMA_signal_10303), .Z0_t (Inst_bSbox_M13), .Z0_f (new_AGEMA_signal_10424), .Z1_t (new_AGEMA_signal_10425), .Z1_f (new_AGEMA_signal_10426) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M14_U1 ( .A0_t (Inst_bSbox_T2), .A0_f (new_AGEMA_signal_9276), .A1_t (new_AGEMA_signal_9277), .A1_f (new_AGEMA_signal_9278), .B0_t (Inst_bSbox_T10), .B0_f (new_AGEMA_signal_10271), .B1_t (new_AGEMA_signal_10272), .B1_f (new_AGEMA_signal_10273), .Z0_t (Inst_bSbox_M14), .Z0_f (new_AGEMA_signal_10427), .Z1_t (new_AGEMA_signal_10428), .Z1_f (new_AGEMA_signal_10429) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M15_U1 ( .A0_t (Inst_bSbox_M14), .A0_f (new_AGEMA_signal_10427), .A1_t (new_AGEMA_signal_10428), .A1_f (new_AGEMA_signal_10429), .B0_t (Inst_bSbox_M11), .B0_f (new_AGEMA_signal_10301), .B1_t (new_AGEMA_signal_10302), .B1_f (new_AGEMA_signal_10303), .Z0_t (Inst_bSbox_M15), .Z0_f (new_AGEMA_signal_10529), .Z1_t (new_AGEMA_signal_10530), .Z1_f (new_AGEMA_signal_10531) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M16_U1 ( .A0_t (Inst_bSbox_M3), .A0_f (new_AGEMA_signal_10412), .A1_t (new_AGEMA_signal_10413), .A1_f (new_AGEMA_signal_10414), .B0_t (Inst_bSbox_M2), .B0_f (new_AGEMA_signal_10409), .B1_t (new_AGEMA_signal_10410), .B1_f (new_AGEMA_signal_10411), .Z0_t (Inst_bSbox_M16), .Z0_f (new_AGEMA_signal_10532), .Z1_t (new_AGEMA_signal_10533), .Z1_f (new_AGEMA_signal_10534) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M17_U1 ( .A0_t (Inst_bSbox_M5), .A0_f (new_AGEMA_signal_10415), .A1_t (new_AGEMA_signal_10416), .A1_f (new_AGEMA_signal_10417), .B0_t (Inst_bSbox_T24), .B0_f (new_AGEMA_signal_10403), .B1_t (new_AGEMA_signal_10404), .B1_f (new_AGEMA_signal_10405), .Z0_t (Inst_bSbox_M17), .Z0_f (new_AGEMA_signal_10535), .Z1_t (new_AGEMA_signal_10536), .Z1_f (new_AGEMA_signal_10537) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M18_U1 ( .A0_t (Inst_bSbox_M8), .A0_f (new_AGEMA_signal_10418), .A1_t (new_AGEMA_signal_10419), .A1_f (new_AGEMA_signal_10420), .B0_t (Inst_bSbox_M7), .B0_f (new_AGEMA_signal_10298), .B1_t (new_AGEMA_signal_10299), .B1_f (new_AGEMA_signal_10300), .Z0_t (Inst_bSbox_M18), .Z0_f (new_AGEMA_signal_10538), .Z1_t (new_AGEMA_signal_10539), .Z1_f (new_AGEMA_signal_10540) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M19_U1 ( .A0_t (Inst_bSbox_M10), .A0_f (new_AGEMA_signal_10526), .A1_t (new_AGEMA_signal_10527), .A1_f (new_AGEMA_signal_10528), .B0_t (Inst_bSbox_M15), .B0_f (new_AGEMA_signal_10529), .B1_t (new_AGEMA_signal_10530), .B1_f (new_AGEMA_signal_10531), .Z0_t (Inst_bSbox_M19), .Z0_f (new_AGEMA_signal_10682), .Z1_t (new_AGEMA_signal_10683), .Z1_f (new_AGEMA_signal_10684) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M20_U1 ( .A0_t (Inst_bSbox_M16), .A0_f (new_AGEMA_signal_10532), .A1_t (new_AGEMA_signal_10533), .A1_f (new_AGEMA_signal_10534), .B0_t (Inst_bSbox_M13), .B0_f (new_AGEMA_signal_10424), .B1_t (new_AGEMA_signal_10425), .B1_f (new_AGEMA_signal_10426), .Z0_t (Inst_bSbox_M20), .Z0_f (new_AGEMA_signal_10685), .Z1_t (new_AGEMA_signal_10686), .Z1_f (new_AGEMA_signal_10687) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M21_U1 ( .A0_t (Inst_bSbox_M17), .A0_f (new_AGEMA_signal_10535), .A1_t (new_AGEMA_signal_10536), .A1_f (new_AGEMA_signal_10537), .B0_t (Inst_bSbox_M15), .B0_f (new_AGEMA_signal_10529), .B1_t (new_AGEMA_signal_10530), .B1_f (new_AGEMA_signal_10531), .Z0_t (Inst_bSbox_M21), .Z0_f (new_AGEMA_signal_10688), .Z1_t (new_AGEMA_signal_10689), .Z1_f (new_AGEMA_signal_10690) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M22_U1 ( .A0_t (Inst_bSbox_M18), .A0_f (new_AGEMA_signal_10538), .A1_t (new_AGEMA_signal_10539), .A1_f (new_AGEMA_signal_10540), .B0_t (Inst_bSbox_M13), .B0_f (new_AGEMA_signal_10424), .B1_t (new_AGEMA_signal_10425), .B1_f (new_AGEMA_signal_10426), .Z0_t (Inst_bSbox_M22), .Z0_f (new_AGEMA_signal_10691), .Z1_t (new_AGEMA_signal_10692), .Z1_f (new_AGEMA_signal_10693) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M23_U1 ( .A0_t (Inst_bSbox_M19), .A0_f (new_AGEMA_signal_10682), .A1_t (new_AGEMA_signal_10683), .A1_f (new_AGEMA_signal_10684), .B0_t (Inst_bSbox_T25), .B0_f (new_AGEMA_signal_10406), .B1_t (new_AGEMA_signal_10407), .B1_f (new_AGEMA_signal_10408), .Z0_t (Inst_bSbox_M23), .Z0_f (new_AGEMA_signal_10817), .Z1_t (new_AGEMA_signal_10818), .Z1_f (new_AGEMA_signal_10819) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M24_U1 ( .A0_t (Inst_bSbox_M22), .A0_f (new_AGEMA_signal_10691), .A1_t (new_AGEMA_signal_10692), .A1_f (new_AGEMA_signal_10693), .B0_t (Inst_bSbox_M23), .B0_f (new_AGEMA_signal_10817), .B1_t (new_AGEMA_signal_10818), .B1_f (new_AGEMA_signal_10819), .Z0_t (Inst_bSbox_M24), .Z0_f (new_AGEMA_signal_10925), .Z1_t (new_AGEMA_signal_10926), .Z1_f (new_AGEMA_signal_10927) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M25_U1 ( .A0_t (Inst_bSbox_M22), .A0_f (new_AGEMA_signal_10691), .A1_t (new_AGEMA_signal_10692), .A1_f (new_AGEMA_signal_10693), .B0_t (Inst_bSbox_M20), .B0_f (new_AGEMA_signal_10685), .B1_t (new_AGEMA_signal_10686), .B1_f (new_AGEMA_signal_10687), .Z0_t (Inst_bSbox_M25), .Z0_f (new_AGEMA_signal_10820), .Z1_t (new_AGEMA_signal_10821), .Z1_f (new_AGEMA_signal_10822) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M26_U1 ( .A0_t (Inst_bSbox_M21), .A0_f (new_AGEMA_signal_10688), .A1_t (new_AGEMA_signal_10689), .A1_f (new_AGEMA_signal_10690), .B0_t (Inst_bSbox_M25), .B0_f (new_AGEMA_signal_10820), .B1_t (new_AGEMA_signal_10821), .B1_f (new_AGEMA_signal_10822), .Z0_t (Inst_bSbox_M26), .Z0_f (new_AGEMA_signal_10928), .Z1_t (new_AGEMA_signal_10929), .Z1_f (new_AGEMA_signal_10930) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M27_U1 ( .A0_t (Inst_bSbox_M20), .A0_f (new_AGEMA_signal_10685), .A1_t (new_AGEMA_signal_10686), .A1_f (new_AGEMA_signal_10687), .B0_t (Inst_bSbox_M21), .B0_f (new_AGEMA_signal_10688), .B1_t (new_AGEMA_signal_10689), .B1_f (new_AGEMA_signal_10690), .Z0_t (Inst_bSbox_M27), .Z0_f (new_AGEMA_signal_10823), .Z1_t (new_AGEMA_signal_10824), .Z1_f (new_AGEMA_signal_10825) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M28_U1 ( .A0_t (Inst_bSbox_M23), .A0_f (new_AGEMA_signal_10817), .A1_t (new_AGEMA_signal_10818), .A1_f (new_AGEMA_signal_10819), .B0_t (Inst_bSbox_M25), .B0_f (new_AGEMA_signal_10820), .B1_t (new_AGEMA_signal_10821), .B1_f (new_AGEMA_signal_10822), .Z0_t (Inst_bSbox_M28), .Z0_f (new_AGEMA_signal_10931), .Z1_t (new_AGEMA_signal_10932), .Z1_f (new_AGEMA_signal_10933) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M29_U1 ( .A0_t (Inst_bSbox_M28), .A0_f (new_AGEMA_signal_10931), .A1_t (new_AGEMA_signal_10932), .A1_f (new_AGEMA_signal_10933), .B0_t (Inst_bSbox_M27), .B0_f (new_AGEMA_signal_10823), .B1_t (new_AGEMA_signal_10824), .B1_f (new_AGEMA_signal_10825), .Z0_t (Inst_bSbox_M29), .Z0_f (new_AGEMA_signal_11036), .Z1_t (new_AGEMA_signal_11037), .Z1_f (new_AGEMA_signal_11038) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M30_U1 ( .A0_t (Inst_bSbox_M26), .A0_f (new_AGEMA_signal_10928), .A1_t (new_AGEMA_signal_10929), .A1_f (new_AGEMA_signal_10930), .B0_t (Inst_bSbox_M24), .B0_f (new_AGEMA_signal_10925), .B1_t (new_AGEMA_signal_10926), .B1_f (new_AGEMA_signal_10927), .Z0_t (Inst_bSbox_M30), .Z0_f (new_AGEMA_signal_11039), .Z1_t (new_AGEMA_signal_11040), .Z1_f (new_AGEMA_signal_11041) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M31_U1 ( .A0_t (Inst_bSbox_M20), .A0_f (new_AGEMA_signal_10685), .A1_t (new_AGEMA_signal_10686), .A1_f (new_AGEMA_signal_10687), .B0_t (Inst_bSbox_M23), .B0_f (new_AGEMA_signal_10817), .B1_t (new_AGEMA_signal_10818), .B1_f (new_AGEMA_signal_10819), .Z0_t (Inst_bSbox_M31), .Z0_f (new_AGEMA_signal_10934), .Z1_t (new_AGEMA_signal_10935), .Z1_f (new_AGEMA_signal_10936) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M32_U1 ( .A0_t (Inst_bSbox_M27), .A0_f (new_AGEMA_signal_10823), .A1_t (new_AGEMA_signal_10824), .A1_f (new_AGEMA_signal_10825), .B0_t (Inst_bSbox_M31), .B0_f (new_AGEMA_signal_10934), .B1_t (new_AGEMA_signal_10935), .B1_f (new_AGEMA_signal_10936), .Z0_t (Inst_bSbox_M32), .Z0_f (new_AGEMA_signal_11042), .Z1_t (new_AGEMA_signal_11043), .Z1_f (new_AGEMA_signal_11044) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M33_U1 ( .A0_t (Inst_bSbox_M27), .A0_f (new_AGEMA_signal_10823), .A1_t (new_AGEMA_signal_10824), .A1_f (new_AGEMA_signal_10825), .B0_t (Inst_bSbox_M25), .B0_f (new_AGEMA_signal_10820), .B1_t (new_AGEMA_signal_10821), .B1_f (new_AGEMA_signal_10822), .Z0_t (Inst_bSbox_M33), .Z0_f (new_AGEMA_signal_10937), .Z1_t (new_AGEMA_signal_10938), .Z1_f (new_AGEMA_signal_10939) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M34_U1 ( .A0_t (Inst_bSbox_M21), .A0_f (new_AGEMA_signal_10688), .A1_t (new_AGEMA_signal_10689), .A1_f (new_AGEMA_signal_10690), .B0_t (Inst_bSbox_M22), .B0_f (new_AGEMA_signal_10691), .B1_t (new_AGEMA_signal_10692), .B1_f (new_AGEMA_signal_10693), .Z0_t (Inst_bSbox_M34), .Z0_f (new_AGEMA_signal_10826), .Z1_t (new_AGEMA_signal_10827), .Z1_f (new_AGEMA_signal_10828) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M35_U1 ( .A0_t (Inst_bSbox_M24), .A0_f (new_AGEMA_signal_10925), .A1_t (new_AGEMA_signal_10926), .A1_f (new_AGEMA_signal_10927), .B0_t (Inst_bSbox_M34), .B0_f (new_AGEMA_signal_10826), .B1_t (new_AGEMA_signal_10827), .B1_f (new_AGEMA_signal_10828), .Z0_t (Inst_bSbox_M35), .Z0_f (new_AGEMA_signal_11045), .Z1_t (new_AGEMA_signal_11046), .Z1_f (new_AGEMA_signal_11047) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M36_U1 ( .A0_t (Inst_bSbox_M24), .A0_f (new_AGEMA_signal_10925), .A1_t (new_AGEMA_signal_10926), .A1_f (new_AGEMA_signal_10927), .B0_t (Inst_bSbox_M25), .B0_f (new_AGEMA_signal_10820), .B1_t (new_AGEMA_signal_10821), .B1_f (new_AGEMA_signal_10822), .Z0_t (Inst_bSbox_M36), .Z0_f (new_AGEMA_signal_11048), .Z1_t (new_AGEMA_signal_11049), .Z1_f (new_AGEMA_signal_11050) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M37_U1 ( .A0_t (Inst_bSbox_M21), .A0_f (new_AGEMA_signal_10688), .A1_t (new_AGEMA_signal_10689), .A1_f (new_AGEMA_signal_10690), .B0_t (Inst_bSbox_M29), .B0_f (new_AGEMA_signal_11036), .B1_t (new_AGEMA_signal_11037), .B1_f (new_AGEMA_signal_11038), .Z0_t (Inst_bSbox_M37), .Z0_f (new_AGEMA_signal_11123), .Z1_t (new_AGEMA_signal_11124), .Z1_f (new_AGEMA_signal_11125) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M38_U1 ( .A0_t (Inst_bSbox_M32), .A0_f (new_AGEMA_signal_11042), .A1_t (new_AGEMA_signal_11043), .A1_f (new_AGEMA_signal_11044), .B0_t (Inst_bSbox_M33), .B0_f (new_AGEMA_signal_10937), .B1_t (new_AGEMA_signal_10938), .B1_f (new_AGEMA_signal_10939), .Z0_t (Inst_bSbox_M38), .Z0_f (new_AGEMA_signal_11126), .Z1_t (new_AGEMA_signal_11127), .Z1_f (new_AGEMA_signal_11128) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M39_U1 ( .A0_t (Inst_bSbox_M23), .A0_f (new_AGEMA_signal_10817), .A1_t (new_AGEMA_signal_10818), .A1_f (new_AGEMA_signal_10819), .B0_t (Inst_bSbox_M30), .B0_f (new_AGEMA_signal_11039), .B1_t (new_AGEMA_signal_11040), .B1_f (new_AGEMA_signal_11041), .Z0_t (Inst_bSbox_M39), .Z0_f (new_AGEMA_signal_11129), .Z1_t (new_AGEMA_signal_11130), .Z1_f (new_AGEMA_signal_11131) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M40_U1 ( .A0_t (Inst_bSbox_M35), .A0_f (new_AGEMA_signal_11045), .A1_t (new_AGEMA_signal_11046), .A1_f (new_AGEMA_signal_11047), .B0_t (Inst_bSbox_M36), .B0_f (new_AGEMA_signal_11048), .B1_t (new_AGEMA_signal_11049), .B1_f (new_AGEMA_signal_11050), .Z0_t (Inst_bSbox_M40), .Z0_f (new_AGEMA_signal_11132), .Z1_t (new_AGEMA_signal_11133), .Z1_f (new_AGEMA_signal_11134) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M41_U1 ( .A0_t (Inst_bSbox_M38), .A0_f (new_AGEMA_signal_11126), .A1_t (new_AGEMA_signal_11127), .A1_f (new_AGEMA_signal_11128), .B0_t (Inst_bSbox_M40), .B0_f (new_AGEMA_signal_11132), .B1_t (new_AGEMA_signal_11133), .B1_f (new_AGEMA_signal_11134), .Z0_t (Inst_bSbox_M41), .Z0_f (new_AGEMA_signal_11162), .Z1_t (new_AGEMA_signal_11163), .Z1_f (new_AGEMA_signal_11164) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M42_U1 ( .A0_t (Inst_bSbox_M37), .A0_f (new_AGEMA_signal_11123), .A1_t (new_AGEMA_signal_11124), .A1_f (new_AGEMA_signal_11125), .B0_t (Inst_bSbox_M39), .B0_f (new_AGEMA_signal_11129), .B1_t (new_AGEMA_signal_11130), .B1_f (new_AGEMA_signal_11131), .Z0_t (Inst_bSbox_M42), .Z0_f (new_AGEMA_signal_11165), .Z1_t (new_AGEMA_signal_11166), .Z1_f (new_AGEMA_signal_11167) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M43_U1 ( .A0_t (Inst_bSbox_M37), .A0_f (new_AGEMA_signal_11123), .A1_t (new_AGEMA_signal_11124), .A1_f (new_AGEMA_signal_11125), .B0_t (Inst_bSbox_M38), .B0_f (new_AGEMA_signal_11126), .B1_t (new_AGEMA_signal_11127), .B1_f (new_AGEMA_signal_11128), .Z0_t (Inst_bSbox_M43), .Z0_f (new_AGEMA_signal_11168), .Z1_t (new_AGEMA_signal_11169), .Z1_f (new_AGEMA_signal_11170) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M44_U1 ( .A0_t (Inst_bSbox_M39), .A0_f (new_AGEMA_signal_11129), .A1_t (new_AGEMA_signal_11130), .A1_f (new_AGEMA_signal_11131), .B0_t (Inst_bSbox_M40), .B0_f (new_AGEMA_signal_11132), .B1_t (new_AGEMA_signal_11133), .B1_f (new_AGEMA_signal_11134), .Z0_t (Inst_bSbox_M44), .Z0_f (new_AGEMA_signal_11171), .Z1_t (new_AGEMA_signal_11172), .Z1_f (new_AGEMA_signal_11173) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M45_U1 ( .A0_t (Inst_bSbox_M42), .A0_f (new_AGEMA_signal_11165), .A1_t (new_AGEMA_signal_11166), .A1_f (new_AGEMA_signal_11167), .B0_t (Inst_bSbox_M41), .B0_f (new_AGEMA_signal_11162), .B1_t (new_AGEMA_signal_11163), .B1_f (new_AGEMA_signal_11164), .Z0_t (Inst_bSbox_M45), .Z0_f (new_AGEMA_signal_11198), .Z1_t (new_AGEMA_signal_11199), .Z1_f (new_AGEMA_signal_11200) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M46_U1 ( .A0_t (Inst_bSbox_M44), .A0_f (new_AGEMA_signal_11171), .A1_t (new_AGEMA_signal_11172), .A1_f (new_AGEMA_signal_11173), .B0_t (Inst_bSbox_T6), .B0_f (new_AGEMA_signal_9771), .B1_t (new_AGEMA_signal_9772), .B1_f (new_AGEMA_signal_9773), .Z0_t (Inst_bSbox_M46), .Z0_f (new_AGEMA_signal_11201), .Z1_t (new_AGEMA_signal_11202), .Z1_f (new_AGEMA_signal_11203) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M47_U1 ( .A0_t (Inst_bSbox_M40), .A0_f (new_AGEMA_signal_11132), .A1_t (new_AGEMA_signal_11133), .A1_f (new_AGEMA_signal_11134), .B0_t (Inst_bSbox_T8), .B0_f (new_AGEMA_signal_10268), .B1_t (new_AGEMA_signal_10269), .B1_f (new_AGEMA_signal_10270), .Z0_t (Inst_bSbox_M47), .Z0_f (new_AGEMA_signal_11174), .Z1_t (new_AGEMA_signal_11175), .Z1_f (new_AGEMA_signal_11176) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M48_U1 ( .A0_t (Inst_bSbox_M39), .A0_f (new_AGEMA_signal_11129), .A1_t (new_AGEMA_signal_11130), .A1_f (new_AGEMA_signal_11131), .B0_t (SboxIn[0]), .B0_f (new_AGEMA_signal_8115), .B1_t (new_AGEMA_signal_8116), .B1_f (new_AGEMA_signal_8117), .Z0_t (Inst_bSbox_M48), .Z0_f (new_AGEMA_signal_11177), .Z1_t (new_AGEMA_signal_11178), .Z1_f (new_AGEMA_signal_11179) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M49_U1 ( .A0_t (Inst_bSbox_M43), .A0_f (new_AGEMA_signal_11168), .A1_t (new_AGEMA_signal_11169), .A1_f (new_AGEMA_signal_11170), .B0_t (Inst_bSbox_T16), .B0_f (new_AGEMA_signal_9783), .B1_t (new_AGEMA_signal_9784), .B1_f (new_AGEMA_signal_9785), .Z0_t (Inst_bSbox_M49), .Z0_f (new_AGEMA_signal_11204), .Z1_t (new_AGEMA_signal_11205), .Z1_f (new_AGEMA_signal_11206) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M50_U1 ( .A0_t (Inst_bSbox_M38), .A0_f (new_AGEMA_signal_11126), .A1_t (new_AGEMA_signal_11127), .A1_f (new_AGEMA_signal_11128), .B0_t (Inst_bSbox_T9), .B0_f (new_AGEMA_signal_9774), .B1_t (new_AGEMA_signal_9775), .B1_f (new_AGEMA_signal_9776), .Z0_t (Inst_bSbox_M50), .Z0_f (new_AGEMA_signal_11180), .Z1_t (new_AGEMA_signal_11181), .Z1_f (new_AGEMA_signal_11182) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M51_U1 ( .A0_t (Inst_bSbox_M37), .A0_f (new_AGEMA_signal_11123), .A1_t (new_AGEMA_signal_11124), .A1_f (new_AGEMA_signal_11125), .B0_t (Inst_bSbox_T17), .B0_f (new_AGEMA_signal_10277), .B1_t (new_AGEMA_signal_10278), .B1_f (new_AGEMA_signal_10279), .Z0_t (Inst_bSbox_M51), .Z0_f (new_AGEMA_signal_11183), .Z1_t (new_AGEMA_signal_11184), .Z1_f (new_AGEMA_signal_11185) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M52_U1 ( .A0_t (Inst_bSbox_M42), .A0_f (new_AGEMA_signal_11165), .A1_t (new_AGEMA_signal_11166), .A1_f (new_AGEMA_signal_11167), .B0_t (Inst_bSbox_T15), .B0_f (new_AGEMA_signal_9780), .B1_t (new_AGEMA_signal_9781), .B1_f (new_AGEMA_signal_9782), .Z0_t (Inst_bSbox_M52), .Z0_f (new_AGEMA_signal_11207), .Z1_t (new_AGEMA_signal_11208), .Z1_f (new_AGEMA_signal_11209) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M53_U1 ( .A0_t (Inst_bSbox_M45), .A0_f (new_AGEMA_signal_11198), .A1_t (new_AGEMA_signal_11199), .A1_f (new_AGEMA_signal_11200), .B0_t (Inst_bSbox_T27), .B0_f (new_AGEMA_signal_9792), .B1_t (new_AGEMA_signal_9793), .B1_f (new_AGEMA_signal_9794), .Z0_t (Inst_bSbox_M53), .Z0_f (new_AGEMA_signal_11234), .Z1_t (new_AGEMA_signal_11235), .Z1_f (new_AGEMA_signal_11236) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M54_U1 ( .A0_t (Inst_bSbox_M41), .A0_f (new_AGEMA_signal_11162), .A1_t (new_AGEMA_signal_11163), .A1_f (new_AGEMA_signal_11164), .B0_t (Inst_bSbox_T10), .B0_f (new_AGEMA_signal_10271), .B1_t (new_AGEMA_signal_10272), .B1_f (new_AGEMA_signal_10273), .Z0_t (Inst_bSbox_M54), .Z0_f (new_AGEMA_signal_11210), .Z1_t (new_AGEMA_signal_11211), .Z1_f (new_AGEMA_signal_11212) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M55_U1 ( .A0_t (Inst_bSbox_M44), .A0_f (new_AGEMA_signal_11171), .A1_t (new_AGEMA_signal_11172), .A1_f (new_AGEMA_signal_11173), .B0_t (Inst_bSbox_T13), .B0_f (new_AGEMA_signal_9777), .B1_t (new_AGEMA_signal_9778), .B1_f (new_AGEMA_signal_9779), .Z0_t (Inst_bSbox_M55), .Z0_f (new_AGEMA_signal_11213), .Z1_t (new_AGEMA_signal_11214), .Z1_f (new_AGEMA_signal_11215) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M56_U1 ( .A0_t (Inst_bSbox_M40), .A0_f (new_AGEMA_signal_11132), .A1_t (new_AGEMA_signal_11133), .A1_f (new_AGEMA_signal_11134), .B0_t (Inst_bSbox_T23), .B0_f (new_AGEMA_signal_10283), .B1_t (new_AGEMA_signal_10284), .B1_f (new_AGEMA_signal_10285), .Z0_t (Inst_bSbox_M56), .Z0_f (new_AGEMA_signal_11186), .Z1_t (new_AGEMA_signal_11187), .Z1_f (new_AGEMA_signal_11188) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M57_U1 ( .A0_t (Inst_bSbox_M39), .A0_f (new_AGEMA_signal_11129), .A1_t (new_AGEMA_signal_11130), .A1_f (new_AGEMA_signal_11131), .B0_t (Inst_bSbox_T19), .B0_f (new_AGEMA_signal_9786), .B1_t (new_AGEMA_signal_9787), .B1_f (new_AGEMA_signal_9788), .Z0_t (Inst_bSbox_M57), .Z0_f (new_AGEMA_signal_11189), .Z1_t (new_AGEMA_signal_11190), .Z1_f (new_AGEMA_signal_11191) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M58_U1 ( .A0_t (Inst_bSbox_M43), .A0_f (new_AGEMA_signal_11168), .A1_t (new_AGEMA_signal_11169), .A1_f (new_AGEMA_signal_11170), .B0_t (Inst_bSbox_T3), .B0_f (new_AGEMA_signal_9279), .B1_t (new_AGEMA_signal_9280), .B1_f (new_AGEMA_signal_9281), .Z0_t (Inst_bSbox_M58), .Z0_f (new_AGEMA_signal_11216), .Z1_t (new_AGEMA_signal_11217), .Z1_f (new_AGEMA_signal_11218) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M59_U1 ( .A0_t (Inst_bSbox_M38), .A0_f (new_AGEMA_signal_11126), .A1_t (new_AGEMA_signal_11127), .A1_f (new_AGEMA_signal_11128), .B0_t (Inst_bSbox_T22), .B0_f (new_AGEMA_signal_9789), .B1_t (new_AGEMA_signal_9790), .B1_f (new_AGEMA_signal_9791), .Z0_t (Inst_bSbox_M59), .Z0_f (new_AGEMA_signal_11192), .Z1_t (new_AGEMA_signal_11193), .Z1_f (new_AGEMA_signal_11194) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M60_U1 ( .A0_t (Inst_bSbox_M37), .A0_f (new_AGEMA_signal_11123), .A1_t (new_AGEMA_signal_11124), .A1_f (new_AGEMA_signal_11125), .B0_t (Inst_bSbox_T20), .B0_f (new_AGEMA_signal_10280), .B1_t (new_AGEMA_signal_10281), .B1_f (new_AGEMA_signal_10282), .Z0_t (Inst_bSbox_M60), .Z0_f (new_AGEMA_signal_11195), .Z1_t (new_AGEMA_signal_11196), .Z1_f (new_AGEMA_signal_11197) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M61_U1 ( .A0_t (Inst_bSbox_M42), .A0_f (new_AGEMA_signal_11165), .A1_t (new_AGEMA_signal_11166), .A1_f (new_AGEMA_signal_11167), .B0_t (Inst_bSbox_T1), .B0_f (new_AGEMA_signal_9273), .B1_t (new_AGEMA_signal_9274), .B1_f (new_AGEMA_signal_9275), .Z0_t (Inst_bSbox_M61), .Z0_f (new_AGEMA_signal_11219), .Z1_t (new_AGEMA_signal_11220), .Z1_f (new_AGEMA_signal_11221) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M62_U1 ( .A0_t (Inst_bSbox_M45), .A0_f (new_AGEMA_signal_11198), .A1_t (new_AGEMA_signal_11199), .A1_f (new_AGEMA_signal_11200), .B0_t (Inst_bSbox_T4), .B0_f (new_AGEMA_signal_9282), .B1_t (new_AGEMA_signal_9283), .B1_f (new_AGEMA_signal_9284), .Z0_t (Inst_bSbox_M62), .Z0_f (new_AGEMA_signal_11237), .Z1_t (new_AGEMA_signal_11238), .Z1_f (new_AGEMA_signal_11239) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M63_U1 ( .A0_t (Inst_bSbox_M41), .A0_f (new_AGEMA_signal_11162), .A1_t (new_AGEMA_signal_11163), .A1_f (new_AGEMA_signal_11164), .B0_t (Inst_bSbox_T2), .B0_f (new_AGEMA_signal_9276), .B1_t (new_AGEMA_signal_9277), .B1_f (new_AGEMA_signal_9278), .Z0_t (Inst_bSbox_M63), .Z0_f (new_AGEMA_signal_11222), .Z1_t (new_AGEMA_signal_11223), .Z1_f (new_AGEMA_signal_11224) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L0_U1 ( .A0_t (Inst_bSbox_M61), .A0_f (new_AGEMA_signal_11219), .A1_t (new_AGEMA_signal_11220), .A1_f (new_AGEMA_signal_11221), .B0_t (Inst_bSbox_M62), .B0_f (new_AGEMA_signal_11237), .B1_t (new_AGEMA_signal_11238), .B1_f (new_AGEMA_signal_11239), .Z0_t (Inst_bSbox_L0), .Z0_f (new_AGEMA_signal_11264), .Z1_t (new_AGEMA_signal_11265), .Z1_f (new_AGEMA_signal_11266) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L1_U1 ( .A0_t (Inst_bSbox_M50), .A0_f (new_AGEMA_signal_11180), .A1_t (new_AGEMA_signal_11181), .A1_f (new_AGEMA_signal_11182), .B0_t (Inst_bSbox_M56), .B0_f (new_AGEMA_signal_11186), .B1_t (new_AGEMA_signal_11187), .B1_f (new_AGEMA_signal_11188), .Z0_t (Inst_bSbox_L1), .Z0_f (new_AGEMA_signal_11225), .Z1_t (new_AGEMA_signal_11226), .Z1_f (new_AGEMA_signal_11227) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L2_U1 ( .A0_t (Inst_bSbox_M46), .A0_f (new_AGEMA_signal_11201), .A1_t (new_AGEMA_signal_11202), .A1_f (new_AGEMA_signal_11203), .B0_t (Inst_bSbox_M48), .B0_f (new_AGEMA_signal_11177), .B1_t (new_AGEMA_signal_11178), .B1_f (new_AGEMA_signal_11179), .Z0_t (Inst_bSbox_L2), .Z0_f (new_AGEMA_signal_11240), .Z1_t (new_AGEMA_signal_11241), .Z1_f (new_AGEMA_signal_11242) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L3_U1 ( .A0_t (Inst_bSbox_M47), .A0_f (new_AGEMA_signal_11174), .A1_t (new_AGEMA_signal_11175), .A1_f (new_AGEMA_signal_11176), .B0_t (Inst_bSbox_M55), .B0_f (new_AGEMA_signal_11213), .B1_t (new_AGEMA_signal_11214), .B1_f (new_AGEMA_signal_11215), .Z0_t (Inst_bSbox_L3), .Z0_f (new_AGEMA_signal_11243), .Z1_t (new_AGEMA_signal_11244), .Z1_f (new_AGEMA_signal_11245) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L4_U1 ( .A0_t (Inst_bSbox_M54), .A0_f (new_AGEMA_signal_11210), .A1_t (new_AGEMA_signal_11211), .A1_f (new_AGEMA_signal_11212), .B0_t (Inst_bSbox_M58), .B0_f (new_AGEMA_signal_11216), .B1_t (new_AGEMA_signal_11217), .B1_f (new_AGEMA_signal_11218), .Z0_t (Inst_bSbox_L4), .Z0_f (new_AGEMA_signal_11246), .Z1_t (new_AGEMA_signal_11247), .Z1_f (new_AGEMA_signal_11248) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L5_U1 ( .A0_t (Inst_bSbox_M49), .A0_f (new_AGEMA_signal_11204), .A1_t (new_AGEMA_signal_11205), .A1_f (new_AGEMA_signal_11206), .B0_t (Inst_bSbox_M61), .B0_f (new_AGEMA_signal_11219), .B1_t (new_AGEMA_signal_11220), .B1_f (new_AGEMA_signal_11221), .Z0_t (Inst_bSbox_L5), .Z0_f (new_AGEMA_signal_11249), .Z1_t (new_AGEMA_signal_11250), .Z1_f (new_AGEMA_signal_11251) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L6_U1 ( .A0_t (Inst_bSbox_M62), .A0_f (new_AGEMA_signal_11237), .A1_t (new_AGEMA_signal_11238), .A1_f (new_AGEMA_signal_11239), .B0_t (Inst_bSbox_L5), .B0_f (new_AGEMA_signal_11249), .B1_t (new_AGEMA_signal_11250), .B1_f (new_AGEMA_signal_11251), .Z0_t (Inst_bSbox_L6), .Z0_f (new_AGEMA_signal_11267), .Z1_t (new_AGEMA_signal_11268), .Z1_f (new_AGEMA_signal_11269) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L7_U1 ( .A0_t (Inst_bSbox_M46), .A0_f (new_AGEMA_signal_11201), .A1_t (new_AGEMA_signal_11202), .A1_f (new_AGEMA_signal_11203), .B0_t (Inst_bSbox_L3), .B0_f (new_AGEMA_signal_11243), .B1_t (new_AGEMA_signal_11244), .B1_f (new_AGEMA_signal_11245), .Z0_t (Inst_bSbox_L7), .Z0_f (new_AGEMA_signal_11270), .Z1_t (new_AGEMA_signal_11271), .Z1_f (new_AGEMA_signal_11272) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L8_U1 ( .A0_t (Inst_bSbox_M51), .A0_f (new_AGEMA_signal_11183), .A1_t (new_AGEMA_signal_11184), .A1_f (new_AGEMA_signal_11185), .B0_t (Inst_bSbox_M59), .B0_f (new_AGEMA_signal_11192), .B1_t (new_AGEMA_signal_11193), .B1_f (new_AGEMA_signal_11194), .Z0_t (Inst_bSbox_L8), .Z0_f (new_AGEMA_signal_11228), .Z1_t (new_AGEMA_signal_11229), .Z1_f (new_AGEMA_signal_11230) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L9_U1 ( .A0_t (Inst_bSbox_M52), .A0_f (new_AGEMA_signal_11207), .A1_t (new_AGEMA_signal_11208), .A1_f (new_AGEMA_signal_11209), .B0_t (Inst_bSbox_M53), .B0_f (new_AGEMA_signal_11234), .B1_t (new_AGEMA_signal_11235), .B1_f (new_AGEMA_signal_11236), .Z0_t (Inst_bSbox_L9), .Z0_f (new_AGEMA_signal_11273), .Z1_t (new_AGEMA_signal_11274), .Z1_f (new_AGEMA_signal_11275) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L10_U1 ( .A0_t (Inst_bSbox_M53), .A0_f (new_AGEMA_signal_11234), .A1_t (new_AGEMA_signal_11235), .A1_f (new_AGEMA_signal_11236), .B0_t (Inst_bSbox_L4), .B0_f (new_AGEMA_signal_11246), .B1_t (new_AGEMA_signal_11247), .B1_f (new_AGEMA_signal_11248), .Z0_t (Inst_bSbox_L10), .Z0_f (new_AGEMA_signal_11276), .Z1_t (new_AGEMA_signal_11277), .Z1_f (new_AGEMA_signal_11278) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L11_U1 ( .A0_t (Inst_bSbox_M60), .A0_f (new_AGEMA_signal_11195), .A1_t (new_AGEMA_signal_11196), .A1_f (new_AGEMA_signal_11197), .B0_t (Inst_bSbox_L2), .B0_f (new_AGEMA_signal_11240), .B1_t (new_AGEMA_signal_11241), .B1_f (new_AGEMA_signal_11242), .Z0_t (Inst_bSbox_L11), .Z0_f (new_AGEMA_signal_11279), .Z1_t (new_AGEMA_signal_11280), .Z1_f (new_AGEMA_signal_11281) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L12_U1 ( .A0_t (Inst_bSbox_M48), .A0_f (new_AGEMA_signal_11177), .A1_t (new_AGEMA_signal_11178), .A1_f (new_AGEMA_signal_11179), .B0_t (Inst_bSbox_M51), .B0_f (new_AGEMA_signal_11183), .B1_t (new_AGEMA_signal_11184), .B1_f (new_AGEMA_signal_11185), .Z0_t (Inst_bSbox_L12), .Z0_f (new_AGEMA_signal_11231), .Z1_t (new_AGEMA_signal_11232), .Z1_f (new_AGEMA_signal_11233) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L13_U1 ( .A0_t (Inst_bSbox_M50), .A0_f (new_AGEMA_signal_11180), .A1_t (new_AGEMA_signal_11181), .A1_f (new_AGEMA_signal_11182), .B0_t (Inst_bSbox_L0), .B0_f (new_AGEMA_signal_11264), .B1_t (new_AGEMA_signal_11265), .B1_f (new_AGEMA_signal_11266), .Z0_t (Inst_bSbox_L13), .Z0_f (new_AGEMA_signal_11291), .Z1_t (new_AGEMA_signal_11292), .Z1_f (new_AGEMA_signal_11293) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L14_U1 ( .A0_t (Inst_bSbox_M52), .A0_f (new_AGEMA_signal_11207), .A1_t (new_AGEMA_signal_11208), .A1_f (new_AGEMA_signal_11209), .B0_t (Inst_bSbox_M61), .B0_f (new_AGEMA_signal_11219), .B1_t (new_AGEMA_signal_11220), .B1_f (new_AGEMA_signal_11221), .Z0_t (Inst_bSbox_L14), .Z0_f (new_AGEMA_signal_11252), .Z1_t (new_AGEMA_signal_11253), .Z1_f (new_AGEMA_signal_11254) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L15_U1 ( .A0_t (Inst_bSbox_M55), .A0_f (new_AGEMA_signal_11213), .A1_t (new_AGEMA_signal_11214), .A1_f (new_AGEMA_signal_11215), .B0_t (Inst_bSbox_L1), .B0_f (new_AGEMA_signal_11225), .B1_t (new_AGEMA_signal_11226), .B1_f (new_AGEMA_signal_11227), .Z0_t (Inst_bSbox_L15), .Z0_f (new_AGEMA_signal_11255), .Z1_t (new_AGEMA_signal_11256), .Z1_f (new_AGEMA_signal_11257) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L16_U1 ( .A0_t (Inst_bSbox_M56), .A0_f (new_AGEMA_signal_11186), .A1_t (new_AGEMA_signal_11187), .A1_f (new_AGEMA_signal_11188), .B0_t (Inst_bSbox_L0), .B0_f (new_AGEMA_signal_11264), .B1_t (new_AGEMA_signal_11265), .B1_f (new_AGEMA_signal_11266), .Z0_t (Inst_bSbox_L16), .Z0_f (new_AGEMA_signal_11294), .Z1_t (new_AGEMA_signal_11295), .Z1_f (new_AGEMA_signal_11296) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L17_U1 ( .A0_t (Inst_bSbox_M57), .A0_f (new_AGEMA_signal_11189), .A1_t (new_AGEMA_signal_11190), .A1_f (new_AGEMA_signal_11191), .B0_t (Inst_bSbox_L1), .B0_f (new_AGEMA_signal_11225), .B1_t (new_AGEMA_signal_11226), .B1_f (new_AGEMA_signal_11227), .Z0_t (Inst_bSbox_L17), .Z0_f (new_AGEMA_signal_11258), .Z1_t (new_AGEMA_signal_11259), .Z1_f (new_AGEMA_signal_11260) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L18_U1 ( .A0_t (Inst_bSbox_M58), .A0_f (new_AGEMA_signal_11216), .A1_t (new_AGEMA_signal_11217), .A1_f (new_AGEMA_signal_11218), .B0_t (Inst_bSbox_L8), .B0_f (new_AGEMA_signal_11228), .B1_t (new_AGEMA_signal_11229), .B1_f (new_AGEMA_signal_11230), .Z0_t (Inst_bSbox_L18), .Z0_f (new_AGEMA_signal_11261), .Z1_t (new_AGEMA_signal_11262), .Z1_f (new_AGEMA_signal_11263) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L19_U1 ( .A0_t (Inst_bSbox_M63), .A0_f (new_AGEMA_signal_11222), .A1_t (new_AGEMA_signal_11223), .A1_f (new_AGEMA_signal_11224), .B0_t (Inst_bSbox_L4), .B0_f (new_AGEMA_signal_11246), .B1_t (new_AGEMA_signal_11247), .B1_f (new_AGEMA_signal_11248), .Z0_t (Inst_bSbox_L19), .Z0_f (new_AGEMA_signal_11282), .Z1_t (new_AGEMA_signal_11283), .Z1_f (new_AGEMA_signal_11284) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L20_U1 ( .A0_t (Inst_bSbox_L0), .A0_f (new_AGEMA_signal_11264), .A1_t (new_AGEMA_signal_11265), .A1_f (new_AGEMA_signal_11266), .B0_t (Inst_bSbox_L1), .B0_f (new_AGEMA_signal_11225), .B1_t (new_AGEMA_signal_11226), .B1_f (new_AGEMA_signal_11227), .Z0_t (Inst_bSbox_L20), .Z0_f (new_AGEMA_signal_11297), .Z1_t (new_AGEMA_signal_11298), .Z1_f (new_AGEMA_signal_11299) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L21_U1 ( .A0_t (Inst_bSbox_L1), .A0_f (new_AGEMA_signal_11225), .A1_t (new_AGEMA_signal_11226), .A1_f (new_AGEMA_signal_11227), .B0_t (Inst_bSbox_L7), .B0_f (new_AGEMA_signal_11270), .B1_t (new_AGEMA_signal_11271), .B1_f (new_AGEMA_signal_11272), .Z0_t (Inst_bSbox_L21), .Z0_f (new_AGEMA_signal_11300), .Z1_t (new_AGEMA_signal_11301), .Z1_f (new_AGEMA_signal_11302) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L22_U1 ( .A0_t (Inst_bSbox_L3), .A0_f (new_AGEMA_signal_11243), .A1_t (new_AGEMA_signal_11244), .A1_f (new_AGEMA_signal_11245), .B0_t (Inst_bSbox_L12), .B0_f (new_AGEMA_signal_11231), .B1_t (new_AGEMA_signal_11232), .B1_f (new_AGEMA_signal_11233), .Z0_t (Inst_bSbox_L22), .Z0_f (new_AGEMA_signal_11285), .Z1_t (new_AGEMA_signal_11286), .Z1_f (new_AGEMA_signal_11287) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L23_U1 ( .A0_t (Inst_bSbox_L18), .A0_f (new_AGEMA_signal_11261), .A1_t (new_AGEMA_signal_11262), .A1_f (new_AGEMA_signal_11263), .B0_t (Inst_bSbox_L2), .B0_f (new_AGEMA_signal_11240), .B1_t (new_AGEMA_signal_11241), .B1_f (new_AGEMA_signal_11242), .Z0_t (Inst_bSbox_L23), .Z0_f (new_AGEMA_signal_11288), .Z1_t (new_AGEMA_signal_11289), .Z1_f (new_AGEMA_signal_11290) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L24_U1 ( .A0_t (Inst_bSbox_L15), .A0_f (new_AGEMA_signal_11255), .A1_t (new_AGEMA_signal_11256), .A1_f (new_AGEMA_signal_11257), .B0_t (Inst_bSbox_L9), .B0_f (new_AGEMA_signal_11273), .B1_t (new_AGEMA_signal_11274), .B1_f (new_AGEMA_signal_11275), .Z0_t (Inst_bSbox_L24), .Z0_f (new_AGEMA_signal_11303), .Z1_t (new_AGEMA_signal_11304), .Z1_f (new_AGEMA_signal_11305) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L25_U1 ( .A0_t (Inst_bSbox_L6), .A0_f (new_AGEMA_signal_11267), .A1_t (new_AGEMA_signal_11268), .A1_f (new_AGEMA_signal_11269), .B0_t (Inst_bSbox_L10), .B0_f (new_AGEMA_signal_11276), .B1_t (new_AGEMA_signal_11277), .B1_f (new_AGEMA_signal_11278), .Z0_t (Inst_bSbox_L25), .Z0_f (new_AGEMA_signal_11306), .Z1_t (new_AGEMA_signal_11307), .Z1_f (new_AGEMA_signal_11308) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L26_U1 ( .A0_t (Inst_bSbox_L7), .A0_f (new_AGEMA_signal_11270), .A1_t (new_AGEMA_signal_11271), .A1_f (new_AGEMA_signal_11272), .B0_t (Inst_bSbox_L9), .B0_f (new_AGEMA_signal_11273), .B1_t (new_AGEMA_signal_11274), .B1_f (new_AGEMA_signal_11275), .Z0_t (Inst_bSbox_L26), .Z0_f (new_AGEMA_signal_11309), .Z1_t (new_AGEMA_signal_11310), .Z1_f (new_AGEMA_signal_11311) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L27_U1 ( .A0_t (Inst_bSbox_L8), .A0_f (new_AGEMA_signal_11228), .A1_t (new_AGEMA_signal_11229), .A1_f (new_AGEMA_signal_11230), .B0_t (Inst_bSbox_L10), .B0_f (new_AGEMA_signal_11276), .B1_t (new_AGEMA_signal_11277), .B1_f (new_AGEMA_signal_11278), .Z0_t (Inst_bSbox_L27), .Z0_f (new_AGEMA_signal_11312), .Z1_t (new_AGEMA_signal_11313), .Z1_f (new_AGEMA_signal_11314) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L28_U1 ( .A0_t (Inst_bSbox_L11), .A0_f (new_AGEMA_signal_11279), .A1_t (new_AGEMA_signal_11280), .A1_f (new_AGEMA_signal_11281), .B0_t (Inst_bSbox_L14), .B0_f (new_AGEMA_signal_11252), .B1_t (new_AGEMA_signal_11253), .B1_f (new_AGEMA_signal_11254), .Z0_t (Inst_bSbox_L28), .Z0_f (new_AGEMA_signal_11315), .Z1_t (new_AGEMA_signal_11316), .Z1_f (new_AGEMA_signal_11317) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L29_U1 ( .A0_t (Inst_bSbox_L11), .A0_f (new_AGEMA_signal_11279), .A1_t (new_AGEMA_signal_11280), .A1_f (new_AGEMA_signal_11281), .B0_t (Inst_bSbox_L17), .B0_f (new_AGEMA_signal_11258), .B1_t (new_AGEMA_signal_11259), .B1_f (new_AGEMA_signal_11260), .Z0_t (Inst_bSbox_L29), .Z0_f (new_AGEMA_signal_11318), .Z1_t (new_AGEMA_signal_11319), .Z1_f (new_AGEMA_signal_11320) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_S0_U1 ( .A0_t (Inst_bSbox_L6), .A0_f (new_AGEMA_signal_11267), .A1_t (new_AGEMA_signal_11268), .A1_f (new_AGEMA_signal_11269), .B0_t (Inst_bSbox_L24), .B0_f (new_AGEMA_signal_11303), .B1_t (new_AGEMA_signal_11304), .B1_f (new_AGEMA_signal_11305), .Z0_t (SboxOut[7]), .Z0_f (new_AGEMA_signal_11330), .Z1_t (new_AGEMA_signal_11331), .Z1_f (new_AGEMA_signal_11332) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Inst_bSbox_XOR_S1_U1 ( .A0_t (Inst_bSbox_L16), .A0_f (new_AGEMA_signal_11294), .A1_t (new_AGEMA_signal_11295), .A1_f (new_AGEMA_signal_11296), .B0_t (Inst_bSbox_L26), .B0_f (new_AGEMA_signal_11309), .B1_t (new_AGEMA_signal_11310), .B1_f (new_AGEMA_signal_11311), .Z0_t (SboxOut[6]), .Z0_f (new_AGEMA_signal_11333), .Z1_t (new_AGEMA_signal_11334), .Z1_f (new_AGEMA_signal_11335) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Inst_bSbox_XOR_S2_U1 ( .A0_t (Inst_bSbox_L19), .A0_f (new_AGEMA_signal_11282), .A1_t (new_AGEMA_signal_11283), .A1_f (new_AGEMA_signal_11284), .B0_t (Inst_bSbox_L28), .B0_f (new_AGEMA_signal_11315), .B1_t (new_AGEMA_signal_11316), .B1_f (new_AGEMA_signal_11317), .Z0_t (SboxOut[5]), .Z0_f (new_AGEMA_signal_11336), .Z1_t (new_AGEMA_signal_11337), .Z1_f (new_AGEMA_signal_11338) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_S3_U1 ( .A0_t (Inst_bSbox_L6), .A0_f (new_AGEMA_signal_11267), .A1_t (new_AGEMA_signal_11268), .A1_f (new_AGEMA_signal_11269), .B0_t (Inst_bSbox_L21), .B0_f (new_AGEMA_signal_11300), .B1_t (new_AGEMA_signal_11301), .B1_f (new_AGEMA_signal_11302), .Z0_t (SboxOut[4]), .Z0_f (new_AGEMA_signal_11339), .Z1_t (new_AGEMA_signal_11340), .Z1_f (new_AGEMA_signal_11341) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_S4_U1 ( .A0_t (Inst_bSbox_L20), .A0_f (new_AGEMA_signal_11297), .A1_t (new_AGEMA_signal_11298), .A1_f (new_AGEMA_signal_11299), .B0_t (Inst_bSbox_L22), .B0_f (new_AGEMA_signal_11285), .B1_t (new_AGEMA_signal_11286), .B1_f (new_AGEMA_signal_11287), .Z0_t (SboxOut[3]), .Z0_f (new_AGEMA_signal_11342), .Z1_t (new_AGEMA_signal_11343), .Z1_f (new_AGEMA_signal_11344) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_S5_U1 ( .A0_t (Inst_bSbox_L25), .A0_f (new_AGEMA_signal_11306), .A1_t (new_AGEMA_signal_11307), .A1_f (new_AGEMA_signal_11308), .B0_t (Inst_bSbox_L29), .B0_f (new_AGEMA_signal_11318), .B1_t (new_AGEMA_signal_11319), .B1_f (new_AGEMA_signal_11320), .Z0_t (SboxOut[2]), .Z0_f (new_AGEMA_signal_11345), .Z1_t (new_AGEMA_signal_11346), .Z1_f (new_AGEMA_signal_11347) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Inst_bSbox_XOR_S6_U1 ( .A0_t (Inst_bSbox_L13), .A0_f (new_AGEMA_signal_11291), .A1_t (new_AGEMA_signal_11292), .A1_f (new_AGEMA_signal_11293), .B0_t (Inst_bSbox_L27), .B0_f (new_AGEMA_signal_11312), .B1_t (new_AGEMA_signal_11313), .B1_f (new_AGEMA_signal_11314), .Z0_t (SboxOut[1]), .Z0_f (new_AGEMA_signal_11348), .Z1_t (new_AGEMA_signal_11349), .Z1_f (new_AGEMA_signal_11350) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Inst_bSbox_XOR_S7_U1 ( .A0_t (Inst_bSbox_L6), .A0_f (new_AGEMA_signal_11267), .A1_t (new_AGEMA_signal_11268), .A1_f (new_AGEMA_signal_11269), .B0_t (Inst_bSbox_L23), .B0_f (new_AGEMA_signal_11288), .B1_t (new_AGEMA_signal_11289), .B1_f (new_AGEMA_signal_11290), .Z0_t (SboxOut[0]), .Z0_f (new_AGEMA_signal_11321), .Z1_t (new_AGEMA_signal_11322), .Z1_f (new_AGEMA_signal_11323) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1), .NL(1'b0)) new_AGEMA_gate_3161 ( .A0_t (ctrl_n9), .A0_f (new_AGEMA_signal_7394), .B0_t (1'b0), .B0_f (1'b1), .Z0_t (enRCon), .Z0_f (new_AGEMA_signal_5791) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1), .NL(1'b0)) new_AGEMA_gate_3162 ( .A0_t (start_t), .A0_f (start_f), .B0_t (1'b0), .B0_f (1'b1), .Z0_t (nReset), .Z0_f (new_AGEMA_signal_3502) ) ;

    /* register cells */
endmodule
