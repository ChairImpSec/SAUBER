/* modified netlist. Source: module LED in file /mnt/c/Users/amirm/Desktop/Papers_in_progress/SAUBER/Design for our FPGA/12-LED_round_based_encryption_PortParallel/4-AGEMA/LED.v */
/* 0 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 1 register stage(s) in total */

module LED_SAUBER_Pipeline_d1 (IN_plaintext, IN_key, IN_reset, OUT_ciphertext, OUT_done);
    input [63:0] IN_plaintext ;
    input [127:0] IN_key ;
    input IN_reset ;
    output [63:0] OUT_ciphertext ;
    output OUT_done ;
    wire n15 ;
    wire n16 ;
    wire n17 ;
    wire n18 ;
    wire n19 ;
    wire n20 ;
    wire LED_128_Instance_n29 ;
    wire LED_128_Instance_n19 ;
    wire LED_128_Instance_n18 ;
    wire LED_128_Instance_n17 ;
    wire LED_128_Instance_n16 ;
    wire LED_128_Instance_n13 ;
    wire LED_128_Instance_n12 ;
    wire LED_128_Instance_n11 ;
    wire LED_128_Instance_n9 ;
    wire LED_128_Instance_n8 ;
    wire LED_128_Instance_n31 ;
    wire LED_128_Instance_n24 ;
    wire LED_128_Instance_ks_0 ;
    wire LED_128_Instance_ks_3_ ;
    wire LED_128_Instance_n23 ;
    wire LED_128_Instance_n22 ;
    wire LED_128_Instance_MUX_state0_mux_inst_0_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_0_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_1_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_1_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_2_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_2_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_3_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_3_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_4_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_4_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_5_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_5_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_6_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_6_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_7_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_7_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_8_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_8_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_9_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_9_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_10_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_10_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_11_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_11_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_12_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_12_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_13_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_13_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_14_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_14_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_15_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_15_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_16_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_16_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_17_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_17_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_18_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_18_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_19_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_19_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_20_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_20_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_21_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_21_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_22_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_22_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_23_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_23_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_24_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_24_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_25_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_25_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_26_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_26_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_27_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_27_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_28_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_28_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_29_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_29_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_30_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_30_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_31_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_31_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_32_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_32_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_33_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_33_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_34_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_34_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_35_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_35_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_36_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_36_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_37_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_37_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_38_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_38_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_39_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_39_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_40_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_40_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_41_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_41_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_42_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_42_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_43_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_43_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_44_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_44_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_45_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_45_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_46_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_46_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_47_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_47_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_48_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_48_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_49_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_49_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_50_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_50_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_51_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_51_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_52_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_52_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_53_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_53_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_54_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_54_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_55_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_55_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_56_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_56_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_57_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_57_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_58_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_58_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_59_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_59_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_60_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_60_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_61_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_61_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_62_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_62_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_63_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_63_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_0_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_0_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_1_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_1_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_2_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_2_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_3_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_3_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_4_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_4_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_5_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_5_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_6_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_6_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_7_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_7_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_8_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_8_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_9_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_9_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_10_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_10_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_11_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_11_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_12_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_12_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_13_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_13_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_14_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_14_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_15_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_15_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_16_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_16_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_17_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_17_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_18_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_18_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_19_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_19_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_20_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_20_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_21_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_21_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_22_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_22_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_23_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_23_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_24_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_24_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_25_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_25_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_26_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_26_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_27_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_27_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_28_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_28_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_29_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_29_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_30_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_30_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_31_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_31_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_32_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_32_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_33_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_33_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_34_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_34_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_35_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_35_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_36_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_36_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_37_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_37_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_38_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_38_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_39_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_39_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_40_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_40_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_41_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_41_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_42_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_42_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_43_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_43_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_44_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_44_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_45_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_45_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_46_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_46_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_47_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_47_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_48_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_48_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_49_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_49_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_50_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_50_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_51_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_51_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_52_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_52_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_53_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_53_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_54_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_54_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_55_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_55_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_56_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_56_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_57_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_57_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_58_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_58_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_59_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_59_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_60_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_60_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_61_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_61_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_62_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_62_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_63_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_63_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_0_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_0_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_1_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_1_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_2_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_2_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_3_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_3_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_4_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_4_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_5_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_5_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_6_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_6_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_7_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_7_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_8_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_8_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_9_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_9_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_10_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_10_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_11_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_11_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_12_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_12_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_13_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_13_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_14_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_14_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_15_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_15_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_16_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_16_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_17_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_17_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_18_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_18_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_19_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_19_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_20_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_20_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_21_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_21_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_22_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_22_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_23_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_23_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_24_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_24_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_25_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_25_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_26_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_26_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_27_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_27_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_28_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_28_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_29_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_29_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_30_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_30_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_31_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_31_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_32_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_32_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_33_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_33_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_34_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_34_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_35_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_35_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_36_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_36_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_37_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_37_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_38_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_38_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_39_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_39_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_40_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_40_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_41_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_41_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_42_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_42_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_43_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_43_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_44_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_44_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_45_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_45_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_46_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_46_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_47_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_47_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_48_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_48_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_49_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_49_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_50_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_50_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_51_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_51_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_52_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_52_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_53_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_53_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_54_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_54_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_55_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_55_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_56_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_56_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_57_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_57_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_58_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_58_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_59_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_59_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_60_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_60_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_61_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_61_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_62_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_62_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_63_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_63_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_0_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_0_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_1_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_1_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_2_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_2_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_3_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_3_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_4_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_4_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_5_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_5_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_6_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_6_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_7_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_7_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_8_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_8_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_9_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_9_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_10_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_10_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_11_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_11_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_12_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_12_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_13_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_13_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_14_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_14_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_15_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_15_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_16_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_16_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_17_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_17_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_18_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_18_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_19_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_19_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_20_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_20_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_21_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_21_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_22_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_22_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_23_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_23_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_24_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_24_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_25_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_25_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_26_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_26_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_27_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_27_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_28_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_28_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_29_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_29_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_30_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_30_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_31_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_31_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_32_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_32_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_33_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_33_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_34_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_34_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_35_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_35_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_36_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_36_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_37_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_37_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_38_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_38_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_39_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_39_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_40_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_40_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_41_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_41_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_42_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_42_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_43_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_43_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_44_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_44_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_45_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_45_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_46_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_46_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_47_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_47_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_48_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_48_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_49_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_49_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_50_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_50_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_51_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_51_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_52_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_52_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_53_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_53_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_54_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_54_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_55_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_55_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_56_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_56_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_57_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_57_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_58_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_58_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_59_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_59_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_60_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_60_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_61_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_61_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_62_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_62_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_63_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_63_U1_X ;
    wire LED_128_Instance_SBox_Instance_0_L8 ;
    wire LED_128_Instance_SBox_Instance_0_L7 ;
    wire LED_128_Instance_SBox_Instance_0_T3 ;
    wire LED_128_Instance_SBox_Instance_0_T1 ;
    wire LED_128_Instance_SBox_Instance_0_Q7 ;
    wire LED_128_Instance_SBox_Instance_0_Q6 ;
    wire LED_128_Instance_SBox_Instance_0_L5 ;
    wire LED_128_Instance_SBox_Instance_0_T2 ;
    wire LED_128_Instance_SBox_Instance_0_L4 ;
    wire LED_128_Instance_SBox_Instance_0_Q3 ;
    wire LED_128_Instance_SBox_Instance_0_L3 ;
    wire LED_128_Instance_SBox_Instance_0_Q2 ;
    wire LED_128_Instance_SBox_Instance_0_T0 ;
    wire LED_128_Instance_SBox_Instance_0_L2 ;
    wire LED_128_Instance_SBox_Instance_0_L1 ;
    wire LED_128_Instance_SBox_Instance_0_L0 ;
    wire LED_128_Instance_SBox_Instance_1_L8 ;
    wire LED_128_Instance_SBox_Instance_1_L7 ;
    wire LED_128_Instance_SBox_Instance_1_T3 ;
    wire LED_128_Instance_SBox_Instance_1_T1 ;
    wire LED_128_Instance_SBox_Instance_1_Q7 ;
    wire LED_128_Instance_SBox_Instance_1_Q6 ;
    wire LED_128_Instance_SBox_Instance_1_L5 ;
    wire LED_128_Instance_SBox_Instance_1_T2 ;
    wire LED_128_Instance_SBox_Instance_1_L4 ;
    wire LED_128_Instance_SBox_Instance_1_Q3 ;
    wire LED_128_Instance_SBox_Instance_1_L3 ;
    wire LED_128_Instance_SBox_Instance_1_Q2 ;
    wire LED_128_Instance_SBox_Instance_1_T0 ;
    wire LED_128_Instance_SBox_Instance_1_L2 ;
    wire LED_128_Instance_SBox_Instance_1_L1 ;
    wire LED_128_Instance_SBox_Instance_1_L0 ;
    wire LED_128_Instance_SBox_Instance_2_L8 ;
    wire LED_128_Instance_SBox_Instance_2_L7 ;
    wire LED_128_Instance_SBox_Instance_2_T3 ;
    wire LED_128_Instance_SBox_Instance_2_T1 ;
    wire LED_128_Instance_SBox_Instance_2_Q7 ;
    wire LED_128_Instance_SBox_Instance_2_Q6 ;
    wire LED_128_Instance_SBox_Instance_2_L5 ;
    wire LED_128_Instance_SBox_Instance_2_T2 ;
    wire LED_128_Instance_SBox_Instance_2_L4 ;
    wire LED_128_Instance_SBox_Instance_2_Q3 ;
    wire LED_128_Instance_SBox_Instance_2_L3 ;
    wire LED_128_Instance_SBox_Instance_2_Q2 ;
    wire LED_128_Instance_SBox_Instance_2_T0 ;
    wire LED_128_Instance_SBox_Instance_2_L2 ;
    wire LED_128_Instance_SBox_Instance_2_L1 ;
    wire LED_128_Instance_SBox_Instance_2_L0 ;
    wire LED_128_Instance_SBox_Instance_3_L8 ;
    wire LED_128_Instance_SBox_Instance_3_L7 ;
    wire LED_128_Instance_SBox_Instance_3_T3 ;
    wire LED_128_Instance_SBox_Instance_3_T1 ;
    wire LED_128_Instance_SBox_Instance_3_Q7 ;
    wire LED_128_Instance_SBox_Instance_3_Q6 ;
    wire LED_128_Instance_SBox_Instance_3_L5 ;
    wire LED_128_Instance_SBox_Instance_3_T2 ;
    wire LED_128_Instance_SBox_Instance_3_L4 ;
    wire LED_128_Instance_SBox_Instance_3_Q3 ;
    wire LED_128_Instance_SBox_Instance_3_L3 ;
    wire LED_128_Instance_SBox_Instance_3_Q2 ;
    wire LED_128_Instance_SBox_Instance_3_T0 ;
    wire LED_128_Instance_SBox_Instance_3_L2 ;
    wire LED_128_Instance_SBox_Instance_3_L1 ;
    wire LED_128_Instance_SBox_Instance_3_L0 ;
    wire LED_128_Instance_SBox_Instance_4_L8 ;
    wire LED_128_Instance_SBox_Instance_4_L7 ;
    wire LED_128_Instance_SBox_Instance_4_T3 ;
    wire LED_128_Instance_SBox_Instance_4_T1 ;
    wire LED_128_Instance_SBox_Instance_4_Q7 ;
    wire LED_128_Instance_SBox_Instance_4_Q6 ;
    wire LED_128_Instance_SBox_Instance_4_L5 ;
    wire LED_128_Instance_SBox_Instance_4_T2 ;
    wire LED_128_Instance_SBox_Instance_4_L4 ;
    wire LED_128_Instance_SBox_Instance_4_Q3 ;
    wire LED_128_Instance_SBox_Instance_4_L3 ;
    wire LED_128_Instance_SBox_Instance_4_Q2 ;
    wire LED_128_Instance_SBox_Instance_4_T0 ;
    wire LED_128_Instance_SBox_Instance_4_L2 ;
    wire LED_128_Instance_SBox_Instance_4_L1 ;
    wire LED_128_Instance_SBox_Instance_4_L0 ;
    wire LED_128_Instance_SBox_Instance_5_L8 ;
    wire LED_128_Instance_SBox_Instance_5_L7 ;
    wire LED_128_Instance_SBox_Instance_5_T3 ;
    wire LED_128_Instance_SBox_Instance_5_T1 ;
    wire LED_128_Instance_SBox_Instance_5_Q7 ;
    wire LED_128_Instance_SBox_Instance_5_Q6 ;
    wire LED_128_Instance_SBox_Instance_5_L5 ;
    wire LED_128_Instance_SBox_Instance_5_T2 ;
    wire LED_128_Instance_SBox_Instance_5_L4 ;
    wire LED_128_Instance_SBox_Instance_5_Q3 ;
    wire LED_128_Instance_SBox_Instance_5_L3 ;
    wire LED_128_Instance_SBox_Instance_5_Q2 ;
    wire LED_128_Instance_SBox_Instance_5_T0 ;
    wire LED_128_Instance_SBox_Instance_5_L2 ;
    wire LED_128_Instance_SBox_Instance_5_L1 ;
    wire LED_128_Instance_SBox_Instance_5_L0 ;
    wire LED_128_Instance_SBox_Instance_6_L8 ;
    wire LED_128_Instance_SBox_Instance_6_L7 ;
    wire LED_128_Instance_SBox_Instance_6_T3 ;
    wire LED_128_Instance_SBox_Instance_6_T1 ;
    wire LED_128_Instance_SBox_Instance_6_Q7 ;
    wire LED_128_Instance_SBox_Instance_6_Q6 ;
    wire LED_128_Instance_SBox_Instance_6_L5 ;
    wire LED_128_Instance_SBox_Instance_6_T2 ;
    wire LED_128_Instance_SBox_Instance_6_L4 ;
    wire LED_128_Instance_SBox_Instance_6_Q3 ;
    wire LED_128_Instance_SBox_Instance_6_L3 ;
    wire LED_128_Instance_SBox_Instance_6_Q2 ;
    wire LED_128_Instance_SBox_Instance_6_T0 ;
    wire LED_128_Instance_SBox_Instance_6_L2 ;
    wire LED_128_Instance_SBox_Instance_6_L1 ;
    wire LED_128_Instance_SBox_Instance_6_L0 ;
    wire LED_128_Instance_SBox_Instance_7_L8 ;
    wire LED_128_Instance_SBox_Instance_7_L7 ;
    wire LED_128_Instance_SBox_Instance_7_T3 ;
    wire LED_128_Instance_SBox_Instance_7_T1 ;
    wire LED_128_Instance_SBox_Instance_7_Q7 ;
    wire LED_128_Instance_SBox_Instance_7_Q6 ;
    wire LED_128_Instance_SBox_Instance_7_L5 ;
    wire LED_128_Instance_SBox_Instance_7_T2 ;
    wire LED_128_Instance_SBox_Instance_7_L4 ;
    wire LED_128_Instance_SBox_Instance_7_Q3 ;
    wire LED_128_Instance_SBox_Instance_7_L3 ;
    wire LED_128_Instance_SBox_Instance_7_Q2 ;
    wire LED_128_Instance_SBox_Instance_7_T0 ;
    wire LED_128_Instance_SBox_Instance_7_L2 ;
    wire LED_128_Instance_SBox_Instance_7_L1 ;
    wire LED_128_Instance_SBox_Instance_7_L0 ;
    wire LED_128_Instance_SBox_Instance_8_L8 ;
    wire LED_128_Instance_SBox_Instance_8_L7 ;
    wire LED_128_Instance_SBox_Instance_8_T3 ;
    wire LED_128_Instance_SBox_Instance_8_T1 ;
    wire LED_128_Instance_SBox_Instance_8_Q7 ;
    wire LED_128_Instance_SBox_Instance_8_Q6 ;
    wire LED_128_Instance_SBox_Instance_8_L5 ;
    wire LED_128_Instance_SBox_Instance_8_T2 ;
    wire LED_128_Instance_SBox_Instance_8_L4 ;
    wire LED_128_Instance_SBox_Instance_8_Q3 ;
    wire LED_128_Instance_SBox_Instance_8_L3 ;
    wire LED_128_Instance_SBox_Instance_8_Q2 ;
    wire LED_128_Instance_SBox_Instance_8_T0 ;
    wire LED_128_Instance_SBox_Instance_8_L2 ;
    wire LED_128_Instance_SBox_Instance_8_L1 ;
    wire LED_128_Instance_SBox_Instance_8_L0 ;
    wire LED_128_Instance_SBox_Instance_9_L8 ;
    wire LED_128_Instance_SBox_Instance_9_L7 ;
    wire LED_128_Instance_SBox_Instance_9_T3 ;
    wire LED_128_Instance_SBox_Instance_9_T1 ;
    wire LED_128_Instance_SBox_Instance_9_Q7 ;
    wire LED_128_Instance_SBox_Instance_9_Q6 ;
    wire LED_128_Instance_SBox_Instance_9_L5 ;
    wire LED_128_Instance_SBox_Instance_9_T2 ;
    wire LED_128_Instance_SBox_Instance_9_L4 ;
    wire LED_128_Instance_SBox_Instance_9_Q3 ;
    wire LED_128_Instance_SBox_Instance_9_L3 ;
    wire LED_128_Instance_SBox_Instance_9_Q2 ;
    wire LED_128_Instance_SBox_Instance_9_T0 ;
    wire LED_128_Instance_SBox_Instance_9_L2 ;
    wire LED_128_Instance_SBox_Instance_9_L1 ;
    wire LED_128_Instance_SBox_Instance_9_L0 ;
    wire LED_128_Instance_SBox_Instance_10_L8 ;
    wire LED_128_Instance_SBox_Instance_10_L7 ;
    wire LED_128_Instance_SBox_Instance_10_T3 ;
    wire LED_128_Instance_SBox_Instance_10_T1 ;
    wire LED_128_Instance_SBox_Instance_10_Q7 ;
    wire LED_128_Instance_SBox_Instance_10_Q6 ;
    wire LED_128_Instance_SBox_Instance_10_L5 ;
    wire LED_128_Instance_SBox_Instance_10_T2 ;
    wire LED_128_Instance_SBox_Instance_10_L4 ;
    wire LED_128_Instance_SBox_Instance_10_Q3 ;
    wire LED_128_Instance_SBox_Instance_10_L3 ;
    wire LED_128_Instance_SBox_Instance_10_Q2 ;
    wire LED_128_Instance_SBox_Instance_10_T0 ;
    wire LED_128_Instance_SBox_Instance_10_L2 ;
    wire LED_128_Instance_SBox_Instance_10_L1 ;
    wire LED_128_Instance_SBox_Instance_10_L0 ;
    wire LED_128_Instance_SBox_Instance_11_L8 ;
    wire LED_128_Instance_SBox_Instance_11_L7 ;
    wire LED_128_Instance_SBox_Instance_11_T3 ;
    wire LED_128_Instance_SBox_Instance_11_T1 ;
    wire LED_128_Instance_SBox_Instance_11_Q7 ;
    wire LED_128_Instance_SBox_Instance_11_Q6 ;
    wire LED_128_Instance_SBox_Instance_11_L5 ;
    wire LED_128_Instance_SBox_Instance_11_T2 ;
    wire LED_128_Instance_SBox_Instance_11_L4 ;
    wire LED_128_Instance_SBox_Instance_11_Q3 ;
    wire LED_128_Instance_SBox_Instance_11_L3 ;
    wire LED_128_Instance_SBox_Instance_11_Q2 ;
    wire LED_128_Instance_SBox_Instance_11_T0 ;
    wire LED_128_Instance_SBox_Instance_11_L2 ;
    wire LED_128_Instance_SBox_Instance_11_L1 ;
    wire LED_128_Instance_SBox_Instance_11_L0 ;
    wire LED_128_Instance_SBox_Instance_12_L8 ;
    wire LED_128_Instance_SBox_Instance_12_L7 ;
    wire LED_128_Instance_SBox_Instance_12_T3 ;
    wire LED_128_Instance_SBox_Instance_12_T1 ;
    wire LED_128_Instance_SBox_Instance_12_Q7 ;
    wire LED_128_Instance_SBox_Instance_12_Q6 ;
    wire LED_128_Instance_SBox_Instance_12_L5 ;
    wire LED_128_Instance_SBox_Instance_12_T2 ;
    wire LED_128_Instance_SBox_Instance_12_L4 ;
    wire LED_128_Instance_SBox_Instance_12_Q3 ;
    wire LED_128_Instance_SBox_Instance_12_L3 ;
    wire LED_128_Instance_SBox_Instance_12_Q2 ;
    wire LED_128_Instance_SBox_Instance_12_T0 ;
    wire LED_128_Instance_SBox_Instance_12_L2 ;
    wire LED_128_Instance_SBox_Instance_12_L1 ;
    wire LED_128_Instance_SBox_Instance_12_L0 ;
    wire LED_128_Instance_SBox_Instance_13_L8 ;
    wire LED_128_Instance_SBox_Instance_13_L7 ;
    wire LED_128_Instance_SBox_Instance_13_T3 ;
    wire LED_128_Instance_SBox_Instance_13_T1 ;
    wire LED_128_Instance_SBox_Instance_13_Q7 ;
    wire LED_128_Instance_SBox_Instance_13_Q6 ;
    wire LED_128_Instance_SBox_Instance_13_L5 ;
    wire LED_128_Instance_SBox_Instance_13_T2 ;
    wire LED_128_Instance_SBox_Instance_13_L4 ;
    wire LED_128_Instance_SBox_Instance_13_Q3 ;
    wire LED_128_Instance_SBox_Instance_13_L3 ;
    wire LED_128_Instance_SBox_Instance_13_Q2 ;
    wire LED_128_Instance_SBox_Instance_13_T0 ;
    wire LED_128_Instance_SBox_Instance_13_L2 ;
    wire LED_128_Instance_SBox_Instance_13_L1 ;
    wire LED_128_Instance_SBox_Instance_13_L0 ;
    wire LED_128_Instance_SBox_Instance_14_L8 ;
    wire LED_128_Instance_SBox_Instance_14_L7 ;
    wire LED_128_Instance_SBox_Instance_14_T3 ;
    wire LED_128_Instance_SBox_Instance_14_T1 ;
    wire LED_128_Instance_SBox_Instance_14_Q7 ;
    wire LED_128_Instance_SBox_Instance_14_Q6 ;
    wire LED_128_Instance_SBox_Instance_14_L5 ;
    wire LED_128_Instance_SBox_Instance_14_T2 ;
    wire LED_128_Instance_SBox_Instance_14_L4 ;
    wire LED_128_Instance_SBox_Instance_14_Q3 ;
    wire LED_128_Instance_SBox_Instance_14_L3 ;
    wire LED_128_Instance_SBox_Instance_14_Q2 ;
    wire LED_128_Instance_SBox_Instance_14_T0 ;
    wire LED_128_Instance_SBox_Instance_14_L2 ;
    wire LED_128_Instance_SBox_Instance_14_L1 ;
    wire LED_128_Instance_SBox_Instance_14_L0 ;
    wire LED_128_Instance_SBox_Instance_15_L8 ;
    wire LED_128_Instance_SBox_Instance_15_L7 ;
    wire LED_128_Instance_SBox_Instance_15_T3 ;
    wire LED_128_Instance_SBox_Instance_15_T1 ;
    wire LED_128_Instance_SBox_Instance_15_Q7 ;
    wire LED_128_Instance_SBox_Instance_15_Q6 ;
    wire LED_128_Instance_SBox_Instance_15_L5 ;
    wire LED_128_Instance_SBox_Instance_15_T2 ;
    wire LED_128_Instance_SBox_Instance_15_L4 ;
    wire LED_128_Instance_SBox_Instance_15_Q3 ;
    wire LED_128_Instance_SBox_Instance_15_L3 ;
    wire LED_128_Instance_SBox_Instance_15_Q2 ;
    wire LED_128_Instance_SBox_Instance_15_T0 ;
    wire LED_128_Instance_SBox_Instance_15_L2 ;
    wire LED_128_Instance_SBox_Instance_15_L1 ;
    wire LED_128_Instance_SBox_Instance_15_L0 ;
    wire LED_128_Instance_MCS_Instance_0_n42 ;
    wire LED_128_Instance_MCS_Instance_0_n41 ;
    wire LED_128_Instance_MCS_Instance_0_n40 ;
    wire LED_128_Instance_MCS_Instance_0_n39 ;
    wire LED_128_Instance_MCS_Instance_0_n38 ;
    wire LED_128_Instance_MCS_Instance_0_n37 ;
    wire LED_128_Instance_MCS_Instance_0_n36 ;
    wire LED_128_Instance_MCS_Instance_0_n35 ;
    wire LED_128_Instance_MCS_Instance_0_n34 ;
    wire LED_128_Instance_MCS_Instance_0_n33 ;
    wire LED_128_Instance_MCS_Instance_0_n32 ;
    wire LED_128_Instance_MCS_Instance_0_n31 ;
    wire LED_128_Instance_MCS_Instance_0_n30 ;
    wire LED_128_Instance_MCS_Instance_0_n29 ;
    wire LED_128_Instance_MCS_Instance_0_n28 ;
    wire LED_128_Instance_MCS_Instance_0_n27 ;
    wire LED_128_Instance_MCS_Instance_0_n26 ;
    wire LED_128_Instance_MCS_Instance_0_n25 ;
    wire LED_128_Instance_MCS_Instance_0_n24 ;
    wire LED_128_Instance_MCS_Instance_0_n23 ;
    wire LED_128_Instance_MCS_Instance_0_n22 ;
    wire LED_128_Instance_MCS_Instance_0_n21 ;
    wire LED_128_Instance_MCS_Instance_0_n20 ;
    wire LED_128_Instance_MCS_Instance_0_n19 ;
    wire LED_128_Instance_MCS_Instance_0_n18 ;
    wire LED_128_Instance_MCS_Instance_0_n17 ;
    wire LED_128_Instance_MCS_Instance_0_n16 ;
    wire LED_128_Instance_MCS_Instance_0_n15 ;
    wire LED_128_Instance_MCS_Instance_0_n14 ;
    wire LED_128_Instance_MCS_Instance_0_n13 ;
    wire LED_128_Instance_MCS_Instance_0_n12 ;
    wire LED_128_Instance_MCS_Instance_0_n11 ;
    wire LED_128_Instance_MCS_Instance_0_n10 ;
    wire LED_128_Instance_MCS_Instance_0_n9 ;
    wire LED_128_Instance_MCS_Instance_0_n8 ;
    wire LED_128_Instance_MCS_Instance_0_n7 ;
    wire LED_128_Instance_MCS_Instance_0_n6 ;
    wire LED_128_Instance_MCS_Instance_0_n5 ;
    wire LED_128_Instance_MCS_Instance_0_n4 ;
    wire LED_128_Instance_MCS_Instance_0_n3 ;
    wire LED_128_Instance_MCS_Instance_0_n2 ;
    wire LED_128_Instance_MCS_Instance_0_n1 ;
    wire LED_128_Instance_MCS_Instance_1_n42 ;
    wire LED_128_Instance_MCS_Instance_1_n41 ;
    wire LED_128_Instance_MCS_Instance_1_n40 ;
    wire LED_128_Instance_MCS_Instance_1_n39 ;
    wire LED_128_Instance_MCS_Instance_1_n38 ;
    wire LED_128_Instance_MCS_Instance_1_n37 ;
    wire LED_128_Instance_MCS_Instance_1_n36 ;
    wire LED_128_Instance_MCS_Instance_1_n35 ;
    wire LED_128_Instance_MCS_Instance_1_n34 ;
    wire LED_128_Instance_MCS_Instance_1_n33 ;
    wire LED_128_Instance_MCS_Instance_1_n32 ;
    wire LED_128_Instance_MCS_Instance_1_n31 ;
    wire LED_128_Instance_MCS_Instance_1_n30 ;
    wire LED_128_Instance_MCS_Instance_1_n29 ;
    wire LED_128_Instance_MCS_Instance_1_n28 ;
    wire LED_128_Instance_MCS_Instance_1_n27 ;
    wire LED_128_Instance_MCS_Instance_1_n26 ;
    wire LED_128_Instance_MCS_Instance_1_n25 ;
    wire LED_128_Instance_MCS_Instance_1_n24 ;
    wire LED_128_Instance_MCS_Instance_1_n23 ;
    wire LED_128_Instance_MCS_Instance_1_n22 ;
    wire LED_128_Instance_MCS_Instance_1_n21 ;
    wire LED_128_Instance_MCS_Instance_1_n20 ;
    wire LED_128_Instance_MCS_Instance_1_n19 ;
    wire LED_128_Instance_MCS_Instance_1_n18 ;
    wire LED_128_Instance_MCS_Instance_1_n17 ;
    wire LED_128_Instance_MCS_Instance_1_n16 ;
    wire LED_128_Instance_MCS_Instance_1_n15 ;
    wire LED_128_Instance_MCS_Instance_1_n14 ;
    wire LED_128_Instance_MCS_Instance_1_n13 ;
    wire LED_128_Instance_MCS_Instance_1_n12 ;
    wire LED_128_Instance_MCS_Instance_1_n11 ;
    wire LED_128_Instance_MCS_Instance_1_n10 ;
    wire LED_128_Instance_MCS_Instance_1_n9 ;
    wire LED_128_Instance_MCS_Instance_1_n8 ;
    wire LED_128_Instance_MCS_Instance_1_n7 ;
    wire LED_128_Instance_MCS_Instance_1_n6 ;
    wire LED_128_Instance_MCS_Instance_1_n5 ;
    wire LED_128_Instance_MCS_Instance_1_n4 ;
    wire LED_128_Instance_MCS_Instance_1_n3 ;
    wire LED_128_Instance_MCS_Instance_1_n2 ;
    wire LED_128_Instance_MCS_Instance_1_n1 ;
    wire LED_128_Instance_MCS_Instance_2_n42 ;
    wire LED_128_Instance_MCS_Instance_2_n41 ;
    wire LED_128_Instance_MCS_Instance_2_n40 ;
    wire LED_128_Instance_MCS_Instance_2_n39 ;
    wire LED_128_Instance_MCS_Instance_2_n38 ;
    wire LED_128_Instance_MCS_Instance_2_n37 ;
    wire LED_128_Instance_MCS_Instance_2_n36 ;
    wire LED_128_Instance_MCS_Instance_2_n35 ;
    wire LED_128_Instance_MCS_Instance_2_n34 ;
    wire LED_128_Instance_MCS_Instance_2_n33 ;
    wire LED_128_Instance_MCS_Instance_2_n32 ;
    wire LED_128_Instance_MCS_Instance_2_n31 ;
    wire LED_128_Instance_MCS_Instance_2_n30 ;
    wire LED_128_Instance_MCS_Instance_2_n29 ;
    wire LED_128_Instance_MCS_Instance_2_n28 ;
    wire LED_128_Instance_MCS_Instance_2_n27 ;
    wire LED_128_Instance_MCS_Instance_2_n26 ;
    wire LED_128_Instance_MCS_Instance_2_n25 ;
    wire LED_128_Instance_MCS_Instance_2_n24 ;
    wire LED_128_Instance_MCS_Instance_2_n23 ;
    wire LED_128_Instance_MCS_Instance_2_n22 ;
    wire LED_128_Instance_MCS_Instance_2_n21 ;
    wire LED_128_Instance_MCS_Instance_2_n20 ;
    wire LED_128_Instance_MCS_Instance_2_n19 ;
    wire LED_128_Instance_MCS_Instance_2_n18 ;
    wire LED_128_Instance_MCS_Instance_2_n17 ;
    wire LED_128_Instance_MCS_Instance_2_n16 ;
    wire LED_128_Instance_MCS_Instance_2_n15 ;
    wire LED_128_Instance_MCS_Instance_2_n14 ;
    wire LED_128_Instance_MCS_Instance_2_n13 ;
    wire LED_128_Instance_MCS_Instance_2_n12 ;
    wire LED_128_Instance_MCS_Instance_2_n11 ;
    wire LED_128_Instance_MCS_Instance_2_n10 ;
    wire LED_128_Instance_MCS_Instance_2_n9 ;
    wire LED_128_Instance_MCS_Instance_2_n8 ;
    wire LED_128_Instance_MCS_Instance_2_n7 ;
    wire LED_128_Instance_MCS_Instance_2_n6 ;
    wire LED_128_Instance_MCS_Instance_2_n5 ;
    wire LED_128_Instance_MCS_Instance_2_n4 ;
    wire LED_128_Instance_MCS_Instance_2_n3 ;
    wire LED_128_Instance_MCS_Instance_2_n2 ;
    wire LED_128_Instance_MCS_Instance_2_n1 ;
    wire LED_128_Instance_MCS_Instance_3_n42 ;
    wire LED_128_Instance_MCS_Instance_3_n41 ;
    wire LED_128_Instance_MCS_Instance_3_n40 ;
    wire LED_128_Instance_MCS_Instance_3_n39 ;
    wire LED_128_Instance_MCS_Instance_3_n38 ;
    wire LED_128_Instance_MCS_Instance_3_n37 ;
    wire LED_128_Instance_MCS_Instance_3_n36 ;
    wire LED_128_Instance_MCS_Instance_3_n35 ;
    wire LED_128_Instance_MCS_Instance_3_n34 ;
    wire LED_128_Instance_MCS_Instance_3_n33 ;
    wire LED_128_Instance_MCS_Instance_3_n32 ;
    wire LED_128_Instance_MCS_Instance_3_n31 ;
    wire LED_128_Instance_MCS_Instance_3_n30 ;
    wire LED_128_Instance_MCS_Instance_3_n29 ;
    wire LED_128_Instance_MCS_Instance_3_n28 ;
    wire LED_128_Instance_MCS_Instance_3_n27 ;
    wire LED_128_Instance_MCS_Instance_3_n26 ;
    wire LED_128_Instance_MCS_Instance_3_n25 ;
    wire LED_128_Instance_MCS_Instance_3_n24 ;
    wire LED_128_Instance_MCS_Instance_3_n23 ;
    wire LED_128_Instance_MCS_Instance_3_n22 ;
    wire LED_128_Instance_MCS_Instance_3_n21 ;
    wire LED_128_Instance_MCS_Instance_3_n20 ;
    wire LED_128_Instance_MCS_Instance_3_n19 ;
    wire LED_128_Instance_MCS_Instance_3_n18 ;
    wire LED_128_Instance_MCS_Instance_3_n17 ;
    wire LED_128_Instance_MCS_Instance_3_n16 ;
    wire LED_128_Instance_MCS_Instance_3_n15 ;
    wire LED_128_Instance_MCS_Instance_3_n14 ;
    wire LED_128_Instance_MCS_Instance_3_n13 ;
    wire LED_128_Instance_MCS_Instance_3_n12 ;
    wire LED_128_Instance_MCS_Instance_3_n11 ;
    wire LED_128_Instance_MCS_Instance_3_n10 ;
    wire LED_128_Instance_MCS_Instance_3_n9 ;
    wire LED_128_Instance_MCS_Instance_3_n8 ;
    wire LED_128_Instance_MCS_Instance_3_n7 ;
    wire LED_128_Instance_MCS_Instance_3_n6 ;
    wire LED_128_Instance_MCS_Instance_3_n5 ;
    wire LED_128_Instance_MCS_Instance_3_n4 ;
    wire LED_128_Instance_MCS_Instance_3_n3 ;
    wire LED_128_Instance_MCS_Instance_3_n2 ;
    wire LED_128_Instance_MCS_Instance_3_n1 ;
    wire LED_128_Instance_ks_reg_2__Q ;
    wire [5:0] roundconstant ;
    wire [63:0] LED_128_Instance_subcells_out ;
    wire [63:0] LED_128_Instance_addconst_out ;
    wire [63:0] LED_128_Instance_addroundkey_tmp ;
    wire [63:0] LED_128_Instance_current_roundkey ;
    wire [63:0] LED_128_Instance_state0 ;
    wire [54:3] LED_128_Instance_addroundkey_out ;
    wire [63:0] LED_128_Instance_mixcolumns_out ;

    /* cells in depth 0 */
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) U16 ( .A0_t (roundconstant[5]), .B0_t (roundconstant[1]), .Z0_t (n15) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) U17 ( .A0_t (roundconstant[0]), .B0_t (n15), .Z0_t (n16) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) U18 ( .A0_t (roundconstant[2]), .B0_t (n16), .Z0_t (n17) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) U19 ( .A0_t (roundconstant[3]), .B0_t (n17), .Z0_t (n18) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) U20 ( .A0_t (roundconstant[4]), .B0_t (n18), .Z0_t (n19) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) U21 ( .A0_t (OUT_done), .B0_t (n19), .Z0_t (n20) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) U22 ( .A0_t (IN_reset), .B0_t (n20), .Z0_t (OUT_done) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) LED_128_Instance_U31 ( .A0_t (roundconstant[3]), .B0_t (IN_reset), .Z0_t (roundconstant[4]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) LED_128_Instance_U30 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_n24), .Z0_t (LED_128_Instance_ks_reg_2__Q) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) LED_128_Instance_U29 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_ks_0), .Z0_t (LED_128_Instance_n24) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) LED_128_Instance_U28 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_ks_3_), .Z0_t (LED_128_Instance_ks_0) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) LED_128_Instance_U27 ( .A0_t (roundconstant[4]), .B0_t (IN_reset), .Z0_t (roundconstant[5]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) LED_128_Instance_U26 ( .A0_t (roundconstant[2]), .B0_t (IN_reset), .Z0_t (roundconstant[3]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) LED_128_Instance_U25 ( .A0_t (roundconstant[1]), .B0_t (IN_reset), .Z0_t (roundconstant[2]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) LED_128_Instance_U24 ( .A0_t (roundconstant[0]), .B0_t (IN_reset), .Z0_t (roundconstant[1]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) LED_128_Instance_U23 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_ks_reg_2__Q), .Z0_t (LED_128_Instance_ks_3_) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b1), .NL(1'b1)) LED_128_Instance_U22 ( .A0_t (LED_128_Instance_n29), .B0_t (IN_reset), .Z0_t (roundconstant[0]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) LED_128_Instance_U20 ( .A0_t (roundconstant[5]), .B0_t (roundconstant[4]), .Z0_t (LED_128_Instance_n29) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) LED_128_Instance_U17 ( .A0_t (roundconstant[0]), .B0_t (LED_128_Instance_n19), .Z0_t (LED_128_Instance_n22) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) LED_128_Instance_U16 ( .A0_t (roundconstant[5]), .B0_t (LED_128_Instance_n18), .Z0_t (LED_128_Instance_n19) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) LED_128_Instance_U15 ( .A0_t (LED_128_Instance_n17), .B0_t (LED_128_Instance_n16), .Z0_t (LED_128_Instance_n18) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) LED_128_Instance_U14 ( .A0_t (roundconstant[2]), .B0_t (roundconstant[1]), .Z0_t (LED_128_Instance_n16) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) LED_128_Instance_U13 ( .A0_t (roundconstant[4]), .B0_t (roundconstant[3]), .Z0_t (LED_128_Instance_n17) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) LED_128_Instance_U11 ( .A0_t (LED_128_Instance_n31), .B0_t (LED_128_Instance_n13), .Z0_t (LED_128_Instance_n23) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) LED_128_Instance_U10 ( .A0_t (LED_128_Instance_ks_0), .B0_t (LED_128_Instance_n12), .Z0_t (LED_128_Instance_n13) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) LED_128_Instance_U9 ( .A0_t (LED_128_Instance_ks_3_), .B0_t (LED_128_Instance_n11), .Z0_t (LED_128_Instance_n12) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) LED_128_Instance_U8 ( .A0_t (LED_128_Instance_n24), .B0_t (LED_128_Instance_ks_reg_2__Q), .Z0_t (LED_128_Instance_n11) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) LED_128_Instance_U6 ( .A0_t (LED_128_Instance_ks_0), .B0_t (LED_128_Instance_n9), .Z0_t (LED_128_Instance_n31) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) LED_128_Instance_U5 ( .A0_t (LED_128_Instance_ks_3_), .B0_t (LED_128_Instance_n8), .Z0_t (LED_128_Instance_n9) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) LED_128_Instance_U4 ( .A0_t (LED_128_Instance_n24), .B0_t (LED_128_Instance_ks_reg_2__Q), .Z0_t (LED_128_Instance_n8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_0_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[0]), .B0_t (LED_128_Instance_addconst_out[0]), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_0_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_0_U1_AND1_U1 ( .A0_t (LED_128_Instance_n22), .B0_t (LED_128_Instance_MUX_state0_mux_inst_0_U1_X), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_0_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_0_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_0_U1_Y), .B0_t (LED_128_Instance_mixcolumns_out[0]), .Z0_t (LED_128_Instance_state0[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_1_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[1]), .B0_t (LED_128_Instance_addconst_out[1]), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_1_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_1_U1_AND1_U1 ( .A0_t (LED_128_Instance_n22), .B0_t (LED_128_Instance_MUX_state0_mux_inst_1_U1_X), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_1_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_1_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_1_U1_Y), .B0_t (LED_128_Instance_mixcolumns_out[1]), .Z0_t (LED_128_Instance_state0[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_2_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[2]), .B0_t (LED_128_Instance_addconst_out[2]), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_2_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_2_U1_AND1_U1 ( .A0_t (LED_128_Instance_n22), .B0_t (LED_128_Instance_MUX_state0_mux_inst_2_U1_X), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_2_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_2_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_2_U1_Y), .B0_t (LED_128_Instance_mixcolumns_out[2]), .Z0_t (LED_128_Instance_state0[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_3_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[3]), .B0_t (LED_128_Instance_addroundkey_out[3]), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_3_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_3_U1_AND1_U1 ( .A0_t (LED_128_Instance_n22), .B0_t (LED_128_Instance_MUX_state0_mux_inst_3_U1_X), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_3_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_3_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_3_U1_Y), .B0_t (LED_128_Instance_mixcolumns_out[3]), .Z0_t (LED_128_Instance_state0[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_4_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[4]), .B0_t (LED_128_Instance_addroundkey_out[4]), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_4_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_4_U1_AND1_U1 ( .A0_t (LED_128_Instance_n22), .B0_t (LED_128_Instance_MUX_state0_mux_inst_4_U1_X), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_4_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_4_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_4_U1_Y), .B0_t (LED_128_Instance_mixcolumns_out[4]), .Z0_t (LED_128_Instance_state0[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_5_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[5]), .B0_t (LED_128_Instance_addroundkey_out[5]), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_5_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_5_U1_AND1_U1 ( .A0_t (LED_128_Instance_n22), .B0_t (LED_128_Instance_MUX_state0_mux_inst_5_U1_X), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_5_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_5_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_5_U1_Y), .B0_t (LED_128_Instance_mixcolumns_out[5]), .Z0_t (LED_128_Instance_state0[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_6_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[6]), .B0_t (LED_128_Instance_addroundkey_out[6]), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_6_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_6_U1_AND1_U1 ( .A0_t (LED_128_Instance_n22), .B0_t (LED_128_Instance_MUX_state0_mux_inst_6_U1_X), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_6_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_6_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_6_U1_Y), .B0_t (LED_128_Instance_mixcolumns_out[6]), .Z0_t (LED_128_Instance_state0[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_7_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[7]), .B0_t (LED_128_Instance_addconst_out[7]), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_7_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_7_U1_AND1_U1 ( .A0_t (LED_128_Instance_n22), .B0_t (LED_128_Instance_MUX_state0_mux_inst_7_U1_X), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_7_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_7_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_7_U1_Y), .B0_t (LED_128_Instance_mixcolumns_out[7]), .Z0_t (LED_128_Instance_state0[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_8_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[8]), .B0_t (LED_128_Instance_addconst_out[8]), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_8_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_8_U1_AND1_U1 ( .A0_t (LED_128_Instance_n22), .B0_t (LED_128_Instance_MUX_state0_mux_inst_8_U1_X), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_8_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_8_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_8_U1_Y), .B0_t (LED_128_Instance_mixcolumns_out[8]), .Z0_t (LED_128_Instance_state0[8]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_9_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[9]), .B0_t (LED_128_Instance_addconst_out[9]), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_9_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_9_U1_AND1_U1 ( .A0_t (LED_128_Instance_n22), .B0_t (LED_128_Instance_MUX_state0_mux_inst_9_U1_X), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_9_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_9_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_9_U1_Y), .B0_t (LED_128_Instance_mixcolumns_out[9]), .Z0_t (LED_128_Instance_state0[9]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_10_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[10]), .B0_t (LED_128_Instance_addconst_out[10]), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_10_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_10_U1_AND1_U1 ( .A0_t (LED_128_Instance_n22), .B0_t (LED_128_Instance_MUX_state0_mux_inst_10_U1_X), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_10_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_10_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_10_U1_Y), .B0_t (LED_128_Instance_mixcolumns_out[10]), .Z0_t (LED_128_Instance_state0[10]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_11_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[11]), .B0_t (LED_128_Instance_addconst_out[11]), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_11_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_11_U1_AND1_U1 ( .A0_t (LED_128_Instance_n22), .B0_t (LED_128_Instance_MUX_state0_mux_inst_11_U1_X), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_11_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_11_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_11_U1_Y), .B0_t (LED_128_Instance_mixcolumns_out[11]), .Z0_t (LED_128_Instance_state0[11]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_12_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[12]), .B0_t (LED_128_Instance_addconst_out[12]), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_12_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_12_U1_AND1_U1 ( .A0_t (LED_128_Instance_n22), .B0_t (LED_128_Instance_MUX_state0_mux_inst_12_U1_X), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_12_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_12_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_12_U1_Y), .B0_t (LED_128_Instance_mixcolumns_out[12]), .Z0_t (LED_128_Instance_state0[12]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_13_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[13]), .B0_t (LED_128_Instance_addconst_out[13]), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_13_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_13_U1_AND1_U1 ( .A0_t (LED_128_Instance_n22), .B0_t (LED_128_Instance_MUX_state0_mux_inst_13_U1_X), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_13_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_13_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_13_U1_Y), .B0_t (LED_128_Instance_mixcolumns_out[13]), .Z0_t (LED_128_Instance_state0[13]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_14_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[14]), .B0_t (LED_128_Instance_addconst_out[14]), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_14_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_14_U1_AND1_U1 ( .A0_t (LED_128_Instance_n22), .B0_t (LED_128_Instance_MUX_state0_mux_inst_14_U1_X), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_14_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_14_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_14_U1_Y), .B0_t (LED_128_Instance_mixcolumns_out[14]), .Z0_t (LED_128_Instance_state0[14]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_15_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[15]), .B0_t (LED_128_Instance_addconst_out[15]), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_15_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_15_U1_AND1_U1 ( .A0_t (LED_128_Instance_n22), .B0_t (LED_128_Instance_MUX_state0_mux_inst_15_U1_X), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_15_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_15_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_15_U1_Y), .B0_t (LED_128_Instance_mixcolumns_out[15]), .Z0_t (LED_128_Instance_state0[15]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_16_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[16]), .B0_t (LED_128_Instance_addroundkey_out[16]), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_16_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_16_U1_AND1_U1 ( .A0_t (LED_128_Instance_n22), .B0_t (LED_128_Instance_MUX_state0_mux_inst_16_U1_X), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_16_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_16_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_16_U1_Y), .B0_t (LED_128_Instance_mixcolumns_out[16]), .Z0_t (LED_128_Instance_state0[16]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_17_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[17]), .B0_t (LED_128_Instance_addconst_out[17]), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_17_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_17_U1_AND1_U1 ( .A0_t (LED_128_Instance_n22), .B0_t (LED_128_Instance_MUX_state0_mux_inst_17_U1_X), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_17_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_17_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_17_U1_Y), .B0_t (LED_128_Instance_mixcolumns_out[17]), .Z0_t (LED_128_Instance_state0[17]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_18_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[18]), .B0_t (LED_128_Instance_addconst_out[18]), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_18_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_18_U1_AND1_U1 ( .A0_t (LED_128_Instance_n22), .B0_t (LED_128_Instance_MUX_state0_mux_inst_18_U1_X), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_18_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_18_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_18_U1_Y), .B0_t (LED_128_Instance_mixcolumns_out[18]), .Z0_t (LED_128_Instance_state0[18]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_19_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[19]), .B0_t (LED_128_Instance_addroundkey_out[19]), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_19_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_19_U1_AND1_U1 ( .A0_t (LED_128_Instance_n22), .B0_t (LED_128_Instance_MUX_state0_mux_inst_19_U1_X), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_19_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_19_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_19_U1_Y), .B0_t (LED_128_Instance_mixcolumns_out[19]), .Z0_t (LED_128_Instance_state0[19]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_20_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[20]), .B0_t (LED_128_Instance_addroundkey_out[20]), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_20_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_20_U1_AND1_U1 ( .A0_t (LED_128_Instance_n22), .B0_t (LED_128_Instance_MUX_state0_mux_inst_20_U1_X), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_20_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_20_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_20_U1_Y), .B0_t (LED_128_Instance_mixcolumns_out[20]), .Z0_t (LED_128_Instance_state0[20]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_21_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[21]), .B0_t (LED_128_Instance_addroundkey_out[21]), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_21_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_21_U1_AND1_U1 ( .A0_t (LED_128_Instance_n22), .B0_t (LED_128_Instance_MUX_state0_mux_inst_21_U1_X), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_21_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_21_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_21_U1_Y), .B0_t (LED_128_Instance_mixcolumns_out[21]), .Z0_t (LED_128_Instance_state0[21]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_22_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[22]), .B0_t (LED_128_Instance_addroundkey_out[22]), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_22_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_22_U1_AND1_U1 ( .A0_t (LED_128_Instance_n22), .B0_t (LED_128_Instance_MUX_state0_mux_inst_22_U1_X), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_22_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_22_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_22_U1_Y), .B0_t (LED_128_Instance_mixcolumns_out[22]), .Z0_t (LED_128_Instance_state0[22]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_23_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[23]), .B0_t (LED_128_Instance_addconst_out[23]), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_23_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_23_U1_AND1_U1 ( .A0_t (LED_128_Instance_n22), .B0_t (LED_128_Instance_MUX_state0_mux_inst_23_U1_X), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_23_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_23_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_23_U1_Y), .B0_t (LED_128_Instance_mixcolumns_out[23]), .Z0_t (LED_128_Instance_state0[23]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_24_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[24]), .B0_t (LED_128_Instance_addconst_out[24]), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_24_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_24_U1_AND1_U1 ( .A0_t (LED_128_Instance_n22), .B0_t (LED_128_Instance_MUX_state0_mux_inst_24_U1_X), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_24_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_24_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_24_U1_Y), .B0_t (LED_128_Instance_mixcolumns_out[24]), .Z0_t (LED_128_Instance_state0[24]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_25_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[25]), .B0_t (LED_128_Instance_addconst_out[25]), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_25_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_25_U1_AND1_U1 ( .A0_t (LED_128_Instance_n22), .B0_t (LED_128_Instance_MUX_state0_mux_inst_25_U1_X), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_25_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_25_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_25_U1_Y), .B0_t (LED_128_Instance_mixcolumns_out[25]), .Z0_t (LED_128_Instance_state0[25]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_26_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[26]), .B0_t (LED_128_Instance_addconst_out[26]), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_26_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_26_U1_AND1_U1 ( .A0_t (LED_128_Instance_n22), .B0_t (LED_128_Instance_MUX_state0_mux_inst_26_U1_X), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_26_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_26_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_26_U1_Y), .B0_t (LED_128_Instance_mixcolumns_out[26]), .Z0_t (LED_128_Instance_state0[26]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_27_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[27]), .B0_t (LED_128_Instance_addconst_out[27]), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_27_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_27_U1_AND1_U1 ( .A0_t (LED_128_Instance_n22), .B0_t (LED_128_Instance_MUX_state0_mux_inst_27_U1_X), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_27_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_27_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_27_U1_Y), .B0_t (LED_128_Instance_mixcolumns_out[27]), .Z0_t (LED_128_Instance_state0[27]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_28_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[28]), .B0_t (LED_128_Instance_addconst_out[28]), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_28_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_28_U1_AND1_U1 ( .A0_t (LED_128_Instance_n22), .B0_t (LED_128_Instance_MUX_state0_mux_inst_28_U1_X), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_28_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_28_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_28_U1_Y), .B0_t (LED_128_Instance_mixcolumns_out[28]), .Z0_t (LED_128_Instance_state0[28]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_29_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[29]), .B0_t (LED_128_Instance_addconst_out[29]), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_29_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_29_U1_AND1_U1 ( .A0_t (LED_128_Instance_n22), .B0_t (LED_128_Instance_MUX_state0_mux_inst_29_U1_X), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_29_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_29_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_29_U1_Y), .B0_t (LED_128_Instance_mixcolumns_out[29]), .Z0_t (LED_128_Instance_state0[29]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_30_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[30]), .B0_t (LED_128_Instance_addconst_out[30]), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_30_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_30_U1_AND1_U1 ( .A0_t (LED_128_Instance_n22), .B0_t (LED_128_Instance_MUX_state0_mux_inst_30_U1_X), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_30_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_30_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_30_U1_Y), .B0_t (LED_128_Instance_mixcolumns_out[30]), .Z0_t (LED_128_Instance_state0[30]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_31_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[31]), .B0_t (LED_128_Instance_addconst_out[31]), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_31_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_31_U1_AND1_U1 ( .A0_t (LED_128_Instance_n22), .B0_t (LED_128_Instance_MUX_state0_mux_inst_31_U1_X), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_31_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_31_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_31_U1_Y), .B0_t (LED_128_Instance_mixcolumns_out[31]), .Z0_t (LED_128_Instance_state0[31]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_32_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[32]), .B0_t (LED_128_Instance_addconst_out[32]), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_32_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_32_U1_AND1_U1 ( .A0_t (LED_128_Instance_n22), .B0_t (LED_128_Instance_MUX_state0_mux_inst_32_U1_X), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_32_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_32_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_32_U1_Y), .B0_t (LED_128_Instance_mixcolumns_out[32]), .Z0_t (LED_128_Instance_state0[32]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_33_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[33]), .B0_t (LED_128_Instance_addroundkey_out[33]), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_33_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_33_U1_AND1_U1 ( .A0_t (LED_128_Instance_n22), .B0_t (LED_128_Instance_MUX_state0_mux_inst_33_U1_X), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_33_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_33_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_33_U1_Y), .B0_t (LED_128_Instance_mixcolumns_out[33]), .Z0_t (LED_128_Instance_state0[33]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_34_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[34]), .B0_t (LED_128_Instance_addconst_out[34]), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_34_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_34_U1_AND1_U1 ( .A0_t (LED_128_Instance_n22), .B0_t (LED_128_Instance_MUX_state0_mux_inst_34_U1_X), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_34_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_34_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_34_U1_Y), .B0_t (LED_128_Instance_mixcolumns_out[34]), .Z0_t (LED_128_Instance_state0[34]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_35_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[35]), .B0_t (LED_128_Instance_addconst_out[35]), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_35_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_35_U1_AND1_U1 ( .A0_t (LED_128_Instance_n22), .B0_t (LED_128_Instance_MUX_state0_mux_inst_35_U1_X), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_35_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_35_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_35_U1_Y), .B0_t (LED_128_Instance_mixcolumns_out[35]), .Z0_t (LED_128_Instance_state0[35]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_36_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[36]), .B0_t (LED_128_Instance_addroundkey_out[36]), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_36_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_36_U1_AND1_U1 ( .A0_t (LED_128_Instance_n22), .B0_t (LED_128_Instance_MUX_state0_mux_inst_36_U1_X), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_36_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_36_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_36_U1_Y), .B0_t (LED_128_Instance_mixcolumns_out[36]), .Z0_t (LED_128_Instance_state0[36]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_37_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[37]), .B0_t (LED_128_Instance_addroundkey_out[37]), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_37_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_37_U1_AND1_U1 ( .A0_t (LED_128_Instance_n22), .B0_t (LED_128_Instance_MUX_state0_mux_inst_37_U1_X), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_37_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_37_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_37_U1_Y), .B0_t (LED_128_Instance_mixcolumns_out[37]), .Z0_t (LED_128_Instance_state0[37]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_38_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[38]), .B0_t (LED_128_Instance_addroundkey_out[38]), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_38_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_38_U1_AND1_U1 ( .A0_t (LED_128_Instance_n22), .B0_t (LED_128_Instance_MUX_state0_mux_inst_38_U1_X), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_38_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_38_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_38_U1_Y), .B0_t (LED_128_Instance_mixcolumns_out[38]), .Z0_t (LED_128_Instance_state0[38]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_39_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[39]), .B0_t (LED_128_Instance_addconst_out[39]), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_39_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_39_U1_AND1_U1 ( .A0_t (LED_128_Instance_n22), .B0_t (LED_128_Instance_MUX_state0_mux_inst_39_U1_X), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_39_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_39_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_39_U1_Y), .B0_t (LED_128_Instance_mixcolumns_out[39]), .Z0_t (LED_128_Instance_state0[39]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_40_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[40]), .B0_t (LED_128_Instance_addconst_out[40]), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_40_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_40_U1_AND1_U1 ( .A0_t (LED_128_Instance_n22), .B0_t (LED_128_Instance_MUX_state0_mux_inst_40_U1_X), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_40_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_40_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_40_U1_Y), .B0_t (LED_128_Instance_mixcolumns_out[40]), .Z0_t (LED_128_Instance_state0[40]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_41_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[41]), .B0_t (LED_128_Instance_addconst_out[41]), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_41_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_41_U1_AND1_U1 ( .A0_t (LED_128_Instance_n22), .B0_t (LED_128_Instance_MUX_state0_mux_inst_41_U1_X), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_41_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_41_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_41_U1_Y), .B0_t (LED_128_Instance_mixcolumns_out[41]), .Z0_t (LED_128_Instance_state0[41]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_42_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[42]), .B0_t (LED_128_Instance_addconst_out[42]), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_42_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_42_U1_AND1_U1 ( .A0_t (LED_128_Instance_n22), .B0_t (LED_128_Instance_MUX_state0_mux_inst_42_U1_X), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_42_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_42_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_42_U1_Y), .B0_t (LED_128_Instance_mixcolumns_out[42]), .Z0_t (LED_128_Instance_state0[42]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_43_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[43]), .B0_t (LED_128_Instance_addconst_out[43]), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_43_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_43_U1_AND1_U1 ( .A0_t (LED_128_Instance_n22), .B0_t (LED_128_Instance_MUX_state0_mux_inst_43_U1_X), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_43_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_43_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_43_U1_Y), .B0_t (LED_128_Instance_mixcolumns_out[43]), .Z0_t (LED_128_Instance_state0[43]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_44_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[44]), .B0_t (LED_128_Instance_addconst_out[44]), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_44_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_44_U1_AND1_U1 ( .A0_t (LED_128_Instance_n22), .B0_t (LED_128_Instance_MUX_state0_mux_inst_44_U1_X), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_44_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_44_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_44_U1_Y), .B0_t (LED_128_Instance_mixcolumns_out[44]), .Z0_t (LED_128_Instance_state0[44]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_45_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[45]), .B0_t (LED_128_Instance_addconst_out[45]), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_45_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_45_U1_AND1_U1 ( .A0_t (LED_128_Instance_n22), .B0_t (LED_128_Instance_MUX_state0_mux_inst_45_U1_X), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_45_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_45_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_45_U1_Y), .B0_t (LED_128_Instance_mixcolumns_out[45]), .Z0_t (LED_128_Instance_state0[45]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_46_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[46]), .B0_t (LED_128_Instance_addconst_out[46]), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_46_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_46_U1_AND1_U1 ( .A0_t (LED_128_Instance_n22), .B0_t (LED_128_Instance_MUX_state0_mux_inst_46_U1_X), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_46_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_46_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_46_U1_Y), .B0_t (LED_128_Instance_mixcolumns_out[46]), .Z0_t (LED_128_Instance_state0[46]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_47_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[47]), .B0_t (LED_128_Instance_addconst_out[47]), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_47_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_47_U1_AND1_U1 ( .A0_t (LED_128_Instance_n22), .B0_t (LED_128_Instance_MUX_state0_mux_inst_47_U1_X), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_47_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_47_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_47_U1_Y), .B0_t (LED_128_Instance_mixcolumns_out[47]), .Z0_t (LED_128_Instance_state0[47]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_48_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[48]), .B0_t (LED_128_Instance_addroundkey_out[48]), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_48_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_48_U1_AND1_U1 ( .A0_t (LED_128_Instance_n22), .B0_t (LED_128_Instance_MUX_state0_mux_inst_48_U1_X), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_48_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_48_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_48_U1_Y), .B0_t (LED_128_Instance_mixcolumns_out[48]), .Z0_t (LED_128_Instance_state0[48]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_49_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[49]), .B0_t (LED_128_Instance_addroundkey_out[49]), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_49_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_49_U1_AND1_U1 ( .A0_t (LED_128_Instance_n22), .B0_t (LED_128_Instance_MUX_state0_mux_inst_49_U1_X), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_49_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_49_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_49_U1_Y), .B0_t (LED_128_Instance_mixcolumns_out[49]), .Z0_t (LED_128_Instance_state0[49]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_50_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[50]), .B0_t (LED_128_Instance_addconst_out[50]), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_50_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_50_U1_AND1_U1 ( .A0_t (LED_128_Instance_n22), .B0_t (LED_128_Instance_MUX_state0_mux_inst_50_U1_X), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_50_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_50_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_50_U1_Y), .B0_t (LED_128_Instance_mixcolumns_out[50]), .Z0_t (LED_128_Instance_state0[50]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_51_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[51]), .B0_t (LED_128_Instance_addconst_out[51]), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_51_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_51_U1_AND1_U1 ( .A0_t (LED_128_Instance_n22), .B0_t (LED_128_Instance_MUX_state0_mux_inst_51_U1_X), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_51_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_51_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_51_U1_Y), .B0_t (LED_128_Instance_mixcolumns_out[51]), .Z0_t (LED_128_Instance_state0[51]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_52_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[52]), .B0_t (LED_128_Instance_addroundkey_out[52]), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_52_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_52_U1_AND1_U1 ( .A0_t (LED_128_Instance_n22), .B0_t (LED_128_Instance_MUX_state0_mux_inst_52_U1_X), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_52_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_52_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_52_U1_Y), .B0_t (LED_128_Instance_mixcolumns_out[52]), .Z0_t (LED_128_Instance_state0[52]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_53_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[53]), .B0_t (LED_128_Instance_addroundkey_out[53]), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_53_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_53_U1_AND1_U1 ( .A0_t (LED_128_Instance_n22), .B0_t (LED_128_Instance_MUX_state0_mux_inst_53_U1_X), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_53_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_53_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_53_U1_Y), .B0_t (LED_128_Instance_mixcolumns_out[53]), .Z0_t (LED_128_Instance_state0[53]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_54_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[54]), .B0_t (LED_128_Instance_addroundkey_out[54]), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_54_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_54_U1_AND1_U1 ( .A0_t (LED_128_Instance_n22), .B0_t (LED_128_Instance_MUX_state0_mux_inst_54_U1_X), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_54_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_54_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_54_U1_Y), .B0_t (LED_128_Instance_mixcolumns_out[54]), .Z0_t (LED_128_Instance_state0[54]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_55_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[55]), .B0_t (LED_128_Instance_addconst_out[55]), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_55_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_55_U1_AND1_U1 ( .A0_t (LED_128_Instance_n22), .B0_t (LED_128_Instance_MUX_state0_mux_inst_55_U1_X), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_55_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_55_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_55_U1_Y), .B0_t (LED_128_Instance_mixcolumns_out[55]), .Z0_t (LED_128_Instance_state0[55]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_56_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[56]), .B0_t (LED_128_Instance_addconst_out[56]), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_56_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_56_U1_AND1_U1 ( .A0_t (LED_128_Instance_n22), .B0_t (LED_128_Instance_MUX_state0_mux_inst_56_U1_X), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_56_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_56_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_56_U1_Y), .B0_t (LED_128_Instance_mixcolumns_out[56]), .Z0_t (LED_128_Instance_state0[56]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_57_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[57]), .B0_t (LED_128_Instance_addconst_out[57]), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_57_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_57_U1_AND1_U1 ( .A0_t (LED_128_Instance_n22), .B0_t (LED_128_Instance_MUX_state0_mux_inst_57_U1_X), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_57_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_57_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_57_U1_Y), .B0_t (LED_128_Instance_mixcolumns_out[57]), .Z0_t (LED_128_Instance_state0[57]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_58_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[58]), .B0_t (LED_128_Instance_addconst_out[58]), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_58_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_58_U1_AND1_U1 ( .A0_t (LED_128_Instance_n22), .B0_t (LED_128_Instance_MUX_state0_mux_inst_58_U1_X), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_58_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_58_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_58_U1_Y), .B0_t (LED_128_Instance_mixcolumns_out[58]), .Z0_t (LED_128_Instance_state0[58]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_59_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[59]), .B0_t (LED_128_Instance_addconst_out[59]), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_59_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_59_U1_AND1_U1 ( .A0_t (LED_128_Instance_n22), .B0_t (LED_128_Instance_MUX_state0_mux_inst_59_U1_X), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_59_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_59_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_59_U1_Y), .B0_t (LED_128_Instance_mixcolumns_out[59]), .Z0_t (LED_128_Instance_state0[59]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_60_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[60]), .B0_t (LED_128_Instance_addconst_out[60]), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_60_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_60_U1_AND1_U1 ( .A0_t (LED_128_Instance_n22), .B0_t (LED_128_Instance_MUX_state0_mux_inst_60_U1_X), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_60_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_60_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_60_U1_Y), .B0_t (LED_128_Instance_mixcolumns_out[60]), .Z0_t (LED_128_Instance_state0[60]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_61_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[61]), .B0_t (LED_128_Instance_addconst_out[61]), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_61_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_61_U1_AND1_U1 ( .A0_t (LED_128_Instance_n22), .B0_t (LED_128_Instance_MUX_state0_mux_inst_61_U1_X), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_61_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_61_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_61_U1_Y), .B0_t (LED_128_Instance_mixcolumns_out[61]), .Z0_t (LED_128_Instance_state0[61]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_62_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[62]), .B0_t (LED_128_Instance_addconst_out[62]), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_62_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_62_U1_AND1_U1 ( .A0_t (LED_128_Instance_n22), .B0_t (LED_128_Instance_MUX_state0_mux_inst_62_U1_X), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_62_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_62_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_62_U1_Y), .B0_t (LED_128_Instance_mixcolumns_out[62]), .Z0_t (LED_128_Instance_state0[62]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_63_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[63]), .B0_t (LED_128_Instance_addconst_out[63]), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_63_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_63_U1_AND1_U1 ( .A0_t (LED_128_Instance_n22), .B0_t (LED_128_Instance_MUX_state0_mux_inst_63_U1_X), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_63_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_63_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_63_U1_Y), .B0_t (LED_128_Instance_mixcolumns_out[63]), .Z0_t (LED_128_Instance_state0[63]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_0_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[0]), .B0_t (IN_plaintext[0]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_0_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_0_U1_AND1_U1 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_MUX_state1_mux_inst_0_U1_X), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_0_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_0_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_0_U1_Y), .B0_t (LED_128_Instance_state0[0]), .Z0_t (OUT_ciphertext[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_1_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[1]), .B0_t (IN_plaintext[1]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_1_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_1_U1_AND1_U1 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_MUX_state1_mux_inst_1_U1_X), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_1_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_1_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_1_U1_Y), .B0_t (LED_128_Instance_state0[1]), .Z0_t (OUT_ciphertext[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_2_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[2]), .B0_t (IN_plaintext[2]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_2_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_2_U1_AND1_U1 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_MUX_state1_mux_inst_2_U1_X), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_2_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_2_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_2_U1_Y), .B0_t (LED_128_Instance_state0[2]), .Z0_t (OUT_ciphertext[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_3_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[3]), .B0_t (IN_plaintext[3]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_3_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_3_U1_AND1_U1 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_MUX_state1_mux_inst_3_U1_X), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_3_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_3_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_3_U1_Y), .B0_t (LED_128_Instance_state0[3]), .Z0_t (OUT_ciphertext[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_4_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[4]), .B0_t (IN_plaintext[4]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_4_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_4_U1_AND1_U1 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_MUX_state1_mux_inst_4_U1_X), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_4_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_4_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_4_U1_Y), .B0_t (LED_128_Instance_state0[4]), .Z0_t (OUT_ciphertext[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_5_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[5]), .B0_t (IN_plaintext[5]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_5_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_5_U1_AND1_U1 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_MUX_state1_mux_inst_5_U1_X), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_5_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_5_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_5_U1_Y), .B0_t (LED_128_Instance_state0[5]), .Z0_t (OUT_ciphertext[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_6_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[6]), .B0_t (IN_plaintext[6]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_6_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_6_U1_AND1_U1 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_MUX_state1_mux_inst_6_U1_X), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_6_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_6_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_6_U1_Y), .B0_t (LED_128_Instance_state0[6]), .Z0_t (OUT_ciphertext[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_7_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[7]), .B0_t (IN_plaintext[7]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_7_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_7_U1_AND1_U1 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_MUX_state1_mux_inst_7_U1_X), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_7_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_7_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_7_U1_Y), .B0_t (LED_128_Instance_state0[7]), .Z0_t (OUT_ciphertext[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_8_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[8]), .B0_t (IN_plaintext[8]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_8_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_8_U1_AND1_U1 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_MUX_state1_mux_inst_8_U1_X), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_8_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_8_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_8_U1_Y), .B0_t (LED_128_Instance_state0[8]), .Z0_t (OUT_ciphertext[8]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_9_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[9]), .B0_t (IN_plaintext[9]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_9_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_9_U1_AND1_U1 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_MUX_state1_mux_inst_9_U1_X), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_9_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_9_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_9_U1_Y), .B0_t (LED_128_Instance_state0[9]), .Z0_t (OUT_ciphertext[9]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_10_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[10]), .B0_t (IN_plaintext[10]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_10_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_10_U1_AND1_U1 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_MUX_state1_mux_inst_10_U1_X), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_10_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_10_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_10_U1_Y), .B0_t (LED_128_Instance_state0[10]), .Z0_t (OUT_ciphertext[10]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_11_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[11]), .B0_t (IN_plaintext[11]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_11_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_11_U1_AND1_U1 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_MUX_state1_mux_inst_11_U1_X), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_11_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_11_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_11_U1_Y), .B0_t (LED_128_Instance_state0[11]), .Z0_t (OUT_ciphertext[11]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_12_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[12]), .B0_t (IN_plaintext[12]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_12_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_12_U1_AND1_U1 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_MUX_state1_mux_inst_12_U1_X), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_12_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_12_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_12_U1_Y), .B0_t (LED_128_Instance_state0[12]), .Z0_t (OUT_ciphertext[12]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_13_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[13]), .B0_t (IN_plaintext[13]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_13_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_13_U1_AND1_U1 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_MUX_state1_mux_inst_13_U1_X), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_13_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_13_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_13_U1_Y), .B0_t (LED_128_Instance_state0[13]), .Z0_t (OUT_ciphertext[13]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_14_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[14]), .B0_t (IN_plaintext[14]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_14_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_14_U1_AND1_U1 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_MUX_state1_mux_inst_14_U1_X), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_14_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_14_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_14_U1_Y), .B0_t (LED_128_Instance_state0[14]), .Z0_t (OUT_ciphertext[14]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_15_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[15]), .B0_t (IN_plaintext[15]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_15_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_15_U1_AND1_U1 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_MUX_state1_mux_inst_15_U1_X), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_15_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_15_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_15_U1_Y), .B0_t (LED_128_Instance_state0[15]), .Z0_t (OUT_ciphertext[15]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_16_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[16]), .B0_t (IN_plaintext[16]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_16_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_16_U1_AND1_U1 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_MUX_state1_mux_inst_16_U1_X), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_16_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_16_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_16_U1_Y), .B0_t (LED_128_Instance_state0[16]), .Z0_t (OUT_ciphertext[16]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_17_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[17]), .B0_t (IN_plaintext[17]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_17_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_17_U1_AND1_U1 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_MUX_state1_mux_inst_17_U1_X), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_17_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_17_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_17_U1_Y), .B0_t (LED_128_Instance_state0[17]), .Z0_t (OUT_ciphertext[17]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_18_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[18]), .B0_t (IN_plaintext[18]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_18_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_18_U1_AND1_U1 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_MUX_state1_mux_inst_18_U1_X), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_18_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_18_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_18_U1_Y), .B0_t (LED_128_Instance_state0[18]), .Z0_t (OUT_ciphertext[18]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_19_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[19]), .B0_t (IN_plaintext[19]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_19_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_19_U1_AND1_U1 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_MUX_state1_mux_inst_19_U1_X), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_19_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_19_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_19_U1_Y), .B0_t (LED_128_Instance_state0[19]), .Z0_t (OUT_ciphertext[19]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_20_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[20]), .B0_t (IN_plaintext[20]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_20_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_20_U1_AND1_U1 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_MUX_state1_mux_inst_20_U1_X), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_20_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_20_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_20_U1_Y), .B0_t (LED_128_Instance_state0[20]), .Z0_t (OUT_ciphertext[20]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_21_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[21]), .B0_t (IN_plaintext[21]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_21_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_21_U1_AND1_U1 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_MUX_state1_mux_inst_21_U1_X), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_21_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_21_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_21_U1_Y), .B0_t (LED_128_Instance_state0[21]), .Z0_t (OUT_ciphertext[21]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_22_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[22]), .B0_t (IN_plaintext[22]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_22_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_22_U1_AND1_U1 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_MUX_state1_mux_inst_22_U1_X), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_22_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_22_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_22_U1_Y), .B0_t (LED_128_Instance_state0[22]), .Z0_t (OUT_ciphertext[22]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_23_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[23]), .B0_t (IN_plaintext[23]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_23_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_23_U1_AND1_U1 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_MUX_state1_mux_inst_23_U1_X), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_23_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_23_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_23_U1_Y), .B0_t (LED_128_Instance_state0[23]), .Z0_t (OUT_ciphertext[23]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_24_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[24]), .B0_t (IN_plaintext[24]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_24_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_24_U1_AND1_U1 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_MUX_state1_mux_inst_24_U1_X), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_24_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_24_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_24_U1_Y), .B0_t (LED_128_Instance_state0[24]), .Z0_t (OUT_ciphertext[24]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_25_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[25]), .B0_t (IN_plaintext[25]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_25_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_25_U1_AND1_U1 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_MUX_state1_mux_inst_25_U1_X), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_25_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_25_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_25_U1_Y), .B0_t (LED_128_Instance_state0[25]), .Z0_t (OUT_ciphertext[25]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_26_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[26]), .B0_t (IN_plaintext[26]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_26_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_26_U1_AND1_U1 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_MUX_state1_mux_inst_26_U1_X), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_26_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_26_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_26_U1_Y), .B0_t (LED_128_Instance_state0[26]), .Z0_t (OUT_ciphertext[26]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_27_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[27]), .B0_t (IN_plaintext[27]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_27_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_27_U1_AND1_U1 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_MUX_state1_mux_inst_27_U1_X), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_27_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_27_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_27_U1_Y), .B0_t (LED_128_Instance_state0[27]), .Z0_t (OUT_ciphertext[27]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_28_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[28]), .B0_t (IN_plaintext[28]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_28_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_28_U1_AND1_U1 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_MUX_state1_mux_inst_28_U1_X), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_28_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_28_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_28_U1_Y), .B0_t (LED_128_Instance_state0[28]), .Z0_t (OUT_ciphertext[28]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_29_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[29]), .B0_t (IN_plaintext[29]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_29_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_29_U1_AND1_U1 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_MUX_state1_mux_inst_29_U1_X), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_29_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_29_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_29_U1_Y), .B0_t (LED_128_Instance_state0[29]), .Z0_t (OUT_ciphertext[29]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_30_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[30]), .B0_t (IN_plaintext[30]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_30_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_30_U1_AND1_U1 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_MUX_state1_mux_inst_30_U1_X), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_30_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_30_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_30_U1_Y), .B0_t (LED_128_Instance_state0[30]), .Z0_t (OUT_ciphertext[30]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_31_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[31]), .B0_t (IN_plaintext[31]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_31_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_31_U1_AND1_U1 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_MUX_state1_mux_inst_31_U1_X), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_31_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_31_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_31_U1_Y), .B0_t (LED_128_Instance_state0[31]), .Z0_t (OUT_ciphertext[31]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_32_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[32]), .B0_t (IN_plaintext[32]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_32_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_32_U1_AND1_U1 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_MUX_state1_mux_inst_32_U1_X), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_32_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_32_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_32_U1_Y), .B0_t (LED_128_Instance_state0[32]), .Z0_t (OUT_ciphertext[32]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_33_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[33]), .B0_t (IN_plaintext[33]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_33_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_33_U1_AND1_U1 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_MUX_state1_mux_inst_33_U1_X), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_33_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_33_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_33_U1_Y), .B0_t (LED_128_Instance_state0[33]), .Z0_t (OUT_ciphertext[33]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_34_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[34]), .B0_t (IN_plaintext[34]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_34_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_34_U1_AND1_U1 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_MUX_state1_mux_inst_34_U1_X), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_34_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_34_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_34_U1_Y), .B0_t (LED_128_Instance_state0[34]), .Z0_t (OUT_ciphertext[34]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_35_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[35]), .B0_t (IN_plaintext[35]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_35_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_35_U1_AND1_U1 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_MUX_state1_mux_inst_35_U1_X), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_35_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_35_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_35_U1_Y), .B0_t (LED_128_Instance_state0[35]), .Z0_t (OUT_ciphertext[35]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_36_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[36]), .B0_t (IN_plaintext[36]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_36_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_36_U1_AND1_U1 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_MUX_state1_mux_inst_36_U1_X), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_36_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_36_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_36_U1_Y), .B0_t (LED_128_Instance_state0[36]), .Z0_t (OUT_ciphertext[36]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_37_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[37]), .B0_t (IN_plaintext[37]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_37_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_37_U1_AND1_U1 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_MUX_state1_mux_inst_37_U1_X), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_37_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_37_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_37_U1_Y), .B0_t (LED_128_Instance_state0[37]), .Z0_t (OUT_ciphertext[37]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_38_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[38]), .B0_t (IN_plaintext[38]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_38_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_38_U1_AND1_U1 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_MUX_state1_mux_inst_38_U1_X), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_38_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_38_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_38_U1_Y), .B0_t (LED_128_Instance_state0[38]), .Z0_t (OUT_ciphertext[38]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_39_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[39]), .B0_t (IN_plaintext[39]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_39_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_39_U1_AND1_U1 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_MUX_state1_mux_inst_39_U1_X), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_39_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_39_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_39_U1_Y), .B0_t (LED_128_Instance_state0[39]), .Z0_t (OUT_ciphertext[39]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_40_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[40]), .B0_t (IN_plaintext[40]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_40_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_40_U1_AND1_U1 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_MUX_state1_mux_inst_40_U1_X), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_40_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_40_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_40_U1_Y), .B0_t (LED_128_Instance_state0[40]), .Z0_t (OUT_ciphertext[40]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_41_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[41]), .B0_t (IN_plaintext[41]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_41_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_41_U1_AND1_U1 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_MUX_state1_mux_inst_41_U1_X), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_41_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_41_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_41_U1_Y), .B0_t (LED_128_Instance_state0[41]), .Z0_t (OUT_ciphertext[41]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_42_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[42]), .B0_t (IN_plaintext[42]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_42_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_42_U1_AND1_U1 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_MUX_state1_mux_inst_42_U1_X), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_42_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_42_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_42_U1_Y), .B0_t (LED_128_Instance_state0[42]), .Z0_t (OUT_ciphertext[42]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_43_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[43]), .B0_t (IN_plaintext[43]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_43_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_43_U1_AND1_U1 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_MUX_state1_mux_inst_43_U1_X), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_43_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_43_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_43_U1_Y), .B0_t (LED_128_Instance_state0[43]), .Z0_t (OUT_ciphertext[43]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_44_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[44]), .B0_t (IN_plaintext[44]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_44_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_44_U1_AND1_U1 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_MUX_state1_mux_inst_44_U1_X), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_44_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_44_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_44_U1_Y), .B0_t (LED_128_Instance_state0[44]), .Z0_t (OUT_ciphertext[44]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_45_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[45]), .B0_t (IN_plaintext[45]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_45_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_45_U1_AND1_U1 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_MUX_state1_mux_inst_45_U1_X), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_45_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_45_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_45_U1_Y), .B0_t (LED_128_Instance_state0[45]), .Z0_t (OUT_ciphertext[45]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_46_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[46]), .B0_t (IN_plaintext[46]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_46_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_46_U1_AND1_U1 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_MUX_state1_mux_inst_46_U1_X), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_46_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_46_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_46_U1_Y), .B0_t (LED_128_Instance_state0[46]), .Z0_t (OUT_ciphertext[46]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_47_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[47]), .B0_t (IN_plaintext[47]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_47_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_47_U1_AND1_U1 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_MUX_state1_mux_inst_47_U1_X), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_47_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_47_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_47_U1_Y), .B0_t (LED_128_Instance_state0[47]), .Z0_t (OUT_ciphertext[47]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_48_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[48]), .B0_t (IN_plaintext[48]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_48_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_48_U1_AND1_U1 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_MUX_state1_mux_inst_48_U1_X), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_48_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_48_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_48_U1_Y), .B0_t (LED_128_Instance_state0[48]), .Z0_t (OUT_ciphertext[48]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_49_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[49]), .B0_t (IN_plaintext[49]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_49_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_49_U1_AND1_U1 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_MUX_state1_mux_inst_49_U1_X), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_49_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_49_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_49_U1_Y), .B0_t (LED_128_Instance_state0[49]), .Z0_t (OUT_ciphertext[49]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_50_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[50]), .B0_t (IN_plaintext[50]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_50_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_50_U1_AND1_U1 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_MUX_state1_mux_inst_50_U1_X), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_50_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_50_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_50_U1_Y), .B0_t (LED_128_Instance_state0[50]), .Z0_t (OUT_ciphertext[50]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_51_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[51]), .B0_t (IN_plaintext[51]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_51_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_51_U1_AND1_U1 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_MUX_state1_mux_inst_51_U1_X), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_51_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_51_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_51_U1_Y), .B0_t (LED_128_Instance_state0[51]), .Z0_t (OUT_ciphertext[51]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_52_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[52]), .B0_t (IN_plaintext[52]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_52_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_52_U1_AND1_U1 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_MUX_state1_mux_inst_52_U1_X), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_52_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_52_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_52_U1_Y), .B0_t (LED_128_Instance_state0[52]), .Z0_t (OUT_ciphertext[52]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_53_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[53]), .B0_t (IN_plaintext[53]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_53_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_53_U1_AND1_U1 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_MUX_state1_mux_inst_53_U1_X), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_53_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_53_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_53_U1_Y), .B0_t (LED_128_Instance_state0[53]), .Z0_t (OUT_ciphertext[53]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_54_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[54]), .B0_t (IN_plaintext[54]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_54_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_54_U1_AND1_U1 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_MUX_state1_mux_inst_54_U1_X), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_54_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_54_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_54_U1_Y), .B0_t (LED_128_Instance_state0[54]), .Z0_t (OUT_ciphertext[54]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_55_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[55]), .B0_t (IN_plaintext[55]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_55_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_55_U1_AND1_U1 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_MUX_state1_mux_inst_55_U1_X), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_55_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_55_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_55_U1_Y), .B0_t (LED_128_Instance_state0[55]), .Z0_t (OUT_ciphertext[55]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_56_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[56]), .B0_t (IN_plaintext[56]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_56_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_56_U1_AND1_U1 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_MUX_state1_mux_inst_56_U1_X), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_56_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_56_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_56_U1_Y), .B0_t (LED_128_Instance_state0[56]), .Z0_t (OUT_ciphertext[56]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_57_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[57]), .B0_t (IN_plaintext[57]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_57_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_57_U1_AND1_U1 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_MUX_state1_mux_inst_57_U1_X), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_57_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_57_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_57_U1_Y), .B0_t (LED_128_Instance_state0[57]), .Z0_t (OUT_ciphertext[57]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_58_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[58]), .B0_t (IN_plaintext[58]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_58_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_58_U1_AND1_U1 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_MUX_state1_mux_inst_58_U1_X), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_58_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_58_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_58_U1_Y), .B0_t (LED_128_Instance_state0[58]), .Z0_t (OUT_ciphertext[58]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_59_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[59]), .B0_t (IN_plaintext[59]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_59_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_59_U1_AND1_U1 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_MUX_state1_mux_inst_59_U1_X), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_59_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_59_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_59_U1_Y), .B0_t (LED_128_Instance_state0[59]), .Z0_t (OUT_ciphertext[59]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_60_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[60]), .B0_t (IN_plaintext[60]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_60_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_60_U1_AND1_U1 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_MUX_state1_mux_inst_60_U1_X), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_60_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_60_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_60_U1_Y), .B0_t (LED_128_Instance_state0[60]), .Z0_t (OUT_ciphertext[60]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_61_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[61]), .B0_t (IN_plaintext[61]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_61_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_61_U1_AND1_U1 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_MUX_state1_mux_inst_61_U1_X), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_61_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_61_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_61_U1_Y), .B0_t (LED_128_Instance_state0[61]), .Z0_t (OUT_ciphertext[61]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_62_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[62]), .B0_t (IN_plaintext[62]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_62_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_62_U1_AND1_U1 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_MUX_state1_mux_inst_62_U1_X), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_62_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_62_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_62_U1_Y), .B0_t (LED_128_Instance_state0[62]), .Z0_t (OUT_ciphertext[62]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_63_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[63]), .B0_t (IN_plaintext[63]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_63_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_63_U1_AND1_U1 ( .A0_t (IN_reset), .B0_t (LED_128_Instance_MUX_state1_mux_inst_63_U1_X), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_63_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_63_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_63_U1_Y), .B0_t (LED_128_Instance_state0[63]), .Z0_t (OUT_ciphertext[63]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_0_U1_XOR1_U1 ( .A0_t (IN_key[64]), .B0_t (IN_key[0]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_0_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_0_U1_AND1_U1 ( .A0_t (LED_128_Instance_n31), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_0_U1_X), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_0_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_0_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_0_U1_Y), .B0_t (IN_key[64]), .Z0_t (LED_128_Instance_current_roundkey[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_1_U1_XOR1_U1 ( .A0_t (IN_key[65]), .B0_t (IN_key[1]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_1_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_1_U1_AND1_U1 ( .A0_t (LED_128_Instance_n31), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_1_U1_X), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_1_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_1_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_1_U1_Y), .B0_t (IN_key[65]), .Z0_t (LED_128_Instance_current_roundkey[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_2_U1_XOR1_U1 ( .A0_t (IN_key[66]), .B0_t (IN_key[2]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_2_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_2_U1_AND1_U1 ( .A0_t (LED_128_Instance_n31), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_2_U1_X), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_2_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_2_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_2_U1_Y), .B0_t (IN_key[66]), .Z0_t (LED_128_Instance_current_roundkey[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_3_U1_XOR1_U1 ( .A0_t (IN_key[67]), .B0_t (IN_key[3]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_3_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_3_U1_AND1_U1 ( .A0_t (LED_128_Instance_n31), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_3_U1_X), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_3_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_3_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_3_U1_Y), .B0_t (IN_key[67]), .Z0_t (LED_128_Instance_current_roundkey[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_4_U1_XOR1_U1 ( .A0_t (IN_key[68]), .B0_t (IN_key[4]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_4_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_4_U1_AND1_U1 ( .A0_t (LED_128_Instance_n31), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_4_U1_X), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_4_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_4_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_4_U1_Y), .B0_t (IN_key[68]), .Z0_t (LED_128_Instance_current_roundkey[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_5_U1_XOR1_U1 ( .A0_t (IN_key[69]), .B0_t (IN_key[5]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_5_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_5_U1_AND1_U1 ( .A0_t (LED_128_Instance_n31), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_5_U1_X), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_5_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_5_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_5_U1_Y), .B0_t (IN_key[69]), .Z0_t (LED_128_Instance_current_roundkey[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_6_U1_XOR1_U1 ( .A0_t (IN_key[70]), .B0_t (IN_key[6]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_6_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_6_U1_AND1_U1 ( .A0_t (LED_128_Instance_n31), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_6_U1_X), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_6_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_6_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_6_U1_Y), .B0_t (IN_key[70]), .Z0_t (LED_128_Instance_current_roundkey[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_7_U1_XOR1_U1 ( .A0_t (IN_key[71]), .B0_t (IN_key[7]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_7_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_7_U1_AND1_U1 ( .A0_t (LED_128_Instance_n31), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_7_U1_X), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_7_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_7_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_7_U1_Y), .B0_t (IN_key[71]), .Z0_t (LED_128_Instance_current_roundkey[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_8_U1_XOR1_U1 ( .A0_t (IN_key[72]), .B0_t (IN_key[8]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_8_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_8_U1_AND1_U1 ( .A0_t (LED_128_Instance_n31), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_8_U1_X), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_8_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_8_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_8_U1_Y), .B0_t (IN_key[72]), .Z0_t (LED_128_Instance_current_roundkey[8]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_9_U1_XOR1_U1 ( .A0_t (IN_key[73]), .B0_t (IN_key[9]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_9_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_9_U1_AND1_U1 ( .A0_t (LED_128_Instance_n31), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_9_U1_X), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_9_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_9_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_9_U1_Y), .B0_t (IN_key[73]), .Z0_t (LED_128_Instance_current_roundkey[9]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_10_U1_XOR1_U1 ( .A0_t (IN_key[74]), .B0_t (IN_key[10]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_10_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_10_U1_AND1_U1 ( .A0_t (LED_128_Instance_n31), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_10_U1_X), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_10_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_10_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_10_U1_Y), .B0_t (IN_key[74]), .Z0_t (LED_128_Instance_current_roundkey[10]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_11_U1_XOR1_U1 ( .A0_t (IN_key[75]), .B0_t (IN_key[11]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_11_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_11_U1_AND1_U1 ( .A0_t (LED_128_Instance_n31), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_11_U1_X), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_11_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_11_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_11_U1_Y), .B0_t (IN_key[75]), .Z0_t (LED_128_Instance_current_roundkey[11]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_12_U1_XOR1_U1 ( .A0_t (IN_key[76]), .B0_t (IN_key[12]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_12_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_12_U1_AND1_U1 ( .A0_t (LED_128_Instance_n31), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_12_U1_X), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_12_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_12_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_12_U1_Y), .B0_t (IN_key[76]), .Z0_t (LED_128_Instance_current_roundkey[12]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_13_U1_XOR1_U1 ( .A0_t (IN_key[77]), .B0_t (IN_key[13]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_13_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_13_U1_AND1_U1 ( .A0_t (LED_128_Instance_n31), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_13_U1_X), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_13_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_13_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_13_U1_Y), .B0_t (IN_key[77]), .Z0_t (LED_128_Instance_current_roundkey[13]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_14_U1_XOR1_U1 ( .A0_t (IN_key[78]), .B0_t (IN_key[14]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_14_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_14_U1_AND1_U1 ( .A0_t (LED_128_Instance_n31), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_14_U1_X), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_14_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_14_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_14_U1_Y), .B0_t (IN_key[78]), .Z0_t (LED_128_Instance_current_roundkey[14]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_15_U1_XOR1_U1 ( .A0_t (IN_key[79]), .B0_t (IN_key[15]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_15_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_15_U1_AND1_U1 ( .A0_t (LED_128_Instance_n31), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_15_U1_X), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_15_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_15_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_15_U1_Y), .B0_t (IN_key[79]), .Z0_t (LED_128_Instance_current_roundkey[15]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_16_U1_XOR1_U1 ( .A0_t (IN_key[80]), .B0_t (IN_key[16]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_16_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_16_U1_AND1_U1 ( .A0_t (LED_128_Instance_n31), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_16_U1_X), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_16_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_16_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_16_U1_Y), .B0_t (IN_key[80]), .Z0_t (LED_128_Instance_current_roundkey[16]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_17_U1_XOR1_U1 ( .A0_t (IN_key[81]), .B0_t (IN_key[17]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_17_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_17_U1_AND1_U1 ( .A0_t (LED_128_Instance_n31), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_17_U1_X), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_17_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_17_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_17_U1_Y), .B0_t (IN_key[81]), .Z0_t (LED_128_Instance_current_roundkey[17]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_18_U1_XOR1_U1 ( .A0_t (IN_key[82]), .B0_t (IN_key[18]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_18_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_18_U1_AND1_U1 ( .A0_t (LED_128_Instance_n31), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_18_U1_X), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_18_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_18_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_18_U1_Y), .B0_t (IN_key[82]), .Z0_t (LED_128_Instance_current_roundkey[18]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_19_U1_XOR1_U1 ( .A0_t (IN_key[83]), .B0_t (IN_key[19]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_19_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_19_U1_AND1_U1 ( .A0_t (LED_128_Instance_n31), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_19_U1_X), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_19_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_19_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_19_U1_Y), .B0_t (IN_key[83]), .Z0_t (LED_128_Instance_current_roundkey[19]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_20_U1_XOR1_U1 ( .A0_t (IN_key[84]), .B0_t (IN_key[20]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_20_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_20_U1_AND1_U1 ( .A0_t (LED_128_Instance_n31), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_20_U1_X), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_20_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_20_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_20_U1_Y), .B0_t (IN_key[84]), .Z0_t (LED_128_Instance_current_roundkey[20]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_21_U1_XOR1_U1 ( .A0_t (IN_key[85]), .B0_t (IN_key[21]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_21_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_21_U1_AND1_U1 ( .A0_t (LED_128_Instance_n31), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_21_U1_X), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_21_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_21_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_21_U1_Y), .B0_t (IN_key[85]), .Z0_t (LED_128_Instance_current_roundkey[21]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_22_U1_XOR1_U1 ( .A0_t (IN_key[86]), .B0_t (IN_key[22]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_22_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_22_U1_AND1_U1 ( .A0_t (LED_128_Instance_n31), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_22_U1_X), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_22_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_22_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_22_U1_Y), .B0_t (IN_key[86]), .Z0_t (LED_128_Instance_current_roundkey[22]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_23_U1_XOR1_U1 ( .A0_t (IN_key[87]), .B0_t (IN_key[23]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_23_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_23_U1_AND1_U1 ( .A0_t (LED_128_Instance_n31), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_23_U1_X), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_23_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_23_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_23_U1_Y), .B0_t (IN_key[87]), .Z0_t (LED_128_Instance_current_roundkey[23]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_24_U1_XOR1_U1 ( .A0_t (IN_key[88]), .B0_t (IN_key[24]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_24_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_24_U1_AND1_U1 ( .A0_t (LED_128_Instance_n31), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_24_U1_X), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_24_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_24_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_24_U1_Y), .B0_t (IN_key[88]), .Z0_t (LED_128_Instance_current_roundkey[24]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_25_U1_XOR1_U1 ( .A0_t (IN_key[89]), .B0_t (IN_key[25]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_25_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_25_U1_AND1_U1 ( .A0_t (LED_128_Instance_n31), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_25_U1_X), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_25_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_25_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_25_U1_Y), .B0_t (IN_key[89]), .Z0_t (LED_128_Instance_current_roundkey[25]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_26_U1_XOR1_U1 ( .A0_t (IN_key[90]), .B0_t (IN_key[26]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_26_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_26_U1_AND1_U1 ( .A0_t (LED_128_Instance_n31), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_26_U1_X), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_26_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_26_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_26_U1_Y), .B0_t (IN_key[90]), .Z0_t (LED_128_Instance_current_roundkey[26]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_27_U1_XOR1_U1 ( .A0_t (IN_key[91]), .B0_t (IN_key[27]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_27_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_27_U1_AND1_U1 ( .A0_t (LED_128_Instance_n31), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_27_U1_X), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_27_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_27_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_27_U1_Y), .B0_t (IN_key[91]), .Z0_t (LED_128_Instance_current_roundkey[27]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_28_U1_XOR1_U1 ( .A0_t (IN_key[92]), .B0_t (IN_key[28]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_28_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_28_U1_AND1_U1 ( .A0_t (LED_128_Instance_n31), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_28_U1_X), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_28_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_28_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_28_U1_Y), .B0_t (IN_key[92]), .Z0_t (LED_128_Instance_current_roundkey[28]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_29_U1_XOR1_U1 ( .A0_t (IN_key[93]), .B0_t (IN_key[29]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_29_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_29_U1_AND1_U1 ( .A0_t (LED_128_Instance_n31), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_29_U1_X), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_29_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_29_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_29_U1_Y), .B0_t (IN_key[93]), .Z0_t (LED_128_Instance_current_roundkey[29]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_30_U1_XOR1_U1 ( .A0_t (IN_key[94]), .B0_t (IN_key[30]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_30_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_30_U1_AND1_U1 ( .A0_t (LED_128_Instance_n31), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_30_U1_X), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_30_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_30_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_30_U1_Y), .B0_t (IN_key[94]), .Z0_t (LED_128_Instance_current_roundkey[30]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_31_U1_XOR1_U1 ( .A0_t (IN_key[95]), .B0_t (IN_key[31]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_31_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_31_U1_AND1_U1 ( .A0_t (LED_128_Instance_n31), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_31_U1_X), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_31_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_31_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_31_U1_Y), .B0_t (IN_key[95]), .Z0_t (LED_128_Instance_current_roundkey[31]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_32_U1_XOR1_U1 ( .A0_t (IN_key[96]), .B0_t (IN_key[32]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_32_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_32_U1_AND1_U1 ( .A0_t (LED_128_Instance_n31), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_32_U1_X), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_32_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_32_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_32_U1_Y), .B0_t (IN_key[96]), .Z0_t (LED_128_Instance_current_roundkey[32]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_33_U1_XOR1_U1 ( .A0_t (IN_key[97]), .B0_t (IN_key[33]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_33_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_33_U1_AND1_U1 ( .A0_t (LED_128_Instance_n31), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_33_U1_X), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_33_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_33_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_33_U1_Y), .B0_t (IN_key[97]), .Z0_t (LED_128_Instance_current_roundkey[33]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_34_U1_XOR1_U1 ( .A0_t (IN_key[98]), .B0_t (IN_key[34]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_34_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_34_U1_AND1_U1 ( .A0_t (LED_128_Instance_n31), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_34_U1_X), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_34_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_34_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_34_U1_Y), .B0_t (IN_key[98]), .Z0_t (LED_128_Instance_current_roundkey[34]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_35_U1_XOR1_U1 ( .A0_t (IN_key[99]), .B0_t (IN_key[35]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_35_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_35_U1_AND1_U1 ( .A0_t (LED_128_Instance_n31), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_35_U1_X), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_35_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_35_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_35_U1_Y), .B0_t (IN_key[99]), .Z0_t (LED_128_Instance_current_roundkey[35]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_36_U1_XOR1_U1 ( .A0_t (IN_key[100]), .B0_t (IN_key[36]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_36_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_36_U1_AND1_U1 ( .A0_t (LED_128_Instance_n31), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_36_U1_X), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_36_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_36_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_36_U1_Y), .B0_t (IN_key[100]), .Z0_t (LED_128_Instance_current_roundkey[36]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_37_U1_XOR1_U1 ( .A0_t (IN_key[101]), .B0_t (IN_key[37]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_37_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_37_U1_AND1_U1 ( .A0_t (LED_128_Instance_n31), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_37_U1_X), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_37_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_37_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_37_U1_Y), .B0_t (IN_key[101]), .Z0_t (LED_128_Instance_current_roundkey[37]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_38_U1_XOR1_U1 ( .A0_t (IN_key[102]), .B0_t (IN_key[38]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_38_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_38_U1_AND1_U1 ( .A0_t (LED_128_Instance_n31), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_38_U1_X), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_38_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_38_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_38_U1_Y), .B0_t (IN_key[102]), .Z0_t (LED_128_Instance_current_roundkey[38]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_39_U1_XOR1_U1 ( .A0_t (IN_key[103]), .B0_t (IN_key[39]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_39_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_39_U1_AND1_U1 ( .A0_t (LED_128_Instance_n31), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_39_U1_X), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_39_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_39_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_39_U1_Y), .B0_t (IN_key[103]), .Z0_t (LED_128_Instance_current_roundkey[39]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_40_U1_XOR1_U1 ( .A0_t (IN_key[104]), .B0_t (IN_key[40]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_40_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_40_U1_AND1_U1 ( .A0_t (LED_128_Instance_n31), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_40_U1_X), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_40_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_40_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_40_U1_Y), .B0_t (IN_key[104]), .Z0_t (LED_128_Instance_current_roundkey[40]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_41_U1_XOR1_U1 ( .A0_t (IN_key[105]), .B0_t (IN_key[41]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_41_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_41_U1_AND1_U1 ( .A0_t (LED_128_Instance_n31), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_41_U1_X), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_41_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_41_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_41_U1_Y), .B0_t (IN_key[105]), .Z0_t (LED_128_Instance_current_roundkey[41]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_42_U1_XOR1_U1 ( .A0_t (IN_key[106]), .B0_t (IN_key[42]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_42_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_42_U1_AND1_U1 ( .A0_t (LED_128_Instance_n31), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_42_U1_X), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_42_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_42_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_42_U1_Y), .B0_t (IN_key[106]), .Z0_t (LED_128_Instance_current_roundkey[42]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_43_U1_XOR1_U1 ( .A0_t (IN_key[107]), .B0_t (IN_key[43]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_43_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_43_U1_AND1_U1 ( .A0_t (LED_128_Instance_n31), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_43_U1_X), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_43_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_43_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_43_U1_Y), .B0_t (IN_key[107]), .Z0_t (LED_128_Instance_current_roundkey[43]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_44_U1_XOR1_U1 ( .A0_t (IN_key[108]), .B0_t (IN_key[44]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_44_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_44_U1_AND1_U1 ( .A0_t (LED_128_Instance_n31), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_44_U1_X), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_44_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_44_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_44_U1_Y), .B0_t (IN_key[108]), .Z0_t (LED_128_Instance_current_roundkey[44]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_45_U1_XOR1_U1 ( .A0_t (IN_key[109]), .B0_t (IN_key[45]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_45_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_45_U1_AND1_U1 ( .A0_t (LED_128_Instance_n31), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_45_U1_X), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_45_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_45_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_45_U1_Y), .B0_t (IN_key[109]), .Z0_t (LED_128_Instance_current_roundkey[45]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_46_U1_XOR1_U1 ( .A0_t (IN_key[110]), .B0_t (IN_key[46]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_46_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_46_U1_AND1_U1 ( .A0_t (LED_128_Instance_n31), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_46_U1_X), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_46_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_46_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_46_U1_Y), .B0_t (IN_key[110]), .Z0_t (LED_128_Instance_current_roundkey[46]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_47_U1_XOR1_U1 ( .A0_t (IN_key[111]), .B0_t (IN_key[47]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_47_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_47_U1_AND1_U1 ( .A0_t (LED_128_Instance_n31), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_47_U1_X), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_47_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_47_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_47_U1_Y), .B0_t (IN_key[111]), .Z0_t (LED_128_Instance_current_roundkey[47]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_48_U1_XOR1_U1 ( .A0_t (IN_key[112]), .B0_t (IN_key[48]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_48_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_48_U1_AND1_U1 ( .A0_t (LED_128_Instance_n31), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_48_U1_X), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_48_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_48_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_48_U1_Y), .B0_t (IN_key[112]), .Z0_t (LED_128_Instance_current_roundkey[48]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_49_U1_XOR1_U1 ( .A0_t (IN_key[113]), .B0_t (IN_key[49]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_49_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_49_U1_AND1_U1 ( .A0_t (LED_128_Instance_n31), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_49_U1_X), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_49_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_49_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_49_U1_Y), .B0_t (IN_key[113]), .Z0_t (LED_128_Instance_current_roundkey[49]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_50_U1_XOR1_U1 ( .A0_t (IN_key[114]), .B0_t (IN_key[50]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_50_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_50_U1_AND1_U1 ( .A0_t (LED_128_Instance_n31), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_50_U1_X), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_50_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_50_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_50_U1_Y), .B0_t (IN_key[114]), .Z0_t (LED_128_Instance_current_roundkey[50]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_51_U1_XOR1_U1 ( .A0_t (IN_key[115]), .B0_t (IN_key[51]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_51_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_51_U1_AND1_U1 ( .A0_t (LED_128_Instance_n31), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_51_U1_X), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_51_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_51_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_51_U1_Y), .B0_t (IN_key[115]), .Z0_t (LED_128_Instance_current_roundkey[51]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_52_U1_XOR1_U1 ( .A0_t (IN_key[116]), .B0_t (IN_key[52]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_52_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_52_U1_AND1_U1 ( .A0_t (LED_128_Instance_n31), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_52_U1_X), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_52_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_52_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_52_U1_Y), .B0_t (IN_key[116]), .Z0_t (LED_128_Instance_current_roundkey[52]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_53_U1_XOR1_U1 ( .A0_t (IN_key[117]), .B0_t (IN_key[53]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_53_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_53_U1_AND1_U1 ( .A0_t (LED_128_Instance_n31), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_53_U1_X), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_53_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_53_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_53_U1_Y), .B0_t (IN_key[117]), .Z0_t (LED_128_Instance_current_roundkey[53]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_54_U1_XOR1_U1 ( .A0_t (IN_key[118]), .B0_t (IN_key[54]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_54_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_54_U1_AND1_U1 ( .A0_t (LED_128_Instance_n31), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_54_U1_X), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_54_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_54_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_54_U1_Y), .B0_t (IN_key[118]), .Z0_t (LED_128_Instance_current_roundkey[54]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_55_U1_XOR1_U1 ( .A0_t (IN_key[119]), .B0_t (IN_key[55]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_55_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_55_U1_AND1_U1 ( .A0_t (LED_128_Instance_n31), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_55_U1_X), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_55_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_55_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_55_U1_Y), .B0_t (IN_key[119]), .Z0_t (LED_128_Instance_current_roundkey[55]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_56_U1_XOR1_U1 ( .A0_t (IN_key[120]), .B0_t (IN_key[56]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_56_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_56_U1_AND1_U1 ( .A0_t (LED_128_Instance_n31), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_56_U1_X), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_56_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_56_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_56_U1_Y), .B0_t (IN_key[120]), .Z0_t (LED_128_Instance_current_roundkey[56]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_57_U1_XOR1_U1 ( .A0_t (IN_key[121]), .B0_t (IN_key[57]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_57_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_57_U1_AND1_U1 ( .A0_t (LED_128_Instance_n31), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_57_U1_X), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_57_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_57_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_57_U1_Y), .B0_t (IN_key[121]), .Z0_t (LED_128_Instance_current_roundkey[57]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_58_U1_XOR1_U1 ( .A0_t (IN_key[122]), .B0_t (IN_key[58]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_58_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_58_U1_AND1_U1 ( .A0_t (LED_128_Instance_n31), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_58_U1_X), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_58_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_58_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_58_U1_Y), .B0_t (IN_key[122]), .Z0_t (LED_128_Instance_current_roundkey[58]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_59_U1_XOR1_U1 ( .A0_t (IN_key[123]), .B0_t (IN_key[59]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_59_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_59_U1_AND1_U1 ( .A0_t (LED_128_Instance_n31), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_59_U1_X), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_59_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_59_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_59_U1_Y), .B0_t (IN_key[123]), .Z0_t (LED_128_Instance_current_roundkey[59]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_60_U1_XOR1_U1 ( .A0_t (IN_key[124]), .B0_t (IN_key[60]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_60_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_60_U1_AND1_U1 ( .A0_t (LED_128_Instance_n31), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_60_U1_X), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_60_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_60_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_60_U1_Y), .B0_t (IN_key[124]), .Z0_t (LED_128_Instance_current_roundkey[60]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_61_U1_XOR1_U1 ( .A0_t (IN_key[125]), .B0_t (IN_key[61]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_61_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_61_U1_AND1_U1 ( .A0_t (LED_128_Instance_n31), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_61_U1_X), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_61_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_61_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_61_U1_Y), .B0_t (IN_key[125]), .Z0_t (LED_128_Instance_current_roundkey[61]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_62_U1_XOR1_U1 ( .A0_t (IN_key[126]), .B0_t (IN_key[62]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_62_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_62_U1_AND1_U1 ( .A0_t (LED_128_Instance_n31), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_62_U1_X), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_62_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_62_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_62_U1_Y), .B0_t (IN_key[126]), .Z0_t (LED_128_Instance_current_roundkey[62]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_63_U1_XOR1_U1 ( .A0_t (IN_key[127]), .B0_t (IN_key[63]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_63_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_63_U1_AND1_U1 ( .A0_t (LED_128_Instance_n31), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_63_U1_X), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_63_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_63_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_63_U1_Y), .B0_t (IN_key[127]), .Z0_t (LED_128_Instance_current_roundkey[63]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U64 ( .A0_t (OUT_ciphertext[28]), .B0_t (LED_128_Instance_current_roundkey[28]), .Z0_t (LED_128_Instance_addroundkey_tmp[28]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U63 ( .A0_t (OUT_ciphertext[24]), .B0_t (LED_128_Instance_current_roundkey[24]), .Z0_t (LED_128_Instance_addroundkey_tmp[24]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U62 ( .A0_t (OUT_ciphertext[12]), .B0_t (LED_128_Instance_current_roundkey[12]), .Z0_t (LED_128_Instance_addroundkey_tmp[12]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U61 ( .A0_t (OUT_ciphertext[8]), .B0_t (LED_128_Instance_current_roundkey[8]), .Z0_t (LED_128_Instance_addroundkey_tmp[8]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U60 ( .A0_t (OUT_ciphertext[0]), .B0_t (LED_128_Instance_current_roundkey[0]), .Z0_t (LED_128_Instance_addroundkey_tmp[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U59 ( .A0_t (OUT_ciphertext[48]), .B0_t (LED_128_Instance_current_roundkey[48]), .Z0_t (LED_128_Instance_addroundkey_tmp[48]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U58 ( .A0_t (OUT_ciphertext[16]), .B0_t (LED_128_Instance_current_roundkey[16]), .Z0_t (LED_128_Instance_addroundkey_tmp[16]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U57 ( .A0_t (OUT_ciphertext[56]), .B0_t (LED_128_Instance_current_roundkey[56]), .Z0_t (LED_128_Instance_addroundkey_tmp[56]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U56 ( .A0_t (OUT_ciphertext[60]), .B0_t (LED_128_Instance_current_roundkey[60]), .Z0_t (LED_128_Instance_addroundkey_tmp[60]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U55 ( .A0_t (OUT_ciphertext[31]), .B0_t (LED_128_Instance_current_roundkey[31]), .Z0_t (LED_128_Instance_addroundkey_tmp[31]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U54 ( .A0_t (OUT_ciphertext[27]), .B0_t (LED_128_Instance_current_roundkey[27]), .Z0_t (LED_128_Instance_addroundkey_tmp[27]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U53 ( .A0_t (OUT_ciphertext[23]), .B0_t (LED_128_Instance_current_roundkey[23]), .Z0_t (LED_128_Instance_addroundkey_tmp[23]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U52 ( .A0_t (OUT_ciphertext[32]), .B0_t (LED_128_Instance_current_roundkey[32]), .Z0_t (LED_128_Instance_addroundkey_tmp[32]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U51 ( .A0_t (OUT_ciphertext[44]), .B0_t (LED_128_Instance_current_roundkey[44]), .Z0_t (LED_128_Instance_addroundkey_tmp[44]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U50 ( .A0_t (OUT_ciphertext[40]), .B0_t (LED_128_Instance_current_roundkey[40]), .Z0_t (LED_128_Instance_addroundkey_tmp[40]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U49 ( .A0_t (OUT_ciphertext[33]), .B0_t (LED_128_Instance_current_roundkey[33]), .Z0_t (LED_128_Instance_addroundkey_tmp[33]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U48 ( .A0_t (OUT_ciphertext[49]), .B0_t (LED_128_Instance_current_roundkey[49]), .Z0_t (LED_128_Instance_addroundkey_tmp[49]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U47 ( .A0_t (OUT_ciphertext[19]), .B0_t (LED_128_Instance_current_roundkey[19]), .Z0_t (LED_128_Instance_addroundkey_tmp[19]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U46 ( .A0_t (OUT_ciphertext[3]), .B0_t (LED_128_Instance_current_roundkey[3]), .Z0_t (LED_128_Instance_addroundkey_tmp[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U45 ( .A0_t (OUT_ciphertext[54]), .B0_t (LED_128_Instance_current_roundkey[54]), .Z0_t (LED_128_Instance_addroundkey_tmp[54]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U44 ( .A0_t (OUT_ciphertext[38]), .B0_t (LED_128_Instance_current_roundkey[38]), .Z0_t (LED_128_Instance_addroundkey_tmp[38]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U43 ( .A0_t (OUT_ciphertext[36]), .B0_t (LED_128_Instance_current_roundkey[36]), .Z0_t (LED_128_Instance_addroundkey_tmp[36]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U42 ( .A0_t (OUT_ciphertext[52]), .B0_t (LED_128_Instance_current_roundkey[52]), .Z0_t (LED_128_Instance_addroundkey_tmp[52]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U41 ( .A0_t (OUT_ciphertext[37]), .B0_t (LED_128_Instance_current_roundkey[37]), .Z0_t (LED_128_Instance_addroundkey_tmp[37]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U40 ( .A0_t (OUT_ciphertext[53]), .B0_t (LED_128_Instance_current_roundkey[53]), .Z0_t (LED_128_Instance_addroundkey_tmp[53]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U39 ( .A0_t (OUT_ciphertext[4]), .B0_t (LED_128_Instance_current_roundkey[4]), .Z0_t (LED_128_Instance_addroundkey_tmp[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U38 ( .A0_t (OUT_ciphertext[6]), .B0_t (LED_128_Instance_current_roundkey[6]), .Z0_t (LED_128_Instance_addroundkey_tmp[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U37 ( .A0_t (OUT_ciphertext[20]), .B0_t (LED_128_Instance_current_roundkey[20]), .Z0_t (LED_128_Instance_addroundkey_tmp[20]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U36 ( .A0_t (OUT_ciphertext[22]), .B0_t (LED_128_Instance_current_roundkey[22]), .Z0_t (LED_128_Instance_addroundkey_tmp[22]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U35 ( .A0_t (OUT_ciphertext[5]), .B0_t (LED_128_Instance_current_roundkey[5]), .Z0_t (LED_128_Instance_addroundkey_tmp[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U34 ( .A0_t (OUT_ciphertext[21]), .B0_t (LED_128_Instance_current_roundkey[21]), .Z0_t (LED_128_Instance_addroundkey_tmp[21]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U33 ( .A0_t (OUT_ciphertext[58]), .B0_t (LED_128_Instance_current_roundkey[58]), .Z0_t (LED_128_Instance_addroundkey_tmp[58]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U32 ( .A0_t (OUT_ciphertext[50]), .B0_t (LED_128_Instance_current_roundkey[50]), .Z0_t (LED_128_Instance_addroundkey_tmp[50]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U31 ( .A0_t (OUT_ciphertext[62]), .B0_t (LED_128_Instance_current_roundkey[62]), .Z0_t (LED_128_Instance_addroundkey_tmp[62]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U30 ( .A0_t (OUT_ciphertext[34]), .B0_t (LED_128_Instance_current_roundkey[34]), .Z0_t (LED_128_Instance_addroundkey_tmp[34]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U29 ( .A0_t (OUT_ciphertext[46]), .B0_t (LED_128_Instance_current_roundkey[46]), .Z0_t (LED_128_Instance_addroundkey_tmp[46]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U28 ( .A0_t (OUT_ciphertext[42]), .B0_t (LED_128_Instance_current_roundkey[42]), .Z0_t (LED_128_Instance_addroundkey_tmp[42]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U27 ( .A0_t (OUT_ciphertext[14]), .B0_t (LED_128_Instance_current_roundkey[14]), .Z0_t (LED_128_Instance_addroundkey_tmp[14]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U26 ( .A0_t (OUT_ciphertext[18]), .B0_t (LED_128_Instance_current_roundkey[18]), .Z0_t (LED_128_Instance_addroundkey_tmp[18]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U25 ( .A0_t (OUT_ciphertext[10]), .B0_t (LED_128_Instance_current_roundkey[10]), .Z0_t (LED_128_Instance_addroundkey_tmp[10]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U24 ( .A0_t (OUT_ciphertext[30]), .B0_t (LED_128_Instance_current_roundkey[30]), .Z0_t (LED_128_Instance_addroundkey_tmp[30]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U23 ( .A0_t (OUT_ciphertext[26]), .B0_t (LED_128_Instance_current_roundkey[26]), .Z0_t (LED_128_Instance_addroundkey_tmp[26]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U22 ( .A0_t (OUT_ciphertext[2]), .B0_t (LED_128_Instance_current_roundkey[2]), .Z0_t (LED_128_Instance_addroundkey_tmp[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U21 ( .A0_t (OUT_ciphertext[45]), .B0_t (LED_128_Instance_current_roundkey[45]), .Z0_t (LED_128_Instance_addroundkey_tmp[45]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U20 ( .A0_t (OUT_ciphertext[41]), .B0_t (LED_128_Instance_current_roundkey[41]), .Z0_t (LED_128_Instance_addroundkey_tmp[41]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U19 ( .A0_t (OUT_ciphertext[57]), .B0_t (LED_128_Instance_current_roundkey[57]), .Z0_t (LED_128_Instance_addroundkey_tmp[57]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U18 ( .A0_t (OUT_ciphertext[61]), .B0_t (LED_128_Instance_current_roundkey[61]), .Z0_t (LED_128_Instance_addroundkey_tmp[61]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U17 ( .A0_t (OUT_ciphertext[13]), .B0_t (LED_128_Instance_current_roundkey[13]), .Z0_t (LED_128_Instance_addroundkey_tmp[13]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U16 ( .A0_t (OUT_ciphertext[17]), .B0_t (LED_128_Instance_current_roundkey[17]), .Z0_t (LED_128_Instance_addroundkey_tmp[17]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U15 ( .A0_t (OUT_ciphertext[9]), .B0_t (LED_128_Instance_current_roundkey[9]), .Z0_t (LED_128_Instance_addroundkey_tmp[9]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U14 ( .A0_t (OUT_ciphertext[29]), .B0_t (LED_128_Instance_current_roundkey[29]), .Z0_t (LED_128_Instance_addroundkey_tmp[29]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U13 ( .A0_t (OUT_ciphertext[25]), .B0_t (LED_128_Instance_current_roundkey[25]), .Z0_t (LED_128_Instance_addroundkey_tmp[25]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U12 ( .A0_t (OUT_ciphertext[1]), .B0_t (LED_128_Instance_current_roundkey[1]), .Z0_t (LED_128_Instance_addroundkey_tmp[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U11 ( .A0_t (OUT_ciphertext[39]), .B0_t (LED_128_Instance_current_roundkey[39]), .Z0_t (LED_128_Instance_addroundkey_tmp[39]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U10 ( .A0_t (OUT_ciphertext[35]), .B0_t (LED_128_Instance_current_roundkey[35]), .Z0_t (LED_128_Instance_addroundkey_tmp[35]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U9 ( .A0_t (OUT_ciphertext[47]), .B0_t (LED_128_Instance_current_roundkey[47]), .Z0_t (LED_128_Instance_addroundkey_tmp[47]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U8 ( .A0_t (OUT_ciphertext[43]), .B0_t (LED_128_Instance_current_roundkey[43]), .Z0_t (LED_128_Instance_addroundkey_tmp[43]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U7 ( .A0_t (OUT_ciphertext[59]), .B0_t (LED_128_Instance_current_roundkey[59]), .Z0_t (LED_128_Instance_addroundkey_tmp[59]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U6 ( .A0_t (OUT_ciphertext[55]), .B0_t (LED_128_Instance_current_roundkey[55]), .Z0_t (LED_128_Instance_addroundkey_tmp[55]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U5 ( .A0_t (OUT_ciphertext[51]), .B0_t (LED_128_Instance_current_roundkey[51]), .Z0_t (LED_128_Instance_addroundkey_tmp[51]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U4 ( .A0_t (OUT_ciphertext[63]), .B0_t (LED_128_Instance_current_roundkey[63]), .Z0_t (LED_128_Instance_addroundkey_tmp[63]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U3 ( .A0_t (OUT_ciphertext[15]), .B0_t (LED_128_Instance_current_roundkey[15]), .Z0_t (LED_128_Instance_addroundkey_tmp[15]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U2 ( .A0_t (OUT_ciphertext[11]), .B0_t (LED_128_Instance_current_roundkey[11]), .Z0_t (LED_128_Instance_addroundkey_tmp[11]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U1 ( .A0_t (OUT_ciphertext[7]), .B0_t (LED_128_Instance_current_roundkey[7]), .Z0_t (LED_128_Instance_addroundkey_tmp[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_0_U1_XOR1_U1 ( .A0_t (OUT_ciphertext[0]), .B0_t (LED_128_Instance_addroundkey_tmp[0]), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_0_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_0_U1_AND1_U1 ( .A0_t (LED_128_Instance_n23), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_0_U1_X), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_0_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_0_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_0_U1_Y), .B0_t (OUT_ciphertext[0]), .Z0_t (LED_128_Instance_addconst_out[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_1_U1_XOR1_U1 ( .A0_t (OUT_ciphertext[1]), .B0_t (LED_128_Instance_addroundkey_tmp[1]), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_1_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_1_U1_AND1_U1 ( .A0_t (LED_128_Instance_n23), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_1_U1_X), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_1_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_1_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_1_U1_Y), .B0_t (OUT_ciphertext[1]), .Z0_t (LED_128_Instance_addconst_out[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_2_U1_XOR1_U1 ( .A0_t (OUT_ciphertext[2]), .B0_t (LED_128_Instance_addroundkey_tmp[2]), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_2_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_2_U1_AND1_U1 ( .A0_t (LED_128_Instance_n23), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_2_U1_X), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_2_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_2_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_2_U1_Y), .B0_t (OUT_ciphertext[2]), .Z0_t (LED_128_Instance_addconst_out[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_3_U1_XOR1_U1 ( .A0_t (OUT_ciphertext[3]), .B0_t (LED_128_Instance_addroundkey_tmp[3]), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_3_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_3_U1_AND1_U1 ( .A0_t (LED_128_Instance_n23), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_3_U1_X), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_3_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_3_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_3_U1_Y), .B0_t (OUT_ciphertext[3]), .Z0_t (LED_128_Instance_addroundkey_out[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_4_U1_XOR1_U1 ( .A0_t (OUT_ciphertext[4]), .B0_t (LED_128_Instance_addroundkey_tmp[4]), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_4_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_4_U1_AND1_U1 ( .A0_t (LED_128_Instance_n23), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_4_U1_X), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_4_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_4_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_4_U1_Y), .B0_t (OUT_ciphertext[4]), .Z0_t (LED_128_Instance_addroundkey_out[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_5_U1_XOR1_U1 ( .A0_t (OUT_ciphertext[5]), .B0_t (LED_128_Instance_addroundkey_tmp[5]), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_5_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_5_U1_AND1_U1 ( .A0_t (LED_128_Instance_n23), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_5_U1_X), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_5_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_5_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_5_U1_Y), .B0_t (OUT_ciphertext[5]), .Z0_t (LED_128_Instance_addroundkey_out[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_6_U1_XOR1_U1 ( .A0_t (OUT_ciphertext[6]), .B0_t (LED_128_Instance_addroundkey_tmp[6]), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_6_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_6_U1_AND1_U1 ( .A0_t (LED_128_Instance_n23), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_6_U1_X), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_6_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_6_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_6_U1_Y), .B0_t (OUT_ciphertext[6]), .Z0_t (LED_128_Instance_addroundkey_out[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_7_U1_XOR1_U1 ( .A0_t (OUT_ciphertext[7]), .B0_t (LED_128_Instance_addroundkey_tmp[7]), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_7_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_7_U1_AND1_U1 ( .A0_t (LED_128_Instance_n23), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_7_U1_X), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_7_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_7_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_7_U1_Y), .B0_t (OUT_ciphertext[7]), .Z0_t (LED_128_Instance_addconst_out[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_8_U1_XOR1_U1 ( .A0_t (OUT_ciphertext[8]), .B0_t (LED_128_Instance_addroundkey_tmp[8]), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_8_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_8_U1_AND1_U1 ( .A0_t (LED_128_Instance_n23), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_8_U1_X), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_8_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_8_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_8_U1_Y), .B0_t (OUT_ciphertext[8]), .Z0_t (LED_128_Instance_addconst_out[8]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_9_U1_XOR1_U1 ( .A0_t (OUT_ciphertext[9]), .B0_t (LED_128_Instance_addroundkey_tmp[9]), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_9_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_9_U1_AND1_U1 ( .A0_t (LED_128_Instance_n23), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_9_U1_X), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_9_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_9_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_9_U1_Y), .B0_t (OUT_ciphertext[9]), .Z0_t (LED_128_Instance_addconst_out[9]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_10_U1_XOR1_U1 ( .A0_t (OUT_ciphertext[10]), .B0_t (LED_128_Instance_addroundkey_tmp[10]), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_10_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_10_U1_AND1_U1 ( .A0_t (LED_128_Instance_n23), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_10_U1_X), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_10_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_10_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_10_U1_Y), .B0_t (OUT_ciphertext[10]), .Z0_t (LED_128_Instance_addconst_out[10]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_11_U1_XOR1_U1 ( .A0_t (OUT_ciphertext[11]), .B0_t (LED_128_Instance_addroundkey_tmp[11]), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_11_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_11_U1_AND1_U1 ( .A0_t (LED_128_Instance_n23), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_11_U1_X), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_11_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_11_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_11_U1_Y), .B0_t (OUT_ciphertext[11]), .Z0_t (LED_128_Instance_addconst_out[11]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_12_U1_XOR1_U1 ( .A0_t (OUT_ciphertext[12]), .B0_t (LED_128_Instance_addroundkey_tmp[12]), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_12_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_12_U1_AND1_U1 ( .A0_t (LED_128_Instance_n23), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_12_U1_X), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_12_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_12_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_12_U1_Y), .B0_t (OUT_ciphertext[12]), .Z0_t (LED_128_Instance_addconst_out[12]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_13_U1_XOR1_U1 ( .A0_t (OUT_ciphertext[13]), .B0_t (LED_128_Instance_addroundkey_tmp[13]), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_13_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_13_U1_AND1_U1 ( .A0_t (LED_128_Instance_n23), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_13_U1_X), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_13_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_13_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_13_U1_Y), .B0_t (OUT_ciphertext[13]), .Z0_t (LED_128_Instance_addconst_out[13]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_14_U1_XOR1_U1 ( .A0_t (OUT_ciphertext[14]), .B0_t (LED_128_Instance_addroundkey_tmp[14]), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_14_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_14_U1_AND1_U1 ( .A0_t (LED_128_Instance_n23), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_14_U1_X), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_14_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_14_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_14_U1_Y), .B0_t (OUT_ciphertext[14]), .Z0_t (LED_128_Instance_addconst_out[14]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_15_U1_XOR1_U1 ( .A0_t (OUT_ciphertext[15]), .B0_t (LED_128_Instance_addroundkey_tmp[15]), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_15_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_15_U1_AND1_U1 ( .A0_t (LED_128_Instance_n23), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_15_U1_X), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_15_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_15_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_15_U1_Y), .B0_t (OUT_ciphertext[15]), .Z0_t (LED_128_Instance_addconst_out[15]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_16_U1_XOR1_U1 ( .A0_t (OUT_ciphertext[16]), .B0_t (LED_128_Instance_addroundkey_tmp[16]), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_16_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_16_U1_AND1_U1 ( .A0_t (LED_128_Instance_n23), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_16_U1_X), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_16_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_16_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_16_U1_Y), .B0_t (OUT_ciphertext[16]), .Z0_t (LED_128_Instance_addroundkey_out[16]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_17_U1_XOR1_U1 ( .A0_t (OUT_ciphertext[17]), .B0_t (LED_128_Instance_addroundkey_tmp[17]), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_17_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_17_U1_AND1_U1 ( .A0_t (LED_128_Instance_n23), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_17_U1_X), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_17_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_17_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_17_U1_Y), .B0_t (OUT_ciphertext[17]), .Z0_t (LED_128_Instance_addconst_out[17]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_18_U1_XOR1_U1 ( .A0_t (OUT_ciphertext[18]), .B0_t (LED_128_Instance_addroundkey_tmp[18]), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_18_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_18_U1_AND1_U1 ( .A0_t (LED_128_Instance_n23), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_18_U1_X), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_18_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_18_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_18_U1_Y), .B0_t (OUT_ciphertext[18]), .Z0_t (LED_128_Instance_addconst_out[18]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_19_U1_XOR1_U1 ( .A0_t (OUT_ciphertext[19]), .B0_t (LED_128_Instance_addroundkey_tmp[19]), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_19_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_19_U1_AND1_U1 ( .A0_t (LED_128_Instance_n23), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_19_U1_X), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_19_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_19_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_19_U1_Y), .B0_t (OUT_ciphertext[19]), .Z0_t (LED_128_Instance_addroundkey_out[19]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_20_U1_XOR1_U1 ( .A0_t (OUT_ciphertext[20]), .B0_t (LED_128_Instance_addroundkey_tmp[20]), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_20_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_20_U1_AND1_U1 ( .A0_t (LED_128_Instance_n23), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_20_U1_X), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_20_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_20_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_20_U1_Y), .B0_t (OUT_ciphertext[20]), .Z0_t (LED_128_Instance_addroundkey_out[20]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_21_U1_XOR1_U1 ( .A0_t (OUT_ciphertext[21]), .B0_t (LED_128_Instance_addroundkey_tmp[21]), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_21_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_21_U1_AND1_U1 ( .A0_t (LED_128_Instance_n23), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_21_U1_X), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_21_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_21_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_21_U1_Y), .B0_t (OUT_ciphertext[21]), .Z0_t (LED_128_Instance_addroundkey_out[21]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_22_U1_XOR1_U1 ( .A0_t (OUT_ciphertext[22]), .B0_t (LED_128_Instance_addroundkey_tmp[22]), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_22_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_22_U1_AND1_U1 ( .A0_t (LED_128_Instance_n23), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_22_U1_X), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_22_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_22_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_22_U1_Y), .B0_t (OUT_ciphertext[22]), .Z0_t (LED_128_Instance_addroundkey_out[22]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_23_U1_XOR1_U1 ( .A0_t (OUT_ciphertext[23]), .B0_t (LED_128_Instance_addroundkey_tmp[23]), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_23_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_23_U1_AND1_U1 ( .A0_t (LED_128_Instance_n23), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_23_U1_X), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_23_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_23_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_23_U1_Y), .B0_t (OUT_ciphertext[23]), .Z0_t (LED_128_Instance_addconst_out[23]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_24_U1_XOR1_U1 ( .A0_t (OUT_ciphertext[24]), .B0_t (LED_128_Instance_addroundkey_tmp[24]), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_24_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_24_U1_AND1_U1 ( .A0_t (LED_128_Instance_n23), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_24_U1_X), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_24_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_24_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_24_U1_Y), .B0_t (OUT_ciphertext[24]), .Z0_t (LED_128_Instance_addconst_out[24]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_25_U1_XOR1_U1 ( .A0_t (OUT_ciphertext[25]), .B0_t (LED_128_Instance_addroundkey_tmp[25]), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_25_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_25_U1_AND1_U1 ( .A0_t (LED_128_Instance_n23), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_25_U1_X), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_25_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_25_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_25_U1_Y), .B0_t (OUT_ciphertext[25]), .Z0_t (LED_128_Instance_addconst_out[25]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_26_U1_XOR1_U1 ( .A0_t (OUT_ciphertext[26]), .B0_t (LED_128_Instance_addroundkey_tmp[26]), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_26_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_26_U1_AND1_U1 ( .A0_t (LED_128_Instance_n23), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_26_U1_X), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_26_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_26_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_26_U1_Y), .B0_t (OUT_ciphertext[26]), .Z0_t (LED_128_Instance_addconst_out[26]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_27_U1_XOR1_U1 ( .A0_t (OUT_ciphertext[27]), .B0_t (LED_128_Instance_addroundkey_tmp[27]), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_27_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_27_U1_AND1_U1 ( .A0_t (LED_128_Instance_n23), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_27_U1_X), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_27_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_27_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_27_U1_Y), .B0_t (OUT_ciphertext[27]), .Z0_t (LED_128_Instance_addconst_out[27]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_28_U1_XOR1_U1 ( .A0_t (OUT_ciphertext[28]), .B0_t (LED_128_Instance_addroundkey_tmp[28]), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_28_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_28_U1_AND1_U1 ( .A0_t (LED_128_Instance_n23), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_28_U1_X), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_28_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_28_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_28_U1_Y), .B0_t (OUT_ciphertext[28]), .Z0_t (LED_128_Instance_addconst_out[28]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_29_U1_XOR1_U1 ( .A0_t (OUT_ciphertext[29]), .B0_t (LED_128_Instance_addroundkey_tmp[29]), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_29_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_29_U1_AND1_U1 ( .A0_t (LED_128_Instance_n23), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_29_U1_X), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_29_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_29_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_29_U1_Y), .B0_t (OUT_ciphertext[29]), .Z0_t (LED_128_Instance_addconst_out[29]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_30_U1_XOR1_U1 ( .A0_t (OUT_ciphertext[30]), .B0_t (LED_128_Instance_addroundkey_tmp[30]), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_30_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_30_U1_AND1_U1 ( .A0_t (LED_128_Instance_n23), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_30_U1_X), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_30_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_30_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_30_U1_Y), .B0_t (OUT_ciphertext[30]), .Z0_t (LED_128_Instance_addconst_out[30]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_31_U1_XOR1_U1 ( .A0_t (OUT_ciphertext[31]), .B0_t (LED_128_Instance_addroundkey_tmp[31]), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_31_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_31_U1_AND1_U1 ( .A0_t (LED_128_Instance_n23), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_31_U1_X), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_31_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_31_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_31_U1_Y), .B0_t (OUT_ciphertext[31]), .Z0_t (LED_128_Instance_addconst_out[31]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_32_U1_XOR1_U1 ( .A0_t (OUT_ciphertext[32]), .B0_t (LED_128_Instance_addroundkey_tmp[32]), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_32_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_32_U1_AND1_U1 ( .A0_t (LED_128_Instance_n23), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_32_U1_X), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_32_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_32_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_32_U1_Y), .B0_t (OUT_ciphertext[32]), .Z0_t (LED_128_Instance_addconst_out[32]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_33_U1_XOR1_U1 ( .A0_t (OUT_ciphertext[33]), .B0_t (LED_128_Instance_addroundkey_tmp[33]), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_33_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_33_U1_AND1_U1 ( .A0_t (LED_128_Instance_n23), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_33_U1_X), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_33_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_33_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_33_U1_Y), .B0_t (OUT_ciphertext[33]), .Z0_t (LED_128_Instance_addroundkey_out[33]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_34_U1_XOR1_U1 ( .A0_t (OUT_ciphertext[34]), .B0_t (LED_128_Instance_addroundkey_tmp[34]), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_34_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_34_U1_AND1_U1 ( .A0_t (LED_128_Instance_n23), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_34_U1_X), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_34_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_34_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_34_U1_Y), .B0_t (OUT_ciphertext[34]), .Z0_t (LED_128_Instance_addconst_out[34]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_35_U1_XOR1_U1 ( .A0_t (OUT_ciphertext[35]), .B0_t (LED_128_Instance_addroundkey_tmp[35]), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_35_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_35_U1_AND1_U1 ( .A0_t (LED_128_Instance_n23), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_35_U1_X), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_35_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_35_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_35_U1_Y), .B0_t (OUT_ciphertext[35]), .Z0_t (LED_128_Instance_addconst_out[35]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_36_U1_XOR1_U1 ( .A0_t (OUT_ciphertext[36]), .B0_t (LED_128_Instance_addroundkey_tmp[36]), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_36_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_36_U1_AND1_U1 ( .A0_t (LED_128_Instance_n23), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_36_U1_X), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_36_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_36_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_36_U1_Y), .B0_t (OUT_ciphertext[36]), .Z0_t (LED_128_Instance_addroundkey_out[36]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_37_U1_XOR1_U1 ( .A0_t (OUT_ciphertext[37]), .B0_t (LED_128_Instance_addroundkey_tmp[37]), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_37_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_37_U1_AND1_U1 ( .A0_t (LED_128_Instance_n23), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_37_U1_X), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_37_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_37_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_37_U1_Y), .B0_t (OUT_ciphertext[37]), .Z0_t (LED_128_Instance_addroundkey_out[37]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_38_U1_XOR1_U1 ( .A0_t (OUT_ciphertext[38]), .B0_t (LED_128_Instance_addroundkey_tmp[38]), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_38_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_38_U1_AND1_U1 ( .A0_t (LED_128_Instance_n23), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_38_U1_X), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_38_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_38_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_38_U1_Y), .B0_t (OUT_ciphertext[38]), .Z0_t (LED_128_Instance_addroundkey_out[38]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_39_U1_XOR1_U1 ( .A0_t (OUT_ciphertext[39]), .B0_t (LED_128_Instance_addroundkey_tmp[39]), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_39_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_39_U1_AND1_U1 ( .A0_t (LED_128_Instance_n23), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_39_U1_X), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_39_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_39_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_39_U1_Y), .B0_t (OUT_ciphertext[39]), .Z0_t (LED_128_Instance_addconst_out[39]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_40_U1_XOR1_U1 ( .A0_t (OUT_ciphertext[40]), .B0_t (LED_128_Instance_addroundkey_tmp[40]), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_40_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_40_U1_AND1_U1 ( .A0_t (LED_128_Instance_n23), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_40_U1_X), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_40_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_40_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_40_U1_Y), .B0_t (OUT_ciphertext[40]), .Z0_t (LED_128_Instance_addconst_out[40]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_41_U1_XOR1_U1 ( .A0_t (OUT_ciphertext[41]), .B0_t (LED_128_Instance_addroundkey_tmp[41]), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_41_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_41_U1_AND1_U1 ( .A0_t (LED_128_Instance_n23), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_41_U1_X), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_41_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_41_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_41_U1_Y), .B0_t (OUT_ciphertext[41]), .Z0_t (LED_128_Instance_addconst_out[41]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_42_U1_XOR1_U1 ( .A0_t (OUT_ciphertext[42]), .B0_t (LED_128_Instance_addroundkey_tmp[42]), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_42_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_42_U1_AND1_U1 ( .A0_t (LED_128_Instance_n23), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_42_U1_X), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_42_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_42_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_42_U1_Y), .B0_t (OUT_ciphertext[42]), .Z0_t (LED_128_Instance_addconst_out[42]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_43_U1_XOR1_U1 ( .A0_t (OUT_ciphertext[43]), .B0_t (LED_128_Instance_addroundkey_tmp[43]), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_43_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_43_U1_AND1_U1 ( .A0_t (LED_128_Instance_n23), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_43_U1_X), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_43_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_43_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_43_U1_Y), .B0_t (OUT_ciphertext[43]), .Z0_t (LED_128_Instance_addconst_out[43]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_44_U1_XOR1_U1 ( .A0_t (OUT_ciphertext[44]), .B0_t (LED_128_Instance_addroundkey_tmp[44]), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_44_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_44_U1_AND1_U1 ( .A0_t (LED_128_Instance_n23), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_44_U1_X), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_44_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_44_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_44_U1_Y), .B0_t (OUT_ciphertext[44]), .Z0_t (LED_128_Instance_addconst_out[44]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_45_U1_XOR1_U1 ( .A0_t (OUT_ciphertext[45]), .B0_t (LED_128_Instance_addroundkey_tmp[45]), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_45_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_45_U1_AND1_U1 ( .A0_t (LED_128_Instance_n23), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_45_U1_X), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_45_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_45_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_45_U1_Y), .B0_t (OUT_ciphertext[45]), .Z0_t (LED_128_Instance_addconst_out[45]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_46_U1_XOR1_U1 ( .A0_t (OUT_ciphertext[46]), .B0_t (LED_128_Instance_addroundkey_tmp[46]), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_46_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_46_U1_AND1_U1 ( .A0_t (LED_128_Instance_n23), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_46_U1_X), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_46_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_46_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_46_U1_Y), .B0_t (OUT_ciphertext[46]), .Z0_t (LED_128_Instance_addconst_out[46]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_47_U1_XOR1_U1 ( .A0_t (OUT_ciphertext[47]), .B0_t (LED_128_Instance_addroundkey_tmp[47]), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_47_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_47_U1_AND1_U1 ( .A0_t (LED_128_Instance_n23), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_47_U1_X), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_47_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_47_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_47_U1_Y), .B0_t (OUT_ciphertext[47]), .Z0_t (LED_128_Instance_addconst_out[47]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_48_U1_XOR1_U1 ( .A0_t (OUT_ciphertext[48]), .B0_t (LED_128_Instance_addroundkey_tmp[48]), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_48_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_48_U1_AND1_U1 ( .A0_t (LED_128_Instance_n23), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_48_U1_X), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_48_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_48_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_48_U1_Y), .B0_t (OUT_ciphertext[48]), .Z0_t (LED_128_Instance_addroundkey_out[48]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_49_U1_XOR1_U1 ( .A0_t (OUT_ciphertext[49]), .B0_t (LED_128_Instance_addroundkey_tmp[49]), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_49_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_49_U1_AND1_U1 ( .A0_t (LED_128_Instance_n23), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_49_U1_X), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_49_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_49_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_49_U1_Y), .B0_t (OUT_ciphertext[49]), .Z0_t (LED_128_Instance_addroundkey_out[49]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_50_U1_XOR1_U1 ( .A0_t (OUT_ciphertext[50]), .B0_t (LED_128_Instance_addroundkey_tmp[50]), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_50_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_50_U1_AND1_U1 ( .A0_t (LED_128_Instance_n23), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_50_U1_X), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_50_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_50_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_50_U1_Y), .B0_t (OUT_ciphertext[50]), .Z0_t (LED_128_Instance_addconst_out[50]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_51_U1_XOR1_U1 ( .A0_t (OUT_ciphertext[51]), .B0_t (LED_128_Instance_addroundkey_tmp[51]), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_51_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_51_U1_AND1_U1 ( .A0_t (LED_128_Instance_n23), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_51_U1_X), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_51_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_51_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_51_U1_Y), .B0_t (OUT_ciphertext[51]), .Z0_t (LED_128_Instance_addconst_out[51]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_52_U1_XOR1_U1 ( .A0_t (OUT_ciphertext[52]), .B0_t (LED_128_Instance_addroundkey_tmp[52]), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_52_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_52_U1_AND1_U1 ( .A0_t (LED_128_Instance_n23), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_52_U1_X), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_52_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_52_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_52_U1_Y), .B0_t (OUT_ciphertext[52]), .Z0_t (LED_128_Instance_addroundkey_out[52]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_53_U1_XOR1_U1 ( .A0_t (OUT_ciphertext[53]), .B0_t (LED_128_Instance_addroundkey_tmp[53]), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_53_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_53_U1_AND1_U1 ( .A0_t (LED_128_Instance_n23), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_53_U1_X), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_53_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_53_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_53_U1_Y), .B0_t (OUT_ciphertext[53]), .Z0_t (LED_128_Instance_addroundkey_out[53]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_54_U1_XOR1_U1 ( .A0_t (OUT_ciphertext[54]), .B0_t (LED_128_Instance_addroundkey_tmp[54]), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_54_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_54_U1_AND1_U1 ( .A0_t (LED_128_Instance_n23), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_54_U1_X), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_54_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_54_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_54_U1_Y), .B0_t (OUT_ciphertext[54]), .Z0_t (LED_128_Instance_addroundkey_out[54]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_55_U1_XOR1_U1 ( .A0_t (OUT_ciphertext[55]), .B0_t (LED_128_Instance_addroundkey_tmp[55]), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_55_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_55_U1_AND1_U1 ( .A0_t (LED_128_Instance_n23), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_55_U1_X), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_55_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_55_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_55_U1_Y), .B0_t (OUT_ciphertext[55]), .Z0_t (LED_128_Instance_addconst_out[55]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_56_U1_XOR1_U1 ( .A0_t (OUT_ciphertext[56]), .B0_t (LED_128_Instance_addroundkey_tmp[56]), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_56_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_56_U1_AND1_U1 ( .A0_t (LED_128_Instance_n23), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_56_U1_X), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_56_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_56_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_56_U1_Y), .B0_t (OUT_ciphertext[56]), .Z0_t (LED_128_Instance_addconst_out[56]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_57_U1_XOR1_U1 ( .A0_t (OUT_ciphertext[57]), .B0_t (LED_128_Instance_addroundkey_tmp[57]), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_57_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_57_U1_AND1_U1 ( .A0_t (LED_128_Instance_n23), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_57_U1_X), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_57_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_57_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_57_U1_Y), .B0_t (OUT_ciphertext[57]), .Z0_t (LED_128_Instance_addconst_out[57]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_58_U1_XOR1_U1 ( .A0_t (OUT_ciphertext[58]), .B0_t (LED_128_Instance_addroundkey_tmp[58]), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_58_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_58_U1_AND1_U1 ( .A0_t (LED_128_Instance_n23), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_58_U1_X), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_58_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_58_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_58_U1_Y), .B0_t (OUT_ciphertext[58]), .Z0_t (LED_128_Instance_addconst_out[58]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_59_U1_XOR1_U1 ( .A0_t (OUT_ciphertext[59]), .B0_t (LED_128_Instance_addroundkey_tmp[59]), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_59_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_59_U1_AND1_U1 ( .A0_t (LED_128_Instance_n23), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_59_U1_X), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_59_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_59_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_59_U1_Y), .B0_t (OUT_ciphertext[59]), .Z0_t (LED_128_Instance_addconst_out[59]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_60_U1_XOR1_U1 ( .A0_t (OUT_ciphertext[60]), .B0_t (LED_128_Instance_addroundkey_tmp[60]), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_60_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_60_U1_AND1_U1 ( .A0_t (LED_128_Instance_n23), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_60_U1_X), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_60_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_60_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_60_U1_Y), .B0_t (OUT_ciphertext[60]), .Z0_t (LED_128_Instance_addconst_out[60]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_61_U1_XOR1_U1 ( .A0_t (OUT_ciphertext[61]), .B0_t (LED_128_Instance_addroundkey_tmp[61]), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_61_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_61_U1_AND1_U1 ( .A0_t (LED_128_Instance_n23), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_61_U1_X), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_61_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_61_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_61_U1_Y), .B0_t (OUT_ciphertext[61]), .Z0_t (LED_128_Instance_addconst_out[61]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_62_U1_XOR1_U1 ( .A0_t (OUT_ciphertext[62]), .B0_t (LED_128_Instance_addroundkey_tmp[62]), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_62_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_62_U1_AND1_U1 ( .A0_t (LED_128_Instance_n23), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_62_U1_X), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_62_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_62_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_62_U1_Y), .B0_t (OUT_ciphertext[62]), .Z0_t (LED_128_Instance_addconst_out[62]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_63_U1_XOR1_U1 ( .A0_t (OUT_ciphertext[63]), .B0_t (LED_128_Instance_addroundkey_tmp[63]), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_63_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_63_U1_AND1_U1 ( .A0_t (LED_128_Instance_n23), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_63_U1_X), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_63_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_63_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_63_U1_Y), .B0_t (OUT_ciphertext[63]), .Z0_t (LED_128_Instance_addconst_out[63]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_AddConstants_instance_U14 ( .A0_t (roundconstant[2]), .B0_t (LED_128_Instance_addroundkey_out[54]), .Z0_t (LED_128_Instance_addconst_out[54]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_AddConstants_instance_U13 ( .A0_t (roundconstant[5]), .B0_t (LED_128_Instance_addroundkey_out[38]), .Z0_t (LED_128_Instance_addconst_out[38]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_AddConstants_instance_U12 ( .A0_t (roundconstant[5]), .B0_t (LED_128_Instance_addroundkey_out[6]), .Z0_t (LED_128_Instance_addconst_out[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_AddConstants_instance_U11 ( .A0_t (roundconstant[2]), .B0_t (LED_128_Instance_addroundkey_out[22]), .Z0_t (LED_128_Instance_addconst_out[22]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_AddConstants_instance_U10 ( .A0_t (roundconstant[3]), .B0_t (LED_128_Instance_addroundkey_out[36]), .Z0_t (LED_128_Instance_addconst_out[36]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_AddConstants_instance_U9 ( .A0_t (roundconstant[3]), .B0_t (LED_128_Instance_addroundkey_out[4]), .Z0_t (LED_128_Instance_addconst_out[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_AddConstants_instance_U8 ( .A0_t (roundconstant[0]), .B0_t (LED_128_Instance_addroundkey_out[52]), .Z0_t (LED_128_Instance_addconst_out[52]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_AddConstants_instance_U7 ( .A0_t (roundconstant[0]), .B0_t (LED_128_Instance_addroundkey_out[20]), .Z0_t (LED_128_Instance_addconst_out[20]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_AddConstants_instance_U6 ( .A0_t (roundconstant[1]), .B0_t (LED_128_Instance_addroundkey_out[53]), .Z0_t (LED_128_Instance_addconst_out[53]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_AddConstants_instance_U5 ( .A0_t (roundconstant[1]), .B0_t (LED_128_Instance_addroundkey_out[21]), .Z0_t (LED_128_Instance_addconst_out[21]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_AddConstants_instance_U4 ( .A0_t (roundconstant[4]), .B0_t (LED_128_Instance_addroundkey_out[37]), .Z0_t (LED_128_Instance_addconst_out[37]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_AddConstants_instance_U3 ( .A0_t (roundconstant[4]), .B0_t (LED_128_Instance_addroundkey_out[5]), .Z0_t (LED_128_Instance_addconst_out[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_0_XOR1_U1 ( .A0_t (LED_128_Instance_addconst_out[2]), .B0_t (LED_128_Instance_addconst_out[1]), .Z0_t (LED_128_Instance_SBox_Instance_0_L0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_0_XOR2_U1 ( .A0_t (LED_128_Instance_addconst_out[1]), .B0_t (LED_128_Instance_addconst_out[0]), .Z0_t (LED_128_Instance_SBox_Instance_0_L1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_0_XOR3_U1 ( .A0_t (LED_128_Instance_SBox_Instance_0_L1), .B0_t (LED_128_Instance_addroundkey_out[3]), .Z0_t (LED_128_Instance_SBox_Instance_0_L2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_SBox_Instance_0_XOR16_U1 ( .A0_t (LED_128_Instance_SBox_Instance_0_T0), .B0_t (LED_128_Instance_SBox_Instance_0_L2), .Z0_t (LED_128_Instance_SBox_Instance_0_Q2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_0_XOR4_U1 ( .A0_t (LED_128_Instance_addroundkey_out[3]), .B0_t (LED_128_Instance_addconst_out[0]), .Z0_t (LED_128_Instance_SBox_Instance_0_L3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_0_XOR5_U1 ( .A0_t (LED_128_Instance_SBox_Instance_0_L3), .B0_t (LED_128_Instance_SBox_Instance_0_L0), .Z0_t (LED_128_Instance_SBox_Instance_0_Q3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_0_XOR6_U1 ( .A0_t (LED_128_Instance_addroundkey_out[3]), .B0_t (LED_128_Instance_addconst_out[1]), .Z0_t (LED_128_Instance_SBox_Instance_0_L4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_0_XOR7_U1 ( .A0_t (LED_128_Instance_SBox_Instance_0_T0), .B0_t (LED_128_Instance_SBox_Instance_0_T2), .Z0_t (LED_128_Instance_SBox_Instance_0_L5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_SBox_Instance_0_XOR8_U1 ( .A0_t (LED_128_Instance_SBox_Instance_0_L4), .B0_t (LED_128_Instance_SBox_Instance_0_L5), .Z0_t (LED_128_Instance_SBox_Instance_0_Q6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_0_XOR9_U1 ( .A0_t (LED_128_Instance_SBox_Instance_0_L1), .B0_t (LED_128_Instance_addconst_out[2]), .Z0_t (LED_128_Instance_SBox_Instance_0_Q7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_0_AND1_U1 ( .A0_t (LED_128_Instance_SBox_Instance_0_L0), .B0_t (LED_128_Instance_addroundkey_out[3]), .Z0_t (LED_128_Instance_SBox_Instance_0_T0) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_0_AND2_U1 ( .A0_t (LED_128_Instance_SBox_Instance_0_Q2), .B0_t (LED_128_Instance_SBox_Instance_0_Q3), .Z0_t (LED_128_Instance_SBox_Instance_0_T1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_0_AND3_U1 ( .A0_t (LED_128_Instance_addconst_out[1]), .B0_t (LED_128_Instance_addconst_out[2]), .Z0_t (LED_128_Instance_SBox_Instance_0_T2) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_0_AND4_U1 ( .A0_t (LED_128_Instance_SBox_Instance_0_Q6), .B0_t (LED_128_Instance_SBox_Instance_0_Q7), .Z0_t (LED_128_Instance_SBox_Instance_0_T3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_0_XOR10_U1 ( .A0_t (LED_128_Instance_SBox_Instance_0_L5), .B0_t (LED_128_Instance_SBox_Instance_0_T3), .Z0_t (LED_128_Instance_SBox_Instance_0_L7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_0_XOR11_U1 ( .A0_t (LED_128_Instance_addconst_out[0]), .B0_t (LED_128_Instance_SBox_Instance_0_L7), .Z0_t (LED_128_Instance_subcells_out[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_0_XOR12_U1 ( .A0_t (LED_128_Instance_SBox_Instance_0_L5), .B0_t (LED_128_Instance_SBox_Instance_0_T1), .Z0_t (LED_128_Instance_SBox_Instance_0_L8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_0_XOR13_U1 ( .A0_t (LED_128_Instance_SBox_Instance_0_L1), .B0_t (LED_128_Instance_SBox_Instance_0_L8), .Z0_t (LED_128_Instance_subcells_out[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_0_XOR14_U1 ( .A0_t (LED_128_Instance_SBox_Instance_0_L4), .B0_t (LED_128_Instance_SBox_Instance_0_T3), .Z0_t (LED_128_Instance_subcells_out[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_0_XOR15_U1 ( .A0_t (LED_128_Instance_SBox_Instance_0_L3), .B0_t (LED_128_Instance_SBox_Instance_0_T2), .Z0_t (LED_128_Instance_subcells_out[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_1_XOR1_U1 ( .A0_t (LED_128_Instance_addconst_out[6]), .B0_t (LED_128_Instance_addconst_out[5]), .Z0_t (LED_128_Instance_SBox_Instance_1_L0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_1_XOR2_U1 ( .A0_t (LED_128_Instance_addconst_out[5]), .B0_t (LED_128_Instance_addconst_out[4]), .Z0_t (LED_128_Instance_SBox_Instance_1_L1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_1_XOR3_U1 ( .A0_t (LED_128_Instance_SBox_Instance_1_L1), .B0_t (LED_128_Instance_addconst_out[7]), .Z0_t (LED_128_Instance_SBox_Instance_1_L2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_SBox_Instance_1_XOR16_U1 ( .A0_t (LED_128_Instance_SBox_Instance_1_T0), .B0_t (LED_128_Instance_SBox_Instance_1_L2), .Z0_t (LED_128_Instance_SBox_Instance_1_Q2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_1_XOR4_U1 ( .A0_t (LED_128_Instance_addconst_out[7]), .B0_t (LED_128_Instance_addconst_out[4]), .Z0_t (LED_128_Instance_SBox_Instance_1_L3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_1_XOR5_U1 ( .A0_t (LED_128_Instance_SBox_Instance_1_L3), .B0_t (LED_128_Instance_SBox_Instance_1_L0), .Z0_t (LED_128_Instance_SBox_Instance_1_Q3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_1_XOR6_U1 ( .A0_t (LED_128_Instance_addconst_out[7]), .B0_t (LED_128_Instance_addconst_out[5]), .Z0_t (LED_128_Instance_SBox_Instance_1_L4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_1_XOR7_U1 ( .A0_t (LED_128_Instance_SBox_Instance_1_T0), .B0_t (LED_128_Instance_SBox_Instance_1_T2), .Z0_t (LED_128_Instance_SBox_Instance_1_L5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_SBox_Instance_1_XOR8_U1 ( .A0_t (LED_128_Instance_SBox_Instance_1_L4), .B0_t (LED_128_Instance_SBox_Instance_1_L5), .Z0_t (LED_128_Instance_SBox_Instance_1_Q6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_1_XOR9_U1 ( .A0_t (LED_128_Instance_SBox_Instance_1_L1), .B0_t (LED_128_Instance_addconst_out[6]), .Z0_t (LED_128_Instance_SBox_Instance_1_Q7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_1_AND1_U1 ( .A0_t (LED_128_Instance_SBox_Instance_1_L0), .B0_t (LED_128_Instance_addconst_out[7]), .Z0_t (LED_128_Instance_SBox_Instance_1_T0) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_1_AND2_U1 ( .A0_t (LED_128_Instance_SBox_Instance_1_Q2), .B0_t (LED_128_Instance_SBox_Instance_1_Q3), .Z0_t (LED_128_Instance_SBox_Instance_1_T1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_1_AND3_U1 ( .A0_t (LED_128_Instance_addconst_out[5]), .B0_t (LED_128_Instance_addconst_out[6]), .Z0_t (LED_128_Instance_SBox_Instance_1_T2) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_1_AND4_U1 ( .A0_t (LED_128_Instance_SBox_Instance_1_Q6), .B0_t (LED_128_Instance_SBox_Instance_1_Q7), .Z0_t (LED_128_Instance_SBox_Instance_1_T3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_1_XOR10_U1 ( .A0_t (LED_128_Instance_SBox_Instance_1_L5), .B0_t (LED_128_Instance_SBox_Instance_1_T3), .Z0_t (LED_128_Instance_SBox_Instance_1_L7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_1_XOR11_U1 ( .A0_t (LED_128_Instance_addconst_out[4]), .B0_t (LED_128_Instance_SBox_Instance_1_L7), .Z0_t (LED_128_Instance_subcells_out[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_1_XOR12_U1 ( .A0_t (LED_128_Instance_SBox_Instance_1_L5), .B0_t (LED_128_Instance_SBox_Instance_1_T1), .Z0_t (LED_128_Instance_SBox_Instance_1_L8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_1_XOR13_U1 ( .A0_t (LED_128_Instance_SBox_Instance_1_L1), .B0_t (LED_128_Instance_SBox_Instance_1_L8), .Z0_t (LED_128_Instance_subcells_out[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_1_XOR14_U1 ( .A0_t (LED_128_Instance_SBox_Instance_1_L4), .B0_t (LED_128_Instance_SBox_Instance_1_T3), .Z0_t (LED_128_Instance_subcells_out[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_1_XOR15_U1 ( .A0_t (LED_128_Instance_SBox_Instance_1_L3), .B0_t (LED_128_Instance_SBox_Instance_1_T2), .Z0_t (LED_128_Instance_subcells_out[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_2_XOR1_U1 ( .A0_t (LED_128_Instance_addconst_out[10]), .B0_t (LED_128_Instance_addconst_out[9]), .Z0_t (LED_128_Instance_SBox_Instance_2_L0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_2_XOR2_U1 ( .A0_t (LED_128_Instance_addconst_out[9]), .B0_t (LED_128_Instance_addconst_out[8]), .Z0_t (LED_128_Instance_SBox_Instance_2_L1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_2_XOR3_U1 ( .A0_t (LED_128_Instance_SBox_Instance_2_L1), .B0_t (LED_128_Instance_addconst_out[11]), .Z0_t (LED_128_Instance_SBox_Instance_2_L2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_SBox_Instance_2_XOR16_U1 ( .A0_t (LED_128_Instance_SBox_Instance_2_T0), .B0_t (LED_128_Instance_SBox_Instance_2_L2), .Z0_t (LED_128_Instance_SBox_Instance_2_Q2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_2_XOR4_U1 ( .A0_t (LED_128_Instance_addconst_out[11]), .B0_t (LED_128_Instance_addconst_out[8]), .Z0_t (LED_128_Instance_SBox_Instance_2_L3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_2_XOR5_U1 ( .A0_t (LED_128_Instance_SBox_Instance_2_L3), .B0_t (LED_128_Instance_SBox_Instance_2_L0), .Z0_t (LED_128_Instance_SBox_Instance_2_Q3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_2_XOR6_U1 ( .A0_t (LED_128_Instance_addconst_out[11]), .B0_t (LED_128_Instance_addconst_out[9]), .Z0_t (LED_128_Instance_SBox_Instance_2_L4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_2_XOR7_U1 ( .A0_t (LED_128_Instance_SBox_Instance_2_T0), .B0_t (LED_128_Instance_SBox_Instance_2_T2), .Z0_t (LED_128_Instance_SBox_Instance_2_L5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_SBox_Instance_2_XOR8_U1 ( .A0_t (LED_128_Instance_SBox_Instance_2_L4), .B0_t (LED_128_Instance_SBox_Instance_2_L5), .Z0_t (LED_128_Instance_SBox_Instance_2_Q6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_2_XOR9_U1 ( .A0_t (LED_128_Instance_SBox_Instance_2_L1), .B0_t (LED_128_Instance_addconst_out[10]), .Z0_t (LED_128_Instance_SBox_Instance_2_Q7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_2_AND1_U1 ( .A0_t (LED_128_Instance_SBox_Instance_2_L0), .B0_t (LED_128_Instance_addconst_out[11]), .Z0_t (LED_128_Instance_SBox_Instance_2_T0) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_2_AND2_U1 ( .A0_t (LED_128_Instance_SBox_Instance_2_Q2), .B0_t (LED_128_Instance_SBox_Instance_2_Q3), .Z0_t (LED_128_Instance_SBox_Instance_2_T1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_2_AND3_U1 ( .A0_t (LED_128_Instance_addconst_out[9]), .B0_t (LED_128_Instance_addconst_out[10]), .Z0_t (LED_128_Instance_SBox_Instance_2_T2) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_2_AND4_U1 ( .A0_t (LED_128_Instance_SBox_Instance_2_Q6), .B0_t (LED_128_Instance_SBox_Instance_2_Q7), .Z0_t (LED_128_Instance_SBox_Instance_2_T3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_2_XOR10_U1 ( .A0_t (LED_128_Instance_SBox_Instance_2_L5), .B0_t (LED_128_Instance_SBox_Instance_2_T3), .Z0_t (LED_128_Instance_SBox_Instance_2_L7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_2_XOR11_U1 ( .A0_t (LED_128_Instance_addconst_out[8]), .B0_t (LED_128_Instance_SBox_Instance_2_L7), .Z0_t (LED_128_Instance_subcells_out[11]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_2_XOR12_U1 ( .A0_t (LED_128_Instance_SBox_Instance_2_L5), .B0_t (LED_128_Instance_SBox_Instance_2_T1), .Z0_t (LED_128_Instance_SBox_Instance_2_L8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_2_XOR13_U1 ( .A0_t (LED_128_Instance_SBox_Instance_2_L1), .B0_t (LED_128_Instance_SBox_Instance_2_L8), .Z0_t (LED_128_Instance_subcells_out[10]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_2_XOR14_U1 ( .A0_t (LED_128_Instance_SBox_Instance_2_L4), .B0_t (LED_128_Instance_SBox_Instance_2_T3), .Z0_t (LED_128_Instance_subcells_out[9]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_2_XOR15_U1 ( .A0_t (LED_128_Instance_SBox_Instance_2_L3), .B0_t (LED_128_Instance_SBox_Instance_2_T2), .Z0_t (LED_128_Instance_subcells_out[8]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_3_XOR1_U1 ( .A0_t (LED_128_Instance_addconst_out[14]), .B0_t (LED_128_Instance_addconst_out[13]), .Z0_t (LED_128_Instance_SBox_Instance_3_L0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_3_XOR2_U1 ( .A0_t (LED_128_Instance_addconst_out[13]), .B0_t (LED_128_Instance_addconst_out[12]), .Z0_t (LED_128_Instance_SBox_Instance_3_L1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_3_XOR3_U1 ( .A0_t (LED_128_Instance_SBox_Instance_3_L1), .B0_t (LED_128_Instance_addconst_out[15]), .Z0_t (LED_128_Instance_SBox_Instance_3_L2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_SBox_Instance_3_XOR16_U1 ( .A0_t (LED_128_Instance_SBox_Instance_3_T0), .B0_t (LED_128_Instance_SBox_Instance_3_L2), .Z0_t (LED_128_Instance_SBox_Instance_3_Q2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_3_XOR4_U1 ( .A0_t (LED_128_Instance_addconst_out[15]), .B0_t (LED_128_Instance_addconst_out[12]), .Z0_t (LED_128_Instance_SBox_Instance_3_L3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_3_XOR5_U1 ( .A0_t (LED_128_Instance_SBox_Instance_3_L3), .B0_t (LED_128_Instance_SBox_Instance_3_L0), .Z0_t (LED_128_Instance_SBox_Instance_3_Q3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_3_XOR6_U1 ( .A0_t (LED_128_Instance_addconst_out[15]), .B0_t (LED_128_Instance_addconst_out[13]), .Z0_t (LED_128_Instance_SBox_Instance_3_L4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_3_XOR7_U1 ( .A0_t (LED_128_Instance_SBox_Instance_3_T0), .B0_t (LED_128_Instance_SBox_Instance_3_T2), .Z0_t (LED_128_Instance_SBox_Instance_3_L5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_SBox_Instance_3_XOR8_U1 ( .A0_t (LED_128_Instance_SBox_Instance_3_L4), .B0_t (LED_128_Instance_SBox_Instance_3_L5), .Z0_t (LED_128_Instance_SBox_Instance_3_Q6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_3_XOR9_U1 ( .A0_t (LED_128_Instance_SBox_Instance_3_L1), .B0_t (LED_128_Instance_addconst_out[14]), .Z0_t (LED_128_Instance_SBox_Instance_3_Q7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_3_AND1_U1 ( .A0_t (LED_128_Instance_SBox_Instance_3_L0), .B0_t (LED_128_Instance_addconst_out[15]), .Z0_t (LED_128_Instance_SBox_Instance_3_T0) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_3_AND2_U1 ( .A0_t (LED_128_Instance_SBox_Instance_3_Q2), .B0_t (LED_128_Instance_SBox_Instance_3_Q3), .Z0_t (LED_128_Instance_SBox_Instance_3_T1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_3_AND3_U1 ( .A0_t (LED_128_Instance_addconst_out[13]), .B0_t (LED_128_Instance_addconst_out[14]), .Z0_t (LED_128_Instance_SBox_Instance_3_T2) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_3_AND4_U1 ( .A0_t (LED_128_Instance_SBox_Instance_3_Q6), .B0_t (LED_128_Instance_SBox_Instance_3_Q7), .Z0_t (LED_128_Instance_SBox_Instance_3_T3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_3_XOR10_U1 ( .A0_t (LED_128_Instance_SBox_Instance_3_L5), .B0_t (LED_128_Instance_SBox_Instance_3_T3), .Z0_t (LED_128_Instance_SBox_Instance_3_L7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_3_XOR11_U1 ( .A0_t (LED_128_Instance_addconst_out[12]), .B0_t (LED_128_Instance_SBox_Instance_3_L7), .Z0_t (LED_128_Instance_subcells_out[15]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_3_XOR12_U1 ( .A0_t (LED_128_Instance_SBox_Instance_3_L5), .B0_t (LED_128_Instance_SBox_Instance_3_T1), .Z0_t (LED_128_Instance_SBox_Instance_3_L8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_3_XOR13_U1 ( .A0_t (LED_128_Instance_SBox_Instance_3_L1), .B0_t (LED_128_Instance_SBox_Instance_3_L8), .Z0_t (LED_128_Instance_subcells_out[14]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_3_XOR14_U1 ( .A0_t (LED_128_Instance_SBox_Instance_3_L4), .B0_t (LED_128_Instance_SBox_Instance_3_T3), .Z0_t (LED_128_Instance_subcells_out[13]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_3_XOR15_U1 ( .A0_t (LED_128_Instance_SBox_Instance_3_L3), .B0_t (LED_128_Instance_SBox_Instance_3_T2), .Z0_t (LED_128_Instance_subcells_out[12]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_4_XOR1_U1 ( .A0_t (LED_128_Instance_addconst_out[18]), .B0_t (LED_128_Instance_addconst_out[17]), .Z0_t (LED_128_Instance_SBox_Instance_4_L0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_4_XOR2_U1 ( .A0_t (LED_128_Instance_addconst_out[17]), .B0_t (LED_128_Instance_addroundkey_out[16]), .Z0_t (LED_128_Instance_SBox_Instance_4_L1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_4_XOR3_U1 ( .A0_t (LED_128_Instance_SBox_Instance_4_L1), .B0_t (LED_128_Instance_addroundkey_out[19]), .Z0_t (LED_128_Instance_SBox_Instance_4_L2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_SBox_Instance_4_XOR16_U1 ( .A0_t (LED_128_Instance_SBox_Instance_4_T0), .B0_t (LED_128_Instance_SBox_Instance_4_L2), .Z0_t (LED_128_Instance_SBox_Instance_4_Q2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_4_XOR4_U1 ( .A0_t (LED_128_Instance_addroundkey_out[19]), .B0_t (LED_128_Instance_addroundkey_out[16]), .Z0_t (LED_128_Instance_SBox_Instance_4_L3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_4_XOR5_U1 ( .A0_t (LED_128_Instance_SBox_Instance_4_L3), .B0_t (LED_128_Instance_SBox_Instance_4_L0), .Z0_t (LED_128_Instance_SBox_Instance_4_Q3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_4_XOR6_U1 ( .A0_t (LED_128_Instance_addroundkey_out[19]), .B0_t (LED_128_Instance_addconst_out[17]), .Z0_t (LED_128_Instance_SBox_Instance_4_L4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_4_XOR7_U1 ( .A0_t (LED_128_Instance_SBox_Instance_4_T0), .B0_t (LED_128_Instance_SBox_Instance_4_T2), .Z0_t (LED_128_Instance_SBox_Instance_4_L5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_SBox_Instance_4_XOR8_U1 ( .A0_t (LED_128_Instance_SBox_Instance_4_L4), .B0_t (LED_128_Instance_SBox_Instance_4_L5), .Z0_t (LED_128_Instance_SBox_Instance_4_Q6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_4_XOR9_U1 ( .A0_t (LED_128_Instance_SBox_Instance_4_L1), .B0_t (LED_128_Instance_addconst_out[18]), .Z0_t (LED_128_Instance_SBox_Instance_4_Q7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_4_AND1_U1 ( .A0_t (LED_128_Instance_SBox_Instance_4_L0), .B0_t (LED_128_Instance_addroundkey_out[19]), .Z0_t (LED_128_Instance_SBox_Instance_4_T0) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_4_AND2_U1 ( .A0_t (LED_128_Instance_SBox_Instance_4_Q2), .B0_t (LED_128_Instance_SBox_Instance_4_Q3), .Z0_t (LED_128_Instance_SBox_Instance_4_T1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_4_AND3_U1 ( .A0_t (LED_128_Instance_addconst_out[17]), .B0_t (LED_128_Instance_addconst_out[18]), .Z0_t (LED_128_Instance_SBox_Instance_4_T2) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_4_AND4_U1 ( .A0_t (LED_128_Instance_SBox_Instance_4_Q6), .B0_t (LED_128_Instance_SBox_Instance_4_Q7), .Z0_t (LED_128_Instance_SBox_Instance_4_T3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_4_XOR10_U1 ( .A0_t (LED_128_Instance_SBox_Instance_4_L5), .B0_t (LED_128_Instance_SBox_Instance_4_T3), .Z0_t (LED_128_Instance_SBox_Instance_4_L7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_4_XOR11_U1 ( .A0_t (LED_128_Instance_addroundkey_out[16]), .B0_t (LED_128_Instance_SBox_Instance_4_L7), .Z0_t (LED_128_Instance_subcells_out[19]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_4_XOR12_U1 ( .A0_t (LED_128_Instance_SBox_Instance_4_L5), .B0_t (LED_128_Instance_SBox_Instance_4_T1), .Z0_t (LED_128_Instance_SBox_Instance_4_L8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_4_XOR13_U1 ( .A0_t (LED_128_Instance_SBox_Instance_4_L1), .B0_t (LED_128_Instance_SBox_Instance_4_L8), .Z0_t (LED_128_Instance_subcells_out[18]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_4_XOR14_U1 ( .A0_t (LED_128_Instance_SBox_Instance_4_L4), .B0_t (LED_128_Instance_SBox_Instance_4_T3), .Z0_t (LED_128_Instance_subcells_out[17]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_4_XOR15_U1 ( .A0_t (LED_128_Instance_SBox_Instance_4_L3), .B0_t (LED_128_Instance_SBox_Instance_4_T2), .Z0_t (LED_128_Instance_subcells_out[16]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_5_XOR1_U1 ( .A0_t (LED_128_Instance_addconst_out[22]), .B0_t (LED_128_Instance_addconst_out[21]), .Z0_t (LED_128_Instance_SBox_Instance_5_L0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_5_XOR2_U1 ( .A0_t (LED_128_Instance_addconst_out[21]), .B0_t (LED_128_Instance_addconst_out[20]), .Z0_t (LED_128_Instance_SBox_Instance_5_L1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_5_XOR3_U1 ( .A0_t (LED_128_Instance_SBox_Instance_5_L1), .B0_t (LED_128_Instance_addconst_out[23]), .Z0_t (LED_128_Instance_SBox_Instance_5_L2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_SBox_Instance_5_XOR16_U1 ( .A0_t (LED_128_Instance_SBox_Instance_5_T0), .B0_t (LED_128_Instance_SBox_Instance_5_L2), .Z0_t (LED_128_Instance_SBox_Instance_5_Q2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_5_XOR4_U1 ( .A0_t (LED_128_Instance_addconst_out[23]), .B0_t (LED_128_Instance_addconst_out[20]), .Z0_t (LED_128_Instance_SBox_Instance_5_L3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_5_XOR5_U1 ( .A0_t (LED_128_Instance_SBox_Instance_5_L3), .B0_t (LED_128_Instance_SBox_Instance_5_L0), .Z0_t (LED_128_Instance_SBox_Instance_5_Q3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_5_XOR6_U1 ( .A0_t (LED_128_Instance_addconst_out[23]), .B0_t (LED_128_Instance_addconst_out[21]), .Z0_t (LED_128_Instance_SBox_Instance_5_L4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_5_XOR7_U1 ( .A0_t (LED_128_Instance_SBox_Instance_5_T0), .B0_t (LED_128_Instance_SBox_Instance_5_T2), .Z0_t (LED_128_Instance_SBox_Instance_5_L5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_SBox_Instance_5_XOR8_U1 ( .A0_t (LED_128_Instance_SBox_Instance_5_L4), .B0_t (LED_128_Instance_SBox_Instance_5_L5), .Z0_t (LED_128_Instance_SBox_Instance_5_Q6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_5_XOR9_U1 ( .A0_t (LED_128_Instance_SBox_Instance_5_L1), .B0_t (LED_128_Instance_addconst_out[22]), .Z0_t (LED_128_Instance_SBox_Instance_5_Q7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_5_AND1_U1 ( .A0_t (LED_128_Instance_SBox_Instance_5_L0), .B0_t (LED_128_Instance_addconst_out[23]), .Z0_t (LED_128_Instance_SBox_Instance_5_T0) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_5_AND2_U1 ( .A0_t (LED_128_Instance_SBox_Instance_5_Q2), .B0_t (LED_128_Instance_SBox_Instance_5_Q3), .Z0_t (LED_128_Instance_SBox_Instance_5_T1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_5_AND3_U1 ( .A0_t (LED_128_Instance_addconst_out[21]), .B0_t (LED_128_Instance_addconst_out[22]), .Z0_t (LED_128_Instance_SBox_Instance_5_T2) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_5_AND4_U1 ( .A0_t (LED_128_Instance_SBox_Instance_5_Q6), .B0_t (LED_128_Instance_SBox_Instance_5_Q7), .Z0_t (LED_128_Instance_SBox_Instance_5_T3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_5_XOR10_U1 ( .A0_t (LED_128_Instance_SBox_Instance_5_L5), .B0_t (LED_128_Instance_SBox_Instance_5_T3), .Z0_t (LED_128_Instance_SBox_Instance_5_L7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_5_XOR11_U1 ( .A0_t (LED_128_Instance_addconst_out[20]), .B0_t (LED_128_Instance_SBox_Instance_5_L7), .Z0_t (LED_128_Instance_subcells_out[23]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_5_XOR12_U1 ( .A0_t (LED_128_Instance_SBox_Instance_5_L5), .B0_t (LED_128_Instance_SBox_Instance_5_T1), .Z0_t (LED_128_Instance_SBox_Instance_5_L8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_5_XOR13_U1 ( .A0_t (LED_128_Instance_SBox_Instance_5_L1), .B0_t (LED_128_Instance_SBox_Instance_5_L8), .Z0_t (LED_128_Instance_subcells_out[22]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_5_XOR14_U1 ( .A0_t (LED_128_Instance_SBox_Instance_5_L4), .B0_t (LED_128_Instance_SBox_Instance_5_T3), .Z0_t (LED_128_Instance_subcells_out[21]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_5_XOR15_U1 ( .A0_t (LED_128_Instance_SBox_Instance_5_L3), .B0_t (LED_128_Instance_SBox_Instance_5_T2), .Z0_t (LED_128_Instance_subcells_out[20]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_6_XOR1_U1 ( .A0_t (LED_128_Instance_addconst_out[26]), .B0_t (LED_128_Instance_addconst_out[25]), .Z0_t (LED_128_Instance_SBox_Instance_6_L0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_6_XOR2_U1 ( .A0_t (LED_128_Instance_addconst_out[25]), .B0_t (LED_128_Instance_addconst_out[24]), .Z0_t (LED_128_Instance_SBox_Instance_6_L1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_6_XOR3_U1 ( .A0_t (LED_128_Instance_SBox_Instance_6_L1), .B0_t (LED_128_Instance_addconst_out[27]), .Z0_t (LED_128_Instance_SBox_Instance_6_L2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_SBox_Instance_6_XOR16_U1 ( .A0_t (LED_128_Instance_SBox_Instance_6_T0), .B0_t (LED_128_Instance_SBox_Instance_6_L2), .Z0_t (LED_128_Instance_SBox_Instance_6_Q2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_6_XOR4_U1 ( .A0_t (LED_128_Instance_addconst_out[27]), .B0_t (LED_128_Instance_addconst_out[24]), .Z0_t (LED_128_Instance_SBox_Instance_6_L3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_6_XOR5_U1 ( .A0_t (LED_128_Instance_SBox_Instance_6_L3), .B0_t (LED_128_Instance_SBox_Instance_6_L0), .Z0_t (LED_128_Instance_SBox_Instance_6_Q3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_6_XOR6_U1 ( .A0_t (LED_128_Instance_addconst_out[27]), .B0_t (LED_128_Instance_addconst_out[25]), .Z0_t (LED_128_Instance_SBox_Instance_6_L4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_6_XOR7_U1 ( .A0_t (LED_128_Instance_SBox_Instance_6_T0), .B0_t (LED_128_Instance_SBox_Instance_6_T2), .Z0_t (LED_128_Instance_SBox_Instance_6_L5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_SBox_Instance_6_XOR8_U1 ( .A0_t (LED_128_Instance_SBox_Instance_6_L4), .B0_t (LED_128_Instance_SBox_Instance_6_L5), .Z0_t (LED_128_Instance_SBox_Instance_6_Q6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_6_XOR9_U1 ( .A0_t (LED_128_Instance_SBox_Instance_6_L1), .B0_t (LED_128_Instance_addconst_out[26]), .Z0_t (LED_128_Instance_SBox_Instance_6_Q7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_6_AND1_U1 ( .A0_t (LED_128_Instance_SBox_Instance_6_L0), .B0_t (LED_128_Instance_addconst_out[27]), .Z0_t (LED_128_Instance_SBox_Instance_6_T0) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_6_AND2_U1 ( .A0_t (LED_128_Instance_SBox_Instance_6_Q2), .B0_t (LED_128_Instance_SBox_Instance_6_Q3), .Z0_t (LED_128_Instance_SBox_Instance_6_T1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_6_AND3_U1 ( .A0_t (LED_128_Instance_addconst_out[25]), .B0_t (LED_128_Instance_addconst_out[26]), .Z0_t (LED_128_Instance_SBox_Instance_6_T2) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_6_AND4_U1 ( .A0_t (LED_128_Instance_SBox_Instance_6_Q6), .B0_t (LED_128_Instance_SBox_Instance_6_Q7), .Z0_t (LED_128_Instance_SBox_Instance_6_T3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_6_XOR10_U1 ( .A0_t (LED_128_Instance_SBox_Instance_6_L5), .B0_t (LED_128_Instance_SBox_Instance_6_T3), .Z0_t (LED_128_Instance_SBox_Instance_6_L7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_6_XOR11_U1 ( .A0_t (LED_128_Instance_addconst_out[24]), .B0_t (LED_128_Instance_SBox_Instance_6_L7), .Z0_t (LED_128_Instance_subcells_out[27]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_6_XOR12_U1 ( .A0_t (LED_128_Instance_SBox_Instance_6_L5), .B0_t (LED_128_Instance_SBox_Instance_6_T1), .Z0_t (LED_128_Instance_SBox_Instance_6_L8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_6_XOR13_U1 ( .A0_t (LED_128_Instance_SBox_Instance_6_L1), .B0_t (LED_128_Instance_SBox_Instance_6_L8), .Z0_t (LED_128_Instance_subcells_out[26]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_6_XOR14_U1 ( .A0_t (LED_128_Instance_SBox_Instance_6_L4), .B0_t (LED_128_Instance_SBox_Instance_6_T3), .Z0_t (LED_128_Instance_subcells_out[25]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_6_XOR15_U1 ( .A0_t (LED_128_Instance_SBox_Instance_6_L3), .B0_t (LED_128_Instance_SBox_Instance_6_T2), .Z0_t (LED_128_Instance_subcells_out[24]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_7_XOR1_U1 ( .A0_t (LED_128_Instance_addconst_out[30]), .B0_t (LED_128_Instance_addconst_out[29]), .Z0_t (LED_128_Instance_SBox_Instance_7_L0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_7_XOR2_U1 ( .A0_t (LED_128_Instance_addconst_out[29]), .B0_t (LED_128_Instance_addconst_out[28]), .Z0_t (LED_128_Instance_SBox_Instance_7_L1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_7_XOR3_U1 ( .A0_t (LED_128_Instance_SBox_Instance_7_L1), .B0_t (LED_128_Instance_addconst_out[31]), .Z0_t (LED_128_Instance_SBox_Instance_7_L2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_SBox_Instance_7_XOR16_U1 ( .A0_t (LED_128_Instance_SBox_Instance_7_T0), .B0_t (LED_128_Instance_SBox_Instance_7_L2), .Z0_t (LED_128_Instance_SBox_Instance_7_Q2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_7_XOR4_U1 ( .A0_t (LED_128_Instance_addconst_out[31]), .B0_t (LED_128_Instance_addconst_out[28]), .Z0_t (LED_128_Instance_SBox_Instance_7_L3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_7_XOR5_U1 ( .A0_t (LED_128_Instance_SBox_Instance_7_L3), .B0_t (LED_128_Instance_SBox_Instance_7_L0), .Z0_t (LED_128_Instance_SBox_Instance_7_Q3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_7_XOR6_U1 ( .A0_t (LED_128_Instance_addconst_out[31]), .B0_t (LED_128_Instance_addconst_out[29]), .Z0_t (LED_128_Instance_SBox_Instance_7_L4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_7_XOR7_U1 ( .A0_t (LED_128_Instance_SBox_Instance_7_T0), .B0_t (LED_128_Instance_SBox_Instance_7_T2), .Z0_t (LED_128_Instance_SBox_Instance_7_L5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_SBox_Instance_7_XOR8_U1 ( .A0_t (LED_128_Instance_SBox_Instance_7_L4), .B0_t (LED_128_Instance_SBox_Instance_7_L5), .Z0_t (LED_128_Instance_SBox_Instance_7_Q6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_7_XOR9_U1 ( .A0_t (LED_128_Instance_SBox_Instance_7_L1), .B0_t (LED_128_Instance_addconst_out[30]), .Z0_t (LED_128_Instance_SBox_Instance_7_Q7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_7_AND1_U1 ( .A0_t (LED_128_Instance_SBox_Instance_7_L0), .B0_t (LED_128_Instance_addconst_out[31]), .Z0_t (LED_128_Instance_SBox_Instance_7_T0) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_7_AND2_U1 ( .A0_t (LED_128_Instance_SBox_Instance_7_Q2), .B0_t (LED_128_Instance_SBox_Instance_7_Q3), .Z0_t (LED_128_Instance_SBox_Instance_7_T1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_7_AND3_U1 ( .A0_t (LED_128_Instance_addconst_out[29]), .B0_t (LED_128_Instance_addconst_out[30]), .Z0_t (LED_128_Instance_SBox_Instance_7_T2) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_7_AND4_U1 ( .A0_t (LED_128_Instance_SBox_Instance_7_Q6), .B0_t (LED_128_Instance_SBox_Instance_7_Q7), .Z0_t (LED_128_Instance_SBox_Instance_7_T3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_7_XOR10_U1 ( .A0_t (LED_128_Instance_SBox_Instance_7_L5), .B0_t (LED_128_Instance_SBox_Instance_7_T3), .Z0_t (LED_128_Instance_SBox_Instance_7_L7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_7_XOR11_U1 ( .A0_t (LED_128_Instance_addconst_out[28]), .B0_t (LED_128_Instance_SBox_Instance_7_L7), .Z0_t (LED_128_Instance_subcells_out[31]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_7_XOR12_U1 ( .A0_t (LED_128_Instance_SBox_Instance_7_L5), .B0_t (LED_128_Instance_SBox_Instance_7_T1), .Z0_t (LED_128_Instance_SBox_Instance_7_L8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_7_XOR13_U1 ( .A0_t (LED_128_Instance_SBox_Instance_7_L1), .B0_t (LED_128_Instance_SBox_Instance_7_L8), .Z0_t (LED_128_Instance_subcells_out[30]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_7_XOR14_U1 ( .A0_t (LED_128_Instance_SBox_Instance_7_L4), .B0_t (LED_128_Instance_SBox_Instance_7_T3), .Z0_t (LED_128_Instance_subcells_out[29]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_7_XOR15_U1 ( .A0_t (LED_128_Instance_SBox_Instance_7_L3), .B0_t (LED_128_Instance_SBox_Instance_7_T2), .Z0_t (LED_128_Instance_subcells_out[28]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_8_XOR1_U1 ( .A0_t (LED_128_Instance_addconst_out[34]), .B0_t (LED_128_Instance_addroundkey_out[33]), .Z0_t (LED_128_Instance_SBox_Instance_8_L0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_8_XOR2_U1 ( .A0_t (LED_128_Instance_addroundkey_out[33]), .B0_t (LED_128_Instance_addconst_out[32]), .Z0_t (LED_128_Instance_SBox_Instance_8_L1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_8_XOR3_U1 ( .A0_t (LED_128_Instance_SBox_Instance_8_L1), .B0_t (LED_128_Instance_addconst_out[35]), .Z0_t (LED_128_Instance_SBox_Instance_8_L2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_SBox_Instance_8_XOR16_U1 ( .A0_t (LED_128_Instance_SBox_Instance_8_T0), .B0_t (LED_128_Instance_SBox_Instance_8_L2), .Z0_t (LED_128_Instance_SBox_Instance_8_Q2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_8_XOR4_U1 ( .A0_t (LED_128_Instance_addconst_out[35]), .B0_t (LED_128_Instance_addconst_out[32]), .Z0_t (LED_128_Instance_SBox_Instance_8_L3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_8_XOR5_U1 ( .A0_t (LED_128_Instance_SBox_Instance_8_L3), .B0_t (LED_128_Instance_SBox_Instance_8_L0), .Z0_t (LED_128_Instance_SBox_Instance_8_Q3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_8_XOR6_U1 ( .A0_t (LED_128_Instance_addconst_out[35]), .B0_t (LED_128_Instance_addroundkey_out[33]), .Z0_t (LED_128_Instance_SBox_Instance_8_L4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_8_XOR7_U1 ( .A0_t (LED_128_Instance_SBox_Instance_8_T0), .B0_t (LED_128_Instance_SBox_Instance_8_T2), .Z0_t (LED_128_Instance_SBox_Instance_8_L5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_SBox_Instance_8_XOR8_U1 ( .A0_t (LED_128_Instance_SBox_Instance_8_L4), .B0_t (LED_128_Instance_SBox_Instance_8_L5), .Z0_t (LED_128_Instance_SBox_Instance_8_Q6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_8_XOR9_U1 ( .A0_t (LED_128_Instance_SBox_Instance_8_L1), .B0_t (LED_128_Instance_addconst_out[34]), .Z0_t (LED_128_Instance_SBox_Instance_8_Q7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_8_AND1_U1 ( .A0_t (LED_128_Instance_SBox_Instance_8_L0), .B0_t (LED_128_Instance_addconst_out[35]), .Z0_t (LED_128_Instance_SBox_Instance_8_T0) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_8_AND2_U1 ( .A0_t (LED_128_Instance_SBox_Instance_8_Q2), .B0_t (LED_128_Instance_SBox_Instance_8_Q3), .Z0_t (LED_128_Instance_SBox_Instance_8_T1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_8_AND3_U1 ( .A0_t (LED_128_Instance_addroundkey_out[33]), .B0_t (LED_128_Instance_addconst_out[34]), .Z0_t (LED_128_Instance_SBox_Instance_8_T2) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_8_AND4_U1 ( .A0_t (LED_128_Instance_SBox_Instance_8_Q6), .B0_t (LED_128_Instance_SBox_Instance_8_Q7), .Z0_t (LED_128_Instance_SBox_Instance_8_T3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_8_XOR10_U1 ( .A0_t (LED_128_Instance_SBox_Instance_8_L5), .B0_t (LED_128_Instance_SBox_Instance_8_T3), .Z0_t (LED_128_Instance_SBox_Instance_8_L7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_8_XOR11_U1 ( .A0_t (LED_128_Instance_addconst_out[32]), .B0_t (LED_128_Instance_SBox_Instance_8_L7), .Z0_t (LED_128_Instance_subcells_out[35]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_8_XOR12_U1 ( .A0_t (LED_128_Instance_SBox_Instance_8_L5), .B0_t (LED_128_Instance_SBox_Instance_8_T1), .Z0_t (LED_128_Instance_SBox_Instance_8_L8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_8_XOR13_U1 ( .A0_t (LED_128_Instance_SBox_Instance_8_L1), .B0_t (LED_128_Instance_SBox_Instance_8_L8), .Z0_t (LED_128_Instance_subcells_out[34]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_8_XOR14_U1 ( .A0_t (LED_128_Instance_SBox_Instance_8_L4), .B0_t (LED_128_Instance_SBox_Instance_8_T3), .Z0_t (LED_128_Instance_subcells_out[33]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_8_XOR15_U1 ( .A0_t (LED_128_Instance_SBox_Instance_8_L3), .B0_t (LED_128_Instance_SBox_Instance_8_T2), .Z0_t (LED_128_Instance_subcells_out[32]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_9_XOR1_U1 ( .A0_t (LED_128_Instance_addconst_out[38]), .B0_t (LED_128_Instance_addconst_out[37]), .Z0_t (LED_128_Instance_SBox_Instance_9_L0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_9_XOR2_U1 ( .A0_t (LED_128_Instance_addconst_out[37]), .B0_t (LED_128_Instance_addconst_out[36]), .Z0_t (LED_128_Instance_SBox_Instance_9_L1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_9_XOR3_U1 ( .A0_t (LED_128_Instance_SBox_Instance_9_L1), .B0_t (LED_128_Instance_addconst_out[39]), .Z0_t (LED_128_Instance_SBox_Instance_9_L2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_SBox_Instance_9_XOR16_U1 ( .A0_t (LED_128_Instance_SBox_Instance_9_T0), .B0_t (LED_128_Instance_SBox_Instance_9_L2), .Z0_t (LED_128_Instance_SBox_Instance_9_Q2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_9_XOR4_U1 ( .A0_t (LED_128_Instance_addconst_out[39]), .B0_t (LED_128_Instance_addconst_out[36]), .Z0_t (LED_128_Instance_SBox_Instance_9_L3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_9_XOR5_U1 ( .A0_t (LED_128_Instance_SBox_Instance_9_L3), .B0_t (LED_128_Instance_SBox_Instance_9_L0), .Z0_t (LED_128_Instance_SBox_Instance_9_Q3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_9_XOR6_U1 ( .A0_t (LED_128_Instance_addconst_out[39]), .B0_t (LED_128_Instance_addconst_out[37]), .Z0_t (LED_128_Instance_SBox_Instance_9_L4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_9_XOR7_U1 ( .A0_t (LED_128_Instance_SBox_Instance_9_T0), .B0_t (LED_128_Instance_SBox_Instance_9_T2), .Z0_t (LED_128_Instance_SBox_Instance_9_L5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_SBox_Instance_9_XOR8_U1 ( .A0_t (LED_128_Instance_SBox_Instance_9_L4), .B0_t (LED_128_Instance_SBox_Instance_9_L5), .Z0_t (LED_128_Instance_SBox_Instance_9_Q6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_9_XOR9_U1 ( .A0_t (LED_128_Instance_SBox_Instance_9_L1), .B0_t (LED_128_Instance_addconst_out[38]), .Z0_t (LED_128_Instance_SBox_Instance_9_Q7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_9_AND1_U1 ( .A0_t (LED_128_Instance_SBox_Instance_9_L0), .B0_t (LED_128_Instance_addconst_out[39]), .Z0_t (LED_128_Instance_SBox_Instance_9_T0) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_9_AND2_U1 ( .A0_t (LED_128_Instance_SBox_Instance_9_Q2), .B0_t (LED_128_Instance_SBox_Instance_9_Q3), .Z0_t (LED_128_Instance_SBox_Instance_9_T1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_9_AND3_U1 ( .A0_t (LED_128_Instance_addconst_out[37]), .B0_t (LED_128_Instance_addconst_out[38]), .Z0_t (LED_128_Instance_SBox_Instance_9_T2) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_9_AND4_U1 ( .A0_t (LED_128_Instance_SBox_Instance_9_Q6), .B0_t (LED_128_Instance_SBox_Instance_9_Q7), .Z0_t (LED_128_Instance_SBox_Instance_9_T3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_9_XOR10_U1 ( .A0_t (LED_128_Instance_SBox_Instance_9_L5), .B0_t (LED_128_Instance_SBox_Instance_9_T3), .Z0_t (LED_128_Instance_SBox_Instance_9_L7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_9_XOR11_U1 ( .A0_t (LED_128_Instance_addconst_out[36]), .B0_t (LED_128_Instance_SBox_Instance_9_L7), .Z0_t (LED_128_Instance_subcells_out[39]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_9_XOR12_U1 ( .A0_t (LED_128_Instance_SBox_Instance_9_L5), .B0_t (LED_128_Instance_SBox_Instance_9_T1), .Z0_t (LED_128_Instance_SBox_Instance_9_L8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_9_XOR13_U1 ( .A0_t (LED_128_Instance_SBox_Instance_9_L1), .B0_t (LED_128_Instance_SBox_Instance_9_L8), .Z0_t (LED_128_Instance_subcells_out[38]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_9_XOR14_U1 ( .A0_t (LED_128_Instance_SBox_Instance_9_L4), .B0_t (LED_128_Instance_SBox_Instance_9_T3), .Z0_t (LED_128_Instance_subcells_out[37]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_9_XOR15_U1 ( .A0_t (LED_128_Instance_SBox_Instance_9_L3), .B0_t (LED_128_Instance_SBox_Instance_9_T2), .Z0_t (LED_128_Instance_subcells_out[36]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_10_XOR1_U1 ( .A0_t (LED_128_Instance_addconst_out[42]), .B0_t (LED_128_Instance_addconst_out[41]), .Z0_t (LED_128_Instance_SBox_Instance_10_L0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_10_XOR2_U1 ( .A0_t (LED_128_Instance_addconst_out[41]), .B0_t (LED_128_Instance_addconst_out[40]), .Z0_t (LED_128_Instance_SBox_Instance_10_L1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_10_XOR3_U1 ( .A0_t (LED_128_Instance_SBox_Instance_10_L1), .B0_t (LED_128_Instance_addconst_out[43]), .Z0_t (LED_128_Instance_SBox_Instance_10_L2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_SBox_Instance_10_XOR16_U1 ( .A0_t (LED_128_Instance_SBox_Instance_10_T0), .B0_t (LED_128_Instance_SBox_Instance_10_L2), .Z0_t (LED_128_Instance_SBox_Instance_10_Q2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_10_XOR4_U1 ( .A0_t (LED_128_Instance_addconst_out[43]), .B0_t (LED_128_Instance_addconst_out[40]), .Z0_t (LED_128_Instance_SBox_Instance_10_L3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_10_XOR5_U1 ( .A0_t (LED_128_Instance_SBox_Instance_10_L3), .B0_t (LED_128_Instance_SBox_Instance_10_L0), .Z0_t (LED_128_Instance_SBox_Instance_10_Q3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_10_XOR6_U1 ( .A0_t (LED_128_Instance_addconst_out[43]), .B0_t (LED_128_Instance_addconst_out[41]), .Z0_t (LED_128_Instance_SBox_Instance_10_L4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_10_XOR7_U1 ( .A0_t (LED_128_Instance_SBox_Instance_10_T0), .B0_t (LED_128_Instance_SBox_Instance_10_T2), .Z0_t (LED_128_Instance_SBox_Instance_10_L5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_SBox_Instance_10_XOR8_U1 ( .A0_t (LED_128_Instance_SBox_Instance_10_L4), .B0_t (LED_128_Instance_SBox_Instance_10_L5), .Z0_t (LED_128_Instance_SBox_Instance_10_Q6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_10_XOR9_U1 ( .A0_t (LED_128_Instance_SBox_Instance_10_L1), .B0_t (LED_128_Instance_addconst_out[42]), .Z0_t (LED_128_Instance_SBox_Instance_10_Q7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_10_AND1_U1 ( .A0_t (LED_128_Instance_SBox_Instance_10_L0), .B0_t (LED_128_Instance_addconst_out[43]), .Z0_t (LED_128_Instance_SBox_Instance_10_T0) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_10_AND2_U1 ( .A0_t (LED_128_Instance_SBox_Instance_10_Q2), .B0_t (LED_128_Instance_SBox_Instance_10_Q3), .Z0_t (LED_128_Instance_SBox_Instance_10_T1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_10_AND3_U1 ( .A0_t (LED_128_Instance_addconst_out[41]), .B0_t (LED_128_Instance_addconst_out[42]), .Z0_t (LED_128_Instance_SBox_Instance_10_T2) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_10_AND4_U1 ( .A0_t (LED_128_Instance_SBox_Instance_10_Q6), .B0_t (LED_128_Instance_SBox_Instance_10_Q7), .Z0_t (LED_128_Instance_SBox_Instance_10_T3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_10_XOR10_U1 ( .A0_t (LED_128_Instance_SBox_Instance_10_L5), .B0_t (LED_128_Instance_SBox_Instance_10_T3), .Z0_t (LED_128_Instance_SBox_Instance_10_L7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_10_XOR11_U1 ( .A0_t (LED_128_Instance_addconst_out[40]), .B0_t (LED_128_Instance_SBox_Instance_10_L7), .Z0_t (LED_128_Instance_subcells_out[43]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_10_XOR12_U1 ( .A0_t (LED_128_Instance_SBox_Instance_10_L5), .B0_t (LED_128_Instance_SBox_Instance_10_T1), .Z0_t (LED_128_Instance_SBox_Instance_10_L8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_10_XOR13_U1 ( .A0_t (LED_128_Instance_SBox_Instance_10_L1), .B0_t (LED_128_Instance_SBox_Instance_10_L8), .Z0_t (LED_128_Instance_subcells_out[42]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_10_XOR14_U1 ( .A0_t (LED_128_Instance_SBox_Instance_10_L4), .B0_t (LED_128_Instance_SBox_Instance_10_T3), .Z0_t (LED_128_Instance_subcells_out[41]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_10_XOR15_U1 ( .A0_t (LED_128_Instance_SBox_Instance_10_L3), .B0_t (LED_128_Instance_SBox_Instance_10_T2), .Z0_t (LED_128_Instance_subcells_out[40]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_11_XOR1_U1 ( .A0_t (LED_128_Instance_addconst_out[46]), .B0_t (LED_128_Instance_addconst_out[45]), .Z0_t (LED_128_Instance_SBox_Instance_11_L0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_11_XOR2_U1 ( .A0_t (LED_128_Instance_addconst_out[45]), .B0_t (LED_128_Instance_addconst_out[44]), .Z0_t (LED_128_Instance_SBox_Instance_11_L1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_11_XOR3_U1 ( .A0_t (LED_128_Instance_SBox_Instance_11_L1), .B0_t (LED_128_Instance_addconst_out[47]), .Z0_t (LED_128_Instance_SBox_Instance_11_L2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_SBox_Instance_11_XOR16_U1 ( .A0_t (LED_128_Instance_SBox_Instance_11_T0), .B0_t (LED_128_Instance_SBox_Instance_11_L2), .Z0_t (LED_128_Instance_SBox_Instance_11_Q2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_11_XOR4_U1 ( .A0_t (LED_128_Instance_addconst_out[47]), .B0_t (LED_128_Instance_addconst_out[44]), .Z0_t (LED_128_Instance_SBox_Instance_11_L3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_11_XOR5_U1 ( .A0_t (LED_128_Instance_SBox_Instance_11_L3), .B0_t (LED_128_Instance_SBox_Instance_11_L0), .Z0_t (LED_128_Instance_SBox_Instance_11_Q3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_11_XOR6_U1 ( .A0_t (LED_128_Instance_addconst_out[47]), .B0_t (LED_128_Instance_addconst_out[45]), .Z0_t (LED_128_Instance_SBox_Instance_11_L4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_11_XOR7_U1 ( .A0_t (LED_128_Instance_SBox_Instance_11_T0), .B0_t (LED_128_Instance_SBox_Instance_11_T2), .Z0_t (LED_128_Instance_SBox_Instance_11_L5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_SBox_Instance_11_XOR8_U1 ( .A0_t (LED_128_Instance_SBox_Instance_11_L4), .B0_t (LED_128_Instance_SBox_Instance_11_L5), .Z0_t (LED_128_Instance_SBox_Instance_11_Q6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_11_XOR9_U1 ( .A0_t (LED_128_Instance_SBox_Instance_11_L1), .B0_t (LED_128_Instance_addconst_out[46]), .Z0_t (LED_128_Instance_SBox_Instance_11_Q7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_11_AND1_U1 ( .A0_t (LED_128_Instance_SBox_Instance_11_L0), .B0_t (LED_128_Instance_addconst_out[47]), .Z0_t (LED_128_Instance_SBox_Instance_11_T0) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_11_AND2_U1 ( .A0_t (LED_128_Instance_SBox_Instance_11_Q2), .B0_t (LED_128_Instance_SBox_Instance_11_Q3), .Z0_t (LED_128_Instance_SBox_Instance_11_T1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_11_AND3_U1 ( .A0_t (LED_128_Instance_addconst_out[45]), .B0_t (LED_128_Instance_addconst_out[46]), .Z0_t (LED_128_Instance_SBox_Instance_11_T2) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_11_AND4_U1 ( .A0_t (LED_128_Instance_SBox_Instance_11_Q6), .B0_t (LED_128_Instance_SBox_Instance_11_Q7), .Z0_t (LED_128_Instance_SBox_Instance_11_T3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_11_XOR10_U1 ( .A0_t (LED_128_Instance_SBox_Instance_11_L5), .B0_t (LED_128_Instance_SBox_Instance_11_T3), .Z0_t (LED_128_Instance_SBox_Instance_11_L7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_11_XOR11_U1 ( .A0_t (LED_128_Instance_addconst_out[44]), .B0_t (LED_128_Instance_SBox_Instance_11_L7), .Z0_t (LED_128_Instance_subcells_out[47]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_11_XOR12_U1 ( .A0_t (LED_128_Instance_SBox_Instance_11_L5), .B0_t (LED_128_Instance_SBox_Instance_11_T1), .Z0_t (LED_128_Instance_SBox_Instance_11_L8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_11_XOR13_U1 ( .A0_t (LED_128_Instance_SBox_Instance_11_L1), .B0_t (LED_128_Instance_SBox_Instance_11_L8), .Z0_t (LED_128_Instance_subcells_out[46]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_11_XOR14_U1 ( .A0_t (LED_128_Instance_SBox_Instance_11_L4), .B0_t (LED_128_Instance_SBox_Instance_11_T3), .Z0_t (LED_128_Instance_subcells_out[45]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_11_XOR15_U1 ( .A0_t (LED_128_Instance_SBox_Instance_11_L3), .B0_t (LED_128_Instance_SBox_Instance_11_T2), .Z0_t (LED_128_Instance_subcells_out[44]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_12_XOR1_U1 ( .A0_t (LED_128_Instance_addconst_out[50]), .B0_t (LED_128_Instance_addroundkey_out[49]), .Z0_t (LED_128_Instance_SBox_Instance_12_L0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_12_XOR2_U1 ( .A0_t (LED_128_Instance_addroundkey_out[49]), .B0_t (LED_128_Instance_addroundkey_out[48]), .Z0_t (LED_128_Instance_SBox_Instance_12_L1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_12_XOR3_U1 ( .A0_t (LED_128_Instance_SBox_Instance_12_L1), .B0_t (LED_128_Instance_addconst_out[51]), .Z0_t (LED_128_Instance_SBox_Instance_12_L2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_SBox_Instance_12_XOR16_U1 ( .A0_t (LED_128_Instance_SBox_Instance_12_T0), .B0_t (LED_128_Instance_SBox_Instance_12_L2), .Z0_t (LED_128_Instance_SBox_Instance_12_Q2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_12_XOR4_U1 ( .A0_t (LED_128_Instance_addconst_out[51]), .B0_t (LED_128_Instance_addroundkey_out[48]), .Z0_t (LED_128_Instance_SBox_Instance_12_L3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_12_XOR5_U1 ( .A0_t (LED_128_Instance_SBox_Instance_12_L3), .B0_t (LED_128_Instance_SBox_Instance_12_L0), .Z0_t (LED_128_Instance_SBox_Instance_12_Q3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_12_XOR6_U1 ( .A0_t (LED_128_Instance_addconst_out[51]), .B0_t (LED_128_Instance_addroundkey_out[49]), .Z0_t (LED_128_Instance_SBox_Instance_12_L4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_12_XOR7_U1 ( .A0_t (LED_128_Instance_SBox_Instance_12_T0), .B0_t (LED_128_Instance_SBox_Instance_12_T2), .Z0_t (LED_128_Instance_SBox_Instance_12_L5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_SBox_Instance_12_XOR8_U1 ( .A0_t (LED_128_Instance_SBox_Instance_12_L4), .B0_t (LED_128_Instance_SBox_Instance_12_L5), .Z0_t (LED_128_Instance_SBox_Instance_12_Q6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_12_XOR9_U1 ( .A0_t (LED_128_Instance_SBox_Instance_12_L1), .B0_t (LED_128_Instance_addconst_out[50]), .Z0_t (LED_128_Instance_SBox_Instance_12_Q7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_12_AND1_U1 ( .A0_t (LED_128_Instance_SBox_Instance_12_L0), .B0_t (LED_128_Instance_addconst_out[51]), .Z0_t (LED_128_Instance_SBox_Instance_12_T0) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_12_AND2_U1 ( .A0_t (LED_128_Instance_SBox_Instance_12_Q2), .B0_t (LED_128_Instance_SBox_Instance_12_Q3), .Z0_t (LED_128_Instance_SBox_Instance_12_T1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_12_AND3_U1 ( .A0_t (LED_128_Instance_addroundkey_out[49]), .B0_t (LED_128_Instance_addconst_out[50]), .Z0_t (LED_128_Instance_SBox_Instance_12_T2) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_12_AND4_U1 ( .A0_t (LED_128_Instance_SBox_Instance_12_Q6), .B0_t (LED_128_Instance_SBox_Instance_12_Q7), .Z0_t (LED_128_Instance_SBox_Instance_12_T3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_12_XOR10_U1 ( .A0_t (LED_128_Instance_SBox_Instance_12_L5), .B0_t (LED_128_Instance_SBox_Instance_12_T3), .Z0_t (LED_128_Instance_SBox_Instance_12_L7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_12_XOR11_U1 ( .A0_t (LED_128_Instance_addroundkey_out[48]), .B0_t (LED_128_Instance_SBox_Instance_12_L7), .Z0_t (LED_128_Instance_subcells_out[51]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_12_XOR12_U1 ( .A0_t (LED_128_Instance_SBox_Instance_12_L5), .B0_t (LED_128_Instance_SBox_Instance_12_T1), .Z0_t (LED_128_Instance_SBox_Instance_12_L8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_12_XOR13_U1 ( .A0_t (LED_128_Instance_SBox_Instance_12_L1), .B0_t (LED_128_Instance_SBox_Instance_12_L8), .Z0_t (LED_128_Instance_subcells_out[50]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_12_XOR14_U1 ( .A0_t (LED_128_Instance_SBox_Instance_12_L4), .B0_t (LED_128_Instance_SBox_Instance_12_T3), .Z0_t (LED_128_Instance_subcells_out[49]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_12_XOR15_U1 ( .A0_t (LED_128_Instance_SBox_Instance_12_L3), .B0_t (LED_128_Instance_SBox_Instance_12_T2), .Z0_t (LED_128_Instance_subcells_out[48]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_13_XOR1_U1 ( .A0_t (LED_128_Instance_addconst_out[54]), .B0_t (LED_128_Instance_addconst_out[53]), .Z0_t (LED_128_Instance_SBox_Instance_13_L0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_13_XOR2_U1 ( .A0_t (LED_128_Instance_addconst_out[53]), .B0_t (LED_128_Instance_addconst_out[52]), .Z0_t (LED_128_Instance_SBox_Instance_13_L1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_13_XOR3_U1 ( .A0_t (LED_128_Instance_SBox_Instance_13_L1), .B0_t (LED_128_Instance_addconst_out[55]), .Z0_t (LED_128_Instance_SBox_Instance_13_L2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_SBox_Instance_13_XOR16_U1 ( .A0_t (LED_128_Instance_SBox_Instance_13_T0), .B0_t (LED_128_Instance_SBox_Instance_13_L2), .Z0_t (LED_128_Instance_SBox_Instance_13_Q2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_13_XOR4_U1 ( .A0_t (LED_128_Instance_addconst_out[55]), .B0_t (LED_128_Instance_addconst_out[52]), .Z0_t (LED_128_Instance_SBox_Instance_13_L3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_13_XOR5_U1 ( .A0_t (LED_128_Instance_SBox_Instance_13_L3), .B0_t (LED_128_Instance_SBox_Instance_13_L0), .Z0_t (LED_128_Instance_SBox_Instance_13_Q3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_13_XOR6_U1 ( .A0_t (LED_128_Instance_addconst_out[55]), .B0_t (LED_128_Instance_addconst_out[53]), .Z0_t (LED_128_Instance_SBox_Instance_13_L4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_13_XOR7_U1 ( .A0_t (LED_128_Instance_SBox_Instance_13_T0), .B0_t (LED_128_Instance_SBox_Instance_13_T2), .Z0_t (LED_128_Instance_SBox_Instance_13_L5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_SBox_Instance_13_XOR8_U1 ( .A0_t (LED_128_Instance_SBox_Instance_13_L4), .B0_t (LED_128_Instance_SBox_Instance_13_L5), .Z0_t (LED_128_Instance_SBox_Instance_13_Q6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_13_XOR9_U1 ( .A0_t (LED_128_Instance_SBox_Instance_13_L1), .B0_t (LED_128_Instance_addconst_out[54]), .Z0_t (LED_128_Instance_SBox_Instance_13_Q7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_13_AND1_U1 ( .A0_t (LED_128_Instance_SBox_Instance_13_L0), .B0_t (LED_128_Instance_addconst_out[55]), .Z0_t (LED_128_Instance_SBox_Instance_13_T0) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_13_AND2_U1 ( .A0_t (LED_128_Instance_SBox_Instance_13_Q2), .B0_t (LED_128_Instance_SBox_Instance_13_Q3), .Z0_t (LED_128_Instance_SBox_Instance_13_T1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_13_AND3_U1 ( .A0_t (LED_128_Instance_addconst_out[53]), .B0_t (LED_128_Instance_addconst_out[54]), .Z0_t (LED_128_Instance_SBox_Instance_13_T2) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_13_AND4_U1 ( .A0_t (LED_128_Instance_SBox_Instance_13_Q6), .B0_t (LED_128_Instance_SBox_Instance_13_Q7), .Z0_t (LED_128_Instance_SBox_Instance_13_T3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_13_XOR10_U1 ( .A0_t (LED_128_Instance_SBox_Instance_13_L5), .B0_t (LED_128_Instance_SBox_Instance_13_T3), .Z0_t (LED_128_Instance_SBox_Instance_13_L7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_13_XOR11_U1 ( .A0_t (LED_128_Instance_addconst_out[52]), .B0_t (LED_128_Instance_SBox_Instance_13_L7), .Z0_t (LED_128_Instance_subcells_out[55]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_13_XOR12_U1 ( .A0_t (LED_128_Instance_SBox_Instance_13_L5), .B0_t (LED_128_Instance_SBox_Instance_13_T1), .Z0_t (LED_128_Instance_SBox_Instance_13_L8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_13_XOR13_U1 ( .A0_t (LED_128_Instance_SBox_Instance_13_L1), .B0_t (LED_128_Instance_SBox_Instance_13_L8), .Z0_t (LED_128_Instance_subcells_out[54]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_13_XOR14_U1 ( .A0_t (LED_128_Instance_SBox_Instance_13_L4), .B0_t (LED_128_Instance_SBox_Instance_13_T3), .Z0_t (LED_128_Instance_subcells_out[53]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_13_XOR15_U1 ( .A0_t (LED_128_Instance_SBox_Instance_13_L3), .B0_t (LED_128_Instance_SBox_Instance_13_T2), .Z0_t (LED_128_Instance_subcells_out[52]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_14_XOR1_U1 ( .A0_t (LED_128_Instance_addconst_out[58]), .B0_t (LED_128_Instance_addconst_out[57]), .Z0_t (LED_128_Instance_SBox_Instance_14_L0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_14_XOR2_U1 ( .A0_t (LED_128_Instance_addconst_out[57]), .B0_t (LED_128_Instance_addconst_out[56]), .Z0_t (LED_128_Instance_SBox_Instance_14_L1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_14_XOR3_U1 ( .A0_t (LED_128_Instance_SBox_Instance_14_L1), .B0_t (LED_128_Instance_addconst_out[59]), .Z0_t (LED_128_Instance_SBox_Instance_14_L2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_SBox_Instance_14_XOR16_U1 ( .A0_t (LED_128_Instance_SBox_Instance_14_T0), .B0_t (LED_128_Instance_SBox_Instance_14_L2), .Z0_t (LED_128_Instance_SBox_Instance_14_Q2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_14_XOR4_U1 ( .A0_t (LED_128_Instance_addconst_out[59]), .B0_t (LED_128_Instance_addconst_out[56]), .Z0_t (LED_128_Instance_SBox_Instance_14_L3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_14_XOR5_U1 ( .A0_t (LED_128_Instance_SBox_Instance_14_L3), .B0_t (LED_128_Instance_SBox_Instance_14_L0), .Z0_t (LED_128_Instance_SBox_Instance_14_Q3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_14_XOR6_U1 ( .A0_t (LED_128_Instance_addconst_out[59]), .B0_t (LED_128_Instance_addconst_out[57]), .Z0_t (LED_128_Instance_SBox_Instance_14_L4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_14_XOR7_U1 ( .A0_t (LED_128_Instance_SBox_Instance_14_T0), .B0_t (LED_128_Instance_SBox_Instance_14_T2), .Z0_t (LED_128_Instance_SBox_Instance_14_L5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_SBox_Instance_14_XOR8_U1 ( .A0_t (LED_128_Instance_SBox_Instance_14_L4), .B0_t (LED_128_Instance_SBox_Instance_14_L5), .Z0_t (LED_128_Instance_SBox_Instance_14_Q6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_14_XOR9_U1 ( .A0_t (LED_128_Instance_SBox_Instance_14_L1), .B0_t (LED_128_Instance_addconst_out[58]), .Z0_t (LED_128_Instance_SBox_Instance_14_Q7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_14_AND1_U1 ( .A0_t (LED_128_Instance_SBox_Instance_14_L0), .B0_t (LED_128_Instance_addconst_out[59]), .Z0_t (LED_128_Instance_SBox_Instance_14_T0) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_14_AND2_U1 ( .A0_t (LED_128_Instance_SBox_Instance_14_Q2), .B0_t (LED_128_Instance_SBox_Instance_14_Q3), .Z0_t (LED_128_Instance_SBox_Instance_14_T1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_14_AND3_U1 ( .A0_t (LED_128_Instance_addconst_out[57]), .B0_t (LED_128_Instance_addconst_out[58]), .Z0_t (LED_128_Instance_SBox_Instance_14_T2) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_14_AND4_U1 ( .A0_t (LED_128_Instance_SBox_Instance_14_Q6), .B0_t (LED_128_Instance_SBox_Instance_14_Q7), .Z0_t (LED_128_Instance_SBox_Instance_14_T3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_14_XOR10_U1 ( .A0_t (LED_128_Instance_SBox_Instance_14_L5), .B0_t (LED_128_Instance_SBox_Instance_14_T3), .Z0_t (LED_128_Instance_SBox_Instance_14_L7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_14_XOR11_U1 ( .A0_t (LED_128_Instance_addconst_out[56]), .B0_t (LED_128_Instance_SBox_Instance_14_L7), .Z0_t (LED_128_Instance_subcells_out[59]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_14_XOR12_U1 ( .A0_t (LED_128_Instance_SBox_Instance_14_L5), .B0_t (LED_128_Instance_SBox_Instance_14_T1), .Z0_t (LED_128_Instance_SBox_Instance_14_L8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_14_XOR13_U1 ( .A0_t (LED_128_Instance_SBox_Instance_14_L1), .B0_t (LED_128_Instance_SBox_Instance_14_L8), .Z0_t (LED_128_Instance_subcells_out[58]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_14_XOR14_U1 ( .A0_t (LED_128_Instance_SBox_Instance_14_L4), .B0_t (LED_128_Instance_SBox_Instance_14_T3), .Z0_t (LED_128_Instance_subcells_out[57]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_14_XOR15_U1 ( .A0_t (LED_128_Instance_SBox_Instance_14_L3), .B0_t (LED_128_Instance_SBox_Instance_14_T2), .Z0_t (LED_128_Instance_subcells_out[56]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_15_XOR1_U1 ( .A0_t (LED_128_Instance_addconst_out[62]), .B0_t (LED_128_Instance_addconst_out[61]), .Z0_t (LED_128_Instance_SBox_Instance_15_L0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_15_XOR2_U1 ( .A0_t (LED_128_Instance_addconst_out[61]), .B0_t (LED_128_Instance_addconst_out[60]), .Z0_t (LED_128_Instance_SBox_Instance_15_L1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_15_XOR3_U1 ( .A0_t (LED_128_Instance_SBox_Instance_15_L1), .B0_t (LED_128_Instance_addconst_out[63]), .Z0_t (LED_128_Instance_SBox_Instance_15_L2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_SBox_Instance_15_XOR16_U1 ( .A0_t (LED_128_Instance_SBox_Instance_15_T0), .B0_t (LED_128_Instance_SBox_Instance_15_L2), .Z0_t (LED_128_Instance_SBox_Instance_15_Q2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_15_XOR4_U1 ( .A0_t (LED_128_Instance_addconst_out[63]), .B0_t (LED_128_Instance_addconst_out[60]), .Z0_t (LED_128_Instance_SBox_Instance_15_L3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_15_XOR5_U1 ( .A0_t (LED_128_Instance_SBox_Instance_15_L3), .B0_t (LED_128_Instance_SBox_Instance_15_L0), .Z0_t (LED_128_Instance_SBox_Instance_15_Q3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_15_XOR6_U1 ( .A0_t (LED_128_Instance_addconst_out[63]), .B0_t (LED_128_Instance_addconst_out[61]), .Z0_t (LED_128_Instance_SBox_Instance_15_L4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_15_XOR7_U1 ( .A0_t (LED_128_Instance_SBox_Instance_15_T0), .B0_t (LED_128_Instance_SBox_Instance_15_T2), .Z0_t (LED_128_Instance_SBox_Instance_15_L5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_SBox_Instance_15_XOR8_U1 ( .A0_t (LED_128_Instance_SBox_Instance_15_L4), .B0_t (LED_128_Instance_SBox_Instance_15_L5), .Z0_t (LED_128_Instance_SBox_Instance_15_Q6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_15_XOR9_U1 ( .A0_t (LED_128_Instance_SBox_Instance_15_L1), .B0_t (LED_128_Instance_addconst_out[62]), .Z0_t (LED_128_Instance_SBox_Instance_15_Q7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_15_AND1_U1 ( .A0_t (LED_128_Instance_SBox_Instance_15_L0), .B0_t (LED_128_Instance_addconst_out[63]), .Z0_t (LED_128_Instance_SBox_Instance_15_T0) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_15_AND2_U1 ( .A0_t (LED_128_Instance_SBox_Instance_15_Q2), .B0_t (LED_128_Instance_SBox_Instance_15_Q3), .Z0_t (LED_128_Instance_SBox_Instance_15_T1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_15_AND3_U1 ( .A0_t (LED_128_Instance_addconst_out[61]), .B0_t (LED_128_Instance_addconst_out[62]), .Z0_t (LED_128_Instance_SBox_Instance_15_T2) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_15_AND4_U1 ( .A0_t (LED_128_Instance_SBox_Instance_15_Q6), .B0_t (LED_128_Instance_SBox_Instance_15_Q7), .Z0_t (LED_128_Instance_SBox_Instance_15_T3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_15_XOR10_U1 ( .A0_t (LED_128_Instance_SBox_Instance_15_L5), .B0_t (LED_128_Instance_SBox_Instance_15_T3), .Z0_t (LED_128_Instance_SBox_Instance_15_L7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_15_XOR11_U1 ( .A0_t (LED_128_Instance_addconst_out[60]), .B0_t (LED_128_Instance_SBox_Instance_15_L7), .Z0_t (LED_128_Instance_subcells_out[63]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_15_XOR12_U1 ( .A0_t (LED_128_Instance_SBox_Instance_15_L5), .B0_t (LED_128_Instance_SBox_Instance_15_T1), .Z0_t (LED_128_Instance_SBox_Instance_15_L8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_15_XOR13_U1 ( .A0_t (LED_128_Instance_SBox_Instance_15_L1), .B0_t (LED_128_Instance_SBox_Instance_15_L8), .Z0_t (LED_128_Instance_subcells_out[62]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_15_XOR14_U1 ( .A0_t (LED_128_Instance_SBox_Instance_15_L4), .B0_t (LED_128_Instance_SBox_Instance_15_T3), .Z0_t (LED_128_Instance_subcells_out[61]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_15_XOR15_U1 ( .A0_t (LED_128_Instance_SBox_Instance_15_L3), .B0_t (LED_128_Instance_SBox_Instance_15_T2), .Z0_t (LED_128_Instance_subcells_out[60]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U58 ( .A0_t (LED_128_Instance_subcells_out[2]), .B0_t (LED_128_Instance_MCS_Instance_0_n42), .Z0_t (LED_128_Instance_mixcolumns_out[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U57 ( .A0_t (LED_128_Instance_MCS_Instance_0_n41), .B0_t (LED_128_Instance_subcells_out[62]), .Z0_t (LED_128_Instance_mixcolumns_out[19]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U56 ( .A0_t (LED_128_Instance_subcells_out[61]), .B0_t (LED_128_Instance_MCS_Instance_0_n40), .Z0_t (LED_128_Instance_mixcolumns_out[18]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U55 ( .A0_t (LED_128_Instance_MCS_Instance_0_n39), .B0_t (LED_128_Instance_MCS_Instance_0_n42), .Z0_t (LED_128_Instance_MCS_Instance_0_n40) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U54 ( .A0_t (LED_128_Instance_MCS_Instance_0_n38), .B0_t (LED_128_Instance_MCS_Instance_0_n37), .Z0_t (LED_128_Instance_MCS_Instance_0_n42) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U53 ( .A0_t (LED_128_Instance_MCS_Instance_0_n36), .B0_t (LED_128_Instance_MCS_Instance_0_n35), .Z0_t (LED_128_Instance_MCS_Instance_0_n39) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U52 ( .A0_t (LED_128_Instance_MCS_Instance_0_n34), .B0_t (LED_128_Instance_MCS_Instance_0_n36), .Z0_t (LED_128_Instance_mixcolumns_out[35]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U51 ( .A0_t (LED_128_Instance_MCS_Instance_0_n33), .B0_t (LED_128_Instance_MCS_Instance_0_n32), .Z0_t (LED_128_Instance_MCS_Instance_0_n34) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U50 ( .A0_t (LED_128_Instance_MCS_Instance_0_n31), .B0_t (LED_128_Instance_subcells_out[22]), .Z0_t (LED_128_Instance_MCS_Instance_0_n32) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U49 ( .A0_t (LED_128_Instance_MCS_Instance_0_n30), .B0_t (LED_128_Instance_MCS_Instance_0_n29), .Z0_t (LED_128_Instance_MCS_Instance_0_n33) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U48 ( .A0_t (LED_128_Instance_MCS_Instance_0_n28), .B0_t (LED_128_Instance_MCS_Instance_0_n27), .Z0_t (LED_128_Instance_mixcolumns_out[34]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U47 ( .A0_t (LED_128_Instance_MCS_Instance_0_n26), .B0_t (LED_128_Instance_MCS_Instance_0_n25), .Z0_t (LED_128_Instance_MCS_Instance_0_n28) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U46 ( .A0_t (LED_128_Instance_subcells_out[42]), .B0_t (LED_128_Instance_subcells_out[20]), .Z0_t (LED_128_Instance_MCS_Instance_0_n25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U45 ( .A0_t (LED_128_Instance_MCS_Instance_0_n24), .B0_t (LED_128_Instance_MCS_Instance_0_n23), .Z0_t (LED_128_Instance_mixcolumns_out[33]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U44 ( .A0_t (LED_128_Instance_MCS_Instance_0_n22), .B0_t (LED_128_Instance_MCS_Instance_0_n21), .Z0_t (LED_128_Instance_MCS_Instance_0_n24) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U43 ( .A0_t (LED_128_Instance_MCS_Instance_0_n38), .B0_t (LED_128_Instance_subcells_out[41]), .Z0_t (LED_128_Instance_MCS_Instance_0_n21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U42 ( .A0_t (LED_128_Instance_MCS_Instance_0_n29), .B0_t (LED_128_Instance_subcells_out[40]), .Z0_t (LED_128_Instance_MCS_Instance_0_n22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U41 ( .A0_t (LED_128_Instance_subcells_out[0]), .B0_t (LED_128_Instance_MCS_Instance_0_n35), .Z0_t (LED_128_Instance_MCS_Instance_0_n29) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U40 ( .A0_t (LED_128_Instance_MCS_Instance_0_n20), .B0_t (LED_128_Instance_MCS_Instance_0_n19), .Z0_t (LED_128_Instance_mixcolumns_out[32]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U39 ( .A0_t (LED_128_Instance_MCS_Instance_0_n41), .B0_t (LED_128_Instance_subcells_out[23]), .Z0_t (LED_128_Instance_MCS_Instance_0_n20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U38 ( .A0_t (LED_128_Instance_MCS_Instance_0_n18), .B0_t (LED_128_Instance_MCS_Instance_0_n27), .Z0_t (LED_128_Instance_MCS_Instance_0_n41) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U37 ( .A0_t (LED_128_Instance_MCS_Instance_0_n38), .B0_t (LED_128_Instance_MCS_Instance_0_n17), .Z0_t (LED_128_Instance_MCS_Instance_0_n27) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U36 ( .A0_t (LED_128_Instance_subcells_out[3]), .B0_t (LED_128_Instance_MCS_Instance_0_n31), .Z0_t (LED_128_Instance_MCS_Instance_0_n38) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U35 ( .A0_t (LED_128_Instance_subcells_out[43]), .B0_t (LED_128_Instance_subcells_out[21]), .Z0_t (LED_128_Instance_MCS_Instance_0_n31) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U34 ( .A0_t (LED_128_Instance_MCS_Instance_0_n16), .B0_t (LED_128_Instance_MCS_Instance_0_n30), .Z0_t (LED_128_Instance_mixcolumns_out[51]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U33 ( .A0_t (LED_128_Instance_MCS_Instance_0_n15), .B0_t (LED_128_Instance_subcells_out[2]), .Z0_t (LED_128_Instance_MCS_Instance_0_n16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U32 ( .A0_t (LED_128_Instance_subcells_out[23]), .B0_t (LED_128_Instance_MCS_Instance_0_n14), .Z0_t (LED_128_Instance_mixcolumns_out[49]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U31 ( .A0_t (LED_128_Instance_MCS_Instance_0_n13), .B0_t (LED_128_Instance_MCS_Instance_0_n12), .Z0_t (LED_128_Instance_MCS_Instance_0_n14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U30 ( .A0_t (LED_128_Instance_subcells_out[0]), .B0_t (LED_128_Instance_subcells_out[62]), .Z0_t (LED_128_Instance_MCS_Instance_0_n12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U29 ( .A0_t (LED_128_Instance_MCS_Instance_0_n11), .B0_t (LED_128_Instance_subcells_out[20]), .Z0_t (LED_128_Instance_MCS_Instance_0_n13) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U28 ( .A0_t (LED_128_Instance_subcells_out[43]), .B0_t (LED_128_Instance_MCS_Instance_0_n10), .Z0_t (LED_128_Instance_mixcolumns_out[48]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U27 ( .A0_t (LED_128_Instance_MCS_Instance_0_n9), .B0_t (LED_128_Instance_MCS_Instance_0_n36), .Z0_t (LED_128_Instance_MCS_Instance_0_n10) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U26 ( .A0_t (LED_128_Instance_MCS_Instance_0_n11), .B0_t (LED_128_Instance_MCS_Instance_0_n8), .Z0_t (LED_128_Instance_MCS_Instance_0_n9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U25 ( .A0_t (LED_128_Instance_subcells_out[3]), .B0_t (LED_128_Instance_MCS_Instance_0_n37), .Z0_t (LED_128_Instance_MCS_Instance_0_n11) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U24 ( .A0_t (LED_128_Instance_subcells_out[63]), .B0_t (LED_128_Instance_MCS_Instance_0_n30), .Z0_t (LED_128_Instance_MCS_Instance_0_n37) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U23 ( .A0_t (LED_128_Instance_subcells_out[60]), .B0_t (LED_128_Instance_subcells_out[40]), .Z0_t (LED_128_Instance_MCS_Instance_0_n30) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U22 ( .A0_t (LED_128_Instance_MCS_Instance_0_n7), .B0_t (LED_128_Instance_MCS_Instance_0_n17), .Z0_t (LED_128_Instance_mixcolumns_out[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U21 ( .A0_t (LED_128_Instance_MCS_Instance_0_n18), .B0_t (LED_128_Instance_subcells_out[3]), .Z0_t (LED_128_Instance_MCS_Instance_0_n7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U20 ( .A0_t (LED_128_Instance_subcells_out[0]), .B0_t (LED_128_Instance_subcells_out[61]), .Z0_t (LED_128_Instance_MCS_Instance_0_n18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U19 ( .A0_t (LED_128_Instance_MCS_Instance_0_n6), .B0_t (LED_128_Instance_MCS_Instance_0_n5), .Z0_t (LED_128_Instance_mixcolumns_out[17]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U18 ( .A0_t (LED_128_Instance_MCS_Instance_0_n19), .B0_t (LED_128_Instance_MCS_Instance_0_n15), .Z0_t (LED_128_Instance_MCS_Instance_0_n6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U17 ( .A0_t (LED_128_Instance_MCS_Instance_0_n17), .B0_t (LED_128_Instance_MCS_Instance_0_n23), .Z0_t (LED_128_Instance_MCS_Instance_0_n15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U16 ( .A0_t (LED_128_Instance_subcells_out[62]), .B0_t (LED_128_Instance_subcells_out[42]), .Z0_t (LED_128_Instance_MCS_Instance_0_n23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U15 ( .A0_t (LED_128_Instance_subcells_out[41]), .B0_t (LED_128_Instance_subcells_out[22]), .Z0_t (LED_128_Instance_MCS_Instance_0_n17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U14 ( .A0_t (LED_128_Instance_subcells_out[60]), .B0_t (LED_128_Instance_subcells_out[1]), .Z0_t (LED_128_Instance_MCS_Instance_0_n19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U13 ( .A0_t (LED_128_Instance_subcells_out[1]), .B0_t (LED_128_Instance_MCS_Instance_0_n4), .Z0_t (LED_128_Instance_mixcolumns_out[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U12 ( .A0_t (LED_128_Instance_MCS_Instance_0_n3), .B0_t (LED_128_Instance_MCS_Instance_0_n2), .Z0_t (LED_128_Instance_mixcolumns_out[16]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U11 ( .A0_t (LED_128_Instance_subcells_out[22]), .B0_t (LED_128_Instance_MCS_Instance_0_n4), .Z0_t (LED_128_Instance_MCS_Instance_0_n3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U10 ( .A0_t (LED_128_Instance_subcells_out[62]), .B0_t (LED_128_Instance_MCS_Instance_0_n36), .Z0_t (LED_128_Instance_MCS_Instance_0_n4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U9 ( .A0_t (LED_128_Instance_subcells_out[23]), .B0_t (LED_128_Instance_subcells_out[42]), .Z0_t (LED_128_Instance_MCS_Instance_0_n36) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U8 ( .A0_t (LED_128_Instance_subcells_out[63]), .B0_t (LED_128_Instance_MCS_Instance_0_n5), .Z0_t (LED_128_Instance_mixcolumns_out[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U7 ( .A0_t (LED_128_Instance_subcells_out[43]), .B0_t (LED_128_Instance_MCS_Instance_0_n35), .Z0_t (LED_128_Instance_MCS_Instance_0_n5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U6 ( .A0_t (LED_128_Instance_subcells_out[2]), .B0_t (LED_128_Instance_subcells_out[20]), .Z0_t (LED_128_Instance_MCS_Instance_0_n35) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U5 ( .A0_t (LED_128_Instance_MCS_Instance_0_n1), .B0_t (LED_128_Instance_MCS_Instance_0_n8), .Z0_t (LED_128_Instance_mixcolumns_out[50]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U4 ( .A0_t (LED_128_Instance_subcells_out[61]), .B0_t (LED_128_Instance_subcells_out[41]), .Z0_t (LED_128_Instance_MCS_Instance_0_n8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U3 ( .A0_t (LED_128_Instance_subcells_out[21]), .B0_t (LED_128_Instance_MCS_Instance_0_n2), .Z0_t (LED_128_Instance_MCS_Instance_0_n1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U2 ( .A0_t (LED_128_Instance_subcells_out[40]), .B0_t (LED_128_Instance_MCS_Instance_0_n26), .Z0_t (LED_128_Instance_MCS_Instance_0_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U1 ( .A0_t (LED_128_Instance_subcells_out[1]), .B0_t (LED_128_Instance_subcells_out[63]), .Z0_t (LED_128_Instance_MCS_Instance_0_n26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U58 ( .A0_t (LED_128_Instance_subcells_out[6]), .B0_t (LED_128_Instance_MCS_Instance_1_n42), .Z0_t (LED_128_Instance_mixcolumns_out[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U57 ( .A0_t (LED_128_Instance_MCS_Instance_1_n41), .B0_t (LED_128_Instance_subcells_out[50]), .Z0_t (LED_128_Instance_mixcolumns_out[23]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U56 ( .A0_t (LED_128_Instance_subcells_out[49]), .B0_t (LED_128_Instance_MCS_Instance_1_n40), .Z0_t (LED_128_Instance_mixcolumns_out[22]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U55 ( .A0_t (LED_128_Instance_MCS_Instance_1_n39), .B0_t (LED_128_Instance_MCS_Instance_1_n42), .Z0_t (LED_128_Instance_MCS_Instance_1_n40) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U54 ( .A0_t (LED_128_Instance_MCS_Instance_1_n38), .B0_t (LED_128_Instance_MCS_Instance_1_n37), .Z0_t (LED_128_Instance_MCS_Instance_1_n42) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U53 ( .A0_t (LED_128_Instance_MCS_Instance_1_n36), .B0_t (LED_128_Instance_MCS_Instance_1_n35), .Z0_t (LED_128_Instance_MCS_Instance_1_n39) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U52 ( .A0_t (LED_128_Instance_MCS_Instance_1_n34), .B0_t (LED_128_Instance_MCS_Instance_1_n36), .Z0_t (LED_128_Instance_mixcolumns_out[39]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U51 ( .A0_t (LED_128_Instance_MCS_Instance_1_n33), .B0_t (LED_128_Instance_MCS_Instance_1_n32), .Z0_t (LED_128_Instance_MCS_Instance_1_n34) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U50 ( .A0_t (LED_128_Instance_MCS_Instance_1_n31), .B0_t (LED_128_Instance_subcells_out[26]), .Z0_t (LED_128_Instance_MCS_Instance_1_n32) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U49 ( .A0_t (LED_128_Instance_MCS_Instance_1_n30), .B0_t (LED_128_Instance_MCS_Instance_1_n29), .Z0_t (LED_128_Instance_MCS_Instance_1_n33) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U48 ( .A0_t (LED_128_Instance_MCS_Instance_1_n28), .B0_t (LED_128_Instance_MCS_Instance_1_n27), .Z0_t (LED_128_Instance_mixcolumns_out[38]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U47 ( .A0_t (LED_128_Instance_MCS_Instance_1_n26), .B0_t (LED_128_Instance_MCS_Instance_1_n25), .Z0_t (LED_128_Instance_MCS_Instance_1_n28) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U46 ( .A0_t (LED_128_Instance_subcells_out[46]), .B0_t (LED_128_Instance_subcells_out[24]), .Z0_t (LED_128_Instance_MCS_Instance_1_n25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U45 ( .A0_t (LED_128_Instance_MCS_Instance_1_n24), .B0_t (LED_128_Instance_MCS_Instance_1_n23), .Z0_t (LED_128_Instance_mixcolumns_out[37]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U44 ( .A0_t (LED_128_Instance_MCS_Instance_1_n22), .B0_t (LED_128_Instance_MCS_Instance_1_n21), .Z0_t (LED_128_Instance_MCS_Instance_1_n24) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U43 ( .A0_t (LED_128_Instance_MCS_Instance_1_n38), .B0_t (LED_128_Instance_subcells_out[45]), .Z0_t (LED_128_Instance_MCS_Instance_1_n21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U42 ( .A0_t (LED_128_Instance_MCS_Instance_1_n29), .B0_t (LED_128_Instance_subcells_out[44]), .Z0_t (LED_128_Instance_MCS_Instance_1_n22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U41 ( .A0_t (LED_128_Instance_subcells_out[4]), .B0_t (LED_128_Instance_MCS_Instance_1_n35), .Z0_t (LED_128_Instance_MCS_Instance_1_n29) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U40 ( .A0_t (LED_128_Instance_MCS_Instance_1_n20), .B0_t (LED_128_Instance_MCS_Instance_1_n19), .Z0_t (LED_128_Instance_mixcolumns_out[36]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U39 ( .A0_t (LED_128_Instance_MCS_Instance_1_n41), .B0_t (LED_128_Instance_subcells_out[27]), .Z0_t (LED_128_Instance_MCS_Instance_1_n20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U38 ( .A0_t (LED_128_Instance_MCS_Instance_1_n18), .B0_t (LED_128_Instance_MCS_Instance_1_n27), .Z0_t (LED_128_Instance_MCS_Instance_1_n41) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U37 ( .A0_t (LED_128_Instance_MCS_Instance_1_n38), .B0_t (LED_128_Instance_MCS_Instance_1_n17), .Z0_t (LED_128_Instance_MCS_Instance_1_n27) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U36 ( .A0_t (LED_128_Instance_subcells_out[7]), .B0_t (LED_128_Instance_MCS_Instance_1_n31), .Z0_t (LED_128_Instance_MCS_Instance_1_n38) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U35 ( .A0_t (LED_128_Instance_subcells_out[47]), .B0_t (LED_128_Instance_subcells_out[25]), .Z0_t (LED_128_Instance_MCS_Instance_1_n31) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U34 ( .A0_t (LED_128_Instance_MCS_Instance_1_n16), .B0_t (LED_128_Instance_MCS_Instance_1_n30), .Z0_t (LED_128_Instance_mixcolumns_out[55]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U33 ( .A0_t (LED_128_Instance_MCS_Instance_1_n15), .B0_t (LED_128_Instance_subcells_out[6]), .Z0_t (LED_128_Instance_MCS_Instance_1_n16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U32 ( .A0_t (LED_128_Instance_subcells_out[27]), .B0_t (LED_128_Instance_MCS_Instance_1_n14), .Z0_t (LED_128_Instance_mixcolumns_out[53]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U31 ( .A0_t (LED_128_Instance_MCS_Instance_1_n13), .B0_t (LED_128_Instance_MCS_Instance_1_n12), .Z0_t (LED_128_Instance_MCS_Instance_1_n14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U30 ( .A0_t (LED_128_Instance_subcells_out[4]), .B0_t (LED_128_Instance_subcells_out[50]), .Z0_t (LED_128_Instance_MCS_Instance_1_n12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U29 ( .A0_t (LED_128_Instance_MCS_Instance_1_n11), .B0_t (LED_128_Instance_subcells_out[24]), .Z0_t (LED_128_Instance_MCS_Instance_1_n13) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U28 ( .A0_t (LED_128_Instance_subcells_out[47]), .B0_t (LED_128_Instance_MCS_Instance_1_n10), .Z0_t (LED_128_Instance_mixcolumns_out[52]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U27 ( .A0_t (LED_128_Instance_MCS_Instance_1_n9), .B0_t (LED_128_Instance_MCS_Instance_1_n36), .Z0_t (LED_128_Instance_MCS_Instance_1_n10) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U26 ( .A0_t (LED_128_Instance_MCS_Instance_1_n11), .B0_t (LED_128_Instance_MCS_Instance_1_n8), .Z0_t (LED_128_Instance_MCS_Instance_1_n9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U25 ( .A0_t (LED_128_Instance_subcells_out[7]), .B0_t (LED_128_Instance_MCS_Instance_1_n37), .Z0_t (LED_128_Instance_MCS_Instance_1_n11) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U24 ( .A0_t (LED_128_Instance_subcells_out[51]), .B0_t (LED_128_Instance_MCS_Instance_1_n30), .Z0_t (LED_128_Instance_MCS_Instance_1_n37) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U23 ( .A0_t (LED_128_Instance_subcells_out[48]), .B0_t (LED_128_Instance_subcells_out[44]), .Z0_t (LED_128_Instance_MCS_Instance_1_n30) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U22 ( .A0_t (LED_128_Instance_MCS_Instance_1_n7), .B0_t (LED_128_Instance_MCS_Instance_1_n17), .Z0_t (LED_128_Instance_mixcolumns_out[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U21 ( .A0_t (LED_128_Instance_MCS_Instance_1_n18), .B0_t (LED_128_Instance_subcells_out[7]), .Z0_t (LED_128_Instance_MCS_Instance_1_n7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U20 ( .A0_t (LED_128_Instance_subcells_out[4]), .B0_t (LED_128_Instance_subcells_out[49]), .Z0_t (LED_128_Instance_MCS_Instance_1_n18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U19 ( .A0_t (LED_128_Instance_MCS_Instance_1_n6), .B0_t (LED_128_Instance_MCS_Instance_1_n5), .Z0_t (LED_128_Instance_mixcolumns_out[21]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U18 ( .A0_t (LED_128_Instance_MCS_Instance_1_n19), .B0_t (LED_128_Instance_MCS_Instance_1_n15), .Z0_t (LED_128_Instance_MCS_Instance_1_n6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U17 ( .A0_t (LED_128_Instance_MCS_Instance_1_n17), .B0_t (LED_128_Instance_MCS_Instance_1_n23), .Z0_t (LED_128_Instance_MCS_Instance_1_n15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U16 ( .A0_t (LED_128_Instance_subcells_out[50]), .B0_t (LED_128_Instance_subcells_out[46]), .Z0_t (LED_128_Instance_MCS_Instance_1_n23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U15 ( .A0_t (LED_128_Instance_subcells_out[45]), .B0_t (LED_128_Instance_subcells_out[26]), .Z0_t (LED_128_Instance_MCS_Instance_1_n17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U14 ( .A0_t (LED_128_Instance_subcells_out[48]), .B0_t (LED_128_Instance_subcells_out[5]), .Z0_t (LED_128_Instance_MCS_Instance_1_n19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U13 ( .A0_t (LED_128_Instance_subcells_out[5]), .B0_t (LED_128_Instance_MCS_Instance_1_n4), .Z0_t (LED_128_Instance_mixcolumns_out[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U12 ( .A0_t (LED_128_Instance_MCS_Instance_1_n3), .B0_t (LED_128_Instance_MCS_Instance_1_n2), .Z0_t (LED_128_Instance_mixcolumns_out[20]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U11 ( .A0_t (LED_128_Instance_subcells_out[26]), .B0_t (LED_128_Instance_MCS_Instance_1_n4), .Z0_t (LED_128_Instance_MCS_Instance_1_n3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U10 ( .A0_t (LED_128_Instance_subcells_out[50]), .B0_t (LED_128_Instance_MCS_Instance_1_n36), .Z0_t (LED_128_Instance_MCS_Instance_1_n4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U9 ( .A0_t (LED_128_Instance_subcells_out[27]), .B0_t (LED_128_Instance_subcells_out[46]), .Z0_t (LED_128_Instance_MCS_Instance_1_n36) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U8 ( .A0_t (LED_128_Instance_subcells_out[51]), .B0_t (LED_128_Instance_MCS_Instance_1_n5), .Z0_t (LED_128_Instance_mixcolumns_out[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U7 ( .A0_t (LED_128_Instance_subcells_out[47]), .B0_t (LED_128_Instance_MCS_Instance_1_n35), .Z0_t (LED_128_Instance_MCS_Instance_1_n5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U6 ( .A0_t (LED_128_Instance_subcells_out[6]), .B0_t (LED_128_Instance_subcells_out[24]), .Z0_t (LED_128_Instance_MCS_Instance_1_n35) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U5 ( .A0_t (LED_128_Instance_MCS_Instance_1_n1), .B0_t (LED_128_Instance_MCS_Instance_1_n8), .Z0_t (LED_128_Instance_mixcolumns_out[54]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U4 ( .A0_t (LED_128_Instance_subcells_out[49]), .B0_t (LED_128_Instance_subcells_out[45]), .Z0_t (LED_128_Instance_MCS_Instance_1_n8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U3 ( .A0_t (LED_128_Instance_subcells_out[25]), .B0_t (LED_128_Instance_MCS_Instance_1_n2), .Z0_t (LED_128_Instance_MCS_Instance_1_n1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U2 ( .A0_t (LED_128_Instance_subcells_out[44]), .B0_t (LED_128_Instance_MCS_Instance_1_n26), .Z0_t (LED_128_Instance_MCS_Instance_1_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U1 ( .A0_t (LED_128_Instance_subcells_out[5]), .B0_t (LED_128_Instance_subcells_out[51]), .Z0_t (LED_128_Instance_MCS_Instance_1_n26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U58 ( .A0_t (LED_128_Instance_subcells_out[10]), .B0_t (LED_128_Instance_MCS_Instance_2_n42), .Z0_t (LED_128_Instance_mixcolumns_out[9]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U57 ( .A0_t (LED_128_Instance_MCS_Instance_2_n41), .B0_t (LED_128_Instance_subcells_out[54]), .Z0_t (LED_128_Instance_mixcolumns_out[27]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U56 ( .A0_t (LED_128_Instance_subcells_out[53]), .B0_t (LED_128_Instance_MCS_Instance_2_n40), .Z0_t (LED_128_Instance_mixcolumns_out[26]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U55 ( .A0_t (LED_128_Instance_MCS_Instance_2_n39), .B0_t (LED_128_Instance_MCS_Instance_2_n42), .Z0_t (LED_128_Instance_MCS_Instance_2_n40) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U54 ( .A0_t (LED_128_Instance_MCS_Instance_2_n38), .B0_t (LED_128_Instance_MCS_Instance_2_n37), .Z0_t (LED_128_Instance_MCS_Instance_2_n42) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U53 ( .A0_t (LED_128_Instance_MCS_Instance_2_n36), .B0_t (LED_128_Instance_MCS_Instance_2_n35), .Z0_t (LED_128_Instance_MCS_Instance_2_n39) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U52 ( .A0_t (LED_128_Instance_MCS_Instance_2_n34), .B0_t (LED_128_Instance_MCS_Instance_2_n36), .Z0_t (LED_128_Instance_mixcolumns_out[43]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U51 ( .A0_t (LED_128_Instance_MCS_Instance_2_n33), .B0_t (LED_128_Instance_MCS_Instance_2_n32), .Z0_t (LED_128_Instance_MCS_Instance_2_n34) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U50 ( .A0_t (LED_128_Instance_MCS_Instance_2_n31), .B0_t (LED_128_Instance_subcells_out[30]), .Z0_t (LED_128_Instance_MCS_Instance_2_n32) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U49 ( .A0_t (LED_128_Instance_MCS_Instance_2_n30), .B0_t (LED_128_Instance_MCS_Instance_2_n29), .Z0_t (LED_128_Instance_MCS_Instance_2_n33) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U48 ( .A0_t (LED_128_Instance_MCS_Instance_2_n28), .B0_t (LED_128_Instance_MCS_Instance_2_n27), .Z0_t (LED_128_Instance_mixcolumns_out[42]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U47 ( .A0_t (LED_128_Instance_MCS_Instance_2_n26), .B0_t (LED_128_Instance_MCS_Instance_2_n25), .Z0_t (LED_128_Instance_MCS_Instance_2_n28) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U46 ( .A0_t (LED_128_Instance_subcells_out[34]), .B0_t (LED_128_Instance_subcells_out[28]), .Z0_t (LED_128_Instance_MCS_Instance_2_n25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U45 ( .A0_t (LED_128_Instance_MCS_Instance_2_n24), .B0_t (LED_128_Instance_MCS_Instance_2_n23), .Z0_t (LED_128_Instance_mixcolumns_out[41]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U44 ( .A0_t (LED_128_Instance_MCS_Instance_2_n22), .B0_t (LED_128_Instance_MCS_Instance_2_n21), .Z0_t (LED_128_Instance_MCS_Instance_2_n24) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U43 ( .A0_t (LED_128_Instance_MCS_Instance_2_n38), .B0_t (LED_128_Instance_subcells_out[33]), .Z0_t (LED_128_Instance_MCS_Instance_2_n21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U42 ( .A0_t (LED_128_Instance_MCS_Instance_2_n29), .B0_t (LED_128_Instance_subcells_out[32]), .Z0_t (LED_128_Instance_MCS_Instance_2_n22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U41 ( .A0_t (LED_128_Instance_subcells_out[8]), .B0_t (LED_128_Instance_MCS_Instance_2_n35), .Z0_t (LED_128_Instance_MCS_Instance_2_n29) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U40 ( .A0_t (LED_128_Instance_MCS_Instance_2_n20), .B0_t (LED_128_Instance_MCS_Instance_2_n19), .Z0_t (LED_128_Instance_mixcolumns_out[40]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U39 ( .A0_t (LED_128_Instance_MCS_Instance_2_n41), .B0_t (LED_128_Instance_subcells_out[31]), .Z0_t (LED_128_Instance_MCS_Instance_2_n20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U38 ( .A0_t (LED_128_Instance_MCS_Instance_2_n18), .B0_t (LED_128_Instance_MCS_Instance_2_n27), .Z0_t (LED_128_Instance_MCS_Instance_2_n41) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U37 ( .A0_t (LED_128_Instance_MCS_Instance_2_n38), .B0_t (LED_128_Instance_MCS_Instance_2_n17), .Z0_t (LED_128_Instance_MCS_Instance_2_n27) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U36 ( .A0_t (LED_128_Instance_subcells_out[11]), .B0_t (LED_128_Instance_MCS_Instance_2_n31), .Z0_t (LED_128_Instance_MCS_Instance_2_n38) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U35 ( .A0_t (LED_128_Instance_subcells_out[35]), .B0_t (LED_128_Instance_subcells_out[29]), .Z0_t (LED_128_Instance_MCS_Instance_2_n31) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U34 ( .A0_t (LED_128_Instance_MCS_Instance_2_n16), .B0_t (LED_128_Instance_MCS_Instance_2_n30), .Z0_t (LED_128_Instance_mixcolumns_out[59]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U33 ( .A0_t (LED_128_Instance_MCS_Instance_2_n15), .B0_t (LED_128_Instance_subcells_out[10]), .Z0_t (LED_128_Instance_MCS_Instance_2_n16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U32 ( .A0_t (LED_128_Instance_subcells_out[31]), .B0_t (LED_128_Instance_MCS_Instance_2_n14), .Z0_t (LED_128_Instance_mixcolumns_out[57]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U31 ( .A0_t (LED_128_Instance_MCS_Instance_2_n13), .B0_t (LED_128_Instance_MCS_Instance_2_n12), .Z0_t (LED_128_Instance_MCS_Instance_2_n14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U30 ( .A0_t (LED_128_Instance_subcells_out[8]), .B0_t (LED_128_Instance_subcells_out[54]), .Z0_t (LED_128_Instance_MCS_Instance_2_n12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U29 ( .A0_t (LED_128_Instance_MCS_Instance_2_n11), .B0_t (LED_128_Instance_subcells_out[28]), .Z0_t (LED_128_Instance_MCS_Instance_2_n13) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U28 ( .A0_t (LED_128_Instance_subcells_out[35]), .B0_t (LED_128_Instance_MCS_Instance_2_n10), .Z0_t (LED_128_Instance_mixcolumns_out[56]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U27 ( .A0_t (LED_128_Instance_MCS_Instance_2_n9), .B0_t (LED_128_Instance_MCS_Instance_2_n36), .Z0_t (LED_128_Instance_MCS_Instance_2_n10) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U26 ( .A0_t (LED_128_Instance_MCS_Instance_2_n11), .B0_t (LED_128_Instance_MCS_Instance_2_n8), .Z0_t (LED_128_Instance_MCS_Instance_2_n9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U25 ( .A0_t (LED_128_Instance_subcells_out[11]), .B0_t (LED_128_Instance_MCS_Instance_2_n37), .Z0_t (LED_128_Instance_MCS_Instance_2_n11) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U24 ( .A0_t (LED_128_Instance_subcells_out[55]), .B0_t (LED_128_Instance_MCS_Instance_2_n30), .Z0_t (LED_128_Instance_MCS_Instance_2_n37) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U23 ( .A0_t (LED_128_Instance_subcells_out[52]), .B0_t (LED_128_Instance_subcells_out[32]), .Z0_t (LED_128_Instance_MCS_Instance_2_n30) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U22 ( .A0_t (LED_128_Instance_MCS_Instance_2_n7), .B0_t (LED_128_Instance_MCS_Instance_2_n17), .Z0_t (LED_128_Instance_mixcolumns_out[10]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U21 ( .A0_t (LED_128_Instance_MCS_Instance_2_n18), .B0_t (LED_128_Instance_subcells_out[11]), .Z0_t (LED_128_Instance_MCS_Instance_2_n7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U20 ( .A0_t (LED_128_Instance_subcells_out[8]), .B0_t (LED_128_Instance_subcells_out[53]), .Z0_t (LED_128_Instance_MCS_Instance_2_n18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U19 ( .A0_t (LED_128_Instance_MCS_Instance_2_n6), .B0_t (LED_128_Instance_MCS_Instance_2_n5), .Z0_t (LED_128_Instance_mixcolumns_out[25]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U18 ( .A0_t (LED_128_Instance_MCS_Instance_2_n19), .B0_t (LED_128_Instance_MCS_Instance_2_n15), .Z0_t (LED_128_Instance_MCS_Instance_2_n6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U17 ( .A0_t (LED_128_Instance_MCS_Instance_2_n17), .B0_t (LED_128_Instance_MCS_Instance_2_n23), .Z0_t (LED_128_Instance_MCS_Instance_2_n15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U16 ( .A0_t (LED_128_Instance_subcells_out[54]), .B0_t (LED_128_Instance_subcells_out[34]), .Z0_t (LED_128_Instance_MCS_Instance_2_n23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U15 ( .A0_t (LED_128_Instance_subcells_out[33]), .B0_t (LED_128_Instance_subcells_out[30]), .Z0_t (LED_128_Instance_MCS_Instance_2_n17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U14 ( .A0_t (LED_128_Instance_subcells_out[52]), .B0_t (LED_128_Instance_subcells_out[9]), .Z0_t (LED_128_Instance_MCS_Instance_2_n19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U13 ( .A0_t (LED_128_Instance_subcells_out[9]), .B0_t (LED_128_Instance_MCS_Instance_2_n4), .Z0_t (LED_128_Instance_mixcolumns_out[11]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U12 ( .A0_t (LED_128_Instance_MCS_Instance_2_n3), .B0_t (LED_128_Instance_MCS_Instance_2_n2), .Z0_t (LED_128_Instance_mixcolumns_out[24]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U11 ( .A0_t (LED_128_Instance_subcells_out[30]), .B0_t (LED_128_Instance_MCS_Instance_2_n4), .Z0_t (LED_128_Instance_MCS_Instance_2_n3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U10 ( .A0_t (LED_128_Instance_subcells_out[54]), .B0_t (LED_128_Instance_MCS_Instance_2_n36), .Z0_t (LED_128_Instance_MCS_Instance_2_n4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U9 ( .A0_t (LED_128_Instance_subcells_out[31]), .B0_t (LED_128_Instance_subcells_out[34]), .Z0_t (LED_128_Instance_MCS_Instance_2_n36) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U8 ( .A0_t (LED_128_Instance_subcells_out[55]), .B0_t (LED_128_Instance_MCS_Instance_2_n5), .Z0_t (LED_128_Instance_mixcolumns_out[8]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U7 ( .A0_t (LED_128_Instance_subcells_out[35]), .B0_t (LED_128_Instance_MCS_Instance_2_n35), .Z0_t (LED_128_Instance_MCS_Instance_2_n5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U6 ( .A0_t (LED_128_Instance_subcells_out[10]), .B0_t (LED_128_Instance_subcells_out[28]), .Z0_t (LED_128_Instance_MCS_Instance_2_n35) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U5 ( .A0_t (LED_128_Instance_MCS_Instance_2_n1), .B0_t (LED_128_Instance_MCS_Instance_2_n8), .Z0_t (LED_128_Instance_mixcolumns_out[58]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U4 ( .A0_t (LED_128_Instance_subcells_out[53]), .B0_t (LED_128_Instance_subcells_out[33]), .Z0_t (LED_128_Instance_MCS_Instance_2_n8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U3 ( .A0_t (LED_128_Instance_subcells_out[29]), .B0_t (LED_128_Instance_MCS_Instance_2_n2), .Z0_t (LED_128_Instance_MCS_Instance_2_n1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U2 ( .A0_t (LED_128_Instance_subcells_out[32]), .B0_t (LED_128_Instance_MCS_Instance_2_n26), .Z0_t (LED_128_Instance_MCS_Instance_2_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U1 ( .A0_t (LED_128_Instance_subcells_out[9]), .B0_t (LED_128_Instance_subcells_out[55]), .Z0_t (LED_128_Instance_MCS_Instance_2_n26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U58 ( .A0_t (LED_128_Instance_subcells_out[14]), .B0_t (LED_128_Instance_MCS_Instance_3_n42), .Z0_t (LED_128_Instance_mixcolumns_out[13]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U57 ( .A0_t (LED_128_Instance_MCS_Instance_3_n41), .B0_t (LED_128_Instance_subcells_out[58]), .Z0_t (LED_128_Instance_mixcolumns_out[31]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U56 ( .A0_t (LED_128_Instance_subcells_out[57]), .B0_t (LED_128_Instance_MCS_Instance_3_n40), .Z0_t (LED_128_Instance_mixcolumns_out[30]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U55 ( .A0_t (LED_128_Instance_MCS_Instance_3_n39), .B0_t (LED_128_Instance_MCS_Instance_3_n42), .Z0_t (LED_128_Instance_MCS_Instance_3_n40) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U54 ( .A0_t (LED_128_Instance_MCS_Instance_3_n38), .B0_t (LED_128_Instance_MCS_Instance_3_n37), .Z0_t (LED_128_Instance_MCS_Instance_3_n42) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U53 ( .A0_t (LED_128_Instance_MCS_Instance_3_n36), .B0_t (LED_128_Instance_MCS_Instance_3_n35), .Z0_t (LED_128_Instance_MCS_Instance_3_n39) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U52 ( .A0_t (LED_128_Instance_MCS_Instance_3_n34), .B0_t (LED_128_Instance_MCS_Instance_3_n36), .Z0_t (LED_128_Instance_mixcolumns_out[47]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U51 ( .A0_t (LED_128_Instance_MCS_Instance_3_n33), .B0_t (LED_128_Instance_MCS_Instance_3_n32), .Z0_t (LED_128_Instance_MCS_Instance_3_n34) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U50 ( .A0_t (LED_128_Instance_MCS_Instance_3_n31), .B0_t (LED_128_Instance_subcells_out[18]), .Z0_t (LED_128_Instance_MCS_Instance_3_n32) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U49 ( .A0_t (LED_128_Instance_MCS_Instance_3_n30), .B0_t (LED_128_Instance_MCS_Instance_3_n29), .Z0_t (LED_128_Instance_MCS_Instance_3_n33) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U48 ( .A0_t (LED_128_Instance_MCS_Instance_3_n28), .B0_t (LED_128_Instance_MCS_Instance_3_n27), .Z0_t (LED_128_Instance_mixcolumns_out[46]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U47 ( .A0_t (LED_128_Instance_MCS_Instance_3_n26), .B0_t (LED_128_Instance_MCS_Instance_3_n25), .Z0_t (LED_128_Instance_MCS_Instance_3_n28) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U46 ( .A0_t (LED_128_Instance_subcells_out[38]), .B0_t (LED_128_Instance_subcells_out[16]), .Z0_t (LED_128_Instance_MCS_Instance_3_n25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U45 ( .A0_t (LED_128_Instance_MCS_Instance_3_n24), .B0_t (LED_128_Instance_MCS_Instance_3_n23), .Z0_t (LED_128_Instance_mixcolumns_out[45]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U44 ( .A0_t (LED_128_Instance_MCS_Instance_3_n22), .B0_t (LED_128_Instance_MCS_Instance_3_n21), .Z0_t (LED_128_Instance_MCS_Instance_3_n24) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U43 ( .A0_t (LED_128_Instance_MCS_Instance_3_n38), .B0_t (LED_128_Instance_subcells_out[37]), .Z0_t (LED_128_Instance_MCS_Instance_3_n21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U42 ( .A0_t (LED_128_Instance_MCS_Instance_3_n29), .B0_t (LED_128_Instance_subcells_out[36]), .Z0_t (LED_128_Instance_MCS_Instance_3_n22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U41 ( .A0_t (LED_128_Instance_subcells_out[12]), .B0_t (LED_128_Instance_MCS_Instance_3_n35), .Z0_t (LED_128_Instance_MCS_Instance_3_n29) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U40 ( .A0_t (LED_128_Instance_MCS_Instance_3_n20), .B0_t (LED_128_Instance_MCS_Instance_3_n19), .Z0_t (LED_128_Instance_mixcolumns_out[44]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U39 ( .A0_t (LED_128_Instance_MCS_Instance_3_n41), .B0_t (LED_128_Instance_subcells_out[19]), .Z0_t (LED_128_Instance_MCS_Instance_3_n20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U38 ( .A0_t (LED_128_Instance_MCS_Instance_3_n18), .B0_t (LED_128_Instance_MCS_Instance_3_n27), .Z0_t (LED_128_Instance_MCS_Instance_3_n41) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U37 ( .A0_t (LED_128_Instance_MCS_Instance_3_n38), .B0_t (LED_128_Instance_MCS_Instance_3_n17), .Z0_t (LED_128_Instance_MCS_Instance_3_n27) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U36 ( .A0_t (LED_128_Instance_subcells_out[15]), .B0_t (LED_128_Instance_MCS_Instance_3_n31), .Z0_t (LED_128_Instance_MCS_Instance_3_n38) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U35 ( .A0_t (LED_128_Instance_subcells_out[39]), .B0_t (LED_128_Instance_subcells_out[17]), .Z0_t (LED_128_Instance_MCS_Instance_3_n31) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U34 ( .A0_t (LED_128_Instance_MCS_Instance_3_n16), .B0_t (LED_128_Instance_MCS_Instance_3_n30), .Z0_t (LED_128_Instance_mixcolumns_out[63]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U33 ( .A0_t (LED_128_Instance_MCS_Instance_3_n15), .B0_t (LED_128_Instance_subcells_out[14]), .Z0_t (LED_128_Instance_MCS_Instance_3_n16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U32 ( .A0_t (LED_128_Instance_subcells_out[19]), .B0_t (LED_128_Instance_MCS_Instance_3_n14), .Z0_t (LED_128_Instance_mixcolumns_out[61]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U31 ( .A0_t (LED_128_Instance_MCS_Instance_3_n13), .B0_t (LED_128_Instance_MCS_Instance_3_n12), .Z0_t (LED_128_Instance_MCS_Instance_3_n14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U30 ( .A0_t (LED_128_Instance_subcells_out[12]), .B0_t (LED_128_Instance_subcells_out[58]), .Z0_t (LED_128_Instance_MCS_Instance_3_n12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U29 ( .A0_t (LED_128_Instance_MCS_Instance_3_n11), .B0_t (LED_128_Instance_subcells_out[16]), .Z0_t (LED_128_Instance_MCS_Instance_3_n13) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U28 ( .A0_t (LED_128_Instance_subcells_out[39]), .B0_t (LED_128_Instance_MCS_Instance_3_n10), .Z0_t (LED_128_Instance_mixcolumns_out[60]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U27 ( .A0_t (LED_128_Instance_MCS_Instance_3_n9), .B0_t (LED_128_Instance_MCS_Instance_3_n36), .Z0_t (LED_128_Instance_MCS_Instance_3_n10) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U26 ( .A0_t (LED_128_Instance_MCS_Instance_3_n11), .B0_t (LED_128_Instance_MCS_Instance_3_n8), .Z0_t (LED_128_Instance_MCS_Instance_3_n9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U25 ( .A0_t (LED_128_Instance_subcells_out[15]), .B0_t (LED_128_Instance_MCS_Instance_3_n37), .Z0_t (LED_128_Instance_MCS_Instance_3_n11) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U24 ( .A0_t (LED_128_Instance_subcells_out[59]), .B0_t (LED_128_Instance_MCS_Instance_3_n30), .Z0_t (LED_128_Instance_MCS_Instance_3_n37) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U23 ( .A0_t (LED_128_Instance_subcells_out[56]), .B0_t (LED_128_Instance_subcells_out[36]), .Z0_t (LED_128_Instance_MCS_Instance_3_n30) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U22 ( .A0_t (LED_128_Instance_MCS_Instance_3_n7), .B0_t (LED_128_Instance_MCS_Instance_3_n17), .Z0_t (LED_128_Instance_mixcolumns_out[14]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U21 ( .A0_t (LED_128_Instance_MCS_Instance_3_n18), .B0_t (LED_128_Instance_subcells_out[15]), .Z0_t (LED_128_Instance_MCS_Instance_3_n7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U20 ( .A0_t (LED_128_Instance_subcells_out[12]), .B0_t (LED_128_Instance_subcells_out[57]), .Z0_t (LED_128_Instance_MCS_Instance_3_n18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U19 ( .A0_t (LED_128_Instance_MCS_Instance_3_n6), .B0_t (LED_128_Instance_MCS_Instance_3_n5), .Z0_t (LED_128_Instance_mixcolumns_out[29]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U18 ( .A0_t (LED_128_Instance_MCS_Instance_3_n19), .B0_t (LED_128_Instance_MCS_Instance_3_n15), .Z0_t (LED_128_Instance_MCS_Instance_3_n6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U17 ( .A0_t (LED_128_Instance_MCS_Instance_3_n17), .B0_t (LED_128_Instance_MCS_Instance_3_n23), .Z0_t (LED_128_Instance_MCS_Instance_3_n15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U16 ( .A0_t (LED_128_Instance_subcells_out[58]), .B0_t (LED_128_Instance_subcells_out[38]), .Z0_t (LED_128_Instance_MCS_Instance_3_n23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U15 ( .A0_t (LED_128_Instance_subcells_out[37]), .B0_t (LED_128_Instance_subcells_out[18]), .Z0_t (LED_128_Instance_MCS_Instance_3_n17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U14 ( .A0_t (LED_128_Instance_subcells_out[56]), .B0_t (LED_128_Instance_subcells_out[13]), .Z0_t (LED_128_Instance_MCS_Instance_3_n19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U13 ( .A0_t (LED_128_Instance_subcells_out[13]), .B0_t (LED_128_Instance_MCS_Instance_3_n4), .Z0_t (LED_128_Instance_mixcolumns_out[15]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U12 ( .A0_t (LED_128_Instance_MCS_Instance_3_n3), .B0_t (LED_128_Instance_MCS_Instance_3_n2), .Z0_t (LED_128_Instance_mixcolumns_out[28]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U11 ( .A0_t (LED_128_Instance_subcells_out[18]), .B0_t (LED_128_Instance_MCS_Instance_3_n4), .Z0_t (LED_128_Instance_MCS_Instance_3_n3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U10 ( .A0_t (LED_128_Instance_subcells_out[58]), .B0_t (LED_128_Instance_MCS_Instance_3_n36), .Z0_t (LED_128_Instance_MCS_Instance_3_n4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U9 ( .A0_t (LED_128_Instance_subcells_out[19]), .B0_t (LED_128_Instance_subcells_out[38]), .Z0_t (LED_128_Instance_MCS_Instance_3_n36) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U8 ( .A0_t (LED_128_Instance_subcells_out[59]), .B0_t (LED_128_Instance_MCS_Instance_3_n5), .Z0_t (LED_128_Instance_mixcolumns_out[12]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U7 ( .A0_t (LED_128_Instance_subcells_out[39]), .B0_t (LED_128_Instance_MCS_Instance_3_n35), .Z0_t (LED_128_Instance_MCS_Instance_3_n5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U6 ( .A0_t (LED_128_Instance_subcells_out[14]), .B0_t (LED_128_Instance_subcells_out[16]), .Z0_t (LED_128_Instance_MCS_Instance_3_n35) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U5 ( .A0_t (LED_128_Instance_MCS_Instance_3_n1), .B0_t (LED_128_Instance_MCS_Instance_3_n8), .Z0_t (LED_128_Instance_mixcolumns_out[62]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U4 ( .A0_t (LED_128_Instance_subcells_out[57]), .B0_t (LED_128_Instance_subcells_out[37]), .Z0_t (LED_128_Instance_MCS_Instance_3_n8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U3 ( .A0_t (LED_128_Instance_subcells_out[17]), .B0_t (LED_128_Instance_MCS_Instance_3_n2), .Z0_t (LED_128_Instance_MCS_Instance_3_n1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U2 ( .A0_t (LED_128_Instance_subcells_out[36]), .B0_t (LED_128_Instance_MCS_Instance_3_n26), .Z0_t (LED_128_Instance_MCS_Instance_3_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U1 ( .A0_t (LED_128_Instance_subcells_out[13]), .B0_t (LED_128_Instance_subcells_out[59]), .Z0_t (LED_128_Instance_MCS_Instance_3_n26) ) ;

    /* register cells */
endmodule
