//-----------------------------------------

module top(input wire [59:0] io_in_0t, io_in_0f, io_in_1t, io_in_1f, ctrl_io_in_0t, ctrl_io_in_0f,  output wire [59:0] io_out_0t, io_out_0f, io_out_1t, io_out_1f, io_oeb, ctrl_io_out_0t, ctrl_io_out_0f, ctrl_io_oeb);


    assign io_oeb      = 60'b11111111000000000000;
    assign ctrl_io_oeb = 60'b10000;

    AES_SAUBER_Pipeline_d1 generated_module (
        .port_in_s0_t(io_in_0t[7:0]),
        .port_in_s0_f(io_in_0f[7:0]),
        .port_in_s1_t(io_in_1t[7:0]),
        .port_in_s1_f(io_in_1f[7:0]),
        .start_t(ctrl_io_in_0t[1]),
        .start_f(ctrl_io_in_0f[1]),
        .done_t(ctrl_io_out_0t[5]),
        .done_f(ctrl_io_out_0f[5]),
        .port_out_s0_t(io_out_0t[19:12]),
        .port_out_s0_f(io_out_0f[19:12]),
        .port_out_s1_t(io_out_1t[19:12]),
        .port_out_s1_f(io_out_1f[19:12])
    );

endmodule


/* modified netlist. Source: module AES in file /mnt/c/Users/amirm/Desktop/Papers_in_progress/SAUBER/Design for our FPGA/6-AES_EncSerial_PortSerial/4-AGEMA/AES.v */
/* 0 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 1 register stage(s) in total */

module AES_SAUBER_Pipeline_d1 (port_in_s0_t, start_t, start_f, port_in_s0_f, port_in_s1_t, port_in_s1_f, port_out_s0_t, done_t, port_out_s0_f, port_out_s1_t, port_out_s1_f, done_f);
    input [7:0] port_in_s0_t ;
    input start_t ;
    input start_f ;
    input [7:0] port_in_s0_f ;
    input [7:0] port_in_s1_t ;
    input [7:0] port_in_s1_f ;
    output [7:0] port_out_s0_t ;
    output done_t ;
    output [7:0] port_out_s0_f ;
    output [7:0] port_out_s1_t ;
    output [7:0] port_out_s1_f ;
    output done_f ;
    wire selMC ;
    wire selXOR ;
    wire enRCon ;
    wire intFinal ;
    wire enKS ;
    wire intselXOR ;
    wire notFirst ;
    wire ctrl_n24 ;
    wire ctrl_n19 ;
    wire ctrl_n18 ;
    wire ctrl_n17 ;
    wire ctrl_n14 ;
    wire ctrl_n13 ;
    wire ctrl_n12 ;
    wire ctrl_n11 ;
    wire ctrl_n10 ;
    wire ctrl_n9 ;
    wire ctrl_n4 ;
    wire ctrl_finalStep ;
    wire ctrl_n5 ;
    wire ctrl_seq4Out_1_ ;
    wire ctrl_seq4In_1_ ;
    wire ctrl_nRstSeq4 ;
    wire ctrl_n22 ;
    wire ctrl_seq6Out_4_ ;
    wire ctrl_seq6In_1_ ;
    wire ctrl_seq6In_2_ ;
    wire ctrl_seq6In_3_ ;
    wire ctrl_seq6In_4_ ;
    wire ctrl_seq6_SFF_0_n2 ;
    wire ctrl_seq6_SFF_0_n1 ;
    wire ctrl_seq6_SFF_0_QD ;
    wire ctrl_seq6_SFF_0_MUXInst_Y ;
    wire ctrl_seq6_SFF_0_MUXInst_X ;
    wire ctrl_seq6_SFF_1_n2 ;
    wire ctrl_seq6_SFF_1_n1 ;
    wire ctrl_seq6_SFF_1_QD ;
    wire ctrl_seq6_SFF_1_MUXInst_Y ;
    wire ctrl_seq6_SFF_1_MUXInst_X ;
    wire ctrl_seq6_SFF_2_n2 ;
    wire ctrl_seq6_SFF_2_n1 ;
    wire ctrl_seq6_SFF_2_QD ;
    wire ctrl_seq6_SFF_2_MUXInst_Y ;
    wire ctrl_seq6_SFF_2_MUXInst_X ;
    wire ctrl_seq6_SFF_3_n2 ;
    wire ctrl_seq6_SFF_3_n1 ;
    wire ctrl_seq6_SFF_3_QD ;
    wire ctrl_seq6_SFF_3_MUXInst_Y ;
    wire ctrl_seq6_SFF_3_MUXInst_X ;
    wire ctrl_seq6_SFF_4_n2 ;
    wire ctrl_seq6_SFF_4_n1 ;
    wire ctrl_seq6_SFF_4_QD ;
    wire ctrl_seq6_SFF_4_MUXInst_Y ;
    wire ctrl_seq6_SFF_4_MUXInst_X ;
    wire ctrl_seq4_SFF_0_n2 ;
    wire ctrl_seq4_SFF_0_n1 ;
    wire ctrl_seq4_SFF_0_QD ;
    wire ctrl_seq4_SFF_0_MUXInst_Y ;
    wire ctrl_seq4_SFF_0_MUXInst_X ;
    wire ctrl_seq4_SFF_1_n2 ;
    wire ctrl_seq4_SFF_1_n1 ;
    wire ctrl_seq4_SFF_1_QD ;
    wire ctrl_seq4_SFF_1_MUXInst_Y ;
    wire ctrl_seq4_SFF_1_MUXInst_X ;
    wire MUX_StateIn_mux_inst_0_Y ;
    wire MUX_StateIn_mux_inst_0_X ;
    wire MUX_StateIn_mux_inst_1_Y ;
    wire MUX_StateIn_mux_inst_1_X ;
    wire MUX_StateIn_mux_inst_2_Y ;
    wire MUX_StateIn_mux_inst_2_X ;
    wire MUX_StateIn_mux_inst_3_Y ;
    wire MUX_StateIn_mux_inst_3_X ;
    wire MUX_StateIn_mux_inst_4_Y ;
    wire MUX_StateIn_mux_inst_4_X ;
    wire MUX_StateIn_mux_inst_5_Y ;
    wire MUX_StateIn_mux_inst_5_X ;
    wire MUX_StateIn_mux_inst_6_Y ;
    wire MUX_StateIn_mux_inst_6_X ;
    wire MUX_StateIn_mux_inst_7_Y ;
    wire MUX_StateIn_mux_inst_7_X ;
    wire stateArray_nReset_selMC ;
    wire stateArray_S00reg_gff_1_SFF_0_MUXInst_Y ;
    wire stateArray_S00reg_gff_1_SFF_0_MUXInst_X ;
    wire stateArray_S00reg_gff_1_SFF_1_MUXInst_Y ;
    wire stateArray_S00reg_gff_1_SFF_1_MUXInst_X ;
    wire stateArray_S00reg_gff_1_SFF_2_MUXInst_Y ;
    wire stateArray_S00reg_gff_1_SFF_2_MUXInst_X ;
    wire stateArray_S00reg_gff_1_SFF_3_MUXInst_Y ;
    wire stateArray_S00reg_gff_1_SFF_3_MUXInst_X ;
    wire stateArray_S00reg_gff_1_SFF_4_MUXInst_Y ;
    wire stateArray_S00reg_gff_1_SFF_4_MUXInst_X ;
    wire stateArray_S00reg_gff_1_SFF_5_MUXInst_Y ;
    wire stateArray_S00reg_gff_1_SFF_5_MUXInst_X ;
    wire stateArray_S00reg_gff_1_SFF_6_MUXInst_Y ;
    wire stateArray_S00reg_gff_1_SFF_6_MUXInst_X ;
    wire stateArray_S00reg_gff_1_SFF_7_MUXInst_Y ;
    wire stateArray_S00reg_gff_1_SFF_7_MUXInst_X ;
    wire stateArray_S01reg_gff_1_SFF_0_MUXInst_Y ;
    wire stateArray_S01reg_gff_1_SFF_0_MUXInst_X ;
    wire stateArray_S01reg_gff_1_SFF_1_MUXInst_Y ;
    wire stateArray_S01reg_gff_1_SFF_1_MUXInst_X ;
    wire stateArray_S01reg_gff_1_SFF_2_MUXInst_Y ;
    wire stateArray_S01reg_gff_1_SFF_2_MUXInst_X ;
    wire stateArray_S01reg_gff_1_SFF_3_MUXInst_Y ;
    wire stateArray_S01reg_gff_1_SFF_3_MUXInst_X ;
    wire stateArray_S01reg_gff_1_SFF_4_MUXInst_Y ;
    wire stateArray_S01reg_gff_1_SFF_4_MUXInst_X ;
    wire stateArray_S01reg_gff_1_SFF_5_MUXInst_Y ;
    wire stateArray_S01reg_gff_1_SFF_5_MUXInst_X ;
    wire stateArray_S01reg_gff_1_SFF_6_MUXInst_Y ;
    wire stateArray_S01reg_gff_1_SFF_6_MUXInst_X ;
    wire stateArray_S01reg_gff_1_SFF_7_MUXInst_Y ;
    wire stateArray_S01reg_gff_1_SFF_7_MUXInst_X ;
    wire stateArray_S02reg_gff_1_SFF_0_MUXInst_Y ;
    wire stateArray_S02reg_gff_1_SFF_0_MUXInst_X ;
    wire stateArray_S02reg_gff_1_SFF_1_MUXInst_Y ;
    wire stateArray_S02reg_gff_1_SFF_1_MUXInst_X ;
    wire stateArray_S02reg_gff_1_SFF_2_MUXInst_Y ;
    wire stateArray_S02reg_gff_1_SFF_2_MUXInst_X ;
    wire stateArray_S02reg_gff_1_SFF_3_MUXInst_Y ;
    wire stateArray_S02reg_gff_1_SFF_3_MUXInst_X ;
    wire stateArray_S02reg_gff_1_SFF_4_MUXInst_Y ;
    wire stateArray_S02reg_gff_1_SFF_4_MUXInst_X ;
    wire stateArray_S02reg_gff_1_SFF_5_MUXInst_Y ;
    wire stateArray_S02reg_gff_1_SFF_5_MUXInst_X ;
    wire stateArray_S02reg_gff_1_SFF_6_MUXInst_Y ;
    wire stateArray_S02reg_gff_1_SFF_6_MUXInst_X ;
    wire stateArray_S02reg_gff_1_SFF_7_MUXInst_Y ;
    wire stateArray_S02reg_gff_1_SFF_7_MUXInst_X ;
    wire stateArray_S03reg_gff_1_SFF_0_MUXInst_Y ;
    wire stateArray_S03reg_gff_1_SFF_0_MUXInst_X ;
    wire stateArray_S03reg_gff_1_SFF_1_MUXInst_Y ;
    wire stateArray_S03reg_gff_1_SFF_1_MUXInst_X ;
    wire stateArray_S03reg_gff_1_SFF_2_MUXInst_Y ;
    wire stateArray_S03reg_gff_1_SFF_2_MUXInst_X ;
    wire stateArray_S03reg_gff_1_SFF_3_MUXInst_Y ;
    wire stateArray_S03reg_gff_1_SFF_3_MUXInst_X ;
    wire stateArray_S03reg_gff_1_SFF_4_MUXInst_Y ;
    wire stateArray_S03reg_gff_1_SFF_4_MUXInst_X ;
    wire stateArray_S03reg_gff_1_SFF_5_MUXInst_Y ;
    wire stateArray_S03reg_gff_1_SFF_5_MUXInst_X ;
    wire stateArray_S03reg_gff_1_SFF_6_MUXInst_Y ;
    wire stateArray_S03reg_gff_1_SFF_6_MUXInst_X ;
    wire stateArray_S03reg_gff_1_SFF_7_MUXInst_Y ;
    wire stateArray_S03reg_gff_1_SFF_7_MUXInst_X ;
    wire stateArray_S10reg_gff_1_SFF_0_MUXInst_Y ;
    wire stateArray_S10reg_gff_1_SFF_0_MUXInst_X ;
    wire stateArray_S10reg_gff_1_SFF_1_MUXInst_Y ;
    wire stateArray_S10reg_gff_1_SFF_1_MUXInst_X ;
    wire stateArray_S10reg_gff_1_SFF_2_MUXInst_Y ;
    wire stateArray_S10reg_gff_1_SFF_2_MUXInst_X ;
    wire stateArray_S10reg_gff_1_SFF_3_MUXInst_Y ;
    wire stateArray_S10reg_gff_1_SFF_3_MUXInst_X ;
    wire stateArray_S10reg_gff_1_SFF_4_MUXInst_Y ;
    wire stateArray_S10reg_gff_1_SFF_4_MUXInst_X ;
    wire stateArray_S10reg_gff_1_SFF_5_MUXInst_Y ;
    wire stateArray_S10reg_gff_1_SFF_5_MUXInst_X ;
    wire stateArray_S10reg_gff_1_SFF_6_MUXInst_Y ;
    wire stateArray_S10reg_gff_1_SFF_6_MUXInst_X ;
    wire stateArray_S10reg_gff_1_SFF_7_MUXInst_Y ;
    wire stateArray_S10reg_gff_1_SFF_7_MUXInst_X ;
    wire stateArray_S11reg_gff_1_SFF_0_MUXInst_Y ;
    wire stateArray_S11reg_gff_1_SFF_0_MUXInst_X ;
    wire stateArray_S11reg_gff_1_SFF_1_MUXInst_Y ;
    wire stateArray_S11reg_gff_1_SFF_1_MUXInst_X ;
    wire stateArray_S11reg_gff_1_SFF_2_MUXInst_Y ;
    wire stateArray_S11reg_gff_1_SFF_2_MUXInst_X ;
    wire stateArray_S11reg_gff_1_SFF_3_MUXInst_Y ;
    wire stateArray_S11reg_gff_1_SFF_3_MUXInst_X ;
    wire stateArray_S11reg_gff_1_SFF_4_MUXInst_Y ;
    wire stateArray_S11reg_gff_1_SFF_4_MUXInst_X ;
    wire stateArray_S11reg_gff_1_SFF_5_MUXInst_Y ;
    wire stateArray_S11reg_gff_1_SFF_5_MUXInst_X ;
    wire stateArray_S11reg_gff_1_SFF_6_MUXInst_Y ;
    wire stateArray_S11reg_gff_1_SFF_6_MUXInst_X ;
    wire stateArray_S11reg_gff_1_SFF_7_MUXInst_Y ;
    wire stateArray_S11reg_gff_1_SFF_7_MUXInst_X ;
    wire stateArray_S12reg_gff_1_SFF_0_MUXInst_Y ;
    wire stateArray_S12reg_gff_1_SFF_0_MUXInst_X ;
    wire stateArray_S12reg_gff_1_SFF_1_MUXInst_Y ;
    wire stateArray_S12reg_gff_1_SFF_1_MUXInst_X ;
    wire stateArray_S12reg_gff_1_SFF_2_MUXInst_Y ;
    wire stateArray_S12reg_gff_1_SFF_2_MUXInst_X ;
    wire stateArray_S12reg_gff_1_SFF_3_MUXInst_Y ;
    wire stateArray_S12reg_gff_1_SFF_3_MUXInst_X ;
    wire stateArray_S12reg_gff_1_SFF_4_MUXInst_Y ;
    wire stateArray_S12reg_gff_1_SFF_4_MUXInst_X ;
    wire stateArray_S12reg_gff_1_SFF_5_MUXInst_Y ;
    wire stateArray_S12reg_gff_1_SFF_5_MUXInst_X ;
    wire stateArray_S12reg_gff_1_SFF_6_MUXInst_Y ;
    wire stateArray_S12reg_gff_1_SFF_6_MUXInst_X ;
    wire stateArray_S12reg_gff_1_SFF_7_MUXInst_Y ;
    wire stateArray_S12reg_gff_1_SFF_7_MUXInst_X ;
    wire stateArray_S13reg_gff_1_SFF_0_MUXInst_Y ;
    wire stateArray_S13reg_gff_1_SFF_0_MUXInst_X ;
    wire stateArray_S13reg_gff_1_SFF_1_MUXInst_Y ;
    wire stateArray_S13reg_gff_1_SFF_1_MUXInst_X ;
    wire stateArray_S13reg_gff_1_SFF_2_MUXInst_Y ;
    wire stateArray_S13reg_gff_1_SFF_2_MUXInst_X ;
    wire stateArray_S13reg_gff_1_SFF_3_MUXInst_Y ;
    wire stateArray_S13reg_gff_1_SFF_3_MUXInst_X ;
    wire stateArray_S13reg_gff_1_SFF_4_MUXInst_Y ;
    wire stateArray_S13reg_gff_1_SFF_4_MUXInst_X ;
    wire stateArray_S13reg_gff_1_SFF_5_MUXInst_Y ;
    wire stateArray_S13reg_gff_1_SFF_5_MUXInst_X ;
    wire stateArray_S13reg_gff_1_SFF_6_MUXInst_Y ;
    wire stateArray_S13reg_gff_1_SFF_6_MUXInst_X ;
    wire stateArray_S13reg_gff_1_SFF_7_MUXInst_Y ;
    wire stateArray_S13reg_gff_1_SFF_7_MUXInst_X ;
    wire stateArray_S20reg_gff_1_SFF_0_MUXInst_Y ;
    wire stateArray_S20reg_gff_1_SFF_0_MUXInst_X ;
    wire stateArray_S20reg_gff_1_SFF_1_MUXInst_Y ;
    wire stateArray_S20reg_gff_1_SFF_1_MUXInst_X ;
    wire stateArray_S20reg_gff_1_SFF_2_MUXInst_Y ;
    wire stateArray_S20reg_gff_1_SFF_2_MUXInst_X ;
    wire stateArray_S20reg_gff_1_SFF_3_MUXInst_Y ;
    wire stateArray_S20reg_gff_1_SFF_3_MUXInst_X ;
    wire stateArray_S20reg_gff_1_SFF_4_MUXInst_Y ;
    wire stateArray_S20reg_gff_1_SFF_4_MUXInst_X ;
    wire stateArray_S20reg_gff_1_SFF_5_MUXInst_Y ;
    wire stateArray_S20reg_gff_1_SFF_5_MUXInst_X ;
    wire stateArray_S20reg_gff_1_SFF_6_MUXInst_Y ;
    wire stateArray_S20reg_gff_1_SFF_6_MUXInst_X ;
    wire stateArray_S20reg_gff_1_SFF_7_MUXInst_Y ;
    wire stateArray_S20reg_gff_1_SFF_7_MUXInst_X ;
    wire stateArray_S21reg_gff_1_SFF_0_MUXInst_Y ;
    wire stateArray_S21reg_gff_1_SFF_0_MUXInst_X ;
    wire stateArray_S21reg_gff_1_SFF_1_MUXInst_Y ;
    wire stateArray_S21reg_gff_1_SFF_1_MUXInst_X ;
    wire stateArray_S21reg_gff_1_SFF_2_MUXInst_Y ;
    wire stateArray_S21reg_gff_1_SFF_2_MUXInst_X ;
    wire stateArray_S21reg_gff_1_SFF_3_MUXInst_Y ;
    wire stateArray_S21reg_gff_1_SFF_3_MUXInst_X ;
    wire stateArray_S21reg_gff_1_SFF_4_MUXInst_Y ;
    wire stateArray_S21reg_gff_1_SFF_4_MUXInst_X ;
    wire stateArray_S21reg_gff_1_SFF_5_MUXInst_Y ;
    wire stateArray_S21reg_gff_1_SFF_5_MUXInst_X ;
    wire stateArray_S21reg_gff_1_SFF_6_MUXInst_Y ;
    wire stateArray_S21reg_gff_1_SFF_6_MUXInst_X ;
    wire stateArray_S21reg_gff_1_SFF_7_MUXInst_Y ;
    wire stateArray_S21reg_gff_1_SFF_7_MUXInst_X ;
    wire stateArray_S22reg_gff_1_SFF_0_MUXInst_Y ;
    wire stateArray_S22reg_gff_1_SFF_0_MUXInst_X ;
    wire stateArray_S22reg_gff_1_SFF_1_MUXInst_Y ;
    wire stateArray_S22reg_gff_1_SFF_1_MUXInst_X ;
    wire stateArray_S22reg_gff_1_SFF_2_MUXInst_Y ;
    wire stateArray_S22reg_gff_1_SFF_2_MUXInst_X ;
    wire stateArray_S22reg_gff_1_SFF_3_MUXInst_Y ;
    wire stateArray_S22reg_gff_1_SFF_3_MUXInst_X ;
    wire stateArray_S22reg_gff_1_SFF_4_MUXInst_Y ;
    wire stateArray_S22reg_gff_1_SFF_4_MUXInst_X ;
    wire stateArray_S22reg_gff_1_SFF_5_MUXInst_Y ;
    wire stateArray_S22reg_gff_1_SFF_5_MUXInst_X ;
    wire stateArray_S22reg_gff_1_SFF_6_MUXInst_Y ;
    wire stateArray_S22reg_gff_1_SFF_6_MUXInst_X ;
    wire stateArray_S22reg_gff_1_SFF_7_MUXInst_Y ;
    wire stateArray_S22reg_gff_1_SFF_7_MUXInst_X ;
    wire stateArray_S23reg_gff_1_SFF_0_MUXInst_Y ;
    wire stateArray_S23reg_gff_1_SFF_0_MUXInst_X ;
    wire stateArray_S23reg_gff_1_SFF_1_MUXInst_Y ;
    wire stateArray_S23reg_gff_1_SFF_1_MUXInst_X ;
    wire stateArray_S23reg_gff_1_SFF_2_MUXInst_Y ;
    wire stateArray_S23reg_gff_1_SFF_2_MUXInst_X ;
    wire stateArray_S23reg_gff_1_SFF_3_MUXInst_Y ;
    wire stateArray_S23reg_gff_1_SFF_3_MUXInst_X ;
    wire stateArray_S23reg_gff_1_SFF_4_MUXInst_Y ;
    wire stateArray_S23reg_gff_1_SFF_4_MUXInst_X ;
    wire stateArray_S23reg_gff_1_SFF_5_MUXInst_Y ;
    wire stateArray_S23reg_gff_1_SFF_5_MUXInst_X ;
    wire stateArray_S23reg_gff_1_SFF_6_MUXInst_Y ;
    wire stateArray_S23reg_gff_1_SFF_6_MUXInst_X ;
    wire stateArray_S23reg_gff_1_SFF_7_MUXInst_Y ;
    wire stateArray_S23reg_gff_1_SFF_7_MUXInst_X ;
    wire stateArray_S30reg_gff_1_SFF_0_MUXInst_Y ;
    wire stateArray_S30reg_gff_1_SFF_0_MUXInst_X ;
    wire stateArray_S30reg_gff_1_SFF_1_MUXInst_Y ;
    wire stateArray_S30reg_gff_1_SFF_1_MUXInst_X ;
    wire stateArray_S30reg_gff_1_SFF_2_MUXInst_Y ;
    wire stateArray_S30reg_gff_1_SFF_2_MUXInst_X ;
    wire stateArray_S30reg_gff_1_SFF_3_MUXInst_Y ;
    wire stateArray_S30reg_gff_1_SFF_3_MUXInst_X ;
    wire stateArray_S30reg_gff_1_SFF_4_MUXInst_Y ;
    wire stateArray_S30reg_gff_1_SFF_4_MUXInst_X ;
    wire stateArray_S30reg_gff_1_SFF_5_MUXInst_Y ;
    wire stateArray_S30reg_gff_1_SFF_5_MUXInst_X ;
    wire stateArray_S30reg_gff_1_SFF_6_MUXInst_Y ;
    wire stateArray_S30reg_gff_1_SFF_6_MUXInst_X ;
    wire stateArray_S30reg_gff_1_SFF_7_MUXInst_Y ;
    wire stateArray_S30reg_gff_1_SFF_7_MUXInst_X ;
    wire stateArray_S31reg_gff_1_SFF_0_MUXInst_Y ;
    wire stateArray_S31reg_gff_1_SFF_0_MUXInst_X ;
    wire stateArray_S31reg_gff_1_SFF_1_MUXInst_Y ;
    wire stateArray_S31reg_gff_1_SFF_1_MUXInst_X ;
    wire stateArray_S31reg_gff_1_SFF_2_MUXInst_Y ;
    wire stateArray_S31reg_gff_1_SFF_2_MUXInst_X ;
    wire stateArray_S31reg_gff_1_SFF_3_MUXInst_Y ;
    wire stateArray_S31reg_gff_1_SFF_3_MUXInst_X ;
    wire stateArray_S31reg_gff_1_SFF_4_MUXInst_Y ;
    wire stateArray_S31reg_gff_1_SFF_4_MUXInst_X ;
    wire stateArray_S31reg_gff_1_SFF_5_MUXInst_Y ;
    wire stateArray_S31reg_gff_1_SFF_5_MUXInst_X ;
    wire stateArray_S31reg_gff_1_SFF_6_MUXInst_Y ;
    wire stateArray_S31reg_gff_1_SFF_6_MUXInst_X ;
    wire stateArray_S31reg_gff_1_SFF_7_MUXInst_Y ;
    wire stateArray_S31reg_gff_1_SFF_7_MUXInst_X ;
    wire stateArray_S32reg_gff_1_SFF_0_MUXInst_Y ;
    wire stateArray_S32reg_gff_1_SFF_0_MUXInst_X ;
    wire stateArray_S32reg_gff_1_SFF_1_MUXInst_Y ;
    wire stateArray_S32reg_gff_1_SFF_1_MUXInst_X ;
    wire stateArray_S32reg_gff_1_SFF_2_MUXInst_Y ;
    wire stateArray_S32reg_gff_1_SFF_2_MUXInst_X ;
    wire stateArray_S32reg_gff_1_SFF_3_MUXInst_Y ;
    wire stateArray_S32reg_gff_1_SFF_3_MUXInst_X ;
    wire stateArray_S32reg_gff_1_SFF_4_MUXInst_Y ;
    wire stateArray_S32reg_gff_1_SFF_4_MUXInst_X ;
    wire stateArray_S32reg_gff_1_SFF_5_MUXInst_Y ;
    wire stateArray_S32reg_gff_1_SFF_5_MUXInst_X ;
    wire stateArray_S32reg_gff_1_SFF_6_MUXInst_Y ;
    wire stateArray_S32reg_gff_1_SFF_6_MUXInst_X ;
    wire stateArray_S32reg_gff_1_SFF_7_MUXInst_Y ;
    wire stateArray_S32reg_gff_1_SFF_7_MUXInst_X ;
    wire stateArray_S33reg_gff_1_SFF_0_MUXInst_Y ;
    wire stateArray_S33reg_gff_1_SFF_0_MUXInst_X ;
    wire stateArray_S33reg_gff_1_SFF_1_MUXInst_Y ;
    wire stateArray_S33reg_gff_1_SFF_1_MUXInst_X ;
    wire stateArray_S33reg_gff_1_SFF_2_MUXInst_Y ;
    wire stateArray_S33reg_gff_1_SFF_2_MUXInst_X ;
    wire stateArray_S33reg_gff_1_SFF_3_MUXInst_Y ;
    wire stateArray_S33reg_gff_1_SFF_3_MUXInst_X ;
    wire stateArray_S33reg_gff_1_SFF_4_MUXInst_Y ;
    wire stateArray_S33reg_gff_1_SFF_4_MUXInst_X ;
    wire stateArray_S33reg_gff_1_SFF_5_MUXInst_Y ;
    wire stateArray_S33reg_gff_1_SFF_5_MUXInst_X ;
    wire stateArray_S33reg_gff_1_SFF_6_MUXInst_Y ;
    wire stateArray_S33reg_gff_1_SFF_6_MUXInst_X ;
    wire stateArray_S33reg_gff_1_SFF_7_MUXInst_Y ;
    wire stateArray_S33reg_gff_1_SFF_7_MUXInst_X ;
    wire stateArray_MUX_inS03ser_mux_inst_0_Y ;
    wire stateArray_MUX_inS03ser_mux_inst_0_X ;
    wire stateArray_MUX_inS03ser_mux_inst_1_Y ;
    wire stateArray_MUX_inS03ser_mux_inst_1_X ;
    wire stateArray_MUX_inS03ser_mux_inst_2_Y ;
    wire stateArray_MUX_inS03ser_mux_inst_2_X ;
    wire stateArray_MUX_inS03ser_mux_inst_3_Y ;
    wire stateArray_MUX_inS03ser_mux_inst_3_X ;
    wire stateArray_MUX_inS03ser_mux_inst_4_Y ;
    wire stateArray_MUX_inS03ser_mux_inst_4_X ;
    wire stateArray_MUX_inS03ser_mux_inst_5_Y ;
    wire stateArray_MUX_inS03ser_mux_inst_5_X ;
    wire stateArray_MUX_inS03ser_mux_inst_6_Y ;
    wire stateArray_MUX_inS03ser_mux_inst_6_X ;
    wire stateArray_MUX_inS03ser_mux_inst_7_Y ;
    wire stateArray_MUX_inS03ser_mux_inst_7_X ;
    wire stateArray_MUX_inS13ser_mux_inst_0_Y ;
    wire stateArray_MUX_inS13ser_mux_inst_0_X ;
    wire stateArray_MUX_inS13ser_mux_inst_1_Y ;
    wire stateArray_MUX_inS13ser_mux_inst_1_X ;
    wire stateArray_MUX_inS13ser_mux_inst_2_Y ;
    wire stateArray_MUX_inS13ser_mux_inst_2_X ;
    wire stateArray_MUX_inS13ser_mux_inst_3_Y ;
    wire stateArray_MUX_inS13ser_mux_inst_3_X ;
    wire stateArray_MUX_inS13ser_mux_inst_4_Y ;
    wire stateArray_MUX_inS13ser_mux_inst_4_X ;
    wire stateArray_MUX_inS13ser_mux_inst_5_Y ;
    wire stateArray_MUX_inS13ser_mux_inst_5_X ;
    wire stateArray_MUX_inS13ser_mux_inst_6_Y ;
    wire stateArray_MUX_inS13ser_mux_inst_6_X ;
    wire stateArray_MUX_inS13ser_mux_inst_7_Y ;
    wire stateArray_MUX_inS13ser_mux_inst_7_X ;
    wire stateArray_MUX_inS23ser_mux_inst_0_Y ;
    wire stateArray_MUX_inS23ser_mux_inst_0_X ;
    wire stateArray_MUX_inS23ser_mux_inst_1_Y ;
    wire stateArray_MUX_inS23ser_mux_inst_1_X ;
    wire stateArray_MUX_inS23ser_mux_inst_2_Y ;
    wire stateArray_MUX_inS23ser_mux_inst_2_X ;
    wire stateArray_MUX_inS23ser_mux_inst_3_Y ;
    wire stateArray_MUX_inS23ser_mux_inst_3_X ;
    wire stateArray_MUX_inS23ser_mux_inst_4_Y ;
    wire stateArray_MUX_inS23ser_mux_inst_4_X ;
    wire stateArray_MUX_inS23ser_mux_inst_5_Y ;
    wire stateArray_MUX_inS23ser_mux_inst_5_X ;
    wire stateArray_MUX_inS23ser_mux_inst_6_Y ;
    wire stateArray_MUX_inS23ser_mux_inst_6_X ;
    wire stateArray_MUX_inS23ser_mux_inst_7_Y ;
    wire stateArray_MUX_inS23ser_mux_inst_7_X ;
    wire stateArray_MUX_input_MC_mux_inst_0_Y ;
    wire stateArray_MUX_input_MC_mux_inst_0_X ;
    wire stateArray_MUX_input_MC_mux_inst_1_Y ;
    wire stateArray_MUX_input_MC_mux_inst_1_X ;
    wire stateArray_MUX_input_MC_mux_inst_2_Y ;
    wire stateArray_MUX_input_MC_mux_inst_2_X ;
    wire stateArray_MUX_input_MC_mux_inst_3_Y ;
    wire stateArray_MUX_input_MC_mux_inst_3_X ;
    wire stateArray_MUX_input_MC_mux_inst_4_Y ;
    wire stateArray_MUX_input_MC_mux_inst_4_X ;
    wire stateArray_MUX_input_MC_mux_inst_5_Y ;
    wire stateArray_MUX_input_MC_mux_inst_5_X ;
    wire stateArray_MUX_input_MC_mux_inst_6_Y ;
    wire stateArray_MUX_input_MC_mux_inst_6_X ;
    wire stateArray_MUX_input_MC_mux_inst_7_Y ;
    wire stateArray_MUX_input_MC_mux_inst_7_X ;
    wire stateArray_MUX_inS33ser_mux_inst_0_Y ;
    wire stateArray_MUX_inS33ser_mux_inst_0_X ;
    wire stateArray_MUX_inS33ser_mux_inst_1_Y ;
    wire stateArray_MUX_inS33ser_mux_inst_1_X ;
    wire stateArray_MUX_inS33ser_mux_inst_2_Y ;
    wire stateArray_MUX_inS33ser_mux_inst_2_X ;
    wire stateArray_MUX_inS33ser_mux_inst_3_Y ;
    wire stateArray_MUX_inS33ser_mux_inst_3_X ;
    wire stateArray_MUX_inS33ser_mux_inst_4_Y ;
    wire stateArray_MUX_inS33ser_mux_inst_4_X ;
    wire stateArray_MUX_inS33ser_mux_inst_5_Y ;
    wire stateArray_MUX_inS33ser_mux_inst_5_X ;
    wire stateArray_MUX_inS33ser_mux_inst_6_Y ;
    wire stateArray_MUX_inS33ser_mux_inst_6_X ;
    wire stateArray_MUX_inS33ser_mux_inst_7_Y ;
    wire stateArray_MUX_inS33ser_mux_inst_7_X ;
    wire MUX_StateInMC_mux_inst_0_Y ;
    wire MUX_StateInMC_mux_inst_0_X ;
    wire MUX_StateInMC_mux_inst_1_Y ;
    wire MUX_StateInMC_mux_inst_1_X ;
    wire MUX_StateInMC_mux_inst_2_Y ;
    wire MUX_StateInMC_mux_inst_2_X ;
    wire MUX_StateInMC_mux_inst_3_Y ;
    wire MUX_StateInMC_mux_inst_3_X ;
    wire MUX_StateInMC_mux_inst_4_Y ;
    wire MUX_StateInMC_mux_inst_4_X ;
    wire MUX_StateInMC_mux_inst_5_Y ;
    wire MUX_StateInMC_mux_inst_5_X ;
    wire MUX_StateInMC_mux_inst_6_Y ;
    wire MUX_StateInMC_mux_inst_6_X ;
    wire MUX_StateInMC_mux_inst_7_Y ;
    wire MUX_StateInMC_mux_inst_7_X ;
    wire MUX_StateInMC_mux_inst_8_Y ;
    wire MUX_StateInMC_mux_inst_8_X ;
    wire MUX_StateInMC_mux_inst_9_Y ;
    wire MUX_StateInMC_mux_inst_9_X ;
    wire MUX_StateInMC_mux_inst_10_Y ;
    wire MUX_StateInMC_mux_inst_10_X ;
    wire MUX_StateInMC_mux_inst_11_Y ;
    wire MUX_StateInMC_mux_inst_11_X ;
    wire MUX_StateInMC_mux_inst_12_Y ;
    wire MUX_StateInMC_mux_inst_12_X ;
    wire MUX_StateInMC_mux_inst_13_Y ;
    wire MUX_StateInMC_mux_inst_13_X ;
    wire MUX_StateInMC_mux_inst_14_Y ;
    wire MUX_StateInMC_mux_inst_14_X ;
    wire MUX_StateInMC_mux_inst_15_Y ;
    wire MUX_StateInMC_mux_inst_15_X ;
    wire MUX_StateInMC_mux_inst_16_Y ;
    wire MUX_StateInMC_mux_inst_16_X ;
    wire MUX_StateInMC_mux_inst_17_Y ;
    wire MUX_StateInMC_mux_inst_17_X ;
    wire MUX_StateInMC_mux_inst_18_Y ;
    wire MUX_StateInMC_mux_inst_18_X ;
    wire MUX_StateInMC_mux_inst_19_Y ;
    wire MUX_StateInMC_mux_inst_19_X ;
    wire MUX_StateInMC_mux_inst_20_Y ;
    wire MUX_StateInMC_mux_inst_20_X ;
    wire MUX_StateInMC_mux_inst_21_Y ;
    wire MUX_StateInMC_mux_inst_21_X ;
    wire MUX_StateInMC_mux_inst_22_Y ;
    wire MUX_StateInMC_mux_inst_22_X ;
    wire MUX_StateInMC_mux_inst_23_Y ;
    wire MUX_StateInMC_mux_inst_23_X ;
    wire MUX_StateInMC_mux_inst_24_Y ;
    wire MUX_StateInMC_mux_inst_24_X ;
    wire MUX_StateInMC_mux_inst_25_Y ;
    wire MUX_StateInMC_mux_inst_25_X ;
    wire MUX_StateInMC_mux_inst_26_Y ;
    wire MUX_StateInMC_mux_inst_26_X ;
    wire MUX_StateInMC_mux_inst_27_Y ;
    wire MUX_StateInMC_mux_inst_27_X ;
    wire MUX_StateInMC_mux_inst_28_Y ;
    wire MUX_StateInMC_mux_inst_28_X ;
    wire MUX_StateInMC_mux_inst_29_Y ;
    wire MUX_StateInMC_mux_inst_29_X ;
    wire MUX_StateInMC_mux_inst_30_Y ;
    wire MUX_StateInMC_mux_inst_30_X ;
    wire MUX_StateInMC_mux_inst_31_Y ;
    wire MUX_StateInMC_mux_inst_31_X ;
    wire KeyArray_n32 ;
    wire KeyArray_n31 ;
    wire KeyArray_n30 ;
    wire KeyArray_n29 ;
    wire KeyArray_n28 ;
    wire KeyArray_n27 ;
    wire KeyArray_n26 ;
    wire KeyArray_n25 ;
    wire KeyArray_nReset_selXOR ;
    wire KeyArray_outS01ser_0_ ;
    wire KeyArray_outS01ser_1_ ;
    wire KeyArray_outS01ser_2_ ;
    wire KeyArray_outS01ser_3_ ;
    wire KeyArray_outS01ser_4_ ;
    wire KeyArray_outS01ser_5_ ;
    wire KeyArray_outS01ser_6_ ;
    wire KeyArray_outS01ser_7_ ;
    wire KeyArray_S00reg_gff_1_SFF_0_n2 ;
    wire KeyArray_S00reg_gff_1_SFF_0_n1 ;
    wire KeyArray_S00reg_gff_1_SFF_0_QD ;
    wire KeyArray_S00reg_gff_1_SFF_0_MUXInst_Y ;
    wire KeyArray_S00reg_gff_1_SFF_0_MUXInst_X ;
    wire KeyArray_S00reg_gff_1_SFF_1_n2 ;
    wire KeyArray_S00reg_gff_1_SFF_1_n1 ;
    wire KeyArray_S00reg_gff_1_SFF_1_QD ;
    wire KeyArray_S00reg_gff_1_SFF_1_MUXInst_Y ;
    wire KeyArray_S00reg_gff_1_SFF_1_MUXInst_X ;
    wire KeyArray_S00reg_gff_1_SFF_2_n2 ;
    wire KeyArray_S00reg_gff_1_SFF_2_n1 ;
    wire KeyArray_S00reg_gff_1_SFF_2_QD ;
    wire KeyArray_S00reg_gff_1_SFF_2_MUXInst_Y ;
    wire KeyArray_S00reg_gff_1_SFF_2_MUXInst_X ;
    wire KeyArray_S00reg_gff_1_SFF_3_n2 ;
    wire KeyArray_S00reg_gff_1_SFF_3_n1 ;
    wire KeyArray_S00reg_gff_1_SFF_3_QD ;
    wire KeyArray_S00reg_gff_1_SFF_3_MUXInst_Y ;
    wire KeyArray_S00reg_gff_1_SFF_3_MUXInst_X ;
    wire KeyArray_S00reg_gff_1_SFF_4_n2 ;
    wire KeyArray_S00reg_gff_1_SFF_4_n1 ;
    wire KeyArray_S00reg_gff_1_SFF_4_QD ;
    wire KeyArray_S00reg_gff_1_SFF_4_MUXInst_Y ;
    wire KeyArray_S00reg_gff_1_SFF_4_MUXInst_X ;
    wire KeyArray_S00reg_gff_1_SFF_5_n2 ;
    wire KeyArray_S00reg_gff_1_SFF_5_n1 ;
    wire KeyArray_S00reg_gff_1_SFF_5_QD ;
    wire KeyArray_S00reg_gff_1_SFF_5_MUXInst_Y ;
    wire KeyArray_S00reg_gff_1_SFF_5_MUXInst_X ;
    wire KeyArray_S00reg_gff_1_SFF_6_n2 ;
    wire KeyArray_S00reg_gff_1_SFF_6_n1 ;
    wire KeyArray_S00reg_gff_1_SFF_6_QD ;
    wire KeyArray_S00reg_gff_1_SFF_6_MUXInst_Y ;
    wire KeyArray_S00reg_gff_1_SFF_6_MUXInst_X ;
    wire KeyArray_S00reg_gff_1_SFF_7_n2 ;
    wire KeyArray_S00reg_gff_1_SFF_7_n1 ;
    wire KeyArray_S00reg_gff_1_SFF_7_QD ;
    wire KeyArray_S00reg_gff_1_SFF_7_MUXInst_Y ;
    wire KeyArray_S00reg_gff_1_SFF_7_MUXInst_X ;
    wire KeyArray_S01reg_gff_1_SFF_0_n2 ;
    wire KeyArray_S01reg_gff_1_SFF_0_n1 ;
    wire KeyArray_S01reg_gff_1_SFF_0_QD ;
    wire KeyArray_S01reg_gff_1_SFF_0_MUXInst_Y ;
    wire KeyArray_S01reg_gff_1_SFF_0_MUXInst_X ;
    wire KeyArray_S01reg_gff_1_SFF_1_n2 ;
    wire KeyArray_S01reg_gff_1_SFF_1_n1 ;
    wire KeyArray_S01reg_gff_1_SFF_1_QD ;
    wire KeyArray_S01reg_gff_1_SFF_1_MUXInst_Y ;
    wire KeyArray_S01reg_gff_1_SFF_1_MUXInst_X ;
    wire KeyArray_S01reg_gff_1_SFF_2_n2 ;
    wire KeyArray_S01reg_gff_1_SFF_2_n1 ;
    wire KeyArray_S01reg_gff_1_SFF_2_QD ;
    wire KeyArray_S01reg_gff_1_SFF_2_MUXInst_Y ;
    wire KeyArray_S01reg_gff_1_SFF_2_MUXInst_X ;
    wire KeyArray_S01reg_gff_1_SFF_3_n2 ;
    wire KeyArray_S01reg_gff_1_SFF_3_n1 ;
    wire KeyArray_S01reg_gff_1_SFF_3_QD ;
    wire KeyArray_S01reg_gff_1_SFF_3_MUXInst_Y ;
    wire KeyArray_S01reg_gff_1_SFF_3_MUXInst_X ;
    wire KeyArray_S01reg_gff_1_SFF_4_n2 ;
    wire KeyArray_S01reg_gff_1_SFF_4_n1 ;
    wire KeyArray_S01reg_gff_1_SFF_4_QD ;
    wire KeyArray_S01reg_gff_1_SFF_4_MUXInst_Y ;
    wire KeyArray_S01reg_gff_1_SFF_4_MUXInst_X ;
    wire KeyArray_S01reg_gff_1_SFF_5_n2 ;
    wire KeyArray_S01reg_gff_1_SFF_5_n1 ;
    wire KeyArray_S01reg_gff_1_SFF_5_QD ;
    wire KeyArray_S01reg_gff_1_SFF_5_MUXInst_Y ;
    wire KeyArray_S01reg_gff_1_SFF_5_MUXInst_X ;
    wire KeyArray_S01reg_gff_1_SFF_6_n2 ;
    wire KeyArray_S01reg_gff_1_SFF_6_n1 ;
    wire KeyArray_S01reg_gff_1_SFF_6_QD ;
    wire KeyArray_S01reg_gff_1_SFF_6_MUXInst_Y ;
    wire KeyArray_S01reg_gff_1_SFF_6_MUXInst_X ;
    wire KeyArray_S01reg_gff_1_SFF_7_n2 ;
    wire KeyArray_S01reg_gff_1_SFF_7_n1 ;
    wire KeyArray_S01reg_gff_1_SFF_7_QD ;
    wire KeyArray_S01reg_gff_1_SFF_7_MUXInst_Y ;
    wire KeyArray_S01reg_gff_1_SFF_7_MUXInst_X ;
    wire KeyArray_S02reg_gff_1_SFF_0_n2 ;
    wire KeyArray_S02reg_gff_1_SFF_0_n1 ;
    wire KeyArray_S02reg_gff_1_SFF_0_QD ;
    wire KeyArray_S02reg_gff_1_SFF_0_MUXInst_Y ;
    wire KeyArray_S02reg_gff_1_SFF_0_MUXInst_X ;
    wire KeyArray_S02reg_gff_1_SFF_1_n2 ;
    wire KeyArray_S02reg_gff_1_SFF_1_n1 ;
    wire KeyArray_S02reg_gff_1_SFF_1_QD ;
    wire KeyArray_S02reg_gff_1_SFF_1_MUXInst_Y ;
    wire KeyArray_S02reg_gff_1_SFF_1_MUXInst_X ;
    wire KeyArray_S02reg_gff_1_SFF_2_n2 ;
    wire KeyArray_S02reg_gff_1_SFF_2_n1 ;
    wire KeyArray_S02reg_gff_1_SFF_2_QD ;
    wire KeyArray_S02reg_gff_1_SFF_2_MUXInst_Y ;
    wire KeyArray_S02reg_gff_1_SFF_2_MUXInst_X ;
    wire KeyArray_S02reg_gff_1_SFF_3_n2 ;
    wire KeyArray_S02reg_gff_1_SFF_3_n1 ;
    wire KeyArray_S02reg_gff_1_SFF_3_QD ;
    wire KeyArray_S02reg_gff_1_SFF_3_MUXInst_Y ;
    wire KeyArray_S02reg_gff_1_SFF_3_MUXInst_X ;
    wire KeyArray_S02reg_gff_1_SFF_4_n2 ;
    wire KeyArray_S02reg_gff_1_SFF_4_n1 ;
    wire KeyArray_S02reg_gff_1_SFF_4_QD ;
    wire KeyArray_S02reg_gff_1_SFF_4_MUXInst_Y ;
    wire KeyArray_S02reg_gff_1_SFF_4_MUXInst_X ;
    wire KeyArray_S02reg_gff_1_SFF_5_n2 ;
    wire KeyArray_S02reg_gff_1_SFF_5_n1 ;
    wire KeyArray_S02reg_gff_1_SFF_5_QD ;
    wire KeyArray_S02reg_gff_1_SFF_5_MUXInst_Y ;
    wire KeyArray_S02reg_gff_1_SFF_5_MUXInst_X ;
    wire KeyArray_S02reg_gff_1_SFF_6_n2 ;
    wire KeyArray_S02reg_gff_1_SFF_6_n1 ;
    wire KeyArray_S02reg_gff_1_SFF_6_QD ;
    wire KeyArray_S02reg_gff_1_SFF_6_MUXInst_Y ;
    wire KeyArray_S02reg_gff_1_SFF_6_MUXInst_X ;
    wire KeyArray_S02reg_gff_1_SFF_7_n2 ;
    wire KeyArray_S02reg_gff_1_SFF_7_n1 ;
    wire KeyArray_S02reg_gff_1_SFF_7_QD ;
    wire KeyArray_S02reg_gff_1_SFF_7_MUXInst_Y ;
    wire KeyArray_S02reg_gff_1_SFF_7_MUXInst_X ;
    wire KeyArray_S03reg_gff_1_SFF_0_n2 ;
    wire KeyArray_S03reg_gff_1_SFF_0_n1 ;
    wire KeyArray_S03reg_gff_1_SFF_0_QD ;
    wire KeyArray_S03reg_gff_1_SFF_0_MUXInst_Y ;
    wire KeyArray_S03reg_gff_1_SFF_0_MUXInst_X ;
    wire KeyArray_S03reg_gff_1_SFF_1_n2 ;
    wire KeyArray_S03reg_gff_1_SFF_1_n1 ;
    wire KeyArray_S03reg_gff_1_SFF_1_QD ;
    wire KeyArray_S03reg_gff_1_SFF_1_MUXInst_Y ;
    wire KeyArray_S03reg_gff_1_SFF_1_MUXInst_X ;
    wire KeyArray_S03reg_gff_1_SFF_2_n2 ;
    wire KeyArray_S03reg_gff_1_SFF_2_n1 ;
    wire KeyArray_S03reg_gff_1_SFF_2_QD ;
    wire KeyArray_S03reg_gff_1_SFF_2_MUXInst_Y ;
    wire KeyArray_S03reg_gff_1_SFF_2_MUXInst_X ;
    wire KeyArray_S03reg_gff_1_SFF_3_n2 ;
    wire KeyArray_S03reg_gff_1_SFF_3_n1 ;
    wire KeyArray_S03reg_gff_1_SFF_3_QD ;
    wire KeyArray_S03reg_gff_1_SFF_3_MUXInst_Y ;
    wire KeyArray_S03reg_gff_1_SFF_3_MUXInst_X ;
    wire KeyArray_S03reg_gff_1_SFF_4_n2 ;
    wire KeyArray_S03reg_gff_1_SFF_4_n1 ;
    wire KeyArray_S03reg_gff_1_SFF_4_QD ;
    wire KeyArray_S03reg_gff_1_SFF_4_MUXInst_Y ;
    wire KeyArray_S03reg_gff_1_SFF_4_MUXInst_X ;
    wire KeyArray_S03reg_gff_1_SFF_5_n2 ;
    wire KeyArray_S03reg_gff_1_SFF_5_n1 ;
    wire KeyArray_S03reg_gff_1_SFF_5_QD ;
    wire KeyArray_S03reg_gff_1_SFF_5_MUXInst_Y ;
    wire KeyArray_S03reg_gff_1_SFF_5_MUXInst_X ;
    wire KeyArray_S03reg_gff_1_SFF_6_n2 ;
    wire KeyArray_S03reg_gff_1_SFF_6_n1 ;
    wire KeyArray_S03reg_gff_1_SFF_6_QD ;
    wire KeyArray_S03reg_gff_1_SFF_6_MUXInst_Y ;
    wire KeyArray_S03reg_gff_1_SFF_6_MUXInst_X ;
    wire KeyArray_S03reg_gff_1_SFF_7_n2 ;
    wire KeyArray_S03reg_gff_1_SFF_7_n1 ;
    wire KeyArray_S03reg_gff_1_SFF_7_QD ;
    wire KeyArray_S03reg_gff_1_SFF_7_MUXInst_Y ;
    wire KeyArray_S03reg_gff_1_SFF_7_MUXInst_X ;
    wire KeyArray_S10reg_gff_1_SFF_0_n2 ;
    wire KeyArray_S10reg_gff_1_SFF_0_n1 ;
    wire KeyArray_S10reg_gff_1_SFF_0_QD ;
    wire KeyArray_S10reg_gff_1_SFF_0_MUXInst_Y ;
    wire KeyArray_S10reg_gff_1_SFF_0_MUXInst_X ;
    wire KeyArray_S10reg_gff_1_SFF_1_n2 ;
    wire KeyArray_S10reg_gff_1_SFF_1_n1 ;
    wire KeyArray_S10reg_gff_1_SFF_1_QD ;
    wire KeyArray_S10reg_gff_1_SFF_1_MUXInst_Y ;
    wire KeyArray_S10reg_gff_1_SFF_1_MUXInst_X ;
    wire KeyArray_S10reg_gff_1_SFF_2_n2 ;
    wire KeyArray_S10reg_gff_1_SFF_2_n1 ;
    wire KeyArray_S10reg_gff_1_SFF_2_QD ;
    wire KeyArray_S10reg_gff_1_SFF_2_MUXInst_Y ;
    wire KeyArray_S10reg_gff_1_SFF_2_MUXInst_X ;
    wire KeyArray_S10reg_gff_1_SFF_3_n2 ;
    wire KeyArray_S10reg_gff_1_SFF_3_n1 ;
    wire KeyArray_S10reg_gff_1_SFF_3_QD ;
    wire KeyArray_S10reg_gff_1_SFF_3_MUXInst_Y ;
    wire KeyArray_S10reg_gff_1_SFF_3_MUXInst_X ;
    wire KeyArray_S10reg_gff_1_SFF_4_n2 ;
    wire KeyArray_S10reg_gff_1_SFF_4_n1 ;
    wire KeyArray_S10reg_gff_1_SFF_4_QD ;
    wire KeyArray_S10reg_gff_1_SFF_4_MUXInst_Y ;
    wire KeyArray_S10reg_gff_1_SFF_4_MUXInst_X ;
    wire KeyArray_S10reg_gff_1_SFF_5_n2 ;
    wire KeyArray_S10reg_gff_1_SFF_5_n1 ;
    wire KeyArray_S10reg_gff_1_SFF_5_QD ;
    wire KeyArray_S10reg_gff_1_SFF_5_MUXInst_Y ;
    wire KeyArray_S10reg_gff_1_SFF_5_MUXInst_X ;
    wire KeyArray_S10reg_gff_1_SFF_6_n2 ;
    wire KeyArray_S10reg_gff_1_SFF_6_n1 ;
    wire KeyArray_S10reg_gff_1_SFF_6_QD ;
    wire KeyArray_S10reg_gff_1_SFF_6_MUXInst_Y ;
    wire KeyArray_S10reg_gff_1_SFF_6_MUXInst_X ;
    wire KeyArray_S10reg_gff_1_SFF_7_n2 ;
    wire KeyArray_S10reg_gff_1_SFF_7_n1 ;
    wire KeyArray_S10reg_gff_1_SFF_7_QD ;
    wire KeyArray_S10reg_gff_1_SFF_7_MUXInst_Y ;
    wire KeyArray_S10reg_gff_1_SFF_7_MUXInst_X ;
    wire KeyArray_S11reg_gff_1_SFF_0_n2 ;
    wire KeyArray_S11reg_gff_1_SFF_0_n1 ;
    wire KeyArray_S11reg_gff_1_SFF_0_QD ;
    wire KeyArray_S11reg_gff_1_SFF_0_MUXInst_Y ;
    wire KeyArray_S11reg_gff_1_SFF_0_MUXInst_X ;
    wire KeyArray_S11reg_gff_1_SFF_1_n2 ;
    wire KeyArray_S11reg_gff_1_SFF_1_n1 ;
    wire KeyArray_S11reg_gff_1_SFF_1_QD ;
    wire KeyArray_S11reg_gff_1_SFF_1_MUXInst_Y ;
    wire KeyArray_S11reg_gff_1_SFF_1_MUXInst_X ;
    wire KeyArray_S11reg_gff_1_SFF_2_n2 ;
    wire KeyArray_S11reg_gff_1_SFF_2_n1 ;
    wire KeyArray_S11reg_gff_1_SFF_2_QD ;
    wire KeyArray_S11reg_gff_1_SFF_2_MUXInst_Y ;
    wire KeyArray_S11reg_gff_1_SFF_2_MUXInst_X ;
    wire KeyArray_S11reg_gff_1_SFF_3_n2 ;
    wire KeyArray_S11reg_gff_1_SFF_3_n1 ;
    wire KeyArray_S11reg_gff_1_SFF_3_QD ;
    wire KeyArray_S11reg_gff_1_SFF_3_MUXInst_Y ;
    wire KeyArray_S11reg_gff_1_SFF_3_MUXInst_X ;
    wire KeyArray_S11reg_gff_1_SFF_4_n2 ;
    wire KeyArray_S11reg_gff_1_SFF_4_n1 ;
    wire KeyArray_S11reg_gff_1_SFF_4_QD ;
    wire KeyArray_S11reg_gff_1_SFF_4_MUXInst_Y ;
    wire KeyArray_S11reg_gff_1_SFF_4_MUXInst_X ;
    wire KeyArray_S11reg_gff_1_SFF_5_n2 ;
    wire KeyArray_S11reg_gff_1_SFF_5_n1 ;
    wire KeyArray_S11reg_gff_1_SFF_5_QD ;
    wire KeyArray_S11reg_gff_1_SFF_5_MUXInst_Y ;
    wire KeyArray_S11reg_gff_1_SFF_5_MUXInst_X ;
    wire KeyArray_S11reg_gff_1_SFF_6_n2 ;
    wire KeyArray_S11reg_gff_1_SFF_6_n1 ;
    wire KeyArray_S11reg_gff_1_SFF_6_QD ;
    wire KeyArray_S11reg_gff_1_SFF_6_MUXInst_Y ;
    wire KeyArray_S11reg_gff_1_SFF_6_MUXInst_X ;
    wire KeyArray_S11reg_gff_1_SFF_7_n2 ;
    wire KeyArray_S11reg_gff_1_SFF_7_n1 ;
    wire KeyArray_S11reg_gff_1_SFF_7_QD ;
    wire KeyArray_S11reg_gff_1_SFF_7_MUXInst_Y ;
    wire KeyArray_S11reg_gff_1_SFF_7_MUXInst_X ;
    wire KeyArray_S12reg_gff_1_SFF_0_n2 ;
    wire KeyArray_S12reg_gff_1_SFF_0_n1 ;
    wire KeyArray_S12reg_gff_1_SFF_0_QD ;
    wire KeyArray_S12reg_gff_1_SFF_0_MUXInst_Y ;
    wire KeyArray_S12reg_gff_1_SFF_0_MUXInst_X ;
    wire KeyArray_S12reg_gff_1_SFF_1_n2 ;
    wire KeyArray_S12reg_gff_1_SFF_1_n1 ;
    wire KeyArray_S12reg_gff_1_SFF_1_QD ;
    wire KeyArray_S12reg_gff_1_SFF_1_MUXInst_Y ;
    wire KeyArray_S12reg_gff_1_SFF_1_MUXInst_X ;
    wire KeyArray_S12reg_gff_1_SFF_2_n2 ;
    wire KeyArray_S12reg_gff_1_SFF_2_n1 ;
    wire KeyArray_S12reg_gff_1_SFF_2_QD ;
    wire KeyArray_S12reg_gff_1_SFF_2_MUXInst_Y ;
    wire KeyArray_S12reg_gff_1_SFF_2_MUXInst_X ;
    wire KeyArray_S12reg_gff_1_SFF_3_n2 ;
    wire KeyArray_S12reg_gff_1_SFF_3_n1 ;
    wire KeyArray_S12reg_gff_1_SFF_3_QD ;
    wire KeyArray_S12reg_gff_1_SFF_3_MUXInst_Y ;
    wire KeyArray_S12reg_gff_1_SFF_3_MUXInst_X ;
    wire KeyArray_S12reg_gff_1_SFF_4_n2 ;
    wire KeyArray_S12reg_gff_1_SFF_4_n1 ;
    wire KeyArray_S12reg_gff_1_SFF_4_QD ;
    wire KeyArray_S12reg_gff_1_SFF_4_MUXInst_Y ;
    wire KeyArray_S12reg_gff_1_SFF_4_MUXInst_X ;
    wire KeyArray_S12reg_gff_1_SFF_5_n2 ;
    wire KeyArray_S12reg_gff_1_SFF_5_n1 ;
    wire KeyArray_S12reg_gff_1_SFF_5_QD ;
    wire KeyArray_S12reg_gff_1_SFF_5_MUXInst_Y ;
    wire KeyArray_S12reg_gff_1_SFF_5_MUXInst_X ;
    wire KeyArray_S12reg_gff_1_SFF_6_n2 ;
    wire KeyArray_S12reg_gff_1_SFF_6_n1 ;
    wire KeyArray_S12reg_gff_1_SFF_6_QD ;
    wire KeyArray_S12reg_gff_1_SFF_6_MUXInst_Y ;
    wire KeyArray_S12reg_gff_1_SFF_6_MUXInst_X ;
    wire KeyArray_S12reg_gff_1_SFF_7_n2 ;
    wire KeyArray_S12reg_gff_1_SFF_7_n1 ;
    wire KeyArray_S12reg_gff_1_SFF_7_QD ;
    wire KeyArray_S12reg_gff_1_SFF_7_MUXInst_Y ;
    wire KeyArray_S12reg_gff_1_SFF_7_MUXInst_X ;
    wire KeyArray_S13reg_gff_1_SFF_0_n2 ;
    wire KeyArray_S13reg_gff_1_SFF_0_n1 ;
    wire KeyArray_S13reg_gff_1_SFF_0_QD ;
    wire KeyArray_S13reg_gff_1_SFF_0_MUXInst_Y ;
    wire KeyArray_S13reg_gff_1_SFF_0_MUXInst_X ;
    wire KeyArray_S13reg_gff_1_SFF_1_n2 ;
    wire KeyArray_S13reg_gff_1_SFF_1_n1 ;
    wire KeyArray_S13reg_gff_1_SFF_1_QD ;
    wire KeyArray_S13reg_gff_1_SFF_1_MUXInst_Y ;
    wire KeyArray_S13reg_gff_1_SFF_1_MUXInst_X ;
    wire KeyArray_S13reg_gff_1_SFF_2_n2 ;
    wire KeyArray_S13reg_gff_1_SFF_2_n1 ;
    wire KeyArray_S13reg_gff_1_SFF_2_QD ;
    wire KeyArray_S13reg_gff_1_SFF_2_MUXInst_Y ;
    wire KeyArray_S13reg_gff_1_SFF_2_MUXInst_X ;
    wire KeyArray_S13reg_gff_1_SFF_3_n2 ;
    wire KeyArray_S13reg_gff_1_SFF_3_n1 ;
    wire KeyArray_S13reg_gff_1_SFF_3_QD ;
    wire KeyArray_S13reg_gff_1_SFF_3_MUXInst_Y ;
    wire KeyArray_S13reg_gff_1_SFF_3_MUXInst_X ;
    wire KeyArray_S13reg_gff_1_SFF_4_n2 ;
    wire KeyArray_S13reg_gff_1_SFF_4_n1 ;
    wire KeyArray_S13reg_gff_1_SFF_4_QD ;
    wire KeyArray_S13reg_gff_1_SFF_4_MUXInst_Y ;
    wire KeyArray_S13reg_gff_1_SFF_4_MUXInst_X ;
    wire KeyArray_S13reg_gff_1_SFF_5_n2 ;
    wire KeyArray_S13reg_gff_1_SFF_5_n1 ;
    wire KeyArray_S13reg_gff_1_SFF_5_QD ;
    wire KeyArray_S13reg_gff_1_SFF_5_MUXInst_Y ;
    wire KeyArray_S13reg_gff_1_SFF_5_MUXInst_X ;
    wire KeyArray_S13reg_gff_1_SFF_6_n2 ;
    wire KeyArray_S13reg_gff_1_SFF_6_n1 ;
    wire KeyArray_S13reg_gff_1_SFF_6_QD ;
    wire KeyArray_S13reg_gff_1_SFF_6_MUXInst_Y ;
    wire KeyArray_S13reg_gff_1_SFF_6_MUXInst_X ;
    wire KeyArray_S13reg_gff_1_SFF_7_n2 ;
    wire KeyArray_S13reg_gff_1_SFF_7_n1 ;
    wire KeyArray_S13reg_gff_1_SFF_7_QD ;
    wire KeyArray_S13reg_gff_1_SFF_7_MUXInst_Y ;
    wire KeyArray_S13reg_gff_1_SFF_7_MUXInst_X ;
    wire KeyArray_S20reg_gff_1_SFF_0_n2 ;
    wire KeyArray_S20reg_gff_1_SFF_0_n1 ;
    wire KeyArray_S20reg_gff_1_SFF_0_QD ;
    wire KeyArray_S20reg_gff_1_SFF_0_MUXInst_Y ;
    wire KeyArray_S20reg_gff_1_SFF_0_MUXInst_X ;
    wire KeyArray_S20reg_gff_1_SFF_1_n2 ;
    wire KeyArray_S20reg_gff_1_SFF_1_n1 ;
    wire KeyArray_S20reg_gff_1_SFF_1_QD ;
    wire KeyArray_S20reg_gff_1_SFF_1_MUXInst_Y ;
    wire KeyArray_S20reg_gff_1_SFF_1_MUXInst_X ;
    wire KeyArray_S20reg_gff_1_SFF_2_n2 ;
    wire KeyArray_S20reg_gff_1_SFF_2_n1 ;
    wire KeyArray_S20reg_gff_1_SFF_2_QD ;
    wire KeyArray_S20reg_gff_1_SFF_2_MUXInst_Y ;
    wire KeyArray_S20reg_gff_1_SFF_2_MUXInst_X ;
    wire KeyArray_S20reg_gff_1_SFF_3_n2 ;
    wire KeyArray_S20reg_gff_1_SFF_3_n1 ;
    wire KeyArray_S20reg_gff_1_SFF_3_QD ;
    wire KeyArray_S20reg_gff_1_SFF_3_MUXInst_Y ;
    wire KeyArray_S20reg_gff_1_SFF_3_MUXInst_X ;
    wire KeyArray_S20reg_gff_1_SFF_4_n2 ;
    wire KeyArray_S20reg_gff_1_SFF_4_n1 ;
    wire KeyArray_S20reg_gff_1_SFF_4_QD ;
    wire KeyArray_S20reg_gff_1_SFF_4_MUXInst_Y ;
    wire KeyArray_S20reg_gff_1_SFF_4_MUXInst_X ;
    wire KeyArray_S20reg_gff_1_SFF_5_n2 ;
    wire KeyArray_S20reg_gff_1_SFF_5_n1 ;
    wire KeyArray_S20reg_gff_1_SFF_5_QD ;
    wire KeyArray_S20reg_gff_1_SFF_5_MUXInst_Y ;
    wire KeyArray_S20reg_gff_1_SFF_5_MUXInst_X ;
    wire KeyArray_S20reg_gff_1_SFF_6_n2 ;
    wire KeyArray_S20reg_gff_1_SFF_6_n1 ;
    wire KeyArray_S20reg_gff_1_SFF_6_QD ;
    wire KeyArray_S20reg_gff_1_SFF_6_MUXInst_Y ;
    wire KeyArray_S20reg_gff_1_SFF_6_MUXInst_X ;
    wire KeyArray_S20reg_gff_1_SFF_7_n2 ;
    wire KeyArray_S20reg_gff_1_SFF_7_n1 ;
    wire KeyArray_S20reg_gff_1_SFF_7_QD ;
    wire KeyArray_S20reg_gff_1_SFF_7_MUXInst_Y ;
    wire KeyArray_S20reg_gff_1_SFF_7_MUXInst_X ;
    wire KeyArray_S21reg_gff_1_SFF_0_n2 ;
    wire KeyArray_S21reg_gff_1_SFF_0_n1 ;
    wire KeyArray_S21reg_gff_1_SFF_0_QD ;
    wire KeyArray_S21reg_gff_1_SFF_0_MUXInst_Y ;
    wire KeyArray_S21reg_gff_1_SFF_0_MUXInst_X ;
    wire KeyArray_S21reg_gff_1_SFF_1_n2 ;
    wire KeyArray_S21reg_gff_1_SFF_1_n1 ;
    wire KeyArray_S21reg_gff_1_SFF_1_QD ;
    wire KeyArray_S21reg_gff_1_SFF_1_MUXInst_Y ;
    wire KeyArray_S21reg_gff_1_SFF_1_MUXInst_X ;
    wire KeyArray_S21reg_gff_1_SFF_2_n2 ;
    wire KeyArray_S21reg_gff_1_SFF_2_n1 ;
    wire KeyArray_S21reg_gff_1_SFF_2_QD ;
    wire KeyArray_S21reg_gff_1_SFF_2_MUXInst_Y ;
    wire KeyArray_S21reg_gff_1_SFF_2_MUXInst_X ;
    wire KeyArray_S21reg_gff_1_SFF_3_n2 ;
    wire KeyArray_S21reg_gff_1_SFF_3_n1 ;
    wire KeyArray_S21reg_gff_1_SFF_3_QD ;
    wire KeyArray_S21reg_gff_1_SFF_3_MUXInst_Y ;
    wire KeyArray_S21reg_gff_1_SFF_3_MUXInst_X ;
    wire KeyArray_S21reg_gff_1_SFF_4_n2 ;
    wire KeyArray_S21reg_gff_1_SFF_4_n1 ;
    wire KeyArray_S21reg_gff_1_SFF_4_QD ;
    wire KeyArray_S21reg_gff_1_SFF_4_MUXInst_Y ;
    wire KeyArray_S21reg_gff_1_SFF_4_MUXInst_X ;
    wire KeyArray_S21reg_gff_1_SFF_5_n2 ;
    wire KeyArray_S21reg_gff_1_SFF_5_n1 ;
    wire KeyArray_S21reg_gff_1_SFF_5_QD ;
    wire KeyArray_S21reg_gff_1_SFF_5_MUXInst_Y ;
    wire KeyArray_S21reg_gff_1_SFF_5_MUXInst_X ;
    wire KeyArray_S21reg_gff_1_SFF_6_n2 ;
    wire KeyArray_S21reg_gff_1_SFF_6_n1 ;
    wire KeyArray_S21reg_gff_1_SFF_6_QD ;
    wire KeyArray_S21reg_gff_1_SFF_6_MUXInst_Y ;
    wire KeyArray_S21reg_gff_1_SFF_6_MUXInst_X ;
    wire KeyArray_S21reg_gff_1_SFF_7_n2 ;
    wire KeyArray_S21reg_gff_1_SFF_7_n1 ;
    wire KeyArray_S21reg_gff_1_SFF_7_QD ;
    wire KeyArray_S21reg_gff_1_SFF_7_MUXInst_Y ;
    wire KeyArray_S21reg_gff_1_SFF_7_MUXInst_X ;
    wire KeyArray_S22reg_gff_1_SFF_0_n2 ;
    wire KeyArray_S22reg_gff_1_SFF_0_n1 ;
    wire KeyArray_S22reg_gff_1_SFF_0_QD ;
    wire KeyArray_S22reg_gff_1_SFF_0_MUXInst_Y ;
    wire KeyArray_S22reg_gff_1_SFF_0_MUXInst_X ;
    wire KeyArray_S22reg_gff_1_SFF_1_n2 ;
    wire KeyArray_S22reg_gff_1_SFF_1_n1 ;
    wire KeyArray_S22reg_gff_1_SFF_1_QD ;
    wire KeyArray_S22reg_gff_1_SFF_1_MUXInst_Y ;
    wire KeyArray_S22reg_gff_1_SFF_1_MUXInst_X ;
    wire KeyArray_S22reg_gff_1_SFF_2_n2 ;
    wire KeyArray_S22reg_gff_1_SFF_2_n1 ;
    wire KeyArray_S22reg_gff_1_SFF_2_QD ;
    wire KeyArray_S22reg_gff_1_SFF_2_MUXInst_Y ;
    wire KeyArray_S22reg_gff_1_SFF_2_MUXInst_X ;
    wire KeyArray_S22reg_gff_1_SFF_3_n2 ;
    wire KeyArray_S22reg_gff_1_SFF_3_n1 ;
    wire KeyArray_S22reg_gff_1_SFF_3_QD ;
    wire KeyArray_S22reg_gff_1_SFF_3_MUXInst_Y ;
    wire KeyArray_S22reg_gff_1_SFF_3_MUXInst_X ;
    wire KeyArray_S22reg_gff_1_SFF_4_n2 ;
    wire KeyArray_S22reg_gff_1_SFF_4_n1 ;
    wire KeyArray_S22reg_gff_1_SFF_4_QD ;
    wire KeyArray_S22reg_gff_1_SFF_4_MUXInst_Y ;
    wire KeyArray_S22reg_gff_1_SFF_4_MUXInst_X ;
    wire KeyArray_S22reg_gff_1_SFF_5_n2 ;
    wire KeyArray_S22reg_gff_1_SFF_5_n1 ;
    wire KeyArray_S22reg_gff_1_SFF_5_QD ;
    wire KeyArray_S22reg_gff_1_SFF_5_MUXInst_Y ;
    wire KeyArray_S22reg_gff_1_SFF_5_MUXInst_X ;
    wire KeyArray_S22reg_gff_1_SFF_6_n2 ;
    wire KeyArray_S22reg_gff_1_SFF_6_n1 ;
    wire KeyArray_S22reg_gff_1_SFF_6_QD ;
    wire KeyArray_S22reg_gff_1_SFF_6_MUXInst_Y ;
    wire KeyArray_S22reg_gff_1_SFF_6_MUXInst_X ;
    wire KeyArray_S22reg_gff_1_SFF_7_n2 ;
    wire KeyArray_S22reg_gff_1_SFF_7_n1 ;
    wire KeyArray_S22reg_gff_1_SFF_7_QD ;
    wire KeyArray_S22reg_gff_1_SFF_7_MUXInst_Y ;
    wire KeyArray_S22reg_gff_1_SFF_7_MUXInst_X ;
    wire KeyArray_S23reg_gff_1_SFF_0_n2 ;
    wire KeyArray_S23reg_gff_1_SFF_0_n1 ;
    wire KeyArray_S23reg_gff_1_SFF_0_QD ;
    wire KeyArray_S23reg_gff_1_SFF_0_MUXInst_Y ;
    wire KeyArray_S23reg_gff_1_SFF_0_MUXInst_X ;
    wire KeyArray_S23reg_gff_1_SFF_1_n2 ;
    wire KeyArray_S23reg_gff_1_SFF_1_n1 ;
    wire KeyArray_S23reg_gff_1_SFF_1_QD ;
    wire KeyArray_S23reg_gff_1_SFF_1_MUXInst_Y ;
    wire KeyArray_S23reg_gff_1_SFF_1_MUXInst_X ;
    wire KeyArray_S23reg_gff_1_SFF_2_n2 ;
    wire KeyArray_S23reg_gff_1_SFF_2_n1 ;
    wire KeyArray_S23reg_gff_1_SFF_2_QD ;
    wire KeyArray_S23reg_gff_1_SFF_2_MUXInst_Y ;
    wire KeyArray_S23reg_gff_1_SFF_2_MUXInst_X ;
    wire KeyArray_S23reg_gff_1_SFF_3_n2 ;
    wire KeyArray_S23reg_gff_1_SFF_3_n1 ;
    wire KeyArray_S23reg_gff_1_SFF_3_QD ;
    wire KeyArray_S23reg_gff_1_SFF_3_MUXInst_Y ;
    wire KeyArray_S23reg_gff_1_SFF_3_MUXInst_X ;
    wire KeyArray_S23reg_gff_1_SFF_4_n2 ;
    wire KeyArray_S23reg_gff_1_SFF_4_n1 ;
    wire KeyArray_S23reg_gff_1_SFF_4_QD ;
    wire KeyArray_S23reg_gff_1_SFF_4_MUXInst_Y ;
    wire KeyArray_S23reg_gff_1_SFF_4_MUXInst_X ;
    wire KeyArray_S23reg_gff_1_SFF_5_n2 ;
    wire KeyArray_S23reg_gff_1_SFF_5_n1 ;
    wire KeyArray_S23reg_gff_1_SFF_5_QD ;
    wire KeyArray_S23reg_gff_1_SFF_5_MUXInst_Y ;
    wire KeyArray_S23reg_gff_1_SFF_5_MUXInst_X ;
    wire KeyArray_S23reg_gff_1_SFF_6_n2 ;
    wire KeyArray_S23reg_gff_1_SFF_6_n1 ;
    wire KeyArray_S23reg_gff_1_SFF_6_QD ;
    wire KeyArray_S23reg_gff_1_SFF_6_MUXInst_Y ;
    wire KeyArray_S23reg_gff_1_SFF_6_MUXInst_X ;
    wire KeyArray_S23reg_gff_1_SFF_7_n2 ;
    wire KeyArray_S23reg_gff_1_SFF_7_n1 ;
    wire KeyArray_S23reg_gff_1_SFF_7_QD ;
    wire KeyArray_S23reg_gff_1_SFF_7_MUXInst_Y ;
    wire KeyArray_S23reg_gff_1_SFF_7_MUXInst_X ;
    wire KeyArray_S30reg_gff_1_SFF_0_n2 ;
    wire KeyArray_S30reg_gff_1_SFF_0_n1 ;
    wire KeyArray_S30reg_gff_1_SFF_0_QD ;
    wire KeyArray_S30reg_gff_1_SFF_0_MUXInst_Y ;
    wire KeyArray_S30reg_gff_1_SFF_0_MUXInst_X ;
    wire KeyArray_S30reg_gff_1_SFF_1_n2 ;
    wire KeyArray_S30reg_gff_1_SFF_1_n1 ;
    wire KeyArray_S30reg_gff_1_SFF_1_QD ;
    wire KeyArray_S30reg_gff_1_SFF_1_MUXInst_Y ;
    wire KeyArray_S30reg_gff_1_SFF_1_MUXInst_X ;
    wire KeyArray_S30reg_gff_1_SFF_2_n2 ;
    wire KeyArray_S30reg_gff_1_SFF_2_n1 ;
    wire KeyArray_S30reg_gff_1_SFF_2_QD ;
    wire KeyArray_S30reg_gff_1_SFF_2_MUXInst_Y ;
    wire KeyArray_S30reg_gff_1_SFF_2_MUXInst_X ;
    wire KeyArray_S30reg_gff_1_SFF_3_n2 ;
    wire KeyArray_S30reg_gff_1_SFF_3_n1 ;
    wire KeyArray_S30reg_gff_1_SFF_3_QD ;
    wire KeyArray_S30reg_gff_1_SFF_3_MUXInst_Y ;
    wire KeyArray_S30reg_gff_1_SFF_3_MUXInst_X ;
    wire KeyArray_S30reg_gff_1_SFF_4_n2 ;
    wire KeyArray_S30reg_gff_1_SFF_4_n1 ;
    wire KeyArray_S30reg_gff_1_SFF_4_QD ;
    wire KeyArray_S30reg_gff_1_SFF_4_MUXInst_Y ;
    wire KeyArray_S30reg_gff_1_SFF_4_MUXInst_X ;
    wire KeyArray_S30reg_gff_1_SFF_5_n2 ;
    wire KeyArray_S30reg_gff_1_SFF_5_n1 ;
    wire KeyArray_S30reg_gff_1_SFF_5_QD ;
    wire KeyArray_S30reg_gff_1_SFF_5_MUXInst_Y ;
    wire KeyArray_S30reg_gff_1_SFF_5_MUXInst_X ;
    wire KeyArray_S30reg_gff_1_SFF_6_n2 ;
    wire KeyArray_S30reg_gff_1_SFF_6_n1 ;
    wire KeyArray_S30reg_gff_1_SFF_6_QD ;
    wire KeyArray_S30reg_gff_1_SFF_6_MUXInst_Y ;
    wire KeyArray_S30reg_gff_1_SFF_6_MUXInst_X ;
    wire KeyArray_S30reg_gff_1_SFF_7_n2 ;
    wire KeyArray_S30reg_gff_1_SFF_7_n1 ;
    wire KeyArray_S30reg_gff_1_SFF_7_QD ;
    wire KeyArray_S30reg_gff_1_SFF_7_MUXInst_Y ;
    wire KeyArray_S30reg_gff_1_SFF_7_MUXInst_X ;
    wire KeyArray_S31reg_gff_1_SFF_0_n2 ;
    wire KeyArray_S31reg_gff_1_SFF_0_n1 ;
    wire KeyArray_S31reg_gff_1_SFF_0_QD ;
    wire KeyArray_S31reg_gff_1_SFF_0_MUXInst_Y ;
    wire KeyArray_S31reg_gff_1_SFF_0_MUXInst_X ;
    wire KeyArray_S31reg_gff_1_SFF_1_n2 ;
    wire KeyArray_S31reg_gff_1_SFF_1_n1 ;
    wire KeyArray_S31reg_gff_1_SFF_1_QD ;
    wire KeyArray_S31reg_gff_1_SFF_1_MUXInst_Y ;
    wire KeyArray_S31reg_gff_1_SFF_1_MUXInst_X ;
    wire KeyArray_S31reg_gff_1_SFF_2_n2 ;
    wire KeyArray_S31reg_gff_1_SFF_2_n1 ;
    wire KeyArray_S31reg_gff_1_SFF_2_QD ;
    wire KeyArray_S31reg_gff_1_SFF_2_MUXInst_Y ;
    wire KeyArray_S31reg_gff_1_SFF_2_MUXInst_X ;
    wire KeyArray_S31reg_gff_1_SFF_3_n2 ;
    wire KeyArray_S31reg_gff_1_SFF_3_n1 ;
    wire KeyArray_S31reg_gff_1_SFF_3_QD ;
    wire KeyArray_S31reg_gff_1_SFF_3_MUXInst_Y ;
    wire KeyArray_S31reg_gff_1_SFF_3_MUXInst_X ;
    wire KeyArray_S31reg_gff_1_SFF_4_n2 ;
    wire KeyArray_S31reg_gff_1_SFF_4_n1 ;
    wire KeyArray_S31reg_gff_1_SFF_4_QD ;
    wire KeyArray_S31reg_gff_1_SFF_4_MUXInst_Y ;
    wire KeyArray_S31reg_gff_1_SFF_4_MUXInst_X ;
    wire KeyArray_S31reg_gff_1_SFF_5_n2 ;
    wire KeyArray_S31reg_gff_1_SFF_5_n1 ;
    wire KeyArray_S31reg_gff_1_SFF_5_QD ;
    wire KeyArray_S31reg_gff_1_SFF_5_MUXInst_Y ;
    wire KeyArray_S31reg_gff_1_SFF_5_MUXInst_X ;
    wire KeyArray_S31reg_gff_1_SFF_6_n2 ;
    wire KeyArray_S31reg_gff_1_SFF_6_n1 ;
    wire KeyArray_S31reg_gff_1_SFF_6_QD ;
    wire KeyArray_S31reg_gff_1_SFF_6_MUXInst_Y ;
    wire KeyArray_S31reg_gff_1_SFF_6_MUXInst_X ;
    wire KeyArray_S31reg_gff_1_SFF_7_n2 ;
    wire KeyArray_S31reg_gff_1_SFF_7_n1 ;
    wire KeyArray_S31reg_gff_1_SFF_7_QD ;
    wire KeyArray_S31reg_gff_1_SFF_7_MUXInst_Y ;
    wire KeyArray_S31reg_gff_1_SFF_7_MUXInst_X ;
    wire KeyArray_S32reg_gff_1_SFF_0_n2 ;
    wire KeyArray_S32reg_gff_1_SFF_0_n1 ;
    wire KeyArray_S32reg_gff_1_SFF_0_QD ;
    wire KeyArray_S32reg_gff_1_SFF_0_MUXInst_Y ;
    wire KeyArray_S32reg_gff_1_SFF_0_MUXInst_X ;
    wire KeyArray_S32reg_gff_1_SFF_1_n2 ;
    wire KeyArray_S32reg_gff_1_SFF_1_n1 ;
    wire KeyArray_S32reg_gff_1_SFF_1_QD ;
    wire KeyArray_S32reg_gff_1_SFF_1_MUXInst_Y ;
    wire KeyArray_S32reg_gff_1_SFF_1_MUXInst_X ;
    wire KeyArray_S32reg_gff_1_SFF_2_n2 ;
    wire KeyArray_S32reg_gff_1_SFF_2_n1 ;
    wire KeyArray_S32reg_gff_1_SFF_2_QD ;
    wire KeyArray_S32reg_gff_1_SFF_2_MUXInst_Y ;
    wire KeyArray_S32reg_gff_1_SFF_2_MUXInst_X ;
    wire KeyArray_S32reg_gff_1_SFF_3_n2 ;
    wire KeyArray_S32reg_gff_1_SFF_3_n1 ;
    wire KeyArray_S32reg_gff_1_SFF_3_QD ;
    wire KeyArray_S32reg_gff_1_SFF_3_MUXInst_Y ;
    wire KeyArray_S32reg_gff_1_SFF_3_MUXInst_X ;
    wire KeyArray_S32reg_gff_1_SFF_4_n2 ;
    wire KeyArray_S32reg_gff_1_SFF_4_n1 ;
    wire KeyArray_S32reg_gff_1_SFF_4_QD ;
    wire KeyArray_S32reg_gff_1_SFF_4_MUXInst_Y ;
    wire KeyArray_S32reg_gff_1_SFF_4_MUXInst_X ;
    wire KeyArray_S32reg_gff_1_SFF_5_n2 ;
    wire KeyArray_S32reg_gff_1_SFF_5_n1 ;
    wire KeyArray_S32reg_gff_1_SFF_5_QD ;
    wire KeyArray_S32reg_gff_1_SFF_5_MUXInst_Y ;
    wire KeyArray_S32reg_gff_1_SFF_5_MUXInst_X ;
    wire KeyArray_S32reg_gff_1_SFF_6_n2 ;
    wire KeyArray_S32reg_gff_1_SFF_6_n1 ;
    wire KeyArray_S32reg_gff_1_SFF_6_QD ;
    wire KeyArray_S32reg_gff_1_SFF_6_MUXInst_Y ;
    wire KeyArray_S32reg_gff_1_SFF_6_MUXInst_X ;
    wire KeyArray_S32reg_gff_1_SFF_7_n2 ;
    wire KeyArray_S32reg_gff_1_SFF_7_n1 ;
    wire KeyArray_S32reg_gff_1_SFF_7_QD ;
    wire KeyArray_S32reg_gff_1_SFF_7_MUXInst_Y ;
    wire KeyArray_S32reg_gff_1_SFF_7_MUXInst_X ;
    wire KeyArray_S33reg_gff_1_SFF_0_n2 ;
    wire KeyArray_S33reg_gff_1_SFF_0_n1 ;
    wire KeyArray_S33reg_gff_1_SFF_0_QD ;
    wire KeyArray_S33reg_gff_1_SFF_0_MUXInst_Y ;
    wire KeyArray_S33reg_gff_1_SFF_0_MUXInst_X ;
    wire KeyArray_S33reg_gff_1_SFF_1_n2 ;
    wire KeyArray_S33reg_gff_1_SFF_1_n1 ;
    wire KeyArray_S33reg_gff_1_SFF_1_QD ;
    wire KeyArray_S33reg_gff_1_SFF_1_MUXInst_Y ;
    wire KeyArray_S33reg_gff_1_SFF_1_MUXInst_X ;
    wire KeyArray_S33reg_gff_1_SFF_2_n2 ;
    wire KeyArray_S33reg_gff_1_SFF_2_n1 ;
    wire KeyArray_S33reg_gff_1_SFF_2_QD ;
    wire KeyArray_S33reg_gff_1_SFF_2_MUXInst_Y ;
    wire KeyArray_S33reg_gff_1_SFF_2_MUXInst_X ;
    wire KeyArray_S33reg_gff_1_SFF_3_n2 ;
    wire KeyArray_S33reg_gff_1_SFF_3_n1 ;
    wire KeyArray_S33reg_gff_1_SFF_3_QD ;
    wire KeyArray_S33reg_gff_1_SFF_3_MUXInst_Y ;
    wire KeyArray_S33reg_gff_1_SFF_3_MUXInst_X ;
    wire KeyArray_S33reg_gff_1_SFF_4_n2 ;
    wire KeyArray_S33reg_gff_1_SFF_4_n1 ;
    wire KeyArray_S33reg_gff_1_SFF_4_QD ;
    wire KeyArray_S33reg_gff_1_SFF_4_MUXInst_Y ;
    wire KeyArray_S33reg_gff_1_SFF_4_MUXInst_X ;
    wire KeyArray_S33reg_gff_1_SFF_5_n2 ;
    wire KeyArray_S33reg_gff_1_SFF_5_n1 ;
    wire KeyArray_S33reg_gff_1_SFF_5_QD ;
    wire KeyArray_S33reg_gff_1_SFF_5_MUXInst_Y ;
    wire KeyArray_S33reg_gff_1_SFF_5_MUXInst_X ;
    wire KeyArray_S33reg_gff_1_SFF_6_n2 ;
    wire KeyArray_S33reg_gff_1_SFF_6_n1 ;
    wire KeyArray_S33reg_gff_1_SFF_6_QD ;
    wire KeyArray_S33reg_gff_1_SFF_6_MUXInst_Y ;
    wire KeyArray_S33reg_gff_1_SFF_6_MUXInst_X ;
    wire KeyArray_S33reg_gff_1_SFF_7_n2 ;
    wire KeyArray_S33reg_gff_1_SFF_7_n1 ;
    wire KeyArray_S33reg_gff_1_SFF_7_QD ;
    wire KeyArray_S33reg_gff_1_SFF_7_MUXInst_Y ;
    wire KeyArray_S33reg_gff_1_SFF_7_MUXInst_X ;
    wire KeyArray_MUX_inS00ser_mux_inst_0_Y ;
    wire KeyArray_MUX_inS00ser_mux_inst_0_X ;
    wire KeyArray_MUX_inS00ser_mux_inst_1_Y ;
    wire KeyArray_MUX_inS00ser_mux_inst_1_X ;
    wire KeyArray_MUX_inS00ser_mux_inst_2_Y ;
    wire KeyArray_MUX_inS00ser_mux_inst_2_X ;
    wire KeyArray_MUX_inS00ser_mux_inst_3_Y ;
    wire KeyArray_MUX_inS00ser_mux_inst_3_X ;
    wire KeyArray_MUX_inS00ser_mux_inst_4_Y ;
    wire KeyArray_MUX_inS00ser_mux_inst_4_X ;
    wire KeyArray_MUX_inS00ser_mux_inst_5_Y ;
    wire KeyArray_MUX_inS00ser_mux_inst_5_X ;
    wire KeyArray_MUX_inS00ser_mux_inst_6_Y ;
    wire KeyArray_MUX_inS00ser_mux_inst_6_X ;
    wire KeyArray_MUX_inS00ser_mux_inst_7_Y ;
    wire KeyArray_MUX_inS00ser_mux_inst_7_X ;
    wire KeyArray_MUX_inS33ser_mux_inst_0_Y ;
    wire KeyArray_MUX_inS33ser_mux_inst_0_X ;
    wire KeyArray_MUX_inS33ser_mux_inst_1_Y ;
    wire KeyArray_MUX_inS33ser_mux_inst_1_X ;
    wire KeyArray_MUX_inS33ser_mux_inst_2_Y ;
    wire KeyArray_MUX_inS33ser_mux_inst_2_X ;
    wire KeyArray_MUX_inS33ser_mux_inst_3_Y ;
    wire KeyArray_MUX_inS33ser_mux_inst_3_X ;
    wire KeyArray_MUX_inS33ser_mux_inst_4_Y ;
    wire KeyArray_MUX_inS33ser_mux_inst_4_X ;
    wire KeyArray_MUX_inS33ser_mux_inst_5_Y ;
    wire KeyArray_MUX_inS33ser_mux_inst_5_X ;
    wire KeyArray_MUX_inS33ser_mux_inst_6_Y ;
    wire KeyArray_MUX_inS33ser_mux_inst_6_X ;
    wire KeyArray_MUX_inS33ser_mux_inst_7_Y ;
    wire KeyArray_MUX_inS33ser_mux_inst_7_X ;
    wire MixColumns_line0_n16 ;
    wire MixColumns_line0_n15 ;
    wire MixColumns_line0_n14 ;
    wire MixColumns_line0_n13 ;
    wire MixColumns_line0_n12 ;
    wire MixColumns_line0_n11 ;
    wire MixColumns_line0_n10 ;
    wire MixColumns_line0_n9 ;
    wire MixColumns_line0_n8 ;
    wire MixColumns_line0_n7 ;
    wire MixColumns_line0_n6 ;
    wire MixColumns_line0_n5 ;
    wire MixColumns_line0_n4 ;
    wire MixColumns_line0_n3 ;
    wire MixColumns_line0_n2 ;
    wire MixColumns_line0_n1 ;
    wire MixColumns_line1_n16 ;
    wire MixColumns_line1_n15 ;
    wire MixColumns_line1_n14 ;
    wire MixColumns_line1_n13 ;
    wire MixColumns_line1_n12 ;
    wire MixColumns_line1_n11 ;
    wire MixColumns_line1_n10 ;
    wire MixColumns_line1_n9 ;
    wire MixColumns_line1_n8 ;
    wire MixColumns_line1_n7 ;
    wire MixColumns_line1_n6 ;
    wire MixColumns_line1_n5 ;
    wire MixColumns_line1_n4 ;
    wire MixColumns_line1_n3 ;
    wire MixColumns_line1_n2 ;
    wire MixColumns_line1_n1 ;
    wire MixColumns_line2_n16 ;
    wire MixColumns_line2_n15 ;
    wire MixColumns_line2_n14 ;
    wire MixColumns_line2_n13 ;
    wire MixColumns_line2_n12 ;
    wire MixColumns_line2_n11 ;
    wire MixColumns_line2_n10 ;
    wire MixColumns_line2_n9 ;
    wire MixColumns_line2_n8 ;
    wire MixColumns_line2_n7 ;
    wire MixColumns_line2_n6 ;
    wire MixColumns_line2_n5 ;
    wire MixColumns_line2_n4 ;
    wire MixColumns_line2_n3 ;
    wire MixColumns_line2_n2 ;
    wire MixColumns_line2_n1 ;
    wire MixColumns_line3_n16 ;
    wire MixColumns_line3_n15 ;
    wire MixColumns_line3_n14 ;
    wire MixColumns_line3_n13 ;
    wire MixColumns_line3_n12 ;
    wire MixColumns_line3_n11 ;
    wire MixColumns_line3_n10 ;
    wire MixColumns_line3_n9 ;
    wire MixColumns_line3_n8 ;
    wire MixColumns_line3_n7 ;
    wire MixColumns_line3_n6 ;
    wire MixColumns_line3_n5 ;
    wire MixColumns_line3_n4 ;
    wire MixColumns_line3_n3 ;
    wire MixColumns_line3_n2 ;
    wire MixColumns_line3_n1 ;
    wire MixColumns_line3_timesTHREE_input2_1_ ;
    wire MixColumns_line3_timesTHREE_input2_3_ ;
    wire MixColumns_line3_timesTHREE_input2_4_ ;
    wire calcRCon_n42 ;
    wire calcRCon_n41 ;
    wire calcRCon_n40 ;
    wire calcRCon_n39 ;
    wire calcRCon_n38 ;
    wire calcRCon_n37 ;
    wire calcRCon_n36 ;
    wire calcRCon_n35 ;
    wire calcRCon_n34 ;
    wire calcRCon_n33 ;
    wire calcRCon_n32 ;
    wire calcRCon_n31 ;
    wire calcRCon_n30 ;
    wire calcRCon_n29 ;
    wire calcRCon_n28 ;
    wire calcRCon_n27 ;
    wire calcRCon_n26 ;
    wire calcRCon_n25 ;
    wire calcRCon_n24 ;
    wire calcRCon_n23 ;
    wire calcRCon_n22 ;
    wire calcRCon_n21 ;
    wire calcRCon_n20 ;
    wire calcRCon_n19 ;
    wire calcRCon_n18 ;
    wire calcRCon_n17 ;
    wire calcRCon_n16 ;
    wire calcRCon_n15 ;
    wire calcRCon_n14 ;
    wire calcRCon_n13 ;
    wire calcRCon_n9 ;
    wire calcRCon_n8 ;
    wire calcRCon_n7 ;
    wire calcRCon_s_current_state_0_ ;
    wire calcRCon_s_current_state_1_ ;
    wire calcRCon_s_current_state_2_ ;
    wire calcRCon_s_current_state_3_ ;
    wire calcRCon_s_current_state_4_ ;
    wire calcRCon_s_current_state_5_ ;
    wire calcRCon_s_current_state_6_ ;
    wire calcRCon_s_current_state_7_ ;
    wire MUX_SboxIn_mux_inst_0_Y ;
    wire MUX_SboxIn_mux_inst_0_X ;
    wire MUX_SboxIn_mux_inst_1_Y ;
    wire MUX_SboxIn_mux_inst_1_X ;
    wire MUX_SboxIn_mux_inst_2_Y ;
    wire MUX_SboxIn_mux_inst_2_X ;
    wire MUX_SboxIn_mux_inst_3_Y ;
    wire MUX_SboxIn_mux_inst_3_X ;
    wire MUX_SboxIn_mux_inst_4_Y ;
    wire MUX_SboxIn_mux_inst_4_X ;
    wire MUX_SboxIn_mux_inst_5_Y ;
    wire MUX_SboxIn_mux_inst_5_X ;
    wire MUX_SboxIn_mux_inst_6_Y ;
    wire MUX_SboxIn_mux_inst_6_X ;
    wire MUX_SboxIn_mux_inst_7_Y ;
    wire MUX_SboxIn_mux_inst_7_X ;
    wire Inst_bSbox_L29 ;
    wire Inst_bSbox_L28 ;
    wire Inst_bSbox_L27 ;
    wire Inst_bSbox_L26 ;
    wire Inst_bSbox_L25 ;
    wire Inst_bSbox_L24 ;
    wire Inst_bSbox_L23 ;
    wire Inst_bSbox_L22 ;
    wire Inst_bSbox_L21 ;
    wire Inst_bSbox_L20 ;
    wire Inst_bSbox_L19 ;
    wire Inst_bSbox_L18 ;
    wire Inst_bSbox_L17 ;
    wire Inst_bSbox_L16 ;
    wire Inst_bSbox_L15 ;
    wire Inst_bSbox_L14 ;
    wire Inst_bSbox_L13 ;
    wire Inst_bSbox_L12 ;
    wire Inst_bSbox_L11 ;
    wire Inst_bSbox_L10 ;
    wire Inst_bSbox_L9 ;
    wire Inst_bSbox_L8 ;
    wire Inst_bSbox_L7 ;
    wire Inst_bSbox_L6 ;
    wire Inst_bSbox_L5 ;
    wire Inst_bSbox_L4 ;
    wire Inst_bSbox_L3 ;
    wire Inst_bSbox_L2 ;
    wire Inst_bSbox_L1 ;
    wire Inst_bSbox_L0 ;
    wire Inst_bSbox_M63 ;
    wire Inst_bSbox_M62 ;
    wire Inst_bSbox_M61 ;
    wire Inst_bSbox_M60 ;
    wire Inst_bSbox_M59 ;
    wire Inst_bSbox_M58 ;
    wire Inst_bSbox_M57 ;
    wire Inst_bSbox_M56 ;
    wire Inst_bSbox_M55 ;
    wire Inst_bSbox_M54 ;
    wire Inst_bSbox_M53 ;
    wire Inst_bSbox_M52 ;
    wire Inst_bSbox_M51 ;
    wire Inst_bSbox_M50 ;
    wire Inst_bSbox_M49 ;
    wire Inst_bSbox_M48 ;
    wire Inst_bSbox_M47 ;
    wire Inst_bSbox_M46 ;
    wire Inst_bSbox_M45 ;
    wire Inst_bSbox_M44 ;
    wire Inst_bSbox_M43 ;
    wire Inst_bSbox_M42 ;
    wire Inst_bSbox_M41 ;
    wire Inst_bSbox_M40 ;
    wire Inst_bSbox_M39 ;
    wire Inst_bSbox_M38 ;
    wire Inst_bSbox_M37 ;
    wire Inst_bSbox_M36 ;
    wire Inst_bSbox_M35 ;
    wire Inst_bSbox_M34 ;
    wire Inst_bSbox_M33 ;
    wire Inst_bSbox_M32 ;
    wire Inst_bSbox_M31 ;
    wire Inst_bSbox_M30 ;
    wire Inst_bSbox_M29 ;
    wire Inst_bSbox_M28 ;
    wire Inst_bSbox_M27 ;
    wire Inst_bSbox_M26 ;
    wire Inst_bSbox_M25 ;
    wire Inst_bSbox_M24 ;
    wire Inst_bSbox_M23 ;
    wire Inst_bSbox_M22 ;
    wire Inst_bSbox_M21 ;
    wire Inst_bSbox_M20 ;
    wire Inst_bSbox_M19 ;
    wire Inst_bSbox_M18 ;
    wire Inst_bSbox_M17 ;
    wire Inst_bSbox_M16 ;
    wire Inst_bSbox_M15 ;
    wire Inst_bSbox_M14 ;
    wire Inst_bSbox_M13 ;
    wire Inst_bSbox_M12 ;
    wire Inst_bSbox_M11 ;
    wire Inst_bSbox_M10 ;
    wire Inst_bSbox_M9 ;
    wire Inst_bSbox_M8 ;
    wire Inst_bSbox_M7 ;
    wire Inst_bSbox_M6 ;
    wire Inst_bSbox_M5 ;
    wire Inst_bSbox_M4 ;
    wire Inst_bSbox_M3 ;
    wire Inst_bSbox_M2 ;
    wire Inst_bSbox_M1 ;
    wire Inst_bSbox_T27 ;
    wire Inst_bSbox_T26 ;
    wire Inst_bSbox_T25 ;
    wire Inst_bSbox_T24 ;
    wire Inst_bSbox_T23 ;
    wire Inst_bSbox_T22 ;
    wire Inst_bSbox_T21 ;
    wire Inst_bSbox_T20 ;
    wire Inst_bSbox_T19 ;
    wire Inst_bSbox_T18 ;
    wire Inst_bSbox_T17 ;
    wire Inst_bSbox_T16 ;
    wire Inst_bSbox_T15 ;
    wire Inst_bSbox_T14 ;
    wire Inst_bSbox_T13 ;
    wire Inst_bSbox_T12 ;
    wire Inst_bSbox_T11 ;
    wire Inst_bSbox_T10 ;
    wire Inst_bSbox_T9 ;
    wire Inst_bSbox_T8 ;
    wire Inst_bSbox_T7 ;
    wire Inst_bSbox_T6 ;
    wire Inst_bSbox_T5 ;
    wire Inst_bSbox_T4 ;
    wire Inst_bSbox_T3 ;
    wire Inst_bSbox_T2 ;
    wire Inst_bSbox_T1 ;
    wire [7:0] SboxOut ;
    wire [7:0] StateOutXORroundKey ;
    wire [7:0] StateIn ;
    wire [31:0] StateInMC ;
    wire [19:0] MCin ;
    wire [31:0] MCout ;
    wire [7:0] keyStateIn ;
    wire [7:0] roundConstant ;
    wire [7:0] keySBIn ;
    wire [7:0] SboxIn ;
    wire [7:0] stateArray_input_MC ;
    wire [7:0] stateArray_inS33ser ;
    wire [7:0] stateArray_outS33ser ;
    wire [7:0] stateArray_outS32ser ;
    wire [7:0] stateArray_outS31ser ;
    wire [7:0] stateArray_inS23ser ;
    wire [7:0] stateArray_outS23ser ;
    wire [7:0] stateArray_outS22ser ;
    wire [7:0] stateArray_outS21ser ;
    wire [7:0] stateArray_inS13ser ;
    wire [7:0] stateArray_outS13ser ;
    wire [7:0] stateArray_outS12ser ;
    wire [7:0] stateArray_outS11ser ;
    wire [7:0] stateArray_inS03ser ;
    wire [7:0] stateArray_outS03ser ;
    wire [7:0] stateArray_outS02ser ;
    wire [7:0] stateArray_outS01ser ;
    wire [7:0] KeyArray_outS01ser_XOR_00 ;
    wire [7:0] KeyArray_inS33ser ;
    wire [7:0] KeyArray_outS33ser ;
    wire [7:0] KeyArray_outS32ser ;
    wire [7:0] KeyArray_inS30par ;
    wire [7:0] KeyArray_outS31ser ;
    wire [7:0] KeyArray_outS30ser ;
    wire [7:0] KeyArray_outS23ser ;
    wire [7:0] KeyArray_outS22ser ;
    wire [7:0] KeyArray_outS21ser ;
    wire [7:0] KeyArray_outS20ser ;
    wire [7:0] KeyArray_outS12ser ;
    wire [7:0] KeyArray_outS11ser ;
    wire [7:0] KeyArray_outS10ser ;
    wire [7:0] KeyArray_outS03ser ;
    wire [7:0] KeyArray_outS02ser ;
    wire [7:0] KeyArray_inS00ser ;
    wire [7:0] MixColumns_line0_S13 ;
    wire [4:1] MixColumns_line0_S02 ;
    wire [4:1] MixColumns_line0_timesTHREE_input2 ;
    wire [7:0] MixColumns_line1_S13 ;
    wire [7:0] MixColumns_line1_S02 ;
    wire [4:1] MixColumns_line1_timesTHREE_input2 ;
    wire [7:0] MixColumns_line2_S13 ;
    wire [7:0] MixColumns_line2_S02 ;
    wire [4:1] MixColumns_line2_timesTHREE_input2 ;
    wire [7:0] MixColumns_line3_S13 ;
    wire [7:0] MixColumns_line3_S02 ;
    wire new_AGEMA_signal_2489 ;
    wire new_AGEMA_signal_2490 ;
    wire new_AGEMA_signal_2491 ;
    wire new_AGEMA_signal_2495 ;
    wire new_AGEMA_signal_2496 ;
    wire new_AGEMA_signal_2497 ;
    wire new_AGEMA_signal_2498 ;
    wire new_AGEMA_signal_2499 ;
    wire new_AGEMA_signal_2500 ;
    wire new_AGEMA_signal_2504 ;
    wire new_AGEMA_signal_2505 ;
    wire new_AGEMA_signal_2506 ;
    wire new_AGEMA_signal_2507 ;
    wire new_AGEMA_signal_2508 ;
    wire new_AGEMA_signal_2509 ;
    wire new_AGEMA_signal_2513 ;
    wire new_AGEMA_signal_2514 ;
    wire new_AGEMA_signal_2515 ;
    wire new_AGEMA_signal_2516 ;
    wire new_AGEMA_signal_2517 ;
    wire new_AGEMA_signal_2518 ;
    wire new_AGEMA_signal_2522 ;
    wire new_AGEMA_signal_2523 ;
    wire new_AGEMA_signal_2524 ;
    wire new_AGEMA_signal_2525 ;
    wire new_AGEMA_signal_2526 ;
    wire new_AGEMA_signal_2527 ;
    wire new_AGEMA_signal_2531 ;
    wire new_AGEMA_signal_2532 ;
    wire new_AGEMA_signal_2533 ;
    wire new_AGEMA_signal_2534 ;
    wire new_AGEMA_signal_2535 ;
    wire new_AGEMA_signal_2536 ;
    wire new_AGEMA_signal_2540 ;
    wire new_AGEMA_signal_2541 ;
    wire new_AGEMA_signal_2542 ;
    wire new_AGEMA_signal_2543 ;
    wire new_AGEMA_signal_2544 ;
    wire new_AGEMA_signal_2545 ;
    wire new_AGEMA_signal_2549 ;
    wire new_AGEMA_signal_2550 ;
    wire new_AGEMA_signal_2551 ;
    wire new_AGEMA_signal_2552 ;
    wire new_AGEMA_signal_2553 ;
    wire new_AGEMA_signal_2554 ;
    wire new_AGEMA_signal_2558 ;
    wire new_AGEMA_signal_2559 ;
    wire new_AGEMA_signal_2560 ;
    wire new_AGEMA_signal_2561 ;
    wire new_AGEMA_signal_2562 ;
    wire new_AGEMA_signal_2563 ;
    wire new_AGEMA_signal_2564 ;
    wire new_AGEMA_signal_2565 ;
    wire new_AGEMA_signal_2566 ;
    wire new_AGEMA_signal_2567 ;
    wire new_AGEMA_signal_2568 ;
    wire new_AGEMA_signal_2569 ;
    wire new_AGEMA_signal_2570 ;
    wire new_AGEMA_signal_2571 ;
    wire new_AGEMA_signal_2573 ;
    wire new_AGEMA_signal_2574 ;
    wire new_AGEMA_signal_2575 ;
    wire new_AGEMA_signal_2576 ;
    wire new_AGEMA_signal_2577 ;
    wire new_AGEMA_signal_2578 ;
    wire new_AGEMA_signal_2579 ;
    wire new_AGEMA_signal_2580 ;
    wire new_AGEMA_signal_2581 ;
    wire new_AGEMA_signal_2582 ;
    wire new_AGEMA_signal_2583 ;
    wire new_AGEMA_signal_2584 ;
    wire new_AGEMA_signal_2585 ;
    wire new_AGEMA_signal_2586 ;
    wire new_AGEMA_signal_2587 ;
    wire new_AGEMA_signal_2588 ;
    wire new_AGEMA_signal_2589 ;
    wire new_AGEMA_signal_2590 ;
    wire new_AGEMA_signal_2591 ;
    wire new_AGEMA_signal_2592 ;
    wire new_AGEMA_signal_2593 ;
    wire new_AGEMA_signal_2594 ;
    wire new_AGEMA_signal_2595 ;
    wire new_AGEMA_signal_2596 ;
    wire new_AGEMA_signal_2597 ;
    wire new_AGEMA_signal_2598 ;
    wire new_AGEMA_signal_2599 ;
    wire new_AGEMA_signal_2600 ;
    wire new_AGEMA_signal_2601 ;
    wire new_AGEMA_signal_2602 ;
    wire new_AGEMA_signal_2603 ;
    wire new_AGEMA_signal_2604 ;
    wire new_AGEMA_signal_2605 ;
    wire new_AGEMA_signal_2606 ;
    wire new_AGEMA_signal_2607 ;
    wire new_AGEMA_signal_2608 ;
    wire new_AGEMA_signal_2609 ;
    wire new_AGEMA_signal_2610 ;
    wire new_AGEMA_signal_2611 ;
    wire new_AGEMA_signal_2612 ;
    wire new_AGEMA_signal_2613 ;
    wire new_AGEMA_signal_2614 ;
    wire new_AGEMA_signal_2615 ;
    wire new_AGEMA_signal_2616 ;
    wire new_AGEMA_signal_2617 ;
    wire new_AGEMA_signal_2618 ;
    wire new_AGEMA_signal_2619 ;
    wire new_AGEMA_signal_2620 ;
    wire new_AGEMA_signal_2621 ;
    wire new_AGEMA_signal_2622 ;
    wire new_AGEMA_signal_2623 ;
    wire new_AGEMA_signal_2624 ;
    wire new_AGEMA_signal_2625 ;
    wire new_AGEMA_signal_2626 ;
    wire new_AGEMA_signal_2627 ;
    wire new_AGEMA_signal_2628 ;
    wire new_AGEMA_signal_2629 ;
    wire new_AGEMA_signal_2630 ;
    wire new_AGEMA_signal_2631 ;
    wire new_AGEMA_signal_2632 ;
    wire new_AGEMA_signal_2633 ;
    wire new_AGEMA_signal_2634 ;
    wire new_AGEMA_signal_2635 ;
    wire new_AGEMA_signal_2636 ;
    wire new_AGEMA_signal_2637 ;
    wire new_AGEMA_signal_2638 ;
    wire new_AGEMA_signal_2639 ;
    wire new_AGEMA_signal_2640 ;
    wire new_AGEMA_signal_2641 ;
    wire new_AGEMA_signal_2642 ;
    wire new_AGEMA_signal_2643 ;
    wire new_AGEMA_signal_2644 ;
    wire new_AGEMA_signal_2645 ;
    wire new_AGEMA_signal_2646 ;
    wire new_AGEMA_signal_2647 ;
    wire new_AGEMA_signal_2648 ;
    wire new_AGEMA_signal_2649 ;
    wire new_AGEMA_signal_2650 ;
    wire new_AGEMA_signal_2651 ;
    wire new_AGEMA_signal_2652 ;
    wire new_AGEMA_signal_2653 ;
    wire new_AGEMA_signal_2654 ;
    wire new_AGEMA_signal_2655 ;
    wire new_AGEMA_signal_2656 ;
    wire new_AGEMA_signal_2657 ;
    wire new_AGEMA_signal_2658 ;
    wire new_AGEMA_signal_2659 ;
    wire new_AGEMA_signal_2660 ;
    wire new_AGEMA_signal_2661 ;
    wire new_AGEMA_signal_2662 ;
    wire new_AGEMA_signal_2663 ;
    wire new_AGEMA_signal_2664 ;
    wire new_AGEMA_signal_2665 ;
    wire new_AGEMA_signal_2666 ;
    wire new_AGEMA_signal_2667 ;
    wire new_AGEMA_signal_2668 ;
    wire new_AGEMA_signal_2669 ;
    wire new_AGEMA_signal_2670 ;
    wire new_AGEMA_signal_2671 ;
    wire new_AGEMA_signal_2672 ;
    wire new_AGEMA_signal_2673 ;
    wire new_AGEMA_signal_2674 ;
    wire new_AGEMA_signal_2675 ;
    wire new_AGEMA_signal_2676 ;
    wire new_AGEMA_signal_2677 ;
    wire new_AGEMA_signal_2678 ;
    wire new_AGEMA_signal_2679 ;
    wire new_AGEMA_signal_2680 ;
    wire new_AGEMA_signal_2681 ;
    wire new_AGEMA_signal_2682 ;
    wire new_AGEMA_signal_2683 ;
    wire new_AGEMA_signal_2684 ;
    wire new_AGEMA_signal_2685 ;
    wire new_AGEMA_signal_2686 ;
    wire new_AGEMA_signal_2687 ;
    wire new_AGEMA_signal_2688 ;
    wire new_AGEMA_signal_2689 ;
    wire new_AGEMA_signal_2690 ;
    wire new_AGEMA_signal_2691 ;
    wire new_AGEMA_signal_2692 ;
    wire new_AGEMA_signal_2693 ;
    wire new_AGEMA_signal_2694 ;
    wire new_AGEMA_signal_2695 ;
    wire new_AGEMA_signal_2696 ;
    wire new_AGEMA_signal_2697 ;
    wire new_AGEMA_signal_2698 ;
    wire new_AGEMA_signal_2699 ;
    wire new_AGEMA_signal_2700 ;
    wire new_AGEMA_signal_2701 ;
    wire new_AGEMA_signal_2702 ;
    wire new_AGEMA_signal_2703 ;
    wire new_AGEMA_signal_2704 ;
    wire new_AGEMA_signal_2705 ;
    wire new_AGEMA_signal_2706 ;
    wire new_AGEMA_signal_2707 ;
    wire new_AGEMA_signal_2708 ;
    wire new_AGEMA_signal_2709 ;
    wire new_AGEMA_signal_2710 ;
    wire new_AGEMA_signal_2711 ;
    wire new_AGEMA_signal_2712 ;
    wire new_AGEMA_signal_2713 ;
    wire new_AGEMA_signal_2714 ;
    wire new_AGEMA_signal_2715 ;
    wire new_AGEMA_signal_2716 ;
    wire new_AGEMA_signal_2717 ;
    wire new_AGEMA_signal_2718 ;
    wire new_AGEMA_signal_2719 ;
    wire new_AGEMA_signal_2720 ;
    wire new_AGEMA_signal_2721 ;
    wire new_AGEMA_signal_2722 ;
    wire new_AGEMA_signal_2723 ;
    wire new_AGEMA_signal_2724 ;
    wire new_AGEMA_signal_2725 ;
    wire new_AGEMA_signal_2726 ;
    wire new_AGEMA_signal_2727 ;
    wire new_AGEMA_signal_2728 ;
    wire new_AGEMA_signal_2729 ;
    wire new_AGEMA_signal_2730 ;
    wire new_AGEMA_signal_2731 ;
    wire new_AGEMA_signal_2732 ;
    wire new_AGEMA_signal_2733 ;
    wire new_AGEMA_signal_2734 ;
    wire new_AGEMA_signal_2735 ;
    wire new_AGEMA_signal_2736 ;
    wire new_AGEMA_signal_2737 ;
    wire new_AGEMA_signal_2738 ;
    wire new_AGEMA_signal_2739 ;
    wire new_AGEMA_signal_2740 ;
    wire new_AGEMA_signal_2741 ;
    wire new_AGEMA_signal_2742 ;
    wire new_AGEMA_signal_2743 ;
    wire new_AGEMA_signal_2744 ;
    wire new_AGEMA_signal_2745 ;
    wire new_AGEMA_signal_2746 ;
    wire new_AGEMA_signal_2747 ;
    wire new_AGEMA_signal_2748 ;
    wire new_AGEMA_signal_2749 ;
    wire new_AGEMA_signal_2750 ;
    wire new_AGEMA_signal_2751 ;
    wire new_AGEMA_signal_2752 ;
    wire new_AGEMA_signal_2753 ;
    wire new_AGEMA_signal_2754 ;
    wire new_AGEMA_signal_2755 ;
    wire new_AGEMA_signal_2756 ;
    wire new_AGEMA_signal_2757 ;
    wire new_AGEMA_signal_2758 ;
    wire new_AGEMA_signal_2759 ;
    wire new_AGEMA_signal_2760 ;
    wire new_AGEMA_signal_2761 ;
    wire new_AGEMA_signal_2762 ;
    wire new_AGEMA_signal_2763 ;
    wire new_AGEMA_signal_2764 ;
    wire new_AGEMA_signal_2765 ;
    wire new_AGEMA_signal_2766 ;
    wire new_AGEMA_signal_2767 ;
    wire new_AGEMA_signal_2768 ;
    wire new_AGEMA_signal_2769 ;
    wire new_AGEMA_signal_2770 ;
    wire new_AGEMA_signal_2771 ;
    wire new_AGEMA_signal_2772 ;
    wire new_AGEMA_signal_2773 ;
    wire new_AGEMA_signal_2774 ;
    wire new_AGEMA_signal_2775 ;
    wire new_AGEMA_signal_2776 ;
    wire new_AGEMA_signal_2777 ;
    wire new_AGEMA_signal_2778 ;
    wire new_AGEMA_signal_2779 ;
    wire new_AGEMA_signal_2780 ;
    wire new_AGEMA_signal_2781 ;
    wire new_AGEMA_signal_2782 ;
    wire new_AGEMA_signal_2783 ;
    wire new_AGEMA_signal_2784 ;
    wire new_AGEMA_signal_2785 ;
    wire new_AGEMA_signal_2786 ;
    wire new_AGEMA_signal_2787 ;
    wire new_AGEMA_signal_2788 ;
    wire new_AGEMA_signal_2789 ;
    wire new_AGEMA_signal_2790 ;
    wire new_AGEMA_signal_2791 ;
    wire new_AGEMA_signal_2792 ;
    wire new_AGEMA_signal_2793 ;
    wire new_AGEMA_signal_2794 ;
    wire new_AGEMA_signal_2795 ;
    wire new_AGEMA_signal_2796 ;
    wire new_AGEMA_signal_2797 ;
    wire new_AGEMA_signal_2798 ;
    wire new_AGEMA_signal_2799 ;
    wire new_AGEMA_signal_2800 ;
    wire new_AGEMA_signal_2801 ;
    wire new_AGEMA_signal_2802 ;
    wire new_AGEMA_signal_2803 ;
    wire new_AGEMA_signal_2804 ;
    wire new_AGEMA_signal_2805 ;
    wire new_AGEMA_signal_2806 ;
    wire new_AGEMA_signal_2807 ;
    wire new_AGEMA_signal_2808 ;
    wire new_AGEMA_signal_2809 ;
    wire new_AGEMA_signal_2810 ;
    wire new_AGEMA_signal_2811 ;
    wire new_AGEMA_signal_2812 ;
    wire new_AGEMA_signal_2813 ;
    wire new_AGEMA_signal_2814 ;
    wire new_AGEMA_signal_2815 ;
    wire new_AGEMA_signal_2816 ;
    wire new_AGEMA_signal_2817 ;
    wire new_AGEMA_signal_2818 ;
    wire new_AGEMA_signal_2819 ;
    wire new_AGEMA_signal_2820 ;
    wire new_AGEMA_signal_2821 ;
    wire new_AGEMA_signal_2822 ;
    wire new_AGEMA_signal_2823 ;
    wire new_AGEMA_signal_2824 ;
    wire new_AGEMA_signal_2825 ;
    wire new_AGEMA_signal_2826 ;
    wire new_AGEMA_signal_2827 ;
    wire new_AGEMA_signal_2828 ;
    wire new_AGEMA_signal_2829 ;
    wire new_AGEMA_signal_2830 ;
    wire new_AGEMA_signal_2831 ;
    wire new_AGEMA_signal_2832 ;
    wire new_AGEMA_signal_2833 ;
    wire new_AGEMA_signal_2834 ;
    wire new_AGEMA_signal_2835 ;
    wire new_AGEMA_signal_2836 ;
    wire new_AGEMA_signal_2837 ;
    wire new_AGEMA_signal_2838 ;
    wire new_AGEMA_signal_2839 ;
    wire new_AGEMA_signal_2840 ;
    wire new_AGEMA_signal_2841 ;
    wire new_AGEMA_signal_2842 ;
    wire new_AGEMA_signal_2843 ;
    wire new_AGEMA_signal_2844 ;
    wire new_AGEMA_signal_2845 ;
    wire new_AGEMA_signal_2846 ;
    wire new_AGEMA_signal_2847 ;
    wire new_AGEMA_signal_2848 ;
    wire new_AGEMA_signal_2849 ;
    wire new_AGEMA_signal_2850 ;
    wire new_AGEMA_signal_2851 ;
    wire new_AGEMA_signal_2852 ;
    wire new_AGEMA_signal_2853 ;
    wire new_AGEMA_signal_2854 ;
    wire new_AGEMA_signal_2855 ;
    wire new_AGEMA_signal_2856 ;
    wire new_AGEMA_signal_2857 ;
    wire new_AGEMA_signal_2858 ;
    wire new_AGEMA_signal_2859 ;
    wire new_AGEMA_signal_2860 ;
    wire new_AGEMA_signal_2861 ;
    wire new_AGEMA_signal_2862 ;
    wire new_AGEMA_signal_2863 ;
    wire new_AGEMA_signal_2864 ;
    wire new_AGEMA_signal_2865 ;
    wire new_AGEMA_signal_2866 ;
    wire new_AGEMA_signal_2867 ;
    wire new_AGEMA_signal_2868 ;
    wire new_AGEMA_signal_2869 ;
    wire new_AGEMA_signal_2870 ;
    wire new_AGEMA_signal_2871 ;
    wire new_AGEMA_signal_2872 ;
    wire new_AGEMA_signal_2873 ;
    wire new_AGEMA_signal_2874 ;
    wire new_AGEMA_signal_2875 ;
    wire new_AGEMA_signal_2876 ;
    wire new_AGEMA_signal_2877 ;
    wire new_AGEMA_signal_2878 ;
    wire new_AGEMA_signal_2879 ;
    wire new_AGEMA_signal_2880 ;
    wire new_AGEMA_signal_2881 ;
    wire new_AGEMA_signal_2882 ;
    wire new_AGEMA_signal_2883 ;
    wire new_AGEMA_signal_2884 ;
    wire new_AGEMA_signal_2885 ;
    wire new_AGEMA_signal_2886 ;
    wire new_AGEMA_signal_2887 ;
    wire new_AGEMA_signal_2888 ;
    wire new_AGEMA_signal_2889 ;
    wire new_AGEMA_signal_2890 ;
    wire new_AGEMA_signal_2891 ;
    wire new_AGEMA_signal_2892 ;
    wire new_AGEMA_signal_2893 ;
    wire new_AGEMA_signal_2894 ;
    wire new_AGEMA_signal_2895 ;
    wire new_AGEMA_signal_2896 ;
    wire new_AGEMA_signal_2897 ;
    wire new_AGEMA_signal_2898 ;
    wire new_AGEMA_signal_2899 ;
    wire new_AGEMA_signal_2900 ;
    wire new_AGEMA_signal_2901 ;
    wire new_AGEMA_signal_2902 ;
    wire new_AGEMA_signal_2903 ;
    wire new_AGEMA_signal_2904 ;
    wire new_AGEMA_signal_2905 ;
    wire new_AGEMA_signal_2906 ;
    wire new_AGEMA_signal_2907 ;
    wire new_AGEMA_signal_2908 ;
    wire new_AGEMA_signal_2909 ;
    wire new_AGEMA_signal_2910 ;
    wire new_AGEMA_signal_2911 ;
    wire new_AGEMA_signal_2912 ;
    wire new_AGEMA_signal_2913 ;
    wire new_AGEMA_signal_2914 ;
    wire new_AGEMA_signal_2915 ;
    wire new_AGEMA_signal_2916 ;
    wire new_AGEMA_signal_2917 ;
    wire new_AGEMA_signal_2918 ;
    wire new_AGEMA_signal_2919 ;
    wire new_AGEMA_signal_2920 ;
    wire new_AGEMA_signal_2921 ;
    wire new_AGEMA_signal_2922 ;
    wire new_AGEMA_signal_2923 ;
    wire new_AGEMA_signal_2924 ;
    wire new_AGEMA_signal_2925 ;
    wire new_AGEMA_signal_2926 ;
    wire new_AGEMA_signal_2927 ;
    wire new_AGEMA_signal_2928 ;
    wire new_AGEMA_signal_2929 ;
    wire new_AGEMA_signal_2930 ;
    wire new_AGEMA_signal_2931 ;
    wire new_AGEMA_signal_2932 ;
    wire new_AGEMA_signal_2933 ;
    wire new_AGEMA_signal_2934 ;
    wire new_AGEMA_signal_2935 ;
    wire new_AGEMA_signal_2936 ;
    wire new_AGEMA_signal_2937 ;
    wire new_AGEMA_signal_2938 ;
    wire new_AGEMA_signal_2939 ;
    wire new_AGEMA_signal_2940 ;
    wire new_AGEMA_signal_2941 ;
    wire new_AGEMA_signal_2942 ;
    wire new_AGEMA_signal_2943 ;
    wire new_AGEMA_signal_2944 ;
    wire new_AGEMA_signal_2945 ;
    wire new_AGEMA_signal_2946 ;
    wire new_AGEMA_signal_2947 ;
    wire new_AGEMA_signal_2948 ;
    wire new_AGEMA_signal_2949 ;
    wire new_AGEMA_signal_2950 ;
    wire new_AGEMA_signal_2951 ;
    wire new_AGEMA_signal_2952 ;
    wire new_AGEMA_signal_2953 ;
    wire new_AGEMA_signal_2954 ;
    wire new_AGEMA_signal_2955 ;
    wire new_AGEMA_signal_2956 ;
    wire new_AGEMA_signal_2957 ;
    wire new_AGEMA_signal_2958 ;
    wire new_AGEMA_signal_2959 ;
    wire new_AGEMA_signal_2960 ;
    wire new_AGEMA_signal_2961 ;
    wire new_AGEMA_signal_2962 ;
    wire new_AGEMA_signal_2963 ;
    wire new_AGEMA_signal_2964 ;
    wire new_AGEMA_signal_2965 ;
    wire new_AGEMA_signal_2966 ;
    wire new_AGEMA_signal_2967 ;
    wire new_AGEMA_signal_2968 ;
    wire new_AGEMA_signal_2969 ;
    wire new_AGEMA_signal_2970 ;
    wire new_AGEMA_signal_2971 ;
    wire new_AGEMA_signal_2972 ;
    wire new_AGEMA_signal_2973 ;
    wire new_AGEMA_signal_2974 ;
    wire new_AGEMA_signal_2975 ;
    wire new_AGEMA_signal_2976 ;
    wire new_AGEMA_signal_2977 ;
    wire new_AGEMA_signal_2978 ;
    wire new_AGEMA_signal_2979 ;
    wire new_AGEMA_signal_2980 ;
    wire new_AGEMA_signal_2981 ;
    wire new_AGEMA_signal_2982 ;
    wire new_AGEMA_signal_2983 ;
    wire new_AGEMA_signal_2984 ;
    wire new_AGEMA_signal_2985 ;
    wire new_AGEMA_signal_2986 ;
    wire new_AGEMA_signal_2987 ;
    wire new_AGEMA_signal_2988 ;
    wire new_AGEMA_signal_2989 ;
    wire new_AGEMA_signal_2990 ;
    wire new_AGEMA_signal_2991 ;
    wire new_AGEMA_signal_2992 ;
    wire new_AGEMA_signal_2993 ;
    wire new_AGEMA_signal_2994 ;
    wire new_AGEMA_signal_2995 ;
    wire new_AGEMA_signal_2996 ;
    wire new_AGEMA_signal_2997 ;
    wire new_AGEMA_signal_2998 ;
    wire new_AGEMA_signal_2999 ;
    wire new_AGEMA_signal_3000 ;
    wire new_AGEMA_signal_3001 ;
    wire new_AGEMA_signal_3002 ;
    wire new_AGEMA_signal_3003 ;
    wire new_AGEMA_signal_3004 ;
    wire new_AGEMA_signal_3005 ;
    wire new_AGEMA_signal_3006 ;
    wire new_AGEMA_signal_3007 ;
    wire new_AGEMA_signal_3008 ;
    wire new_AGEMA_signal_3009 ;
    wire new_AGEMA_signal_3010 ;
    wire new_AGEMA_signal_3011 ;
    wire new_AGEMA_signal_3012 ;
    wire new_AGEMA_signal_3013 ;
    wire new_AGEMA_signal_3014 ;
    wire new_AGEMA_signal_3015 ;
    wire new_AGEMA_signal_3016 ;
    wire new_AGEMA_signal_3017 ;
    wire new_AGEMA_signal_3018 ;
    wire new_AGEMA_signal_3019 ;
    wire new_AGEMA_signal_3020 ;
    wire new_AGEMA_signal_3021 ;
    wire new_AGEMA_signal_3022 ;
    wire new_AGEMA_signal_3023 ;
    wire new_AGEMA_signal_3024 ;
    wire new_AGEMA_signal_3025 ;
    wire new_AGEMA_signal_3026 ;
    wire new_AGEMA_signal_3027 ;
    wire new_AGEMA_signal_3028 ;
    wire new_AGEMA_signal_3029 ;
    wire new_AGEMA_signal_3030 ;
    wire new_AGEMA_signal_3031 ;
    wire new_AGEMA_signal_3032 ;
    wire new_AGEMA_signal_3033 ;
    wire new_AGEMA_signal_3034 ;
    wire new_AGEMA_signal_3035 ;
    wire new_AGEMA_signal_3036 ;
    wire new_AGEMA_signal_3037 ;
    wire new_AGEMA_signal_3038 ;
    wire new_AGEMA_signal_3039 ;
    wire new_AGEMA_signal_3040 ;
    wire new_AGEMA_signal_3041 ;
    wire new_AGEMA_signal_3042 ;
    wire new_AGEMA_signal_3043 ;
    wire new_AGEMA_signal_3044 ;
    wire new_AGEMA_signal_3045 ;
    wire new_AGEMA_signal_3046 ;
    wire new_AGEMA_signal_3047 ;
    wire new_AGEMA_signal_3048 ;
    wire new_AGEMA_signal_3049 ;
    wire new_AGEMA_signal_3050 ;
    wire new_AGEMA_signal_3051 ;
    wire new_AGEMA_signal_3052 ;
    wire new_AGEMA_signal_3053 ;
    wire new_AGEMA_signal_3054 ;
    wire new_AGEMA_signal_3055 ;
    wire new_AGEMA_signal_3056 ;
    wire new_AGEMA_signal_3057 ;
    wire new_AGEMA_signal_3058 ;
    wire new_AGEMA_signal_3059 ;
    wire new_AGEMA_signal_3060 ;
    wire new_AGEMA_signal_3061 ;
    wire new_AGEMA_signal_3062 ;
    wire new_AGEMA_signal_3063 ;
    wire new_AGEMA_signal_3064 ;
    wire new_AGEMA_signal_3065 ;
    wire new_AGEMA_signal_3066 ;
    wire new_AGEMA_signal_3067 ;
    wire new_AGEMA_signal_3068 ;
    wire new_AGEMA_signal_3069 ;
    wire new_AGEMA_signal_3070 ;
    wire new_AGEMA_signal_3071 ;
    wire new_AGEMA_signal_3072 ;
    wire new_AGEMA_signal_3073 ;
    wire new_AGEMA_signal_3074 ;
    wire new_AGEMA_signal_3075 ;
    wire new_AGEMA_signal_3076 ;
    wire new_AGEMA_signal_3077 ;
    wire new_AGEMA_signal_3078 ;
    wire new_AGEMA_signal_3079 ;
    wire new_AGEMA_signal_3080 ;
    wire new_AGEMA_signal_3081 ;
    wire new_AGEMA_signal_3082 ;
    wire new_AGEMA_signal_3083 ;
    wire new_AGEMA_signal_3084 ;
    wire new_AGEMA_signal_3085 ;
    wire new_AGEMA_signal_3086 ;
    wire new_AGEMA_signal_3087 ;
    wire new_AGEMA_signal_3088 ;
    wire new_AGEMA_signal_3089 ;
    wire new_AGEMA_signal_3090 ;
    wire new_AGEMA_signal_3091 ;
    wire new_AGEMA_signal_3092 ;
    wire new_AGEMA_signal_3093 ;
    wire new_AGEMA_signal_3094 ;
    wire new_AGEMA_signal_3095 ;
    wire new_AGEMA_signal_3096 ;
    wire new_AGEMA_signal_3097 ;
    wire new_AGEMA_signal_3098 ;
    wire new_AGEMA_signal_3099 ;
    wire new_AGEMA_signal_3100 ;
    wire new_AGEMA_signal_3101 ;
    wire new_AGEMA_signal_3102 ;
    wire new_AGEMA_signal_3103 ;
    wire new_AGEMA_signal_3104 ;
    wire new_AGEMA_signal_3105 ;
    wire new_AGEMA_signal_3106 ;
    wire new_AGEMA_signal_3107 ;
    wire new_AGEMA_signal_3108 ;
    wire new_AGEMA_signal_3109 ;
    wire new_AGEMA_signal_3110 ;
    wire new_AGEMA_signal_3111 ;
    wire new_AGEMA_signal_3112 ;
    wire new_AGEMA_signal_3113 ;
    wire new_AGEMA_signal_3114 ;
    wire new_AGEMA_signal_3115 ;
    wire new_AGEMA_signal_3116 ;
    wire new_AGEMA_signal_3117 ;
    wire new_AGEMA_signal_3118 ;
    wire new_AGEMA_signal_3119 ;
    wire new_AGEMA_signal_3120 ;
    wire new_AGEMA_signal_3121 ;
    wire new_AGEMA_signal_3122 ;
    wire new_AGEMA_signal_3123 ;
    wire new_AGEMA_signal_3124 ;
    wire new_AGEMA_signal_3125 ;
    wire new_AGEMA_signal_3126 ;
    wire new_AGEMA_signal_3127 ;
    wire new_AGEMA_signal_3128 ;
    wire new_AGEMA_signal_3129 ;
    wire new_AGEMA_signal_3130 ;
    wire new_AGEMA_signal_3131 ;
    wire new_AGEMA_signal_3132 ;
    wire new_AGEMA_signal_3133 ;
    wire new_AGEMA_signal_3134 ;
    wire new_AGEMA_signal_3135 ;
    wire new_AGEMA_signal_3136 ;
    wire new_AGEMA_signal_3137 ;
    wire new_AGEMA_signal_3138 ;
    wire new_AGEMA_signal_3139 ;
    wire new_AGEMA_signal_3140 ;
    wire new_AGEMA_signal_3141 ;
    wire new_AGEMA_signal_3142 ;
    wire new_AGEMA_signal_3143 ;
    wire new_AGEMA_signal_3144 ;
    wire new_AGEMA_signal_3145 ;
    wire new_AGEMA_signal_3146 ;
    wire new_AGEMA_signal_3147 ;
    wire new_AGEMA_signal_3148 ;
    wire new_AGEMA_signal_3149 ;
    wire new_AGEMA_signal_3150 ;
    wire new_AGEMA_signal_3151 ;
    wire new_AGEMA_signal_3152 ;
    wire new_AGEMA_signal_3153 ;
    wire new_AGEMA_signal_3154 ;
    wire new_AGEMA_signal_3155 ;
    wire new_AGEMA_signal_3156 ;
    wire new_AGEMA_signal_3157 ;
    wire new_AGEMA_signal_3158 ;
    wire new_AGEMA_signal_3159 ;
    wire new_AGEMA_signal_3160 ;
    wire new_AGEMA_signal_3161 ;
    wire new_AGEMA_signal_3162 ;
    wire new_AGEMA_signal_3163 ;
    wire new_AGEMA_signal_3164 ;
    wire new_AGEMA_signal_3165 ;
    wire new_AGEMA_signal_3166 ;
    wire new_AGEMA_signal_3167 ;
    wire new_AGEMA_signal_3168 ;
    wire new_AGEMA_signal_3169 ;
    wire new_AGEMA_signal_3170 ;
    wire new_AGEMA_signal_3171 ;
    wire new_AGEMA_signal_3172 ;
    wire new_AGEMA_signal_3173 ;
    wire new_AGEMA_signal_3174 ;
    wire new_AGEMA_signal_3175 ;
    wire new_AGEMA_signal_3176 ;
    wire new_AGEMA_signal_3177 ;
    wire new_AGEMA_signal_3178 ;
    wire new_AGEMA_signal_3179 ;
    wire new_AGEMA_signal_3180 ;
    wire new_AGEMA_signal_3181 ;
    wire new_AGEMA_signal_3182 ;
    wire new_AGEMA_signal_3183 ;
    wire new_AGEMA_signal_3184 ;
    wire new_AGEMA_signal_3185 ;
    wire new_AGEMA_signal_3186 ;
    wire new_AGEMA_signal_3187 ;
    wire new_AGEMA_signal_3188 ;
    wire new_AGEMA_signal_3189 ;
    wire new_AGEMA_signal_3190 ;
    wire new_AGEMA_signal_3191 ;
    wire new_AGEMA_signal_3192 ;
    wire new_AGEMA_signal_3193 ;
    wire new_AGEMA_signal_3194 ;
    wire new_AGEMA_signal_3195 ;
    wire new_AGEMA_signal_3196 ;
    wire new_AGEMA_signal_3197 ;
    wire new_AGEMA_signal_3198 ;
    wire new_AGEMA_signal_3199 ;
    wire new_AGEMA_signal_3200 ;
    wire new_AGEMA_signal_3201 ;
    wire new_AGEMA_signal_3202 ;
    wire new_AGEMA_signal_3203 ;
    wire new_AGEMA_signal_3204 ;
    wire new_AGEMA_signal_3205 ;
    wire new_AGEMA_signal_3206 ;
    wire new_AGEMA_signal_3207 ;
    wire new_AGEMA_signal_3208 ;
    wire new_AGEMA_signal_3209 ;
    wire new_AGEMA_signal_3210 ;
    wire new_AGEMA_signal_3211 ;
    wire new_AGEMA_signal_3212 ;
    wire new_AGEMA_signal_3213 ;
    wire new_AGEMA_signal_3214 ;
    wire new_AGEMA_signal_3215 ;
    wire new_AGEMA_signal_3216 ;
    wire new_AGEMA_signal_3217 ;
    wire new_AGEMA_signal_3218 ;
    wire new_AGEMA_signal_3219 ;
    wire new_AGEMA_signal_3220 ;
    wire new_AGEMA_signal_3221 ;
    wire new_AGEMA_signal_3222 ;
    wire new_AGEMA_signal_3223 ;
    wire new_AGEMA_signal_3224 ;
    wire new_AGEMA_signal_3225 ;
    wire new_AGEMA_signal_3226 ;
    wire new_AGEMA_signal_3227 ;
    wire new_AGEMA_signal_3228 ;
    wire new_AGEMA_signal_3229 ;
    wire new_AGEMA_signal_3230 ;
    wire new_AGEMA_signal_3231 ;
    wire new_AGEMA_signal_3232 ;
    wire new_AGEMA_signal_3233 ;
    wire new_AGEMA_signal_3234 ;
    wire new_AGEMA_signal_3235 ;
    wire new_AGEMA_signal_3236 ;
    wire new_AGEMA_signal_3237 ;
    wire new_AGEMA_signal_3238 ;
    wire new_AGEMA_signal_3239 ;
    wire new_AGEMA_signal_3240 ;
    wire new_AGEMA_signal_3241 ;
    wire new_AGEMA_signal_3242 ;
    wire new_AGEMA_signal_3243 ;
    wire new_AGEMA_signal_3244 ;
    wire new_AGEMA_signal_3245 ;
    wire new_AGEMA_signal_3246 ;
    wire new_AGEMA_signal_3247 ;
    wire new_AGEMA_signal_3248 ;
    wire new_AGEMA_signal_3249 ;
    wire new_AGEMA_signal_3250 ;
    wire new_AGEMA_signal_3251 ;
    wire new_AGEMA_signal_3252 ;
    wire new_AGEMA_signal_3253 ;
    wire new_AGEMA_signal_3254 ;
    wire new_AGEMA_signal_3255 ;
    wire new_AGEMA_signal_3256 ;
    wire new_AGEMA_signal_3257 ;
    wire new_AGEMA_signal_3258 ;
    wire new_AGEMA_signal_3259 ;
    wire new_AGEMA_signal_3260 ;
    wire new_AGEMA_signal_3261 ;
    wire new_AGEMA_signal_3262 ;
    wire new_AGEMA_signal_3263 ;
    wire new_AGEMA_signal_3264 ;
    wire new_AGEMA_signal_3265 ;
    wire new_AGEMA_signal_3266 ;
    wire new_AGEMA_signal_3267 ;
    wire new_AGEMA_signal_3268 ;
    wire new_AGEMA_signal_3269 ;
    wire new_AGEMA_signal_3270 ;
    wire new_AGEMA_signal_3271 ;
    wire new_AGEMA_signal_3272 ;
    wire new_AGEMA_signal_3273 ;
    wire new_AGEMA_signal_3274 ;
    wire new_AGEMA_signal_3275 ;
    wire new_AGEMA_signal_3276 ;
    wire new_AGEMA_signal_3277 ;
    wire new_AGEMA_signal_3278 ;
    wire new_AGEMA_signal_3279 ;
    wire new_AGEMA_signal_3280 ;
    wire new_AGEMA_signal_3281 ;
    wire new_AGEMA_signal_3282 ;
    wire new_AGEMA_signal_3283 ;
    wire new_AGEMA_signal_3284 ;
    wire new_AGEMA_signal_3285 ;
    wire new_AGEMA_signal_3286 ;
    wire new_AGEMA_signal_3287 ;
    wire new_AGEMA_signal_3288 ;
    wire new_AGEMA_signal_3289 ;
    wire new_AGEMA_signal_3290 ;
    wire new_AGEMA_signal_3291 ;
    wire new_AGEMA_signal_3292 ;
    wire new_AGEMA_signal_3293 ;
    wire new_AGEMA_signal_3294 ;
    wire new_AGEMA_signal_3295 ;
    wire new_AGEMA_signal_3296 ;
    wire new_AGEMA_signal_3297 ;
    wire new_AGEMA_signal_3298 ;
    wire new_AGEMA_signal_3299 ;
    wire new_AGEMA_signal_3300 ;
    wire new_AGEMA_signal_3301 ;
    wire new_AGEMA_signal_3302 ;
    wire new_AGEMA_signal_3303 ;
    wire new_AGEMA_signal_3304 ;
    wire new_AGEMA_signal_3305 ;
    wire new_AGEMA_signal_3306 ;
    wire new_AGEMA_signal_3307 ;
    wire new_AGEMA_signal_3308 ;
    wire new_AGEMA_signal_3309 ;
    wire new_AGEMA_signal_3310 ;
    wire new_AGEMA_signal_3311 ;
    wire new_AGEMA_signal_3312 ;
    wire new_AGEMA_signal_3313 ;
    wire new_AGEMA_signal_3314 ;
    wire new_AGEMA_signal_3315 ;
    wire new_AGEMA_signal_3316 ;
    wire new_AGEMA_signal_3317 ;
    wire new_AGEMA_signal_3318 ;
    wire new_AGEMA_signal_3319 ;
    wire new_AGEMA_signal_3320 ;
    wire new_AGEMA_signal_3321 ;
    wire new_AGEMA_signal_3322 ;
    wire new_AGEMA_signal_3323 ;
    wire new_AGEMA_signal_3324 ;
    wire new_AGEMA_signal_3325 ;
    wire new_AGEMA_signal_3326 ;
    wire new_AGEMA_signal_3327 ;
    wire new_AGEMA_signal_3328 ;
    wire new_AGEMA_signal_3329 ;
    wire new_AGEMA_signal_3330 ;
    wire new_AGEMA_signal_3331 ;
    wire new_AGEMA_signal_3332 ;
    wire new_AGEMA_signal_3333 ;
    wire new_AGEMA_signal_3334 ;
    wire new_AGEMA_signal_3335 ;
    wire new_AGEMA_signal_3336 ;
    wire new_AGEMA_signal_3337 ;
    wire new_AGEMA_signal_3338 ;
    wire new_AGEMA_signal_3339 ;
    wire new_AGEMA_signal_3340 ;
    wire new_AGEMA_signal_3341 ;
    wire new_AGEMA_signal_3342 ;
    wire new_AGEMA_signal_3343 ;
    wire new_AGEMA_signal_3344 ;
    wire new_AGEMA_signal_3345 ;
    wire new_AGEMA_signal_3346 ;
    wire new_AGEMA_signal_3347 ;
    wire new_AGEMA_signal_3348 ;
    wire new_AGEMA_signal_3349 ;
    wire new_AGEMA_signal_3350 ;
    wire new_AGEMA_signal_3351 ;
    wire new_AGEMA_signal_3352 ;
    wire new_AGEMA_signal_3353 ;
    wire new_AGEMA_signal_3354 ;
    wire new_AGEMA_signal_3355 ;
    wire new_AGEMA_signal_3356 ;
    wire new_AGEMA_signal_3357 ;
    wire new_AGEMA_signal_3358 ;
    wire new_AGEMA_signal_3359 ;
    wire new_AGEMA_signal_3360 ;
    wire new_AGEMA_signal_3361 ;
    wire new_AGEMA_signal_3362 ;
    wire new_AGEMA_signal_3363 ;
    wire new_AGEMA_signal_3364 ;
    wire new_AGEMA_signal_3365 ;
    wire new_AGEMA_signal_3366 ;
    wire new_AGEMA_signal_3367 ;
    wire new_AGEMA_signal_3368 ;
    wire new_AGEMA_signal_3369 ;
    wire new_AGEMA_signal_3370 ;
    wire new_AGEMA_signal_3371 ;
    wire new_AGEMA_signal_3372 ;
    wire new_AGEMA_signal_3373 ;
    wire new_AGEMA_signal_3374 ;
    wire new_AGEMA_signal_3375 ;
    wire new_AGEMA_signal_3376 ;
    wire new_AGEMA_signal_3377 ;
    wire new_AGEMA_signal_3378 ;
    wire new_AGEMA_signal_3379 ;
    wire new_AGEMA_signal_3380 ;
    wire new_AGEMA_signal_3381 ;
    wire new_AGEMA_signal_3382 ;
    wire new_AGEMA_signal_3383 ;
    wire new_AGEMA_signal_3384 ;
    wire new_AGEMA_signal_3385 ;
    wire new_AGEMA_signal_3386 ;
    wire new_AGEMA_signal_3387 ;
    wire new_AGEMA_signal_3388 ;
    wire new_AGEMA_signal_3389 ;
    wire new_AGEMA_signal_3390 ;
    wire new_AGEMA_signal_3391 ;
    wire new_AGEMA_signal_3392 ;
    wire new_AGEMA_signal_3393 ;
    wire new_AGEMA_signal_3394 ;
    wire new_AGEMA_signal_3395 ;
    wire new_AGEMA_signal_3396 ;
    wire new_AGEMA_signal_3397 ;
    wire new_AGEMA_signal_3398 ;
    wire new_AGEMA_signal_3399 ;
    wire new_AGEMA_signal_3400 ;
    wire new_AGEMA_signal_3401 ;
    wire new_AGEMA_signal_3402 ;
    wire new_AGEMA_signal_3403 ;
    wire new_AGEMA_signal_3404 ;
    wire new_AGEMA_signal_3405 ;
    wire new_AGEMA_signal_3406 ;
    wire new_AGEMA_signal_3407 ;
    wire new_AGEMA_signal_3408 ;
    wire new_AGEMA_signal_3409 ;
    wire new_AGEMA_signal_3410 ;
    wire new_AGEMA_signal_3411 ;
    wire new_AGEMA_signal_3412 ;
    wire new_AGEMA_signal_3413 ;
    wire new_AGEMA_signal_3414 ;
    wire new_AGEMA_signal_3415 ;
    wire new_AGEMA_signal_3416 ;
    wire new_AGEMA_signal_3417 ;
    wire new_AGEMA_signal_3418 ;
    wire new_AGEMA_signal_3419 ;
    wire new_AGEMA_signal_3420 ;
    wire new_AGEMA_signal_3421 ;
    wire new_AGEMA_signal_3422 ;
    wire new_AGEMA_signal_3423 ;
    wire new_AGEMA_signal_3424 ;
    wire new_AGEMA_signal_3425 ;
    wire new_AGEMA_signal_3426 ;
    wire new_AGEMA_signal_3427 ;
    wire new_AGEMA_signal_3428 ;
    wire new_AGEMA_signal_3429 ;
    wire new_AGEMA_signal_3430 ;
    wire new_AGEMA_signal_3431 ;
    wire new_AGEMA_signal_3432 ;
    wire new_AGEMA_signal_3433 ;
    wire new_AGEMA_signal_3434 ;
    wire new_AGEMA_signal_3435 ;
    wire new_AGEMA_signal_3436 ;
    wire new_AGEMA_signal_3437 ;
    wire new_AGEMA_signal_3438 ;
    wire new_AGEMA_signal_3439 ;
    wire new_AGEMA_signal_3440 ;
    wire new_AGEMA_signal_3441 ;
    wire new_AGEMA_signal_3442 ;
    wire new_AGEMA_signal_3443 ;
    wire new_AGEMA_signal_3444 ;
    wire new_AGEMA_signal_3445 ;
    wire new_AGEMA_signal_3446 ;
    wire new_AGEMA_signal_3447 ;
    wire new_AGEMA_signal_3448 ;
    wire new_AGEMA_signal_3449 ;
    wire new_AGEMA_signal_3450 ;
    wire new_AGEMA_signal_3451 ;
    wire new_AGEMA_signal_3452 ;
    wire new_AGEMA_signal_3453 ;
    wire new_AGEMA_signal_3454 ;
    wire new_AGEMA_signal_3455 ;
    wire new_AGEMA_signal_3456 ;
    wire new_AGEMA_signal_3457 ;
    wire new_AGEMA_signal_3458 ;
    wire new_AGEMA_signal_3459 ;
    wire new_AGEMA_signal_3460 ;
    wire new_AGEMA_signal_3461 ;
    wire new_AGEMA_signal_3462 ;
    wire new_AGEMA_signal_3463 ;
    wire new_AGEMA_signal_3464 ;
    wire new_AGEMA_signal_3465 ;
    wire new_AGEMA_signal_3466 ;
    wire new_AGEMA_signal_3467 ;
    wire new_AGEMA_signal_3468 ;
    wire new_AGEMA_signal_3469 ;
    wire new_AGEMA_signal_3470 ;
    wire new_AGEMA_signal_3471 ;
    wire new_AGEMA_signal_3472 ;
    wire new_AGEMA_signal_3473 ;
    wire new_AGEMA_signal_3474 ;
    wire new_AGEMA_signal_3475 ;
    wire new_AGEMA_signal_3476 ;
    wire new_AGEMA_signal_3477 ;
    wire new_AGEMA_signal_3478 ;
    wire new_AGEMA_signal_3479 ;
    wire new_AGEMA_signal_3480 ;
    wire new_AGEMA_signal_3481 ;
    wire new_AGEMA_signal_3482 ;
    wire new_AGEMA_signal_3483 ;
    wire new_AGEMA_signal_3484 ;
    wire new_AGEMA_signal_3485 ;
    wire new_AGEMA_signal_3486 ;
    wire new_AGEMA_signal_3487 ;
    wire new_AGEMA_signal_3488 ;
    wire new_AGEMA_signal_3489 ;
    wire new_AGEMA_signal_3490 ;
    wire new_AGEMA_signal_3491 ;
    wire new_AGEMA_signal_3492 ;
    wire new_AGEMA_signal_3493 ;
    wire new_AGEMA_signal_3494 ;
    wire new_AGEMA_signal_3495 ;
    wire new_AGEMA_signal_3496 ;
    wire new_AGEMA_signal_3497 ;
    wire new_AGEMA_signal_3498 ;
    wire new_AGEMA_signal_3499 ;
    wire new_AGEMA_signal_3500 ;
    wire new_AGEMA_signal_3501 ;
    wire new_AGEMA_signal_3502 ;
    wire new_AGEMA_signal_3503 ;
    wire new_AGEMA_signal_3504 ;
    wire new_AGEMA_signal_3505 ;
    wire new_AGEMA_signal_3506 ;
    wire new_AGEMA_signal_3507 ;
    wire new_AGEMA_signal_3508 ;
    wire new_AGEMA_signal_3509 ;
    wire new_AGEMA_signal_3510 ;
    wire new_AGEMA_signal_3511 ;
    wire new_AGEMA_signal_3512 ;
    wire new_AGEMA_signal_3513 ;
    wire new_AGEMA_signal_3514 ;
    wire new_AGEMA_signal_3515 ;
    wire new_AGEMA_signal_3516 ;
    wire new_AGEMA_signal_3517 ;
    wire new_AGEMA_signal_3518 ;
    wire new_AGEMA_signal_3519 ;
    wire new_AGEMA_signal_3520 ;
    wire new_AGEMA_signal_3521 ;
    wire new_AGEMA_signal_3522 ;
    wire new_AGEMA_signal_3523 ;
    wire new_AGEMA_signal_3524 ;
    wire new_AGEMA_signal_3525 ;
    wire new_AGEMA_signal_3526 ;
    wire new_AGEMA_signal_3527 ;
    wire new_AGEMA_signal_3528 ;
    wire new_AGEMA_signal_3529 ;
    wire new_AGEMA_signal_3530 ;
    wire new_AGEMA_signal_3531 ;
    wire new_AGEMA_signal_3532 ;
    wire new_AGEMA_signal_3533 ;
    wire new_AGEMA_signal_3534 ;
    wire new_AGEMA_signal_3535 ;
    wire new_AGEMA_signal_3536 ;
    wire new_AGEMA_signal_3537 ;
    wire new_AGEMA_signal_3538 ;
    wire new_AGEMA_signal_3539 ;
    wire new_AGEMA_signal_3540 ;
    wire new_AGEMA_signal_3541 ;
    wire new_AGEMA_signal_3542 ;
    wire new_AGEMA_signal_3543 ;
    wire new_AGEMA_signal_3544 ;
    wire new_AGEMA_signal_3545 ;
    wire new_AGEMA_signal_3546 ;
    wire new_AGEMA_signal_3547 ;
    wire new_AGEMA_signal_3548 ;
    wire new_AGEMA_signal_3549 ;
    wire new_AGEMA_signal_3550 ;
    wire new_AGEMA_signal_3551 ;
    wire new_AGEMA_signal_3552 ;
    wire new_AGEMA_signal_3553 ;
    wire new_AGEMA_signal_3554 ;
    wire new_AGEMA_signal_3555 ;
    wire new_AGEMA_signal_3556 ;
    wire new_AGEMA_signal_3557 ;
    wire new_AGEMA_signal_3558 ;
    wire new_AGEMA_signal_3559 ;
    wire new_AGEMA_signal_3560 ;
    wire new_AGEMA_signal_3561 ;
    wire new_AGEMA_signal_3562 ;
    wire new_AGEMA_signal_3563 ;
    wire new_AGEMA_signal_3564 ;
    wire new_AGEMA_signal_3565 ;
    wire new_AGEMA_signal_3566 ;
    wire new_AGEMA_signal_3567 ;
    wire new_AGEMA_signal_3568 ;
    wire new_AGEMA_signal_3569 ;
    wire new_AGEMA_signal_3570 ;
    wire new_AGEMA_signal_3571 ;
    wire new_AGEMA_signal_3572 ;
    wire new_AGEMA_signal_3573 ;
    wire new_AGEMA_signal_3574 ;
    wire new_AGEMA_signal_3575 ;
    wire new_AGEMA_signal_3576 ;
    wire new_AGEMA_signal_3577 ;
    wire new_AGEMA_signal_3578 ;
    wire new_AGEMA_signal_3579 ;
    wire new_AGEMA_signal_3580 ;
    wire new_AGEMA_signal_3581 ;
    wire new_AGEMA_signal_3582 ;
    wire new_AGEMA_signal_3583 ;
    wire new_AGEMA_signal_3584 ;
    wire new_AGEMA_signal_3585 ;
    wire new_AGEMA_signal_3586 ;
    wire new_AGEMA_signal_3587 ;
    wire new_AGEMA_signal_3588 ;
    wire new_AGEMA_signal_3589 ;
    wire new_AGEMA_signal_3590 ;
    wire new_AGEMA_signal_3591 ;
    wire new_AGEMA_signal_3592 ;
    wire new_AGEMA_signal_3593 ;
    wire new_AGEMA_signal_3594 ;
    wire new_AGEMA_signal_3595 ;
    wire new_AGEMA_signal_3596 ;
    wire new_AGEMA_signal_3597 ;
    wire new_AGEMA_signal_3598 ;
    wire new_AGEMA_signal_3599 ;
    wire new_AGEMA_signal_3600 ;
    wire new_AGEMA_signal_3601 ;
    wire new_AGEMA_signal_3602 ;
    wire new_AGEMA_signal_3603 ;
    wire new_AGEMA_signal_3604 ;
    wire new_AGEMA_signal_3605 ;
    wire new_AGEMA_signal_3606 ;
    wire new_AGEMA_signal_3607 ;
    wire new_AGEMA_signal_3608 ;
    wire new_AGEMA_signal_3609 ;
    wire new_AGEMA_signal_3610 ;
    wire new_AGEMA_signal_3611 ;
    wire new_AGEMA_signal_3612 ;
    wire new_AGEMA_signal_3613 ;
    wire new_AGEMA_signal_3614 ;
    wire new_AGEMA_signal_3615 ;
    wire new_AGEMA_signal_3616 ;
    wire new_AGEMA_signal_3617 ;
    wire new_AGEMA_signal_3618 ;
    wire new_AGEMA_signal_3619 ;
    wire new_AGEMA_signal_3620 ;
    wire new_AGEMA_signal_3621 ;
    wire new_AGEMA_signal_3622 ;
    wire new_AGEMA_signal_3623 ;
    wire new_AGEMA_signal_3624 ;
    wire new_AGEMA_signal_3625 ;
    wire new_AGEMA_signal_3626 ;
    wire new_AGEMA_signal_3627 ;
    wire new_AGEMA_signal_3628 ;
    wire new_AGEMA_signal_3629 ;
    wire new_AGEMA_signal_3630 ;
    wire new_AGEMA_signal_3631 ;
    wire new_AGEMA_signal_3632 ;
    wire new_AGEMA_signal_3633 ;
    wire new_AGEMA_signal_3634 ;
    wire new_AGEMA_signal_3635 ;
    wire new_AGEMA_signal_3636 ;
    wire new_AGEMA_signal_3637 ;
    wire new_AGEMA_signal_3638 ;
    wire new_AGEMA_signal_3639 ;
    wire new_AGEMA_signal_3640 ;
    wire new_AGEMA_signal_3641 ;
    wire new_AGEMA_signal_3642 ;
    wire new_AGEMA_signal_3643 ;
    wire new_AGEMA_signal_3644 ;
    wire new_AGEMA_signal_3645 ;
    wire new_AGEMA_signal_3646 ;
    wire new_AGEMA_signal_3647 ;
    wire new_AGEMA_signal_3648 ;
    wire new_AGEMA_signal_3649 ;
    wire new_AGEMA_signal_3650 ;
    wire new_AGEMA_signal_3651 ;
    wire new_AGEMA_signal_3652 ;
    wire new_AGEMA_signal_3653 ;
    wire new_AGEMA_signal_3654 ;
    wire new_AGEMA_signal_3655 ;
    wire new_AGEMA_signal_3656 ;
    wire new_AGEMA_signal_3657 ;
    wire new_AGEMA_signal_3658 ;
    wire new_AGEMA_signal_3659 ;
    wire new_AGEMA_signal_3660 ;
    wire new_AGEMA_signal_3661 ;
    wire new_AGEMA_signal_3662 ;
    wire new_AGEMA_signal_3663 ;
    wire new_AGEMA_signal_3664 ;
    wire new_AGEMA_signal_3665 ;
    wire new_AGEMA_signal_3666 ;
    wire new_AGEMA_signal_3667 ;
    wire new_AGEMA_signal_3668 ;
    wire new_AGEMA_signal_3669 ;
    wire new_AGEMA_signal_3670 ;
    wire new_AGEMA_signal_3671 ;
    wire new_AGEMA_signal_3672 ;
    wire new_AGEMA_signal_3673 ;
    wire new_AGEMA_signal_3674 ;
    wire new_AGEMA_signal_3675 ;
    wire new_AGEMA_signal_3676 ;
    wire new_AGEMA_signal_3677 ;
    wire new_AGEMA_signal_3678 ;
    wire new_AGEMA_signal_3679 ;
    wire new_AGEMA_signal_3680 ;
    wire new_AGEMA_signal_3681 ;
    wire new_AGEMA_signal_3682 ;
    wire new_AGEMA_signal_3683 ;
    wire new_AGEMA_signal_3684 ;
    wire new_AGEMA_signal_3685 ;
    wire new_AGEMA_signal_3686 ;
    wire new_AGEMA_signal_3687 ;
    wire new_AGEMA_signal_3688 ;
    wire new_AGEMA_signal_3689 ;
    wire new_AGEMA_signal_3690 ;
    wire new_AGEMA_signal_3691 ;
    wire new_AGEMA_signal_3692 ;
    wire new_AGEMA_signal_3693 ;
    wire new_AGEMA_signal_3694 ;
    wire new_AGEMA_signal_3695 ;
    wire new_AGEMA_signal_3696 ;
    wire new_AGEMA_signal_3697 ;
    wire new_AGEMA_signal_3698 ;
    wire new_AGEMA_signal_3699 ;
    wire new_AGEMA_signal_3700 ;
    wire new_AGEMA_signal_3701 ;
    wire new_AGEMA_signal_3702 ;
    wire new_AGEMA_signal_3703 ;
    wire new_AGEMA_signal_3704 ;
    wire new_AGEMA_signal_3705 ;
    wire new_AGEMA_signal_3706 ;
    wire new_AGEMA_signal_3707 ;
    wire new_AGEMA_signal_3708 ;
    wire new_AGEMA_signal_3709 ;
    wire new_AGEMA_signal_3710 ;
    wire new_AGEMA_signal_3711 ;
    wire new_AGEMA_signal_3712 ;
    wire new_AGEMA_signal_3713 ;
    wire new_AGEMA_signal_3714 ;
    wire new_AGEMA_signal_3715 ;
    wire new_AGEMA_signal_3716 ;
    wire new_AGEMA_signal_3717 ;
    wire new_AGEMA_signal_3718 ;
    wire new_AGEMA_signal_3719 ;
    wire new_AGEMA_signal_3720 ;
    wire new_AGEMA_signal_3721 ;
    wire new_AGEMA_signal_3722 ;
    wire new_AGEMA_signal_3723 ;
    wire new_AGEMA_signal_3724 ;
    wire new_AGEMA_signal_3725 ;
    wire new_AGEMA_signal_3726 ;
    wire new_AGEMA_signal_3727 ;
    wire new_AGEMA_signal_3728 ;
    wire new_AGEMA_signal_3729 ;
    wire new_AGEMA_signal_3730 ;
    wire new_AGEMA_signal_3731 ;
    wire new_AGEMA_signal_3732 ;
    wire new_AGEMA_signal_3733 ;
    wire new_AGEMA_signal_3734 ;
    wire new_AGEMA_signal_3735 ;
    wire new_AGEMA_signal_3736 ;
    wire new_AGEMA_signal_3737 ;
    wire new_AGEMA_signal_3738 ;
    wire new_AGEMA_signal_3739 ;
    wire new_AGEMA_signal_3740 ;
    wire new_AGEMA_signal_3741 ;
    wire new_AGEMA_signal_3742 ;
    wire new_AGEMA_signal_3743 ;
    wire new_AGEMA_signal_3744 ;
    wire new_AGEMA_signal_3745 ;
    wire new_AGEMA_signal_3746 ;
    wire new_AGEMA_signal_3747 ;
    wire new_AGEMA_signal_3748 ;
    wire new_AGEMA_signal_3749 ;
    wire new_AGEMA_signal_3750 ;
    wire new_AGEMA_signal_3751 ;
    wire new_AGEMA_signal_3752 ;
    wire new_AGEMA_signal_3753 ;
    wire new_AGEMA_signal_3754 ;
    wire new_AGEMA_signal_3755 ;
    wire new_AGEMA_signal_3756 ;
    wire new_AGEMA_signal_3757 ;
    wire new_AGEMA_signal_3758 ;
    wire new_AGEMA_signal_3759 ;
    wire new_AGEMA_signal_3760 ;
    wire new_AGEMA_signal_3761 ;
    wire new_AGEMA_signal_3762 ;
    wire new_AGEMA_signal_3763 ;
    wire new_AGEMA_signal_3764 ;
    wire new_AGEMA_signal_3765 ;
    wire new_AGEMA_signal_3766 ;
    wire new_AGEMA_signal_3767 ;
    wire new_AGEMA_signal_3768 ;
    wire new_AGEMA_signal_3769 ;
    wire new_AGEMA_signal_3770 ;
    wire new_AGEMA_signal_3771 ;
    wire new_AGEMA_signal_3772 ;
    wire new_AGEMA_signal_3773 ;
    wire new_AGEMA_signal_3774 ;
    wire new_AGEMA_signal_3775 ;
    wire new_AGEMA_signal_3776 ;
    wire new_AGEMA_signal_3777 ;
    wire new_AGEMA_signal_3778 ;
    wire new_AGEMA_signal_3779 ;
    wire new_AGEMA_signal_3780 ;
    wire new_AGEMA_signal_3781 ;
    wire new_AGEMA_signal_3782 ;
    wire new_AGEMA_signal_3783 ;
    wire new_AGEMA_signal_3784 ;
    wire new_AGEMA_signal_3785 ;
    wire new_AGEMA_signal_3786 ;
    wire new_AGEMA_signal_3787 ;
    wire new_AGEMA_signal_3788 ;
    wire new_AGEMA_signal_3789 ;
    wire new_AGEMA_signal_3790 ;
    wire new_AGEMA_signal_3791 ;
    wire new_AGEMA_signal_3792 ;
    wire new_AGEMA_signal_3793 ;
    wire new_AGEMA_signal_3794 ;
    wire new_AGEMA_signal_3795 ;
    wire new_AGEMA_signal_3796 ;
    wire new_AGEMA_signal_3797 ;
    wire new_AGEMA_signal_3798 ;
    wire new_AGEMA_signal_3799 ;
    wire new_AGEMA_signal_3800 ;
    wire new_AGEMA_signal_3801 ;
    wire new_AGEMA_signal_3802 ;
    wire new_AGEMA_signal_3803 ;
    wire new_AGEMA_signal_3804 ;
    wire new_AGEMA_signal_3805 ;
    wire new_AGEMA_signal_3806 ;
    wire new_AGEMA_signal_3807 ;
    wire new_AGEMA_signal_3808 ;
    wire new_AGEMA_signal_3809 ;
    wire new_AGEMA_signal_3810 ;
    wire new_AGEMA_signal_3811 ;
    wire new_AGEMA_signal_3812 ;
    wire new_AGEMA_signal_3813 ;
    wire new_AGEMA_signal_3814 ;
    wire new_AGEMA_signal_3815 ;
    wire new_AGEMA_signal_3816 ;
    wire new_AGEMA_signal_3817 ;
    wire new_AGEMA_signal_3818 ;
    wire new_AGEMA_signal_3819 ;
    wire new_AGEMA_signal_3820 ;
    wire new_AGEMA_signal_3821 ;
    wire new_AGEMA_signal_3822 ;
    wire new_AGEMA_signal_3823 ;
    wire new_AGEMA_signal_3824 ;
    wire new_AGEMA_signal_3825 ;
    wire new_AGEMA_signal_3826 ;
    wire new_AGEMA_signal_3827 ;
    wire new_AGEMA_signal_3828 ;
    wire new_AGEMA_signal_3829 ;
    wire new_AGEMA_signal_3830 ;
    wire new_AGEMA_signal_3831 ;
    wire new_AGEMA_signal_3832 ;
    wire new_AGEMA_signal_3833 ;
    wire new_AGEMA_signal_3834 ;
    wire new_AGEMA_signal_3835 ;
    wire new_AGEMA_signal_3836 ;
    wire new_AGEMA_signal_3837 ;
    wire new_AGEMA_signal_3838 ;
    wire new_AGEMA_signal_3839 ;
    wire new_AGEMA_signal_3840 ;
    wire new_AGEMA_signal_3841 ;
    wire new_AGEMA_signal_3842 ;
    wire new_AGEMA_signal_3843 ;
    wire new_AGEMA_signal_3844 ;
    wire new_AGEMA_signal_3845 ;
    wire new_AGEMA_signal_3846 ;
    wire new_AGEMA_signal_3847 ;
    wire new_AGEMA_signal_3848 ;
    wire new_AGEMA_signal_3849 ;
    wire new_AGEMA_signal_3850 ;
    wire new_AGEMA_signal_3851 ;
    wire new_AGEMA_signal_3852 ;
    wire new_AGEMA_signal_3853 ;
    wire new_AGEMA_signal_3854 ;
    wire new_AGEMA_signal_3855 ;
    wire new_AGEMA_signal_3856 ;
    wire new_AGEMA_signal_3857 ;
    wire new_AGEMA_signal_3858 ;
    wire new_AGEMA_signal_3859 ;
    wire new_AGEMA_signal_3860 ;
    wire new_AGEMA_signal_3861 ;
    wire new_AGEMA_signal_3862 ;
    wire new_AGEMA_signal_3863 ;
    wire new_AGEMA_signal_3864 ;
    wire new_AGEMA_signal_3865 ;
    wire new_AGEMA_signal_3866 ;
    wire new_AGEMA_signal_3867 ;
    wire new_AGEMA_signal_3868 ;
    wire new_AGEMA_signal_3869 ;
    wire new_AGEMA_signal_3870 ;
    wire new_AGEMA_signal_3871 ;
    wire new_AGEMA_signal_3872 ;
    wire new_AGEMA_signal_3873 ;
    wire new_AGEMA_signal_3874 ;
    wire new_AGEMA_signal_3875 ;
    wire new_AGEMA_signal_3876 ;
    wire new_AGEMA_signal_3877 ;
    wire new_AGEMA_signal_3878 ;
    wire new_AGEMA_signal_3879 ;
    wire new_AGEMA_signal_3880 ;
    wire new_AGEMA_signal_3881 ;
    wire new_AGEMA_signal_3882 ;
    wire new_AGEMA_signal_3883 ;
    wire new_AGEMA_signal_3884 ;
    wire new_AGEMA_signal_3885 ;
    wire new_AGEMA_signal_3886 ;
    wire new_AGEMA_signal_3887 ;
    wire new_AGEMA_signal_3888 ;
    wire new_AGEMA_signal_3889 ;
    wire new_AGEMA_signal_3890 ;
    wire new_AGEMA_signal_3891 ;
    wire new_AGEMA_signal_3892 ;
    wire new_AGEMA_signal_3893 ;
    wire new_AGEMA_signal_3894 ;
    wire new_AGEMA_signal_3895 ;
    wire new_AGEMA_signal_3896 ;
    wire new_AGEMA_signal_3897 ;
    wire new_AGEMA_signal_3898 ;
    wire new_AGEMA_signal_3899 ;
    wire new_AGEMA_signal_3900 ;
    wire new_AGEMA_signal_3901 ;
    wire new_AGEMA_signal_3902 ;
    wire new_AGEMA_signal_3903 ;
    wire new_AGEMA_signal_3904 ;
    wire new_AGEMA_signal_3905 ;
    wire new_AGEMA_signal_3906 ;
    wire new_AGEMA_signal_3907 ;
    wire new_AGEMA_signal_3908 ;
    wire new_AGEMA_signal_3909 ;
    wire new_AGEMA_signal_3910 ;
    wire new_AGEMA_signal_3911 ;
    wire new_AGEMA_signal_3912 ;
    wire new_AGEMA_signal_3913 ;
    wire new_AGEMA_signal_3914 ;
    wire new_AGEMA_signal_3915 ;
    wire new_AGEMA_signal_3916 ;
    wire new_AGEMA_signal_3917 ;
    wire new_AGEMA_signal_3918 ;
    wire new_AGEMA_signal_3919 ;
    wire new_AGEMA_signal_3920 ;
    wire new_AGEMA_signal_3921 ;
    wire new_AGEMA_signal_3922 ;
    wire new_AGEMA_signal_3923 ;
    wire new_AGEMA_signal_3924 ;
    wire new_AGEMA_signal_3925 ;
    wire new_AGEMA_signal_3926 ;
    wire new_AGEMA_signal_3927 ;
    wire new_AGEMA_signal_3928 ;
    wire new_AGEMA_signal_3929 ;
    wire new_AGEMA_signal_3930 ;
    wire new_AGEMA_signal_3931 ;
    wire new_AGEMA_signal_3932 ;
    wire new_AGEMA_signal_3933 ;
    wire new_AGEMA_signal_3934 ;
    wire new_AGEMA_signal_3935 ;
    wire new_AGEMA_signal_3936 ;
    wire new_AGEMA_signal_3937 ;
    wire new_AGEMA_signal_3938 ;
    wire new_AGEMA_signal_3939 ;
    wire new_AGEMA_signal_3940 ;
    wire new_AGEMA_signal_3941 ;
    wire new_AGEMA_signal_3942 ;
    wire new_AGEMA_signal_3943 ;
    wire new_AGEMA_signal_3944 ;
    wire new_AGEMA_signal_3945 ;
    wire new_AGEMA_signal_3946 ;
    wire new_AGEMA_signal_3947 ;
    wire new_AGEMA_signal_3948 ;
    wire new_AGEMA_signal_3949 ;
    wire new_AGEMA_signal_3950 ;
    wire new_AGEMA_signal_3951 ;
    wire new_AGEMA_signal_3952 ;
    wire new_AGEMA_signal_3953 ;
    wire new_AGEMA_signal_3954 ;
    wire new_AGEMA_signal_3955 ;
    wire new_AGEMA_signal_3956 ;
    wire new_AGEMA_signal_3957 ;
    wire new_AGEMA_signal_3958 ;
    wire new_AGEMA_signal_3959 ;
    wire new_AGEMA_signal_3960 ;
    wire new_AGEMA_signal_3961 ;
    wire new_AGEMA_signal_3962 ;
    wire new_AGEMA_signal_3963 ;
    wire new_AGEMA_signal_3964 ;
    wire new_AGEMA_signal_3965 ;
    wire new_AGEMA_signal_3966 ;
    wire new_AGEMA_signal_3967 ;
    wire new_AGEMA_signal_3968 ;
    wire new_AGEMA_signal_3969 ;
    wire new_AGEMA_signal_3970 ;
    wire new_AGEMA_signal_3971 ;
    wire new_AGEMA_signal_3972 ;
    wire new_AGEMA_signal_3973 ;
    wire new_AGEMA_signal_3974 ;
    wire new_AGEMA_signal_3975 ;
    wire new_AGEMA_signal_3976 ;
    wire new_AGEMA_signal_3977 ;
    wire new_AGEMA_signal_3978 ;
    wire new_AGEMA_signal_3979 ;
    wire new_AGEMA_signal_3980 ;
    wire new_AGEMA_signal_3981 ;
    wire new_AGEMA_signal_3982 ;
    wire new_AGEMA_signal_3983 ;
    wire new_AGEMA_signal_3984 ;
    wire new_AGEMA_signal_3985 ;
    wire new_AGEMA_signal_3986 ;
    wire new_AGEMA_signal_3987 ;
    wire new_AGEMA_signal_3988 ;
    wire new_AGEMA_signal_3989 ;
    wire new_AGEMA_signal_3990 ;
    wire new_AGEMA_signal_3991 ;
    wire new_AGEMA_signal_3992 ;
    wire new_AGEMA_signal_3993 ;
    wire new_AGEMA_signal_3994 ;
    wire new_AGEMA_signal_3995 ;
    wire new_AGEMA_signal_3996 ;
    wire new_AGEMA_signal_3997 ;
    wire new_AGEMA_signal_3998 ;
    wire new_AGEMA_signal_3999 ;
    wire new_AGEMA_signal_4000 ;
    wire new_AGEMA_signal_4001 ;
    wire new_AGEMA_signal_4002 ;
    wire new_AGEMA_signal_4003 ;
    wire new_AGEMA_signal_4004 ;
    wire new_AGEMA_signal_4005 ;
    wire new_AGEMA_signal_4006 ;
    wire new_AGEMA_signal_4007 ;
    wire new_AGEMA_signal_4008 ;
    wire new_AGEMA_signal_4009 ;
    wire new_AGEMA_signal_4010 ;
    wire new_AGEMA_signal_4011 ;
    wire new_AGEMA_signal_4012 ;
    wire new_AGEMA_signal_4013 ;
    wire new_AGEMA_signal_4014 ;
    wire new_AGEMA_signal_4015 ;
    wire new_AGEMA_signal_4016 ;
    wire new_AGEMA_signal_4017 ;
    wire new_AGEMA_signal_4018 ;
    wire new_AGEMA_signal_4019 ;
    wire new_AGEMA_signal_4020 ;
    wire new_AGEMA_signal_4021 ;
    wire new_AGEMA_signal_4022 ;
    wire new_AGEMA_signal_4023 ;
    wire new_AGEMA_signal_4024 ;
    wire new_AGEMA_signal_4025 ;
    wire new_AGEMA_signal_4026 ;
    wire new_AGEMA_signal_4027 ;
    wire new_AGEMA_signal_4028 ;
    wire new_AGEMA_signal_4029 ;
    wire new_AGEMA_signal_4030 ;
    wire new_AGEMA_signal_4031 ;
    wire new_AGEMA_signal_4032 ;
    wire new_AGEMA_signal_4033 ;
    wire new_AGEMA_signal_4034 ;
    wire new_AGEMA_signal_4035 ;
    wire new_AGEMA_signal_4036 ;
    wire new_AGEMA_signal_4037 ;
    wire new_AGEMA_signal_4038 ;
    wire new_AGEMA_signal_4039 ;
    wire new_AGEMA_signal_4040 ;
    wire new_AGEMA_signal_4041 ;
    wire new_AGEMA_signal_4042 ;
    wire new_AGEMA_signal_4043 ;
    wire new_AGEMA_signal_4044 ;
    wire new_AGEMA_signal_4045 ;
    wire new_AGEMA_signal_4046 ;
    wire new_AGEMA_signal_4047 ;
    wire new_AGEMA_signal_4048 ;
    wire new_AGEMA_signal_4049 ;
    wire new_AGEMA_signal_4050 ;
    wire new_AGEMA_signal_4051 ;
    wire new_AGEMA_signal_4052 ;
    wire new_AGEMA_signal_4053 ;
    wire new_AGEMA_signal_4054 ;
    wire new_AGEMA_signal_4055 ;
    wire new_AGEMA_signal_4056 ;
    wire new_AGEMA_signal_4057 ;
    wire new_AGEMA_signal_4058 ;
    wire new_AGEMA_signal_4059 ;
    wire new_AGEMA_signal_4060 ;
    wire new_AGEMA_signal_4061 ;
    wire new_AGEMA_signal_4062 ;
    wire new_AGEMA_signal_4063 ;
    wire new_AGEMA_signal_4064 ;
    wire new_AGEMA_signal_4065 ;
    wire new_AGEMA_signal_4066 ;
    wire new_AGEMA_signal_4067 ;
    wire new_AGEMA_signal_4068 ;
    wire new_AGEMA_signal_4069 ;
    wire new_AGEMA_signal_4070 ;
    wire new_AGEMA_signal_4071 ;
    wire new_AGEMA_signal_4072 ;
    wire new_AGEMA_signal_4073 ;
    wire new_AGEMA_signal_4074 ;
    wire new_AGEMA_signal_4075 ;
    wire new_AGEMA_signal_4076 ;
    wire new_AGEMA_signal_4077 ;
    wire new_AGEMA_signal_4078 ;
    wire new_AGEMA_signal_4079 ;
    wire new_AGEMA_signal_4080 ;
    wire new_AGEMA_signal_4081 ;
    wire new_AGEMA_signal_4082 ;
    wire new_AGEMA_signal_4083 ;
    wire new_AGEMA_signal_4084 ;
    wire new_AGEMA_signal_4085 ;
    wire new_AGEMA_signal_4086 ;
    wire new_AGEMA_signal_4087 ;
    wire new_AGEMA_signal_4088 ;
    wire new_AGEMA_signal_4089 ;
    wire new_AGEMA_signal_4090 ;
    wire new_AGEMA_signal_4091 ;
    wire new_AGEMA_signal_4092 ;
    wire new_AGEMA_signal_4093 ;
    wire new_AGEMA_signal_4094 ;
    wire new_AGEMA_signal_4095 ;
    wire new_AGEMA_signal_4096 ;
    wire new_AGEMA_signal_4097 ;
    wire new_AGEMA_signal_4098 ;
    wire new_AGEMA_signal_4099 ;
    wire new_AGEMA_signal_4100 ;
    wire new_AGEMA_signal_4101 ;
    wire new_AGEMA_signal_4102 ;
    wire new_AGEMA_signal_4103 ;
    wire new_AGEMA_signal_4104 ;
    wire new_AGEMA_signal_4105 ;
    wire new_AGEMA_signal_4106 ;
    wire new_AGEMA_signal_4107 ;
    wire new_AGEMA_signal_4108 ;
    wire new_AGEMA_signal_4109 ;
    wire new_AGEMA_signal_4110 ;
    wire new_AGEMA_signal_4111 ;
    wire new_AGEMA_signal_4112 ;
    wire new_AGEMA_signal_4113 ;
    wire new_AGEMA_signal_4114 ;
    wire new_AGEMA_signal_4115 ;
    wire new_AGEMA_signal_4116 ;
    wire new_AGEMA_signal_4117 ;
    wire new_AGEMA_signal_4118 ;
    wire new_AGEMA_signal_4119 ;
    wire new_AGEMA_signal_4120 ;
    wire new_AGEMA_signal_4121 ;
    wire new_AGEMA_signal_4122 ;
    wire new_AGEMA_signal_4123 ;
    wire new_AGEMA_signal_4124 ;
    wire new_AGEMA_signal_4125 ;
    wire new_AGEMA_signal_4126 ;
    wire new_AGEMA_signal_4127 ;
    wire new_AGEMA_signal_4128 ;
    wire new_AGEMA_signal_4129 ;
    wire new_AGEMA_signal_4130 ;
    wire new_AGEMA_signal_4131 ;
    wire new_AGEMA_signal_4132 ;
    wire new_AGEMA_signal_4133 ;
    wire new_AGEMA_signal_4134 ;
    wire new_AGEMA_signal_4135 ;
    wire new_AGEMA_signal_4136 ;
    wire new_AGEMA_signal_4137 ;
    wire new_AGEMA_signal_4138 ;
    wire new_AGEMA_signal_4139 ;
    wire new_AGEMA_signal_4140 ;
    wire new_AGEMA_signal_4141 ;
    wire new_AGEMA_signal_4142 ;
    wire new_AGEMA_signal_4143 ;
    wire new_AGEMA_signal_4144 ;
    wire new_AGEMA_signal_4145 ;
    wire new_AGEMA_signal_4146 ;
    wire new_AGEMA_signal_4147 ;
    wire new_AGEMA_signal_4148 ;
    wire new_AGEMA_signal_4149 ;
    wire new_AGEMA_signal_4150 ;
    wire new_AGEMA_signal_4151 ;
    wire new_AGEMA_signal_4152 ;
    wire new_AGEMA_signal_4153 ;
    wire new_AGEMA_signal_4154 ;
    wire new_AGEMA_signal_4155 ;
    wire new_AGEMA_signal_4156 ;
    wire new_AGEMA_signal_4157 ;
    wire new_AGEMA_signal_4158 ;
    wire new_AGEMA_signal_4159 ;
    wire new_AGEMA_signal_4160 ;
    wire new_AGEMA_signal_4161 ;
    wire new_AGEMA_signal_4162 ;
    wire new_AGEMA_signal_4163 ;
    wire new_AGEMA_signal_4164 ;
    wire new_AGEMA_signal_4165 ;
    wire new_AGEMA_signal_4166 ;
    wire new_AGEMA_signal_4167 ;
    wire new_AGEMA_signal_4168 ;
    wire new_AGEMA_signal_4169 ;
    wire new_AGEMA_signal_4170 ;
    wire new_AGEMA_signal_4171 ;
    wire new_AGEMA_signal_4172 ;
    wire new_AGEMA_signal_4173 ;
    wire new_AGEMA_signal_4174 ;
    wire new_AGEMA_signal_4175 ;
    wire new_AGEMA_signal_4176 ;
    wire new_AGEMA_signal_4177 ;
    wire new_AGEMA_signal_4178 ;
    wire new_AGEMA_signal_4179 ;
    wire new_AGEMA_signal_4180 ;
    wire new_AGEMA_signal_4181 ;
    wire new_AGEMA_signal_4182 ;
    wire new_AGEMA_signal_4183 ;
    wire new_AGEMA_signal_4184 ;
    wire new_AGEMA_signal_4185 ;
    wire new_AGEMA_signal_4186 ;
    wire new_AGEMA_signal_4187 ;
    wire new_AGEMA_signal_4188 ;
    wire new_AGEMA_signal_4189 ;
    wire new_AGEMA_signal_4190 ;
    wire new_AGEMA_signal_4191 ;
    wire new_AGEMA_signal_4192 ;
    wire new_AGEMA_signal_4193 ;
    wire new_AGEMA_signal_4194 ;
    wire new_AGEMA_signal_4195 ;
    wire new_AGEMA_signal_4196 ;
    wire new_AGEMA_signal_4197 ;
    wire new_AGEMA_signal_4198 ;
    wire new_AGEMA_signal_4199 ;
    wire new_AGEMA_signal_4200 ;
    wire new_AGEMA_signal_4201 ;
    wire new_AGEMA_signal_4202 ;
    wire new_AGEMA_signal_4203 ;
    wire new_AGEMA_signal_4204 ;
    wire new_AGEMA_signal_4205 ;
    wire new_AGEMA_signal_4206 ;
    wire new_AGEMA_signal_4207 ;
    wire new_AGEMA_signal_4208 ;
    wire new_AGEMA_signal_4209 ;
    wire new_AGEMA_signal_4210 ;
    wire new_AGEMA_signal_4211 ;
    wire new_AGEMA_signal_4212 ;
    wire new_AGEMA_signal_4213 ;
    wire new_AGEMA_signal_4214 ;
    wire new_AGEMA_signal_4215 ;
    wire new_AGEMA_signal_4216 ;
    wire new_AGEMA_signal_4217 ;
    wire new_AGEMA_signal_4218 ;
    wire new_AGEMA_signal_4219 ;
    wire new_AGEMA_signal_4220 ;
    wire new_AGEMA_signal_4221 ;
    wire new_AGEMA_signal_4222 ;
    wire new_AGEMA_signal_4223 ;
    wire new_AGEMA_signal_4224 ;
    wire new_AGEMA_signal_4225 ;
    wire new_AGEMA_signal_4226 ;
    wire new_AGEMA_signal_4227 ;
    wire new_AGEMA_signal_4228 ;
    wire new_AGEMA_signal_4229 ;
    wire new_AGEMA_signal_4230 ;
    wire new_AGEMA_signal_4231 ;
    wire new_AGEMA_signal_4232 ;
    wire new_AGEMA_signal_4233 ;
    wire new_AGEMA_signal_4234 ;
    wire new_AGEMA_signal_4235 ;
    wire new_AGEMA_signal_4236 ;
    wire new_AGEMA_signal_4237 ;
    wire new_AGEMA_signal_4238 ;
    wire new_AGEMA_signal_4239 ;
    wire new_AGEMA_signal_4240 ;
    wire new_AGEMA_signal_4241 ;
    wire new_AGEMA_signal_4242 ;
    wire new_AGEMA_signal_4243 ;
    wire new_AGEMA_signal_4244 ;
    wire new_AGEMA_signal_4245 ;
    wire new_AGEMA_signal_4246 ;
    wire new_AGEMA_signal_4247 ;
    wire new_AGEMA_signal_4248 ;
    wire new_AGEMA_signal_4249 ;
    wire new_AGEMA_signal_4250 ;
    wire new_AGEMA_signal_4251 ;
    wire new_AGEMA_signal_4252 ;
    wire new_AGEMA_signal_4253 ;
    wire new_AGEMA_signal_4254 ;
    wire new_AGEMA_signal_4255 ;
    wire new_AGEMA_signal_4256 ;
    wire new_AGEMA_signal_4257 ;
    wire new_AGEMA_signal_4258 ;
    wire new_AGEMA_signal_4259 ;
    wire new_AGEMA_signal_4260 ;
    wire new_AGEMA_signal_4261 ;
    wire new_AGEMA_signal_4262 ;
    wire new_AGEMA_signal_4263 ;
    wire new_AGEMA_signal_4264 ;
    wire new_AGEMA_signal_4265 ;
    wire new_AGEMA_signal_4266 ;
    wire new_AGEMA_signal_4267 ;
    wire new_AGEMA_signal_4268 ;
    wire new_AGEMA_signal_4269 ;
    wire new_AGEMA_signal_4270 ;
    wire new_AGEMA_signal_4271 ;
    wire new_AGEMA_signal_4272 ;
    wire new_AGEMA_signal_4273 ;
    wire new_AGEMA_signal_4274 ;
    wire new_AGEMA_signal_4275 ;
    wire new_AGEMA_signal_4276 ;
    wire new_AGEMA_signal_4277 ;
    wire new_AGEMA_signal_4278 ;
    wire new_AGEMA_signal_4279 ;
    wire new_AGEMA_signal_4280 ;
    wire new_AGEMA_signal_4281 ;
    wire new_AGEMA_signal_4282 ;
    wire new_AGEMA_signal_4283 ;
    wire new_AGEMA_signal_4284 ;
    wire new_AGEMA_signal_4285 ;
    wire new_AGEMA_signal_4286 ;
    wire new_AGEMA_signal_4287 ;
    wire new_AGEMA_signal_4288 ;
    wire new_AGEMA_signal_4289 ;
    wire new_AGEMA_signal_4290 ;
    wire new_AGEMA_signal_4291 ;
    wire new_AGEMA_signal_4292 ;
    wire new_AGEMA_signal_4293 ;
    wire new_AGEMA_signal_4294 ;
    wire new_AGEMA_signal_4295 ;
    wire new_AGEMA_signal_4296 ;
    wire new_AGEMA_signal_4297 ;
    wire new_AGEMA_signal_4298 ;
    wire new_AGEMA_signal_4299 ;
    wire new_AGEMA_signal_4300 ;
    wire new_AGEMA_signal_4301 ;
    wire new_AGEMA_signal_4302 ;
    wire new_AGEMA_signal_4303 ;
    wire new_AGEMA_signal_4304 ;
    wire new_AGEMA_signal_4305 ;
    wire new_AGEMA_signal_4306 ;
    wire new_AGEMA_signal_4307 ;
    wire new_AGEMA_signal_4308 ;
    wire new_AGEMA_signal_4309 ;
    wire new_AGEMA_signal_4310 ;
    wire new_AGEMA_signal_4311 ;
    wire new_AGEMA_signal_4312 ;
    wire new_AGEMA_signal_4313 ;
    wire new_AGEMA_signal_4314 ;
    wire new_AGEMA_signal_4315 ;
    wire new_AGEMA_signal_4316 ;
    wire new_AGEMA_signal_4317 ;
    wire new_AGEMA_signal_4318 ;
    wire new_AGEMA_signal_4319 ;
    wire new_AGEMA_signal_4320 ;
    wire new_AGEMA_signal_4321 ;
    wire new_AGEMA_signal_4322 ;
    wire new_AGEMA_signal_4323 ;
    wire new_AGEMA_signal_4324 ;
    wire new_AGEMA_signal_4325 ;
    wire new_AGEMA_signal_4326 ;
    wire new_AGEMA_signal_4327 ;
    wire new_AGEMA_signal_4328 ;
    wire new_AGEMA_signal_4329 ;
    wire new_AGEMA_signal_4330 ;
    wire new_AGEMA_signal_4331 ;
    wire new_AGEMA_signal_4332 ;
    wire new_AGEMA_signal_4333 ;
    wire new_AGEMA_signal_4334 ;
    wire new_AGEMA_signal_4335 ;
    wire new_AGEMA_signal_4336 ;
    wire new_AGEMA_signal_4337 ;
    wire new_AGEMA_signal_4338 ;
    wire new_AGEMA_signal_4339 ;
    wire new_AGEMA_signal_4340 ;
    wire new_AGEMA_signal_4341 ;
    wire new_AGEMA_signal_4342 ;
    wire new_AGEMA_signal_4343 ;
    wire new_AGEMA_signal_4344 ;
    wire new_AGEMA_signal_4345 ;
    wire new_AGEMA_signal_4346 ;
    wire new_AGEMA_signal_4347 ;
    wire new_AGEMA_signal_4348 ;
    wire new_AGEMA_signal_4349 ;
    wire new_AGEMA_signal_4350 ;
    wire new_AGEMA_signal_4351 ;
    wire new_AGEMA_signal_4352 ;
    wire new_AGEMA_signal_4353 ;
    wire new_AGEMA_signal_4354 ;
    wire new_AGEMA_signal_4355 ;
    wire new_AGEMA_signal_4356 ;
    wire new_AGEMA_signal_4357 ;
    wire new_AGEMA_signal_4358 ;
    wire new_AGEMA_signal_4359 ;
    wire new_AGEMA_signal_4360 ;
    wire new_AGEMA_signal_4361 ;
    wire new_AGEMA_signal_4362 ;
    wire new_AGEMA_signal_4363 ;
    wire new_AGEMA_signal_4364 ;
    wire new_AGEMA_signal_4365 ;
    wire new_AGEMA_signal_4366 ;
    wire new_AGEMA_signal_4367 ;
    wire new_AGEMA_signal_4368 ;
    wire new_AGEMA_signal_4369 ;
    wire new_AGEMA_signal_4370 ;
    wire new_AGEMA_signal_4371 ;
    wire new_AGEMA_signal_4372 ;
    wire new_AGEMA_signal_4373 ;
    wire new_AGEMA_signal_4374 ;
    wire new_AGEMA_signal_4375 ;
    wire new_AGEMA_signal_4376 ;
    wire new_AGEMA_signal_4377 ;
    wire new_AGEMA_signal_4378 ;
    wire new_AGEMA_signal_4379 ;
    wire new_AGEMA_signal_4380 ;
    wire new_AGEMA_signal_4381 ;
    wire new_AGEMA_signal_4382 ;
    wire new_AGEMA_signal_4383 ;
    wire new_AGEMA_signal_4384 ;
    wire new_AGEMA_signal_4385 ;
    wire new_AGEMA_signal_4386 ;
    wire new_AGEMA_signal_4387 ;
    wire new_AGEMA_signal_4388 ;
    wire new_AGEMA_signal_4389 ;
    wire new_AGEMA_signal_4390 ;
    wire new_AGEMA_signal_4391 ;
    wire new_AGEMA_signal_4392 ;
    wire new_AGEMA_signal_4393 ;
    wire new_AGEMA_signal_4394 ;
    wire new_AGEMA_signal_4395 ;
    wire new_AGEMA_signal_4396 ;
    wire new_AGEMA_signal_4397 ;
    wire new_AGEMA_signal_4398 ;
    wire new_AGEMA_signal_4399 ;
    wire new_AGEMA_signal_4400 ;
    wire new_AGEMA_signal_4401 ;
    wire new_AGEMA_signal_4402 ;
    wire new_AGEMA_signal_4403 ;
    wire new_AGEMA_signal_4404 ;
    wire new_AGEMA_signal_4405 ;
    wire new_AGEMA_signal_4406 ;
    wire new_AGEMA_signal_4407 ;
    wire new_AGEMA_signal_4408 ;
    wire new_AGEMA_signal_4409 ;
    wire new_AGEMA_signal_4410 ;
    wire new_AGEMA_signal_4411 ;
    wire new_AGEMA_signal_4412 ;
    wire new_AGEMA_signal_4413 ;
    wire new_AGEMA_signal_4414 ;
    wire new_AGEMA_signal_4415 ;
    wire new_AGEMA_signal_4416 ;
    wire new_AGEMA_signal_4417 ;
    wire new_AGEMA_signal_4418 ;
    wire new_AGEMA_signal_4419 ;
    wire new_AGEMA_signal_4420 ;
    wire new_AGEMA_signal_4421 ;
    wire new_AGEMA_signal_4422 ;
    wire new_AGEMA_signal_4423 ;
    wire new_AGEMA_signal_4424 ;
    wire new_AGEMA_signal_4425 ;
    wire new_AGEMA_signal_4426 ;
    wire new_AGEMA_signal_4427 ;
    wire new_AGEMA_signal_4428 ;
    wire new_AGEMA_signal_4429 ;
    wire new_AGEMA_signal_4430 ;
    wire new_AGEMA_signal_4431 ;
    wire new_AGEMA_signal_4432 ;
    wire new_AGEMA_signal_4433 ;
    wire new_AGEMA_signal_4434 ;
    wire new_AGEMA_signal_4435 ;
    wire new_AGEMA_signal_4436 ;
    wire new_AGEMA_signal_4437 ;
    wire new_AGEMA_signal_4438 ;
    wire new_AGEMA_signal_4439 ;
    wire new_AGEMA_signal_4440 ;
    wire new_AGEMA_signal_4441 ;
    wire new_AGEMA_signal_4442 ;
    wire new_AGEMA_signal_4443 ;
    wire new_AGEMA_signal_4444 ;
    wire new_AGEMA_signal_4445 ;
    wire new_AGEMA_signal_4446 ;
    wire new_AGEMA_signal_4447 ;
    wire new_AGEMA_signal_4448 ;
    wire new_AGEMA_signal_4449 ;
    wire new_AGEMA_signal_4450 ;
    wire new_AGEMA_signal_4451 ;
    wire new_AGEMA_signal_4452 ;
    wire new_AGEMA_signal_4453 ;
    wire new_AGEMA_signal_4454 ;
    wire new_AGEMA_signal_4455 ;
    wire new_AGEMA_signal_4456 ;
    wire new_AGEMA_signal_4457 ;
    wire new_AGEMA_signal_4458 ;
    wire new_AGEMA_signal_4459 ;
    wire new_AGEMA_signal_4460 ;
    wire new_AGEMA_signal_4461 ;
    wire new_AGEMA_signal_4462 ;
    wire new_AGEMA_signal_4463 ;
    wire new_AGEMA_signal_4464 ;
    wire new_AGEMA_signal_4465 ;
    wire new_AGEMA_signal_4466 ;
    wire new_AGEMA_signal_4467 ;
    wire new_AGEMA_signal_4468 ;
    wire new_AGEMA_signal_4469 ;
    wire new_AGEMA_signal_4470 ;
    wire new_AGEMA_signal_4471 ;
    wire new_AGEMA_signal_4472 ;
    wire new_AGEMA_signal_4473 ;
    wire new_AGEMA_signal_4474 ;
    wire new_AGEMA_signal_4475 ;
    wire new_AGEMA_signal_4476 ;
    wire new_AGEMA_signal_4477 ;
    wire new_AGEMA_signal_4478 ;
    wire new_AGEMA_signal_4479 ;
    wire new_AGEMA_signal_4480 ;
    wire new_AGEMA_signal_4481 ;
    wire new_AGEMA_signal_4482 ;
    wire new_AGEMA_signal_4483 ;
    wire new_AGEMA_signal_4484 ;
    wire new_AGEMA_signal_4485 ;
    wire new_AGEMA_signal_4486 ;
    wire new_AGEMA_signal_4487 ;
    wire new_AGEMA_signal_4488 ;
    wire new_AGEMA_signal_4489 ;
    wire new_AGEMA_signal_4490 ;
    wire new_AGEMA_signal_4491 ;
    wire new_AGEMA_signal_4492 ;
    wire new_AGEMA_signal_4493 ;
    wire new_AGEMA_signal_4494 ;
    wire new_AGEMA_signal_4495 ;
    wire new_AGEMA_signal_4496 ;
    wire new_AGEMA_signal_4497 ;
    wire new_AGEMA_signal_4498 ;
    wire new_AGEMA_signal_4499 ;
    wire new_AGEMA_signal_4500 ;
    wire new_AGEMA_signal_4501 ;
    wire new_AGEMA_signal_4502 ;
    wire new_AGEMA_signal_4503 ;
    wire new_AGEMA_signal_4504 ;
    wire new_AGEMA_signal_4505 ;
    wire new_AGEMA_signal_4506 ;
    wire new_AGEMA_signal_4507 ;
    wire new_AGEMA_signal_4508 ;
    wire new_AGEMA_signal_4509 ;
    wire new_AGEMA_signal_4510 ;
    wire new_AGEMA_signal_4511 ;
    wire new_AGEMA_signal_4512 ;
    wire new_AGEMA_signal_4513 ;
    wire new_AGEMA_signal_4514 ;
    wire new_AGEMA_signal_4515 ;
    wire new_AGEMA_signal_4516 ;
    wire new_AGEMA_signal_4517 ;
    wire new_AGEMA_signal_4518 ;
    wire new_AGEMA_signal_4519 ;
    wire new_AGEMA_signal_4520 ;
    wire new_AGEMA_signal_4521 ;
    wire new_AGEMA_signal_4522 ;
    wire new_AGEMA_signal_4523 ;
    wire new_AGEMA_signal_4524 ;
    wire new_AGEMA_signal_4525 ;
    wire new_AGEMA_signal_4526 ;
    wire new_AGEMA_signal_4527 ;
    wire new_AGEMA_signal_4528 ;
    wire new_AGEMA_signal_4529 ;
    wire new_AGEMA_signal_4530 ;
    wire new_AGEMA_signal_4531 ;
    wire new_AGEMA_signal_4532 ;
    wire new_AGEMA_signal_4533 ;
    wire new_AGEMA_signal_4534 ;
    wire new_AGEMA_signal_4535 ;
    wire new_AGEMA_signal_4536 ;
    wire new_AGEMA_signal_4537 ;
    wire new_AGEMA_signal_4538 ;
    wire new_AGEMA_signal_4539 ;
    wire new_AGEMA_signal_4540 ;
    wire new_AGEMA_signal_4541 ;
    wire new_AGEMA_signal_4542 ;
    wire new_AGEMA_signal_4543 ;
    wire new_AGEMA_signal_4544 ;
    wire new_AGEMA_signal_4545 ;
    wire new_AGEMA_signal_4546 ;
    wire new_AGEMA_signal_4547 ;
    wire new_AGEMA_signal_4548 ;
    wire new_AGEMA_signal_4549 ;
    wire new_AGEMA_signal_4550 ;
    wire new_AGEMA_signal_4551 ;
    wire new_AGEMA_signal_4552 ;
    wire new_AGEMA_signal_4553 ;
    wire new_AGEMA_signal_4554 ;
    wire new_AGEMA_signal_4555 ;
    wire new_AGEMA_signal_4556 ;
    wire new_AGEMA_signal_4557 ;
    wire new_AGEMA_signal_4558 ;
    wire new_AGEMA_signal_4559 ;
    wire new_AGEMA_signal_4560 ;
    wire new_AGEMA_signal_4561 ;
    wire new_AGEMA_signal_4562 ;
    wire new_AGEMA_signal_4563 ;
    wire new_AGEMA_signal_4564 ;
    wire new_AGEMA_signal_4565 ;
    wire new_AGEMA_signal_4566 ;
    wire new_AGEMA_signal_4567 ;
    wire new_AGEMA_signal_4568 ;
    wire new_AGEMA_signal_4569 ;
    wire new_AGEMA_signal_4570 ;
    wire new_AGEMA_signal_4571 ;
    wire new_AGEMA_signal_4572 ;
    wire new_AGEMA_signal_4573 ;
    wire new_AGEMA_signal_4574 ;
    wire new_AGEMA_signal_4575 ;
    wire new_AGEMA_signal_4576 ;
    wire new_AGEMA_signal_4577 ;
    wire new_AGEMA_signal_4578 ;
    wire new_AGEMA_signal_4579 ;
    wire new_AGEMA_signal_4580 ;
    wire new_AGEMA_signal_4581 ;
    wire new_AGEMA_signal_4582 ;
    wire new_AGEMA_signal_4583 ;
    wire new_AGEMA_signal_4584 ;
    wire new_AGEMA_signal_4585 ;
    wire new_AGEMA_signal_4586 ;
    wire new_AGEMA_signal_4587 ;
    wire new_AGEMA_signal_4588 ;
    wire new_AGEMA_signal_4589 ;
    wire new_AGEMA_signal_4590 ;
    wire new_AGEMA_signal_4591 ;
    wire new_AGEMA_signal_4592 ;
    wire new_AGEMA_signal_4593 ;
    wire new_AGEMA_signal_4594 ;
    wire new_AGEMA_signal_4595 ;
    wire new_AGEMA_signal_4596 ;
    wire new_AGEMA_signal_4597 ;
    wire new_AGEMA_signal_4598 ;
    wire new_AGEMA_signal_4599 ;
    wire new_AGEMA_signal_4600 ;
    wire new_AGEMA_signal_4601 ;
    wire new_AGEMA_signal_4602 ;
    wire new_AGEMA_signal_4603 ;
    wire new_AGEMA_signal_4604 ;
    wire new_AGEMA_signal_4605 ;
    wire new_AGEMA_signal_4606 ;
    wire new_AGEMA_signal_4607 ;
    wire new_AGEMA_signal_4608 ;
    wire new_AGEMA_signal_4609 ;
    wire new_AGEMA_signal_4610 ;
    wire new_AGEMA_signal_4611 ;
    wire new_AGEMA_signal_4612 ;
    wire new_AGEMA_signal_4613 ;
    wire new_AGEMA_signal_4614 ;
    wire new_AGEMA_signal_4615 ;
    wire new_AGEMA_signal_4616 ;
    wire new_AGEMA_signal_4617 ;
    wire new_AGEMA_signal_4618 ;
    wire new_AGEMA_signal_4619 ;
    wire new_AGEMA_signal_4620 ;
    wire new_AGEMA_signal_4621 ;
    wire new_AGEMA_signal_4622 ;
    wire new_AGEMA_signal_4623 ;
    wire new_AGEMA_signal_4624 ;
    wire new_AGEMA_signal_4625 ;
    wire new_AGEMA_signal_4626 ;
    wire new_AGEMA_signal_4627 ;
    wire new_AGEMA_signal_4628 ;
    wire new_AGEMA_signal_4629 ;
    wire new_AGEMA_signal_4630 ;
    wire new_AGEMA_signal_4631 ;
    wire new_AGEMA_signal_4632 ;
    wire new_AGEMA_signal_4633 ;
    wire new_AGEMA_signal_4634 ;
    wire new_AGEMA_signal_4635 ;
    wire new_AGEMA_signal_4636 ;
    wire new_AGEMA_signal_4637 ;
    wire new_AGEMA_signal_4638 ;
    wire new_AGEMA_signal_4639 ;
    wire new_AGEMA_signal_4640 ;
    wire new_AGEMA_signal_4641 ;
    wire new_AGEMA_signal_4642 ;
    wire new_AGEMA_signal_4643 ;
    wire new_AGEMA_signal_4644 ;
    wire new_AGEMA_signal_4645 ;
    wire new_AGEMA_signal_4646 ;
    wire new_AGEMA_signal_4647 ;
    wire new_AGEMA_signal_4648 ;
    wire new_AGEMA_signal_4649 ;
    wire new_AGEMA_signal_4650 ;
    wire new_AGEMA_signal_4651 ;
    wire new_AGEMA_signal_4652 ;
    wire new_AGEMA_signal_4653 ;
    wire new_AGEMA_signal_4654 ;
    wire new_AGEMA_signal_4655 ;
    wire new_AGEMA_signal_4656 ;
    wire new_AGEMA_signal_4657 ;
    wire new_AGEMA_signal_4658 ;
    wire new_AGEMA_signal_4659 ;
    wire new_AGEMA_signal_4660 ;
    wire new_AGEMA_signal_4661 ;
    wire new_AGEMA_signal_4662 ;
    wire new_AGEMA_signal_4663 ;
    wire new_AGEMA_signal_4664 ;
    wire new_AGEMA_signal_4665 ;
    wire new_AGEMA_signal_4666 ;
    wire new_AGEMA_signal_4667 ;
    wire new_AGEMA_signal_4668 ;
    wire new_AGEMA_signal_4669 ;
    wire new_AGEMA_signal_4670 ;
    wire new_AGEMA_signal_4671 ;
    wire new_AGEMA_signal_4672 ;
    wire new_AGEMA_signal_4673 ;
    wire new_AGEMA_signal_4674 ;
    wire new_AGEMA_signal_4675 ;
    wire new_AGEMA_signal_4676 ;
    wire new_AGEMA_signal_4677 ;
    wire new_AGEMA_signal_4678 ;
    wire new_AGEMA_signal_4679 ;
    wire new_AGEMA_signal_4680 ;
    wire new_AGEMA_signal_4681 ;
    wire new_AGEMA_signal_4682 ;
    wire new_AGEMA_signal_4683 ;
    wire new_AGEMA_signal_4684 ;
    wire new_AGEMA_signal_4685 ;
    wire new_AGEMA_signal_4686 ;
    wire new_AGEMA_signal_4687 ;
    wire new_AGEMA_signal_4688 ;
    wire new_AGEMA_signal_4689 ;
    wire new_AGEMA_signal_4690 ;
    wire new_AGEMA_signal_4691 ;
    wire new_AGEMA_signal_4692 ;
    wire new_AGEMA_signal_4693 ;
    wire new_AGEMA_signal_4694 ;
    wire new_AGEMA_signal_4695 ;
    wire new_AGEMA_signal_4696 ;
    wire new_AGEMA_signal_4697 ;
    wire new_AGEMA_signal_4698 ;
    wire new_AGEMA_signal_4699 ;
    wire new_AGEMA_signal_4700 ;
    wire new_AGEMA_signal_4701 ;
    wire new_AGEMA_signal_4702 ;
    wire new_AGEMA_signal_4703 ;
    wire new_AGEMA_signal_4704 ;
    wire new_AGEMA_signal_4705 ;
    wire new_AGEMA_signal_4706 ;
    wire new_AGEMA_signal_4707 ;
    wire new_AGEMA_signal_4708 ;
    wire new_AGEMA_signal_4709 ;
    wire new_AGEMA_signal_4710 ;
    wire new_AGEMA_signal_4711 ;
    wire new_AGEMA_signal_4712 ;
    wire new_AGEMA_signal_4713 ;
    wire new_AGEMA_signal_4714 ;
    wire new_AGEMA_signal_4715 ;
    wire new_AGEMA_signal_4716 ;
    wire new_AGEMA_signal_4717 ;
    wire new_AGEMA_signal_4718 ;
    wire new_AGEMA_signal_4719 ;
    wire new_AGEMA_signal_4720 ;
    wire new_AGEMA_signal_4721 ;
    wire new_AGEMA_signal_4722 ;
    wire new_AGEMA_signal_4723 ;
    wire new_AGEMA_signal_4724 ;
    wire new_AGEMA_signal_4725 ;
    wire new_AGEMA_signal_4726 ;
    wire new_AGEMA_signal_4727 ;
    wire new_AGEMA_signal_4728 ;
    wire new_AGEMA_signal_4729 ;
    wire new_AGEMA_signal_4730 ;
    wire new_AGEMA_signal_4731 ;
    wire new_AGEMA_signal_4732 ;
    wire new_AGEMA_signal_4733 ;
    wire new_AGEMA_signal_4734 ;
    wire new_AGEMA_signal_4735 ;
    wire new_AGEMA_signal_4736 ;
    wire new_AGEMA_signal_4737 ;
    wire new_AGEMA_signal_4738 ;
    wire new_AGEMA_signal_4739 ;
    wire new_AGEMA_signal_4740 ;
    wire new_AGEMA_signal_4741 ;
    wire new_AGEMA_signal_4742 ;
    wire new_AGEMA_signal_4743 ;
    wire new_AGEMA_signal_4744 ;
    wire new_AGEMA_signal_4745 ;
    wire new_AGEMA_signal_4746 ;
    wire new_AGEMA_signal_4747 ;
    wire new_AGEMA_signal_4748 ;
    wire new_AGEMA_signal_4749 ;
    wire new_AGEMA_signal_4750 ;
    wire new_AGEMA_signal_4751 ;
    wire new_AGEMA_signal_4752 ;
    wire new_AGEMA_signal_4753 ;
    wire new_AGEMA_signal_4754 ;
    wire new_AGEMA_signal_4755 ;
    wire new_AGEMA_signal_4756 ;
    wire new_AGEMA_signal_4757 ;
    wire new_AGEMA_signal_4758 ;
    wire new_AGEMA_signal_4759 ;
    wire new_AGEMA_signal_4760 ;
    wire new_AGEMA_signal_4761 ;
    wire new_AGEMA_signal_4762 ;
    wire new_AGEMA_signal_4763 ;
    wire new_AGEMA_signal_4764 ;
    wire new_AGEMA_signal_4765 ;
    wire new_AGEMA_signal_4766 ;
    wire new_AGEMA_signal_4767 ;
    wire new_AGEMA_signal_4768 ;
    wire new_AGEMA_signal_4769 ;
    wire new_AGEMA_signal_4770 ;
    wire new_AGEMA_signal_4771 ;
    wire new_AGEMA_signal_4772 ;
    wire new_AGEMA_signal_4773 ;
    wire new_AGEMA_signal_4774 ;
    wire new_AGEMA_signal_4775 ;
    wire new_AGEMA_signal_4776 ;
    wire new_AGEMA_signal_4777 ;
    wire new_AGEMA_signal_4778 ;
    wire new_AGEMA_signal_4779 ;
    wire new_AGEMA_signal_4780 ;
    wire new_AGEMA_signal_4781 ;
    wire new_AGEMA_signal_4782 ;
    wire new_AGEMA_signal_4783 ;
    wire new_AGEMA_signal_4784 ;
    wire new_AGEMA_signal_4785 ;
    wire new_AGEMA_signal_4786 ;
    wire new_AGEMA_signal_4787 ;
    wire new_AGEMA_signal_4788 ;
    wire new_AGEMA_signal_4789 ;
    wire new_AGEMA_signal_4790 ;
    wire new_AGEMA_signal_4791 ;
    wire new_AGEMA_signal_4792 ;
    wire new_AGEMA_signal_4793 ;
    wire new_AGEMA_signal_4794 ;
    wire new_AGEMA_signal_4795 ;
    wire new_AGEMA_signal_4796 ;
    wire new_AGEMA_signal_4797 ;
    wire new_AGEMA_signal_4798 ;
    wire new_AGEMA_signal_4799 ;
    wire new_AGEMA_signal_4800 ;
    wire new_AGEMA_signal_4801 ;
    wire new_AGEMA_signal_4802 ;
    wire new_AGEMA_signal_4803 ;
    wire new_AGEMA_signal_4804 ;
    wire new_AGEMA_signal_4805 ;
    wire new_AGEMA_signal_4806 ;
    wire new_AGEMA_signal_4807 ;
    wire new_AGEMA_signal_4808 ;
    wire new_AGEMA_signal_4809 ;
    wire new_AGEMA_signal_4810 ;
    wire new_AGEMA_signal_4811 ;
    wire new_AGEMA_signal_4812 ;
    wire new_AGEMA_signal_4813 ;
    wire new_AGEMA_signal_4814 ;
    wire new_AGEMA_signal_4815 ;
    wire new_AGEMA_signal_4816 ;
    wire new_AGEMA_signal_4817 ;
    wire new_AGEMA_signal_4818 ;
    wire new_AGEMA_signal_4819 ;
    wire new_AGEMA_signal_4820 ;
    wire new_AGEMA_signal_4821 ;
    wire new_AGEMA_signal_4822 ;
    wire new_AGEMA_signal_4823 ;
    wire new_AGEMA_signal_4824 ;
    wire new_AGEMA_signal_4825 ;
    wire new_AGEMA_signal_4826 ;
    wire new_AGEMA_signal_4827 ;
    wire new_AGEMA_signal_4828 ;
    wire new_AGEMA_signal_4829 ;
    wire new_AGEMA_signal_4830 ;
    wire new_AGEMA_signal_4831 ;
    wire new_AGEMA_signal_4832 ;
    wire new_AGEMA_signal_4833 ;
    wire new_AGEMA_signal_4834 ;
    wire new_AGEMA_signal_4835 ;
    wire new_AGEMA_signal_4836 ;
    wire new_AGEMA_signal_4837 ;
    wire new_AGEMA_signal_4838 ;
    wire new_AGEMA_signal_4839 ;
    wire new_AGEMA_signal_4840 ;
    wire new_AGEMA_signal_4841 ;
    wire new_AGEMA_signal_4842 ;
    wire new_AGEMA_signal_4843 ;
    wire new_AGEMA_signal_4844 ;
    wire new_AGEMA_signal_4845 ;
    wire new_AGEMA_signal_4846 ;
    wire new_AGEMA_signal_4847 ;
    wire new_AGEMA_signal_4848 ;
    wire new_AGEMA_signal_4849 ;
    wire new_AGEMA_signal_4850 ;
    wire new_AGEMA_signal_4851 ;
    wire new_AGEMA_signal_4852 ;
    wire new_AGEMA_signal_4853 ;
    wire new_AGEMA_signal_4854 ;
    wire new_AGEMA_signal_4855 ;
    wire new_AGEMA_signal_4856 ;
    wire new_AGEMA_signal_4857 ;
    wire new_AGEMA_signal_4858 ;
    wire new_AGEMA_signal_4859 ;
    wire new_AGEMA_signal_4860 ;
    wire new_AGEMA_signal_4861 ;
    wire new_AGEMA_signal_4862 ;
    wire new_AGEMA_signal_4863 ;
    wire new_AGEMA_signal_4864 ;
    wire new_AGEMA_signal_4865 ;
    wire new_AGEMA_signal_4866 ;
    wire new_AGEMA_signal_4867 ;
    wire new_AGEMA_signal_4868 ;
    wire new_AGEMA_signal_4869 ;
    wire new_AGEMA_signal_4870 ;
    wire new_AGEMA_signal_4871 ;
    wire new_AGEMA_signal_4872 ;
    wire new_AGEMA_signal_4873 ;
    wire new_AGEMA_signal_4874 ;
    wire new_AGEMA_signal_4875 ;
    wire new_AGEMA_signal_4876 ;
    wire new_AGEMA_signal_4877 ;
    wire new_AGEMA_signal_4878 ;
    wire new_AGEMA_signal_4879 ;
    wire new_AGEMA_signal_4880 ;
    wire new_AGEMA_signal_4881 ;
    wire new_AGEMA_signal_4882 ;
    wire new_AGEMA_signal_4883 ;
    wire new_AGEMA_signal_4884 ;
    wire new_AGEMA_signal_4885 ;
    wire new_AGEMA_signal_4886 ;
    wire new_AGEMA_signal_4887 ;
    wire new_AGEMA_signal_4888 ;
    wire new_AGEMA_signal_4889 ;
    wire new_AGEMA_signal_4890 ;
    wire new_AGEMA_signal_4891 ;
    wire new_AGEMA_signal_4892 ;
    wire new_AGEMA_signal_4893 ;
    wire new_AGEMA_signal_4894 ;
    wire new_AGEMA_signal_4895 ;
    wire new_AGEMA_signal_4896 ;
    wire new_AGEMA_signal_4897 ;
    wire new_AGEMA_signal_4898 ;
    wire new_AGEMA_signal_4899 ;
    wire new_AGEMA_signal_4900 ;
    wire new_AGEMA_signal_4901 ;
    wire new_AGEMA_signal_4902 ;
    wire new_AGEMA_signal_4903 ;
    wire new_AGEMA_signal_4904 ;
    wire new_AGEMA_signal_4905 ;
    wire new_AGEMA_signal_4906 ;
    wire new_AGEMA_signal_4907 ;
    wire new_AGEMA_signal_4908 ;
    wire new_AGEMA_signal_4909 ;
    wire new_AGEMA_signal_4910 ;
    wire new_AGEMA_signal_4911 ;
    wire new_AGEMA_signal_4912 ;
    wire new_AGEMA_signal_4913 ;
    wire new_AGEMA_signal_4914 ;
    wire new_AGEMA_signal_4915 ;
    wire new_AGEMA_signal_4916 ;
    wire new_AGEMA_signal_4917 ;
    wire new_AGEMA_signal_4918 ;
    wire new_AGEMA_signal_4919 ;
    wire new_AGEMA_signal_4920 ;
    wire new_AGEMA_signal_4921 ;
    wire new_AGEMA_signal_4922 ;
    wire new_AGEMA_signal_4923 ;
    wire new_AGEMA_signal_4924 ;
    wire new_AGEMA_signal_4925 ;
    wire new_AGEMA_signal_4926 ;
    wire new_AGEMA_signal_4927 ;
    wire new_AGEMA_signal_4928 ;
    wire new_AGEMA_signal_4929 ;
    wire new_AGEMA_signal_4930 ;
    wire new_AGEMA_signal_4931 ;
    wire new_AGEMA_signal_4932 ;
    wire new_AGEMA_signal_4933 ;
    wire new_AGEMA_signal_4934 ;
    wire new_AGEMA_signal_4935 ;
    wire new_AGEMA_signal_4936 ;
    wire new_AGEMA_signal_4937 ;
    wire new_AGEMA_signal_4938 ;
    wire new_AGEMA_signal_4939 ;
    wire new_AGEMA_signal_4940 ;
    wire new_AGEMA_signal_4941 ;
    wire new_AGEMA_signal_4942 ;
    wire new_AGEMA_signal_4943 ;
    wire new_AGEMA_signal_4944 ;
    wire new_AGEMA_signal_4945 ;
    wire new_AGEMA_signal_4946 ;
    wire new_AGEMA_signal_4947 ;
    wire new_AGEMA_signal_4948 ;
    wire new_AGEMA_signal_4949 ;
    wire new_AGEMA_signal_4950 ;
    wire new_AGEMA_signal_4951 ;
    wire new_AGEMA_signal_4952 ;
    wire new_AGEMA_signal_4953 ;
    wire new_AGEMA_signal_4954 ;
    wire new_AGEMA_signal_4955 ;
    wire new_AGEMA_signal_4956 ;
    wire new_AGEMA_signal_4957 ;
    wire new_AGEMA_signal_4958 ;
    wire new_AGEMA_signal_4959 ;
    wire new_AGEMA_signal_4960 ;
    wire new_AGEMA_signal_4961 ;
    wire new_AGEMA_signal_4962 ;
    wire new_AGEMA_signal_4963 ;
    wire new_AGEMA_signal_4964 ;
    wire new_AGEMA_signal_4965 ;
    wire new_AGEMA_signal_4966 ;
    wire new_AGEMA_signal_4967 ;
    wire new_AGEMA_signal_4968 ;
    wire new_AGEMA_signal_4969 ;
    wire new_AGEMA_signal_4970 ;
    wire new_AGEMA_signal_4971 ;
    wire new_AGEMA_signal_4972 ;
    wire new_AGEMA_signal_4973 ;
    wire new_AGEMA_signal_4974 ;
    wire new_AGEMA_signal_4975 ;
    wire new_AGEMA_signal_4976 ;
    wire new_AGEMA_signal_4977 ;
    wire new_AGEMA_signal_4978 ;
    wire new_AGEMA_signal_4979 ;
    wire new_AGEMA_signal_4980 ;
    wire new_AGEMA_signal_4981 ;
    wire new_AGEMA_signal_4982 ;
    wire new_AGEMA_signal_4983 ;
    wire new_AGEMA_signal_4984 ;
    wire new_AGEMA_signal_4985 ;
    wire new_AGEMA_signal_4986 ;
    wire new_AGEMA_signal_4987 ;
    wire new_AGEMA_signal_4988 ;
    wire new_AGEMA_signal_4989 ;
    wire new_AGEMA_signal_4990 ;
    wire new_AGEMA_signal_4991 ;
    wire new_AGEMA_signal_4992 ;
    wire new_AGEMA_signal_4993 ;
    wire new_AGEMA_signal_4994 ;
    wire new_AGEMA_signal_4995 ;
    wire new_AGEMA_signal_4996 ;
    wire new_AGEMA_signal_4997 ;
    wire new_AGEMA_signal_4998 ;
    wire new_AGEMA_signal_4999 ;
    wire new_AGEMA_signal_5000 ;
    wire new_AGEMA_signal_5001 ;
    wire new_AGEMA_signal_5002 ;
    wire new_AGEMA_signal_5003 ;
    wire new_AGEMA_signal_5004 ;
    wire new_AGEMA_signal_5005 ;
    wire new_AGEMA_signal_5006 ;
    wire new_AGEMA_signal_5007 ;
    wire new_AGEMA_signal_5008 ;
    wire new_AGEMA_signal_5009 ;
    wire new_AGEMA_signal_5010 ;
    wire new_AGEMA_signal_5011 ;
    wire new_AGEMA_signal_5012 ;
    wire new_AGEMA_signal_5013 ;
    wire new_AGEMA_signal_5014 ;
    wire new_AGEMA_signal_5015 ;
    wire new_AGEMA_signal_5016 ;
    wire new_AGEMA_signal_5017 ;
    wire new_AGEMA_signal_5018 ;
    wire new_AGEMA_signal_5019 ;
    wire new_AGEMA_signal_5020 ;
    wire new_AGEMA_signal_5021 ;
    wire new_AGEMA_signal_5022 ;
    wire new_AGEMA_signal_5023 ;
    wire new_AGEMA_signal_5024 ;
    wire new_AGEMA_signal_5025 ;
    wire new_AGEMA_signal_5026 ;
    wire new_AGEMA_signal_5027 ;
    wire new_AGEMA_signal_5028 ;
    wire new_AGEMA_signal_5029 ;
    wire new_AGEMA_signal_5030 ;
    wire new_AGEMA_signal_5031 ;
    wire new_AGEMA_signal_5032 ;
    wire new_AGEMA_signal_5033 ;
    wire new_AGEMA_signal_5034 ;
    wire new_AGEMA_signal_5035 ;
    wire new_AGEMA_signal_5036 ;
    wire new_AGEMA_signal_5037 ;
    wire new_AGEMA_signal_5038 ;
    wire new_AGEMA_signal_5039 ;
    wire new_AGEMA_signal_5040 ;
    wire new_AGEMA_signal_5041 ;
    wire new_AGEMA_signal_5042 ;
    wire new_AGEMA_signal_5043 ;
    wire new_AGEMA_signal_5044 ;
    wire new_AGEMA_signal_5045 ;
    wire new_AGEMA_signal_5046 ;
    wire new_AGEMA_signal_5047 ;
    wire new_AGEMA_signal_5048 ;
    wire new_AGEMA_signal_5049 ;
    wire new_AGEMA_signal_5050 ;
    wire new_AGEMA_signal_5051 ;
    wire new_AGEMA_signal_5052 ;
    wire new_AGEMA_signal_5053 ;
    wire new_AGEMA_signal_5054 ;
    wire new_AGEMA_signal_5055 ;
    wire new_AGEMA_signal_5056 ;
    wire new_AGEMA_signal_5057 ;
    wire new_AGEMA_signal_5058 ;
    wire new_AGEMA_signal_5059 ;
    wire new_AGEMA_signal_5060 ;
    wire new_AGEMA_signal_5061 ;
    wire new_AGEMA_signal_5062 ;
    wire new_AGEMA_signal_5063 ;
    wire new_AGEMA_signal_5064 ;
    wire new_AGEMA_signal_5065 ;
    wire new_AGEMA_signal_5066 ;
    wire new_AGEMA_signal_5067 ;
    wire new_AGEMA_signal_5068 ;
    wire new_AGEMA_signal_5069 ;
    wire new_AGEMA_signal_5070 ;
    wire new_AGEMA_signal_5071 ;
    wire new_AGEMA_signal_5072 ;
    wire new_AGEMA_signal_5073 ;
    wire new_AGEMA_signal_5074 ;
    wire new_AGEMA_signal_5075 ;
    wire new_AGEMA_signal_5076 ;
    wire new_AGEMA_signal_5077 ;
    wire new_AGEMA_signal_5078 ;
    wire new_AGEMA_signal_5079 ;
    wire new_AGEMA_signal_5080 ;
    wire new_AGEMA_signal_5081 ;
    wire new_AGEMA_signal_5082 ;
    wire new_AGEMA_signal_5083 ;
    wire new_AGEMA_signal_5084 ;
    wire new_AGEMA_signal_5085 ;
    wire new_AGEMA_signal_5086 ;
    wire new_AGEMA_signal_5087 ;
    wire new_AGEMA_signal_5088 ;
    wire new_AGEMA_signal_5089 ;
    wire new_AGEMA_signal_5090 ;
    wire new_AGEMA_signal_5091 ;
    wire new_AGEMA_signal_5092 ;
    wire new_AGEMA_signal_5093 ;
    wire new_AGEMA_signal_5094 ;
    wire new_AGEMA_signal_5095 ;
    wire new_AGEMA_signal_5096 ;
    wire new_AGEMA_signal_5097 ;
    wire new_AGEMA_signal_5098 ;
    wire new_AGEMA_signal_5099 ;
    wire new_AGEMA_signal_5100 ;
    wire new_AGEMA_signal_5101 ;
    wire new_AGEMA_signal_5102 ;
    wire new_AGEMA_signal_5103 ;
    wire new_AGEMA_signal_5104 ;
    wire new_AGEMA_signal_5105 ;
    wire new_AGEMA_signal_5106 ;
    wire new_AGEMA_signal_5107 ;
    wire new_AGEMA_signal_5108 ;
    wire new_AGEMA_signal_5109 ;
    wire new_AGEMA_signal_5110 ;
    wire new_AGEMA_signal_5111 ;
    wire new_AGEMA_signal_5112 ;
    wire new_AGEMA_signal_5113 ;
    wire new_AGEMA_signal_5114 ;
    wire new_AGEMA_signal_5115 ;
    wire new_AGEMA_signal_5116 ;
    wire new_AGEMA_signal_5117 ;
    wire new_AGEMA_signal_5118 ;
    wire new_AGEMA_signal_5119 ;
    wire new_AGEMA_signal_5120 ;
    wire new_AGEMA_signal_5121 ;
    wire new_AGEMA_signal_5122 ;
    wire new_AGEMA_signal_5123 ;
    wire new_AGEMA_signal_5124 ;
    wire new_AGEMA_signal_5125 ;
    wire new_AGEMA_signal_5126 ;
    wire new_AGEMA_signal_5127 ;
    wire new_AGEMA_signal_5128 ;
    wire new_AGEMA_signal_5129 ;
    wire new_AGEMA_signal_5130 ;
    wire new_AGEMA_signal_5131 ;
    wire new_AGEMA_signal_5132 ;
    wire new_AGEMA_signal_5133 ;
    wire new_AGEMA_signal_5134 ;
    wire new_AGEMA_signal_5135 ;
    wire new_AGEMA_signal_5136 ;
    wire new_AGEMA_signal_5137 ;
    wire new_AGEMA_signal_5138 ;
    wire new_AGEMA_signal_5139 ;
    wire new_AGEMA_signal_5140 ;
    wire new_AGEMA_signal_5141 ;
    wire new_AGEMA_signal_5142 ;
    wire new_AGEMA_signal_5143 ;
    wire new_AGEMA_signal_5144 ;
    wire new_AGEMA_signal_5145 ;
    wire new_AGEMA_signal_5146 ;
    wire new_AGEMA_signal_5147 ;
    wire new_AGEMA_signal_5148 ;
    wire new_AGEMA_signal_5149 ;
    wire new_AGEMA_signal_5150 ;
    wire new_AGEMA_signal_5151 ;
    wire new_AGEMA_signal_5152 ;
    wire new_AGEMA_signal_5153 ;
    wire new_AGEMA_signal_5154 ;
    wire new_AGEMA_signal_5155 ;
    wire new_AGEMA_signal_5156 ;
    wire new_AGEMA_signal_5157 ;
    wire new_AGEMA_signal_5158 ;
    wire new_AGEMA_signal_5159 ;
    wire new_AGEMA_signal_5160 ;
    wire new_AGEMA_signal_5161 ;
    wire new_AGEMA_signal_5162 ;
    wire new_AGEMA_signal_5163 ;
    wire new_AGEMA_signal_5164 ;
    wire new_AGEMA_signal_5165 ;
    wire new_AGEMA_signal_5166 ;
    wire new_AGEMA_signal_5167 ;
    wire new_AGEMA_signal_5168 ;
    wire new_AGEMA_signal_5169 ;
    wire new_AGEMA_signal_5170 ;
    wire new_AGEMA_signal_5171 ;
    wire new_AGEMA_signal_5172 ;
    wire new_AGEMA_signal_5173 ;
    wire new_AGEMA_signal_5174 ;
    wire new_AGEMA_signal_5175 ;
    wire new_AGEMA_signal_5176 ;
    wire new_AGEMA_signal_5177 ;
    wire new_AGEMA_signal_5178 ;
    wire new_AGEMA_signal_5179 ;
    wire new_AGEMA_signal_5180 ;
    wire new_AGEMA_signal_5181 ;
    wire new_AGEMA_signal_5182 ;
    wire new_AGEMA_signal_5183 ;
    wire new_AGEMA_signal_5184 ;
    wire new_AGEMA_signal_5185 ;
    wire new_AGEMA_signal_5186 ;
    wire new_AGEMA_signal_5187 ;
    wire new_AGEMA_signal_5188 ;
    wire new_AGEMA_signal_5189 ;
    wire new_AGEMA_signal_5190 ;
    wire new_AGEMA_signal_5191 ;
    wire new_AGEMA_signal_5192 ;
    wire new_AGEMA_signal_5193 ;
    wire new_AGEMA_signal_5194 ;
    wire new_AGEMA_signal_5195 ;
    wire new_AGEMA_signal_5196 ;
    wire new_AGEMA_signal_5197 ;
    wire new_AGEMA_signal_5198 ;
    wire new_AGEMA_signal_5199 ;
    wire new_AGEMA_signal_5200 ;
    wire new_AGEMA_signal_5201 ;
    wire new_AGEMA_signal_5202 ;
    wire new_AGEMA_signal_5203 ;
    wire new_AGEMA_signal_5204 ;
    wire new_AGEMA_signal_5205 ;
    wire new_AGEMA_signal_5206 ;
    wire new_AGEMA_signal_5207 ;
    wire new_AGEMA_signal_5208 ;
    wire new_AGEMA_signal_5209 ;
    wire new_AGEMA_signal_5210 ;
    wire new_AGEMA_signal_5211 ;
    wire new_AGEMA_signal_5212 ;
    wire new_AGEMA_signal_5213 ;
    wire new_AGEMA_signal_5214 ;
    wire new_AGEMA_signal_5215 ;
    wire new_AGEMA_signal_5216 ;
    wire new_AGEMA_signal_5217 ;
    wire new_AGEMA_signal_5218 ;
    wire new_AGEMA_signal_5219 ;
    wire new_AGEMA_signal_5220 ;
    wire new_AGEMA_signal_5221 ;
    wire new_AGEMA_signal_5222 ;
    wire new_AGEMA_signal_5223 ;
    wire new_AGEMA_signal_5224 ;
    wire new_AGEMA_signal_5225 ;
    wire new_AGEMA_signal_5226 ;
    wire new_AGEMA_signal_5227 ;
    wire new_AGEMA_signal_5228 ;
    wire new_AGEMA_signal_5229 ;
    wire new_AGEMA_signal_5230 ;
    wire new_AGEMA_signal_5231 ;
    wire new_AGEMA_signal_5232 ;
    wire new_AGEMA_signal_5233 ;
    wire new_AGEMA_signal_5234 ;
    wire new_AGEMA_signal_5235 ;
    wire new_AGEMA_signal_5236 ;
    wire new_AGEMA_signal_5237 ;
    wire new_AGEMA_signal_5238 ;
    wire new_AGEMA_signal_5239 ;
    wire new_AGEMA_signal_5240 ;
    wire new_AGEMA_signal_5241 ;
    wire new_AGEMA_signal_5242 ;
    wire new_AGEMA_signal_5243 ;
    wire new_AGEMA_signal_5244 ;
    wire new_AGEMA_signal_5245 ;
    wire new_AGEMA_signal_5246 ;
    wire new_AGEMA_signal_5247 ;
    wire new_AGEMA_signal_5248 ;
    wire new_AGEMA_signal_5249 ;
    wire new_AGEMA_signal_5250 ;
    wire new_AGEMA_signal_5251 ;
    wire new_AGEMA_signal_5252 ;
    wire new_AGEMA_signal_5253 ;
    wire new_AGEMA_signal_5254 ;
    wire new_AGEMA_signal_5255 ;
    wire new_AGEMA_signal_5256 ;
    wire new_AGEMA_signal_5257 ;
    wire new_AGEMA_signal_5258 ;
    wire new_AGEMA_signal_5259 ;
    wire new_AGEMA_signal_5260 ;
    wire new_AGEMA_signal_5261 ;
    wire new_AGEMA_signal_5262 ;
    wire new_AGEMA_signal_5263 ;
    wire new_AGEMA_signal_5264 ;
    wire new_AGEMA_signal_5265 ;
    wire new_AGEMA_signal_5266 ;
    wire new_AGEMA_signal_5267 ;
    wire new_AGEMA_signal_5268 ;
    wire new_AGEMA_signal_5269 ;
    wire new_AGEMA_signal_5270 ;
    wire new_AGEMA_signal_5271 ;
    wire new_AGEMA_signal_5272 ;
    wire new_AGEMA_signal_5273 ;
    wire new_AGEMA_signal_5274 ;
    wire new_AGEMA_signal_5275 ;
    wire new_AGEMA_signal_5276 ;
    wire new_AGEMA_signal_5277 ;
    wire new_AGEMA_signal_5278 ;
    wire new_AGEMA_signal_5279 ;
    wire new_AGEMA_signal_5280 ;
    wire new_AGEMA_signal_5281 ;
    wire new_AGEMA_signal_5282 ;
    wire new_AGEMA_signal_5283 ;
    wire new_AGEMA_signal_5284 ;
    wire new_AGEMA_signal_5285 ;
    wire new_AGEMA_signal_5286 ;
    wire new_AGEMA_signal_5287 ;
    wire new_AGEMA_signal_5288 ;
    wire new_AGEMA_signal_5289 ;
    wire new_AGEMA_signal_5290 ;
    wire new_AGEMA_signal_5291 ;
    wire new_AGEMA_signal_5292 ;
    wire new_AGEMA_signal_5293 ;
    wire new_AGEMA_signal_5294 ;
    wire new_AGEMA_signal_5295 ;
    wire new_AGEMA_signal_5296 ;
    wire new_AGEMA_signal_5297 ;
    wire new_AGEMA_signal_5298 ;
    wire new_AGEMA_signal_5299 ;
    wire new_AGEMA_signal_5300 ;
    wire new_AGEMA_signal_5301 ;
    wire new_AGEMA_signal_5302 ;
    wire new_AGEMA_signal_5303 ;
    wire new_AGEMA_signal_5304 ;
    wire new_AGEMA_signal_5305 ;
    wire new_AGEMA_signal_5306 ;
    wire new_AGEMA_signal_5307 ;
    wire new_AGEMA_signal_5308 ;
    wire new_AGEMA_signal_5309 ;
    wire new_AGEMA_signal_5310 ;
    wire new_AGEMA_signal_5311 ;
    wire new_AGEMA_signal_5312 ;
    wire new_AGEMA_signal_5313 ;
    wire new_AGEMA_signal_5314 ;
    wire new_AGEMA_signal_5315 ;
    wire new_AGEMA_signal_5316 ;
    wire new_AGEMA_signal_5317 ;
    wire new_AGEMA_signal_5318 ;
    wire new_AGEMA_signal_5319 ;
    wire new_AGEMA_signal_5320 ;
    wire new_AGEMA_signal_5321 ;
    wire new_AGEMA_signal_5322 ;
    wire new_AGEMA_signal_5323 ;
    wire new_AGEMA_signal_5324 ;
    wire new_AGEMA_signal_5325 ;
    wire new_AGEMA_signal_5326 ;
    wire new_AGEMA_signal_5327 ;
    wire new_AGEMA_signal_5328 ;
    wire new_AGEMA_signal_5329 ;
    wire new_AGEMA_signal_5330 ;
    wire new_AGEMA_signal_5331 ;
    wire new_AGEMA_signal_5332 ;
    wire new_AGEMA_signal_5333 ;
    wire new_AGEMA_signal_5334 ;
    wire new_AGEMA_signal_5335 ;
    wire new_AGEMA_signal_5336 ;
    wire new_AGEMA_signal_5337 ;
    wire new_AGEMA_signal_5338 ;
    wire new_AGEMA_signal_5339 ;
    wire new_AGEMA_signal_5340 ;
    wire new_AGEMA_signal_5341 ;
    wire new_AGEMA_signal_5342 ;
    wire new_AGEMA_signal_5343 ;
    wire new_AGEMA_signal_5344 ;
    wire new_AGEMA_signal_5345 ;
    wire new_AGEMA_signal_5346 ;
    wire new_AGEMA_signal_5347 ;
    wire new_AGEMA_signal_5348 ;
    wire new_AGEMA_signal_5349 ;
    wire new_AGEMA_signal_5350 ;
    wire new_AGEMA_signal_5351 ;
    wire new_AGEMA_signal_5352 ;
    wire new_AGEMA_signal_5353 ;
    wire new_AGEMA_signal_5354 ;
    wire new_AGEMA_signal_5355 ;
    wire new_AGEMA_signal_5356 ;
    wire new_AGEMA_signal_5357 ;
    wire new_AGEMA_signal_5358 ;
    wire new_AGEMA_signal_5359 ;
    wire new_AGEMA_signal_5360 ;
    wire new_AGEMA_signal_5361 ;
    wire new_AGEMA_signal_5362 ;
    wire new_AGEMA_signal_5363 ;
    wire new_AGEMA_signal_5364 ;
    wire new_AGEMA_signal_5365 ;
    wire new_AGEMA_signal_5366 ;
    wire new_AGEMA_signal_5367 ;
    wire new_AGEMA_signal_5368 ;
    wire new_AGEMA_signal_5369 ;
    wire new_AGEMA_signal_5370 ;
    wire new_AGEMA_signal_5371 ;
    wire new_AGEMA_signal_5372 ;
    wire new_AGEMA_signal_5373 ;
    wire new_AGEMA_signal_5374 ;
    wire new_AGEMA_signal_5375 ;
    wire new_AGEMA_signal_5376 ;
    wire new_AGEMA_signal_5377 ;
    wire new_AGEMA_signal_5378 ;
    wire new_AGEMA_signal_5379 ;
    wire new_AGEMA_signal_5380 ;
    wire new_AGEMA_signal_5381 ;
    wire new_AGEMA_signal_5382 ;
    wire new_AGEMA_signal_5383 ;
    wire new_AGEMA_signal_5384 ;
    wire new_AGEMA_signal_5385 ;
    wire new_AGEMA_signal_5386 ;
    wire new_AGEMA_signal_5387 ;
    wire new_AGEMA_signal_5388 ;
    wire new_AGEMA_signal_5389 ;
    wire new_AGEMA_signal_5390 ;
    wire new_AGEMA_signal_5391 ;
    wire new_AGEMA_signal_5392 ;
    wire new_AGEMA_signal_5393 ;
    wire new_AGEMA_signal_5394 ;
    wire new_AGEMA_signal_5395 ;
    wire new_AGEMA_signal_5396 ;
    wire new_AGEMA_signal_5397 ;
    wire new_AGEMA_signal_5398 ;
    wire new_AGEMA_signal_5399 ;
    wire new_AGEMA_signal_5400 ;
    wire new_AGEMA_signal_5401 ;
    wire new_AGEMA_signal_5402 ;
    wire new_AGEMA_signal_5403 ;
    wire new_AGEMA_signal_5404 ;
    wire new_AGEMA_signal_5405 ;
    wire new_AGEMA_signal_5406 ;
    wire new_AGEMA_signal_5407 ;
    wire new_AGEMA_signal_5408 ;
    wire new_AGEMA_signal_5409 ;
    wire new_AGEMA_signal_5410 ;
    wire new_AGEMA_signal_5411 ;
    wire new_AGEMA_signal_5412 ;
    wire new_AGEMA_signal_5413 ;
    wire new_AGEMA_signal_5414 ;
    wire new_AGEMA_signal_5415 ;
    wire new_AGEMA_signal_5416 ;
    wire new_AGEMA_signal_5417 ;
    wire new_AGEMA_signal_5418 ;
    wire new_AGEMA_signal_5419 ;
    wire new_AGEMA_signal_5420 ;
    wire new_AGEMA_signal_5421 ;
    wire new_AGEMA_signal_5422 ;
    wire new_AGEMA_signal_5423 ;
    wire new_AGEMA_signal_5424 ;
    wire new_AGEMA_signal_5425 ;
    wire new_AGEMA_signal_5426 ;
    wire new_AGEMA_signal_5427 ;
    wire new_AGEMA_signal_5428 ;
    wire new_AGEMA_signal_5429 ;
    wire new_AGEMA_signal_5430 ;
    wire new_AGEMA_signal_5431 ;
    wire new_AGEMA_signal_5432 ;
    wire new_AGEMA_signal_5433 ;
    wire new_AGEMA_signal_5434 ;
    wire new_AGEMA_signal_5435 ;
    wire new_AGEMA_signal_5436 ;
    wire new_AGEMA_signal_5437 ;
    wire new_AGEMA_signal_5438 ;
    wire new_AGEMA_signal_5439 ;
    wire new_AGEMA_signal_5440 ;
    wire new_AGEMA_signal_5441 ;
    wire new_AGEMA_signal_5442 ;
    wire new_AGEMA_signal_5443 ;
    wire new_AGEMA_signal_5444 ;
    wire new_AGEMA_signal_5445 ;
    wire new_AGEMA_signal_5446 ;
    wire new_AGEMA_signal_5447 ;
    wire new_AGEMA_signal_5448 ;
    wire new_AGEMA_signal_5449 ;
    wire new_AGEMA_signal_5450 ;
    wire new_AGEMA_signal_5451 ;
    wire new_AGEMA_signal_5452 ;
    wire new_AGEMA_signal_5453 ;
    wire new_AGEMA_signal_5454 ;
    wire new_AGEMA_signal_5455 ;
    wire new_AGEMA_signal_5456 ;
    wire new_AGEMA_signal_5457 ;
    wire new_AGEMA_signal_5458 ;
    wire new_AGEMA_signal_5459 ;
    wire new_AGEMA_signal_5460 ;
    wire new_AGEMA_signal_5461 ;
    wire new_AGEMA_signal_5462 ;
    wire new_AGEMA_signal_5463 ;
    wire new_AGEMA_signal_5464 ;
    wire new_AGEMA_signal_5465 ;
    wire new_AGEMA_signal_5466 ;
    wire new_AGEMA_signal_5467 ;
    wire new_AGEMA_signal_5468 ;
    wire new_AGEMA_signal_5469 ;
    wire new_AGEMA_signal_5470 ;
    wire new_AGEMA_signal_5471 ;
    wire new_AGEMA_signal_5472 ;
    wire new_AGEMA_signal_5473 ;
    wire new_AGEMA_signal_5474 ;
    wire new_AGEMA_signal_5475 ;
    wire new_AGEMA_signal_5476 ;
    wire new_AGEMA_signal_5477 ;
    wire new_AGEMA_signal_5478 ;
    wire new_AGEMA_signal_5479 ;
    wire new_AGEMA_signal_5480 ;
    wire new_AGEMA_signal_5481 ;
    wire new_AGEMA_signal_5482 ;
    wire new_AGEMA_signal_5483 ;
    wire new_AGEMA_signal_5484 ;
    wire new_AGEMA_signal_5485 ;
    wire new_AGEMA_signal_5486 ;
    wire new_AGEMA_signal_5487 ;
    wire new_AGEMA_signal_5488 ;
    wire new_AGEMA_signal_5489 ;
    wire new_AGEMA_signal_5490 ;
    wire new_AGEMA_signal_5491 ;
    wire new_AGEMA_signal_5492 ;
    wire new_AGEMA_signal_5493 ;
    wire new_AGEMA_signal_5494 ;
    wire new_AGEMA_signal_5495 ;
    wire new_AGEMA_signal_5496 ;
    wire new_AGEMA_signal_5497 ;
    wire new_AGEMA_signal_5498 ;
    wire new_AGEMA_signal_5499 ;
    wire new_AGEMA_signal_5500 ;
    wire new_AGEMA_signal_5501 ;
    wire new_AGEMA_signal_5502 ;
    wire new_AGEMA_signal_5503 ;
    wire new_AGEMA_signal_5504 ;
    wire new_AGEMA_signal_5505 ;
    wire new_AGEMA_signal_5506 ;
    wire new_AGEMA_signal_5507 ;
    wire new_AGEMA_signal_5508 ;
    wire new_AGEMA_signal_5509 ;
    wire new_AGEMA_signal_5510 ;
    wire new_AGEMA_signal_5511 ;
    wire new_AGEMA_signal_5512 ;
    wire new_AGEMA_signal_5513 ;
    wire new_AGEMA_signal_5514 ;
    wire new_AGEMA_signal_5515 ;
    wire new_AGEMA_signal_5516 ;
    wire new_AGEMA_signal_5517 ;
    wire new_AGEMA_signal_5518 ;
    wire new_AGEMA_signal_5519 ;
    wire new_AGEMA_signal_5520 ;
    wire new_AGEMA_signal_5521 ;
    wire new_AGEMA_signal_5522 ;
    wire new_AGEMA_signal_5523 ;
    wire new_AGEMA_signal_5524 ;
    wire new_AGEMA_signal_5525 ;
    wire new_AGEMA_signal_5526 ;
    wire new_AGEMA_signal_5527 ;
    wire new_AGEMA_signal_5528 ;
    wire new_AGEMA_signal_5529 ;
    wire new_AGEMA_signal_5530 ;
    wire new_AGEMA_signal_5531 ;
    wire new_AGEMA_signal_5532 ;
    wire new_AGEMA_signal_5533 ;
    wire new_AGEMA_signal_5534 ;
    wire new_AGEMA_signal_5535 ;
    wire new_AGEMA_signal_5536 ;
    wire new_AGEMA_signal_5537 ;
    wire new_AGEMA_signal_5538 ;
    wire new_AGEMA_signal_5539 ;
    wire new_AGEMA_signal_5540 ;
    wire new_AGEMA_signal_5541 ;
    wire new_AGEMA_signal_5542 ;
    wire new_AGEMA_signal_5543 ;
    wire new_AGEMA_signal_5544 ;
    wire new_AGEMA_signal_5545 ;
    wire new_AGEMA_signal_5546 ;
    wire new_AGEMA_signal_5547 ;
    wire new_AGEMA_signal_5548 ;
    wire new_AGEMA_signal_5549 ;
    wire new_AGEMA_signal_5550 ;
    wire new_AGEMA_signal_5551 ;
    wire new_AGEMA_signal_5552 ;
    wire new_AGEMA_signal_5553 ;
    wire new_AGEMA_signal_5554 ;
    wire new_AGEMA_signal_5555 ;
    wire new_AGEMA_signal_5556 ;
    wire new_AGEMA_signal_5557 ;
    wire new_AGEMA_signal_5558 ;
    wire new_AGEMA_signal_5559 ;
    wire new_AGEMA_signal_5560 ;
    wire new_AGEMA_signal_5561 ;
    wire new_AGEMA_signal_5562 ;
    wire new_AGEMA_signal_5563 ;
    wire new_AGEMA_signal_5564 ;
    wire new_AGEMA_signal_5565 ;
    wire new_AGEMA_signal_5566 ;
    wire new_AGEMA_signal_5567 ;
    wire new_AGEMA_signal_5568 ;
    wire new_AGEMA_signal_5569 ;
    wire new_AGEMA_signal_5570 ;
    wire new_AGEMA_signal_5571 ;
    wire new_AGEMA_signal_5572 ;
    wire new_AGEMA_signal_5573 ;
    wire new_AGEMA_signal_5574 ;
    wire new_AGEMA_signal_5575 ;
    wire new_AGEMA_signal_5576 ;
    wire new_AGEMA_signal_5577 ;
    wire new_AGEMA_signal_5578 ;
    wire new_AGEMA_signal_5579 ;
    wire new_AGEMA_signal_5580 ;
    wire new_AGEMA_signal_5581 ;
    wire new_AGEMA_signal_5582 ;
    wire new_AGEMA_signal_5583 ;
    wire new_AGEMA_signal_5584 ;
    wire new_AGEMA_signal_5585 ;
    wire new_AGEMA_signal_5586 ;
    wire new_AGEMA_signal_5587 ;
    wire new_AGEMA_signal_5588 ;
    wire new_AGEMA_signal_5589 ;
    wire new_AGEMA_signal_5590 ;
    wire new_AGEMA_signal_5591 ;
    wire new_AGEMA_signal_5592 ;
    wire new_AGEMA_signal_5593 ;
    wire new_AGEMA_signal_5594 ;
    wire new_AGEMA_signal_5595 ;
    wire new_AGEMA_signal_5596 ;
    wire new_AGEMA_signal_5597 ;
    wire new_AGEMA_signal_5598 ;
    wire new_AGEMA_signal_5599 ;
    wire new_AGEMA_signal_5600 ;
    wire new_AGEMA_signal_5601 ;
    wire new_AGEMA_signal_5602 ;
    wire new_AGEMA_signal_5603 ;
    wire new_AGEMA_signal_5604 ;
    wire new_AGEMA_signal_5605 ;
    wire new_AGEMA_signal_5606 ;
    wire new_AGEMA_signal_5607 ;
    wire new_AGEMA_signal_5608 ;
    wire new_AGEMA_signal_5609 ;
    wire new_AGEMA_signal_5610 ;
    wire new_AGEMA_signal_5611 ;
    wire new_AGEMA_signal_5612 ;
    wire new_AGEMA_signal_5613 ;
    wire new_AGEMA_signal_5614 ;
    wire new_AGEMA_signal_5615 ;
    wire new_AGEMA_signal_5616 ;
    wire new_AGEMA_signal_5617 ;
    wire new_AGEMA_signal_5618 ;
    wire new_AGEMA_signal_5619 ;
    wire new_AGEMA_signal_5620 ;
    wire new_AGEMA_signal_5621 ;
    wire new_AGEMA_signal_5622 ;
    wire new_AGEMA_signal_5623 ;
    wire new_AGEMA_signal_5624 ;
    wire new_AGEMA_signal_5625 ;
    wire new_AGEMA_signal_5626 ;
    wire new_AGEMA_signal_5627 ;
    wire new_AGEMA_signal_5628 ;
    wire new_AGEMA_signal_5629 ;
    wire new_AGEMA_signal_5630 ;
    wire new_AGEMA_signal_5631 ;
    wire new_AGEMA_signal_5633 ;
    wire new_AGEMA_signal_5634 ;
    wire new_AGEMA_signal_5635 ;
    wire new_AGEMA_signal_5636 ;
    wire new_AGEMA_signal_5637 ;
    wire new_AGEMA_signal_5638 ;
    wire new_AGEMA_signal_5639 ;
    wire new_AGEMA_signal_5640 ;
    wire new_AGEMA_signal_5641 ;
    wire new_AGEMA_signal_5642 ;
    wire new_AGEMA_signal_5643 ;
    wire new_AGEMA_signal_5644 ;
    wire new_AGEMA_signal_5645 ;
    wire new_AGEMA_signal_5646 ;
    wire new_AGEMA_signal_5647 ;
    wire new_AGEMA_signal_5648 ;
    wire new_AGEMA_signal_5649 ;
    wire new_AGEMA_signal_5650 ;
    wire new_AGEMA_signal_5651 ;
    wire new_AGEMA_signal_5652 ;
    wire new_AGEMA_signal_5653 ;
    wire new_AGEMA_signal_5654 ;
    wire new_AGEMA_signal_5655 ;
    wire new_AGEMA_signal_5656 ;
    wire new_AGEMA_signal_5657 ;
    wire new_AGEMA_signal_5658 ;
    wire new_AGEMA_signal_5659 ;
    wire new_AGEMA_signal_5660 ;
    wire new_AGEMA_signal_5661 ;
    wire new_AGEMA_signal_5662 ;
    wire new_AGEMA_signal_5663 ;
    wire new_AGEMA_signal_5664 ;
    wire new_AGEMA_signal_5665 ;
    wire new_AGEMA_signal_5666 ;
    wire new_AGEMA_signal_5667 ;
    wire new_AGEMA_signal_5668 ;
    wire new_AGEMA_signal_5669 ;
    wire new_AGEMA_signal_5670 ;
    wire new_AGEMA_signal_5671 ;
    wire new_AGEMA_signal_5672 ;
    wire new_AGEMA_signal_5673 ;
    wire new_AGEMA_signal_5674 ;
    wire new_AGEMA_signal_5675 ;
    wire new_AGEMA_signal_5676 ;
    wire new_AGEMA_signal_5677 ;
    wire new_AGEMA_signal_5678 ;
    wire new_AGEMA_signal_5679 ;
    wire new_AGEMA_signal_5680 ;
    wire new_AGEMA_signal_5681 ;
    wire new_AGEMA_signal_5682 ;
    wire new_AGEMA_signal_5683 ;
    wire new_AGEMA_signal_5684 ;
    wire new_AGEMA_signal_5685 ;
    wire new_AGEMA_signal_5686 ;
    wire new_AGEMA_signal_5687 ;
    wire new_AGEMA_signal_5688 ;
    wire new_AGEMA_signal_5689 ;
    wire new_AGEMA_signal_5690 ;
    wire new_AGEMA_signal_5691 ;
    wire new_AGEMA_signal_5692 ;
    wire new_AGEMA_signal_5693 ;
    wire new_AGEMA_signal_5694 ;
    wire new_AGEMA_signal_5695 ;
    wire new_AGEMA_signal_5696 ;
    wire new_AGEMA_signal_5697 ;
    wire new_AGEMA_signal_5698 ;
    wire new_AGEMA_signal_5699 ;
    wire new_AGEMA_signal_5700 ;
    wire new_AGEMA_signal_5701 ;
    wire new_AGEMA_signal_5702 ;
    wire new_AGEMA_signal_5703 ;
    wire new_AGEMA_signal_5704 ;
    wire new_AGEMA_signal_5705 ;
    wire new_AGEMA_signal_5706 ;
    wire new_AGEMA_signal_5707 ;
    wire new_AGEMA_signal_5708 ;
    wire new_AGEMA_signal_5709 ;
    wire new_AGEMA_signal_5710 ;
    wire new_AGEMA_signal_5711 ;
    wire new_AGEMA_signal_5712 ;
    wire new_AGEMA_signal_5713 ;
    wire new_AGEMA_signal_5714 ;
    wire new_AGEMA_signal_5715 ;
    wire new_AGEMA_signal_5716 ;
    wire new_AGEMA_signal_5717 ;
    wire new_AGEMA_signal_5718 ;
    wire new_AGEMA_signal_5719 ;
    wire new_AGEMA_signal_5720 ;
    wire new_AGEMA_signal_5721 ;
    wire new_AGEMA_signal_5722 ;
    wire new_AGEMA_signal_5723 ;
    wire new_AGEMA_signal_5724 ;
    wire new_AGEMA_signal_5725 ;
    wire new_AGEMA_signal_5726 ;
    wire new_AGEMA_signal_5727 ;
    wire new_AGEMA_signal_5728 ;
    wire new_AGEMA_signal_5729 ;
    wire new_AGEMA_signal_5730 ;
    wire new_AGEMA_signal_5731 ;
    wire new_AGEMA_signal_5732 ;
    wire new_AGEMA_signal_5733 ;
    wire new_AGEMA_signal_5734 ;
    wire new_AGEMA_signal_5735 ;
    wire new_AGEMA_signal_5736 ;
    wire new_AGEMA_signal_5737 ;
    wire new_AGEMA_signal_5738 ;
    wire new_AGEMA_signal_5739 ;
    wire new_AGEMA_signal_5740 ;
    wire new_AGEMA_signal_5741 ;
    wire new_AGEMA_signal_5742 ;
    wire new_AGEMA_signal_5743 ;
    wire new_AGEMA_signal_5744 ;
    wire new_AGEMA_signal_5745 ;
    wire new_AGEMA_signal_5746 ;
    wire new_AGEMA_signal_5747 ;
    wire new_AGEMA_signal_5748 ;
    wire new_AGEMA_signal_5749 ;
    wire new_AGEMA_signal_5750 ;
    wire new_AGEMA_signal_5751 ;
    wire new_AGEMA_signal_5752 ;
    wire new_AGEMA_signal_5753 ;
    wire new_AGEMA_signal_5754 ;
    wire new_AGEMA_signal_5755 ;
    wire new_AGEMA_signal_5756 ;
    wire new_AGEMA_signal_5757 ;
    wire new_AGEMA_signal_5758 ;
    wire new_AGEMA_signal_5759 ;
    wire new_AGEMA_signal_5760 ;
    wire new_AGEMA_signal_5761 ;
    wire new_AGEMA_signal_5762 ;
    wire new_AGEMA_signal_5763 ;
    wire new_AGEMA_signal_5764 ;
    wire new_AGEMA_signal_5765 ;
    wire new_AGEMA_signal_5766 ;
    wire new_AGEMA_signal_5767 ;
    wire new_AGEMA_signal_5768 ;
    wire new_AGEMA_signal_5769 ;
    wire new_AGEMA_signal_5770 ;
    wire new_AGEMA_signal_5771 ;
    wire new_AGEMA_signal_5772 ;
    wire new_AGEMA_signal_5773 ;
    wire new_AGEMA_signal_5774 ;
    wire new_AGEMA_signal_5775 ;
    wire new_AGEMA_signal_5776 ;
    wire new_AGEMA_signal_5777 ;
    wire new_AGEMA_signal_5778 ;
    wire new_AGEMA_signal_5779 ;
    wire new_AGEMA_signal_5780 ;
    wire new_AGEMA_signal_5781 ;
    wire new_AGEMA_signal_5782 ;
    wire new_AGEMA_signal_5783 ;
    wire new_AGEMA_signal_5784 ;
    wire new_AGEMA_signal_5785 ;
    wire new_AGEMA_signal_5786 ;
    wire new_AGEMA_signal_5787 ;
    wire new_AGEMA_signal_5788 ;
    wire new_AGEMA_signal_5789 ;
    wire new_AGEMA_signal_5790 ;
    wire new_AGEMA_signal_5791 ;
    wire new_AGEMA_signal_5792 ;
    wire new_AGEMA_signal_5793 ;
    wire new_AGEMA_signal_5794 ;
    wire new_AGEMA_signal_5795 ;
    wire new_AGEMA_signal_5796 ;
    wire new_AGEMA_signal_5797 ;
    wire new_AGEMA_signal_5798 ;
    wire new_AGEMA_signal_5799 ;
    wire new_AGEMA_signal_5800 ;
    wire new_AGEMA_signal_5801 ;
    wire new_AGEMA_signal_5802 ;
    wire new_AGEMA_signal_5803 ;
    wire new_AGEMA_signal_5804 ;
    wire new_AGEMA_signal_5805 ;
    wire new_AGEMA_signal_5806 ;
    wire new_AGEMA_signal_5807 ;
    wire new_AGEMA_signal_5808 ;
    wire new_AGEMA_signal_5809 ;
    wire new_AGEMA_signal_5810 ;
    wire new_AGEMA_signal_5811 ;
    wire new_AGEMA_signal_5812 ;
    wire new_AGEMA_signal_5813 ;
    wire new_AGEMA_signal_5814 ;
    wire new_AGEMA_signal_5815 ;
    wire new_AGEMA_signal_5816 ;
    wire new_AGEMA_signal_5817 ;
    wire new_AGEMA_signal_5818 ;
    wire new_AGEMA_signal_5819 ;
    wire new_AGEMA_signal_5820 ;
    wire new_AGEMA_signal_5821 ;
    wire new_AGEMA_signal_5822 ;
    wire new_AGEMA_signal_5823 ;
    wire new_AGEMA_signal_5824 ;
    wire new_AGEMA_signal_5825 ;
    wire new_AGEMA_signal_5826 ;
    wire new_AGEMA_signal_5827 ;
    wire new_AGEMA_signal_5828 ;
    wire new_AGEMA_signal_5829 ;
    wire new_AGEMA_signal_5830 ;
    wire new_AGEMA_signal_5831 ;
    wire new_AGEMA_signal_5832 ;
    wire new_AGEMA_signal_5833 ;
    wire new_AGEMA_signal_5834 ;
    wire new_AGEMA_signal_5835 ;
    wire new_AGEMA_signal_5836 ;
    wire new_AGEMA_signal_5837 ;
    wire new_AGEMA_signal_5838 ;
    wire new_AGEMA_signal_5839 ;
    wire new_AGEMA_signal_5840 ;
    wire new_AGEMA_signal_5841 ;
    wire new_AGEMA_signal_5842 ;
    wire new_AGEMA_signal_5843 ;
    wire new_AGEMA_signal_5844 ;
    wire new_AGEMA_signal_5845 ;
    wire new_AGEMA_signal_5846 ;
    wire new_AGEMA_signal_5847 ;
    wire new_AGEMA_signal_5848 ;
    wire new_AGEMA_signal_5849 ;
    wire new_AGEMA_signal_5850 ;
    wire new_AGEMA_signal_5851 ;
    wire new_AGEMA_signal_5852 ;
    wire new_AGEMA_signal_5853 ;
    wire new_AGEMA_signal_5854 ;
    wire new_AGEMA_signal_5855 ;
    wire new_AGEMA_signal_5856 ;
    wire new_AGEMA_signal_5857 ;
    wire new_AGEMA_signal_5858 ;
    wire new_AGEMA_signal_5859 ;
    wire new_AGEMA_signal_5860 ;
    wire new_AGEMA_signal_5861 ;
    wire new_AGEMA_signal_5862 ;
    wire new_AGEMA_signal_5863 ;
    wire new_AGEMA_signal_5864 ;
    wire new_AGEMA_signal_5865 ;
    wire new_AGEMA_signal_5866 ;
    wire new_AGEMA_signal_5867 ;
    wire new_AGEMA_signal_5868 ;
    wire new_AGEMA_signal_5869 ;
    wire new_AGEMA_signal_5870 ;
    wire new_AGEMA_signal_5871 ;
    wire new_AGEMA_signal_5872 ;
    wire new_AGEMA_signal_5873 ;
    wire new_AGEMA_signal_5874 ;
    wire new_AGEMA_signal_5875 ;
    wire new_AGEMA_signal_5876 ;
    wire new_AGEMA_signal_5877 ;
    wire new_AGEMA_signal_5878 ;
    wire new_AGEMA_signal_5879 ;
    wire new_AGEMA_signal_5880 ;
    wire new_AGEMA_signal_5881 ;
    wire new_AGEMA_signal_5882 ;
    wire new_AGEMA_signal_5883 ;
    wire new_AGEMA_signal_5884 ;
    wire new_AGEMA_signal_5885 ;
    wire new_AGEMA_signal_5886 ;
    wire new_AGEMA_signal_5887 ;
    wire new_AGEMA_signal_5888 ;
    wire new_AGEMA_signal_5889 ;
    wire new_AGEMA_signal_5890 ;
    wire new_AGEMA_signal_5891 ;
    wire new_AGEMA_signal_5892 ;
    wire new_AGEMA_signal_5893 ;
    wire new_AGEMA_signal_5894 ;
    wire new_AGEMA_signal_5895 ;
    wire new_AGEMA_signal_5896 ;
    wire new_AGEMA_signal_5897 ;
    wire new_AGEMA_signal_5898 ;
    wire new_AGEMA_signal_5899 ;
    wire new_AGEMA_signal_5900 ;
    wire new_AGEMA_signal_5901 ;
    wire new_AGEMA_signal_5902 ;
    wire new_AGEMA_signal_5903 ;
    wire new_AGEMA_signal_5904 ;
    wire new_AGEMA_signal_5905 ;
    wire new_AGEMA_signal_5906 ;
    wire new_AGEMA_signal_5907 ;
    wire new_AGEMA_signal_5908 ;
    wire new_AGEMA_signal_5909 ;
    wire new_AGEMA_signal_5910 ;
    wire new_AGEMA_signal_5911 ;
    wire new_AGEMA_signal_5912 ;
    wire new_AGEMA_signal_5913 ;
    wire new_AGEMA_signal_5914 ;
    wire new_AGEMA_signal_5915 ;
    wire new_AGEMA_signal_5916 ;
    wire new_AGEMA_signal_5917 ;
    wire new_AGEMA_signal_5918 ;
    wire new_AGEMA_signal_5919 ;
    wire new_AGEMA_signal_5920 ;
    wire new_AGEMA_signal_5921 ;
    wire new_AGEMA_signal_5922 ;
    wire new_AGEMA_signal_5923 ;
    wire new_AGEMA_signal_5924 ;
    wire new_AGEMA_signal_5925 ;
    wire new_AGEMA_signal_5926 ;
    wire new_AGEMA_signal_5927 ;
    wire new_AGEMA_signal_5928 ;
    wire new_AGEMA_signal_5929 ;
    wire new_AGEMA_signal_5930 ;
    wire new_AGEMA_signal_5931 ;
    wire new_AGEMA_signal_5932 ;
    wire new_AGEMA_signal_5933 ;
    wire new_AGEMA_signal_5934 ;
    wire new_AGEMA_signal_5935 ;
    wire new_AGEMA_signal_5936 ;
    wire new_AGEMA_signal_5937 ;
    wire new_AGEMA_signal_5938 ;
    wire new_AGEMA_signal_5939 ;
    wire new_AGEMA_signal_5940 ;
    wire new_AGEMA_signal_5941 ;
    wire new_AGEMA_signal_5942 ;
    wire new_AGEMA_signal_5943 ;
    wire new_AGEMA_signal_5944 ;
    wire new_AGEMA_signal_5945 ;
    wire new_AGEMA_signal_5946 ;
    wire new_AGEMA_signal_5947 ;
    wire new_AGEMA_signal_5948 ;
    wire new_AGEMA_signal_5949 ;
    wire new_AGEMA_signal_5950 ;
    wire new_AGEMA_signal_5951 ;
    wire new_AGEMA_signal_5952 ;
    wire new_AGEMA_signal_5953 ;
    wire new_AGEMA_signal_5954 ;
    wire new_AGEMA_signal_5955 ;
    wire new_AGEMA_signal_5956 ;
    wire new_AGEMA_signal_5957 ;
    wire new_AGEMA_signal_5958 ;
    wire new_AGEMA_signal_5959 ;
    wire new_AGEMA_signal_5960 ;
    wire new_AGEMA_signal_5961 ;
    wire new_AGEMA_signal_5962 ;
    wire new_AGEMA_signal_5963 ;
    wire new_AGEMA_signal_5964 ;
    wire new_AGEMA_signal_5965 ;
    wire new_AGEMA_signal_5966 ;
    wire new_AGEMA_signal_5967 ;
    wire new_AGEMA_signal_5968 ;
    wire new_AGEMA_signal_5969 ;
    wire new_AGEMA_signal_5970 ;
    wire new_AGEMA_signal_5971 ;
    wire new_AGEMA_signal_5972 ;
    wire new_AGEMA_signal_5973 ;
    wire new_AGEMA_signal_5974 ;
    wire new_AGEMA_signal_5975 ;
    wire new_AGEMA_signal_5976 ;
    wire new_AGEMA_signal_5977 ;
    wire new_AGEMA_signal_5978 ;
    wire new_AGEMA_signal_5979 ;
    wire new_AGEMA_signal_5980 ;
    wire new_AGEMA_signal_5981 ;
    wire new_AGEMA_signal_5982 ;
    wire new_AGEMA_signal_5983 ;
    wire new_AGEMA_signal_5984 ;
    wire new_AGEMA_signal_5985 ;
    wire new_AGEMA_signal_5986 ;
    wire new_AGEMA_signal_5987 ;
    wire new_AGEMA_signal_5988 ;
    wire new_AGEMA_signal_5989 ;
    wire new_AGEMA_signal_5990 ;
    wire new_AGEMA_signal_5991 ;
    wire new_AGEMA_signal_5992 ;
    wire new_AGEMA_signal_5993 ;
    wire new_AGEMA_signal_5994 ;
    wire new_AGEMA_signal_5995 ;
    wire new_AGEMA_signal_5996 ;
    wire new_AGEMA_signal_5997 ;
    wire new_AGEMA_signal_5998 ;
    wire new_AGEMA_signal_5999 ;
    wire new_AGEMA_signal_6000 ;
    wire new_AGEMA_signal_6001 ;
    wire new_AGEMA_signal_6002 ;
    wire new_AGEMA_signal_6003 ;
    wire new_AGEMA_signal_6004 ;
    wire new_AGEMA_signal_6005 ;
    wire new_AGEMA_signal_6006 ;
    wire new_AGEMA_signal_6007 ;
    wire new_AGEMA_signal_6008 ;
    wire new_AGEMA_signal_6009 ;
    wire new_AGEMA_signal_6010 ;
    wire new_AGEMA_signal_6011 ;
    wire new_AGEMA_signal_6012 ;
    wire new_AGEMA_signal_6013 ;
    wire new_AGEMA_signal_6014 ;
    wire new_AGEMA_signal_6015 ;
    wire new_AGEMA_signal_6016 ;
    wire new_AGEMA_signal_6017 ;
    wire new_AGEMA_signal_6018 ;
    wire new_AGEMA_signal_6019 ;
    wire new_AGEMA_signal_6020 ;
    wire new_AGEMA_signal_6021 ;
    wire new_AGEMA_signal_6022 ;
    wire new_AGEMA_signal_6023 ;
    wire new_AGEMA_signal_6024 ;
    wire new_AGEMA_signal_6025 ;
    wire new_AGEMA_signal_6026 ;
    wire new_AGEMA_signal_6027 ;
    wire new_AGEMA_signal_6028 ;
    wire new_AGEMA_signal_6029 ;
    wire new_AGEMA_signal_6030 ;
    wire new_AGEMA_signal_6031 ;
    wire new_AGEMA_signal_6032 ;
    wire new_AGEMA_signal_6033 ;
    wire new_AGEMA_signal_6034 ;
    wire new_AGEMA_signal_6035 ;
    wire new_AGEMA_signal_6036 ;
    wire new_AGEMA_signal_6037 ;
    wire new_AGEMA_signal_6038 ;
    wire new_AGEMA_signal_6039 ;
    wire new_AGEMA_signal_6040 ;
    wire new_AGEMA_signal_6041 ;
    wire new_AGEMA_signal_6042 ;
    wire new_AGEMA_signal_6043 ;
    wire new_AGEMA_signal_6044 ;
    wire new_AGEMA_signal_6045 ;
    wire new_AGEMA_signal_6046 ;
    wire new_AGEMA_signal_6047 ;
    wire new_AGEMA_signal_6048 ;
    wire new_AGEMA_signal_6049 ;
    wire new_AGEMA_signal_6050 ;
    wire new_AGEMA_signal_6051 ;
    wire new_AGEMA_signal_6052 ;
    wire new_AGEMA_signal_6053 ;
    wire new_AGEMA_signal_6054 ;
    wire new_AGEMA_signal_6055 ;
    wire new_AGEMA_signal_6056 ;
    wire new_AGEMA_signal_6057 ;
    wire new_AGEMA_signal_6058 ;
    wire new_AGEMA_signal_6059 ;
    wire new_AGEMA_signal_6060 ;
    wire new_AGEMA_signal_6061 ;
    wire new_AGEMA_signal_6062 ;
    wire new_AGEMA_signal_6063 ;
    wire new_AGEMA_signal_6064 ;
    wire new_AGEMA_signal_6065 ;
    wire new_AGEMA_signal_6066 ;
    wire new_AGEMA_signal_6067 ;
    wire new_AGEMA_signal_6068 ;
    wire new_AGEMA_signal_6069 ;
    wire new_AGEMA_signal_6070 ;
    wire new_AGEMA_signal_6071 ;
    wire new_AGEMA_signal_6072 ;
    wire new_AGEMA_signal_6073 ;
    wire new_AGEMA_signal_6074 ;
    wire new_AGEMA_signal_6075 ;
    wire new_AGEMA_signal_6076 ;
    wire new_AGEMA_signal_6077 ;
    wire new_AGEMA_signal_6078 ;
    wire new_AGEMA_signal_6079 ;
    wire new_AGEMA_signal_6080 ;
    wire new_AGEMA_signal_6081 ;
    wire new_AGEMA_signal_6082 ;
    wire new_AGEMA_signal_6083 ;
    wire new_AGEMA_signal_6084 ;
    wire new_AGEMA_signal_6085 ;
    wire new_AGEMA_signal_6086 ;
    wire new_AGEMA_signal_6087 ;
    wire new_AGEMA_signal_6088 ;
    wire new_AGEMA_signal_6089 ;
    wire new_AGEMA_signal_6090 ;
    wire new_AGEMA_signal_6091 ;
    wire new_AGEMA_signal_6092 ;
    wire new_AGEMA_signal_6093 ;
    wire new_AGEMA_signal_6094 ;
    wire new_AGEMA_signal_6095 ;
    wire new_AGEMA_signal_6096 ;
    wire new_AGEMA_signal_6097 ;
    wire new_AGEMA_signal_6098 ;
    wire new_AGEMA_signal_6099 ;
    wire new_AGEMA_signal_6100 ;
    wire new_AGEMA_signal_6101 ;
    wire new_AGEMA_signal_6102 ;
    wire new_AGEMA_signal_6103 ;
    wire new_AGEMA_signal_6104 ;
    wire new_AGEMA_signal_6105 ;
    wire new_AGEMA_signal_6106 ;
    wire new_AGEMA_signal_6107 ;
    wire new_AGEMA_signal_6108 ;
    wire new_AGEMA_signal_6109 ;
    wire new_AGEMA_signal_6110 ;
    wire new_AGEMA_signal_6111 ;
    wire new_AGEMA_signal_6112 ;
    wire new_AGEMA_signal_6113 ;
    wire new_AGEMA_signal_6114 ;
    wire new_AGEMA_signal_6115 ;
    wire new_AGEMA_signal_6116 ;
    wire new_AGEMA_signal_6117 ;
    wire new_AGEMA_signal_6118 ;
    wire new_AGEMA_signal_6119 ;
    wire new_AGEMA_signal_6120 ;
    wire new_AGEMA_signal_6121 ;
    wire new_AGEMA_signal_6122 ;
    wire new_AGEMA_signal_6123 ;
    wire new_AGEMA_signal_6124 ;
    wire new_AGEMA_signal_6125 ;
    wire new_AGEMA_signal_6126 ;
    wire new_AGEMA_signal_6127 ;
    wire new_AGEMA_signal_6128 ;
    wire new_AGEMA_signal_6129 ;
    wire new_AGEMA_signal_6130 ;
    wire new_AGEMA_signal_6131 ;
    wire new_AGEMA_signal_6132 ;
    wire new_AGEMA_signal_6133 ;
    wire new_AGEMA_signal_6134 ;
    wire new_AGEMA_signal_6135 ;
    wire new_AGEMA_signal_6136 ;
    wire new_AGEMA_signal_6137 ;
    wire new_AGEMA_signal_6138 ;
    wire new_AGEMA_signal_6139 ;
    wire new_AGEMA_signal_6140 ;
    wire new_AGEMA_signal_6141 ;
    wire new_AGEMA_signal_6142 ;
    wire new_AGEMA_signal_6143 ;
    wire new_AGEMA_signal_6144 ;
    wire new_AGEMA_signal_6145 ;
    wire new_AGEMA_signal_6146 ;
    wire new_AGEMA_signal_6147 ;
    wire new_AGEMA_signal_6148 ;
    wire new_AGEMA_signal_6149 ;
    wire new_AGEMA_signal_6150 ;
    wire new_AGEMA_signal_6151 ;
    wire new_AGEMA_signal_6152 ;
    wire new_AGEMA_signal_6153 ;
    wire new_AGEMA_signal_6154 ;
    wire new_AGEMA_signal_6155 ;
    wire new_AGEMA_signal_6156 ;
    wire new_AGEMA_signal_6157 ;
    wire new_AGEMA_signal_6158 ;
    wire new_AGEMA_signal_6159 ;
    wire new_AGEMA_signal_6160 ;
    wire new_AGEMA_signal_6161 ;
    wire new_AGEMA_signal_6162 ;
    wire new_AGEMA_signal_6163 ;
    wire new_AGEMA_signal_6164 ;
    wire new_AGEMA_signal_6165 ;
    wire new_AGEMA_signal_6166 ;
    wire new_AGEMA_signal_6167 ;
    wire new_AGEMA_signal_6168 ;
    wire new_AGEMA_signal_6169 ;
    wire new_AGEMA_signal_6170 ;
    wire new_AGEMA_signal_6171 ;
    wire new_AGEMA_signal_6172 ;
    wire new_AGEMA_signal_6173 ;
    wire new_AGEMA_signal_6174 ;
    wire new_AGEMA_signal_6175 ;
    wire new_AGEMA_signal_6176 ;
    wire new_AGEMA_signal_6177 ;
    wire new_AGEMA_signal_6178 ;
    wire new_AGEMA_signal_6179 ;
    wire new_AGEMA_signal_6180 ;
    wire new_AGEMA_signal_6181 ;
    wire new_AGEMA_signal_6182 ;
    wire new_AGEMA_signal_6183 ;
    wire new_AGEMA_signal_6184 ;
    wire new_AGEMA_signal_6185 ;
    wire new_AGEMA_signal_6186 ;
    wire new_AGEMA_signal_6187 ;
    wire new_AGEMA_signal_6188 ;
    wire new_AGEMA_signal_6189 ;
    wire new_AGEMA_signal_6190 ;
    wire new_AGEMA_signal_6191 ;
    wire new_AGEMA_signal_6192 ;
    wire new_AGEMA_signal_6193 ;
    wire new_AGEMA_signal_6194 ;
    wire new_AGEMA_signal_6195 ;
    wire new_AGEMA_signal_6196 ;
    wire new_AGEMA_signal_6197 ;
    wire new_AGEMA_signal_6198 ;
    wire new_AGEMA_signal_6199 ;
    wire new_AGEMA_signal_6200 ;
    wire new_AGEMA_signal_6201 ;
    wire new_AGEMA_signal_6202 ;
    wire new_AGEMA_signal_6203 ;
    wire new_AGEMA_signal_6204 ;
    wire new_AGEMA_signal_6205 ;
    wire new_AGEMA_signal_6206 ;
    wire new_AGEMA_signal_6207 ;
    wire new_AGEMA_signal_6208 ;
    wire new_AGEMA_signal_6209 ;
    wire new_AGEMA_signal_6210 ;
    wire new_AGEMA_signal_6211 ;
    wire new_AGEMA_signal_6212 ;
    wire new_AGEMA_signal_6213 ;
    wire new_AGEMA_signal_6214 ;
    wire new_AGEMA_signal_6215 ;
    wire new_AGEMA_signal_6216 ;
    wire new_AGEMA_signal_6217 ;
    wire new_AGEMA_signal_6218 ;
    wire new_AGEMA_signal_6219 ;
    wire new_AGEMA_signal_6220 ;
    wire new_AGEMA_signal_6221 ;
    wire new_AGEMA_signal_6222 ;
    wire new_AGEMA_signal_6223 ;
    wire new_AGEMA_signal_6224 ;
    wire new_AGEMA_signal_6225 ;
    wire new_AGEMA_signal_6226 ;
    wire new_AGEMA_signal_6227 ;
    wire new_AGEMA_signal_6228 ;
    wire new_AGEMA_signal_6229 ;
    wire new_AGEMA_signal_6230 ;
    wire new_AGEMA_signal_6231 ;
    wire new_AGEMA_signal_6232 ;
    wire new_AGEMA_signal_6233 ;
    wire new_AGEMA_signal_6234 ;
    wire new_AGEMA_signal_6235 ;
    wire new_AGEMA_signal_6236 ;
    wire new_AGEMA_signal_6237 ;
    wire new_AGEMA_signal_6238 ;
    wire new_AGEMA_signal_6239 ;
    wire new_AGEMA_signal_6240 ;
    wire new_AGEMA_signal_6241 ;
    wire new_AGEMA_signal_6242 ;
    wire new_AGEMA_signal_6243 ;
    wire new_AGEMA_signal_6244 ;
    wire new_AGEMA_signal_6245 ;
    wire new_AGEMA_signal_6246 ;
    wire new_AGEMA_signal_6247 ;
    wire new_AGEMA_signal_6248 ;
    wire new_AGEMA_signal_6249 ;
    wire new_AGEMA_signal_6250 ;
    wire new_AGEMA_signal_6251 ;
    wire new_AGEMA_signal_6252 ;
    wire new_AGEMA_signal_6253 ;
    wire new_AGEMA_signal_6254 ;
    wire new_AGEMA_signal_6255 ;
    wire new_AGEMA_signal_6256 ;
    wire new_AGEMA_signal_6257 ;
    wire new_AGEMA_signal_6258 ;
    wire new_AGEMA_signal_6259 ;
    wire new_AGEMA_signal_6260 ;
    wire new_AGEMA_signal_6261 ;
    wire new_AGEMA_signal_6262 ;
    wire new_AGEMA_signal_6263 ;
    wire new_AGEMA_signal_6264 ;
    wire new_AGEMA_signal_6265 ;
    wire new_AGEMA_signal_6266 ;
    wire new_AGEMA_signal_6267 ;
    wire new_AGEMA_signal_6268 ;
    wire new_AGEMA_signal_6269 ;
    wire new_AGEMA_signal_6270 ;
    wire new_AGEMA_signal_6271 ;
    wire new_AGEMA_signal_6272 ;
    wire new_AGEMA_signal_6273 ;
    wire new_AGEMA_signal_6274 ;
    wire new_AGEMA_signal_6275 ;
    wire new_AGEMA_signal_6276 ;
    wire new_AGEMA_signal_6277 ;
    wire new_AGEMA_signal_6278 ;
    wire new_AGEMA_signal_6279 ;
    wire new_AGEMA_signal_6280 ;
    wire new_AGEMA_signal_6281 ;
    wire new_AGEMA_signal_6282 ;
    wire new_AGEMA_signal_6283 ;
    wire new_AGEMA_signal_6284 ;
    wire new_AGEMA_signal_6285 ;
    wire new_AGEMA_signal_6286 ;
    wire new_AGEMA_signal_6287 ;
    wire new_AGEMA_signal_6288 ;
    wire new_AGEMA_signal_6289 ;
    wire new_AGEMA_signal_6290 ;
    wire new_AGEMA_signal_6291 ;
    wire new_AGEMA_signal_6292 ;
    wire new_AGEMA_signal_6293 ;
    wire new_AGEMA_signal_6294 ;
    wire new_AGEMA_signal_6295 ;
    wire new_AGEMA_signal_6296 ;
    wire new_AGEMA_signal_6297 ;
    wire new_AGEMA_signal_6298 ;
    wire new_AGEMA_signal_6299 ;
    wire new_AGEMA_signal_6300 ;
    wire new_AGEMA_signal_6301 ;
    wire new_AGEMA_signal_6302 ;
    wire new_AGEMA_signal_6303 ;
    wire new_AGEMA_signal_6304 ;
    wire new_AGEMA_signal_6305 ;
    wire new_AGEMA_signal_6306 ;
    wire new_AGEMA_signal_6307 ;
    wire new_AGEMA_signal_6308 ;
    wire new_AGEMA_signal_6309 ;
    wire new_AGEMA_signal_6310 ;
    wire new_AGEMA_signal_6311 ;
    wire new_AGEMA_signal_6312 ;
    wire new_AGEMA_signal_6313 ;
    wire new_AGEMA_signal_6314 ;
    wire new_AGEMA_signal_6315 ;
    wire new_AGEMA_signal_6316 ;
    wire new_AGEMA_signal_6317 ;
    wire new_AGEMA_signal_6318 ;
    wire new_AGEMA_signal_6319 ;
    wire new_AGEMA_signal_6320 ;
    wire new_AGEMA_signal_6321 ;
    wire new_AGEMA_signal_6322 ;
    wire new_AGEMA_signal_6323 ;
    wire new_AGEMA_signal_6324 ;
    wire new_AGEMA_signal_6325 ;
    wire new_AGEMA_signal_6326 ;
    wire new_AGEMA_signal_6327 ;
    wire new_AGEMA_signal_6328 ;
    wire new_AGEMA_signal_6329 ;
    wire new_AGEMA_signal_6330 ;
    wire new_AGEMA_signal_6331 ;
    wire new_AGEMA_signal_6332 ;
    wire new_AGEMA_signal_6333 ;
    wire new_AGEMA_signal_6334 ;
    wire new_AGEMA_signal_6335 ;
    wire new_AGEMA_signal_6336 ;
    wire new_AGEMA_signal_6337 ;
    wire new_AGEMA_signal_6338 ;
    wire new_AGEMA_signal_6339 ;
    wire new_AGEMA_signal_6340 ;
    wire new_AGEMA_signal_6341 ;
    wire new_AGEMA_signal_6342 ;
    wire new_AGEMA_signal_6343 ;
    wire new_AGEMA_signal_6344 ;
    wire new_AGEMA_signal_6345 ;
    wire new_AGEMA_signal_6346 ;
    wire new_AGEMA_signal_6347 ;
    wire new_AGEMA_signal_6348 ;
    wire new_AGEMA_signal_6349 ;
    wire new_AGEMA_signal_6350 ;
    wire new_AGEMA_signal_6351 ;
    wire new_AGEMA_signal_6352 ;
    wire new_AGEMA_signal_6353 ;
    wire new_AGEMA_signal_6354 ;
    wire new_AGEMA_signal_6355 ;
    wire new_AGEMA_signal_6356 ;
    wire new_AGEMA_signal_6357 ;
    wire new_AGEMA_signal_6358 ;
    wire new_AGEMA_signal_6359 ;
    wire new_AGEMA_signal_6360 ;
    wire new_AGEMA_signal_6361 ;
    wire new_AGEMA_signal_6362 ;
    wire new_AGEMA_signal_6363 ;
    wire new_AGEMA_signal_6364 ;
    wire new_AGEMA_signal_6365 ;
    wire new_AGEMA_signal_6366 ;
    wire new_AGEMA_signal_6367 ;
    wire new_AGEMA_signal_6368 ;
    wire new_AGEMA_signal_6369 ;
    wire new_AGEMA_signal_6370 ;
    wire new_AGEMA_signal_6371 ;
    wire new_AGEMA_signal_6372 ;
    wire new_AGEMA_signal_6373 ;
    wire new_AGEMA_signal_6374 ;
    wire new_AGEMA_signal_6375 ;
    wire new_AGEMA_signal_6376 ;
    wire new_AGEMA_signal_6377 ;
    wire new_AGEMA_signal_6378 ;
    wire new_AGEMA_signal_6379 ;
    wire new_AGEMA_signal_6380 ;
    wire new_AGEMA_signal_6381 ;
    wire new_AGEMA_signal_6382 ;
    wire new_AGEMA_signal_6383 ;
    wire new_AGEMA_signal_6384 ;
    wire new_AGEMA_signal_6385 ;
    wire new_AGEMA_signal_6386 ;
    wire new_AGEMA_signal_6387 ;
    wire new_AGEMA_signal_6388 ;
    wire new_AGEMA_signal_6389 ;
    wire new_AGEMA_signal_6390 ;
    wire new_AGEMA_signal_6391 ;
    wire new_AGEMA_signal_6392 ;
    wire new_AGEMA_signal_6393 ;
    wire new_AGEMA_signal_6394 ;
    wire new_AGEMA_signal_6395 ;
    wire new_AGEMA_signal_6396 ;
    wire new_AGEMA_signal_6397 ;
    wire new_AGEMA_signal_6398 ;
    wire new_AGEMA_signal_6399 ;
    wire new_AGEMA_signal_6400 ;
    wire new_AGEMA_signal_6401 ;
    wire new_AGEMA_signal_6402 ;
    wire new_AGEMA_signal_6403 ;
    wire new_AGEMA_signal_6404 ;
    wire new_AGEMA_signal_6405 ;
    wire new_AGEMA_signal_6406 ;
    wire new_AGEMA_signal_6407 ;
    wire new_AGEMA_signal_6408 ;
    wire new_AGEMA_signal_6409 ;
    wire new_AGEMA_signal_6410 ;
    wire new_AGEMA_signal_6411 ;
    wire new_AGEMA_signal_6412 ;
    wire new_AGEMA_signal_6413 ;
    wire new_AGEMA_signal_6414 ;
    wire new_AGEMA_signal_6415 ;
    wire new_AGEMA_signal_6416 ;
    wire new_AGEMA_signal_6417 ;
    wire new_AGEMA_signal_6418 ;
    wire new_AGEMA_signal_6419 ;
    wire new_AGEMA_signal_6420 ;
    wire new_AGEMA_signal_6421 ;
    wire new_AGEMA_signal_6422 ;
    wire new_AGEMA_signal_6423 ;
    wire new_AGEMA_signal_6424 ;
    wire new_AGEMA_signal_6425 ;
    wire new_AGEMA_signal_6426 ;
    wire new_AGEMA_signal_6427 ;
    wire new_AGEMA_signal_6428 ;
    wire new_AGEMA_signal_6429 ;
    wire new_AGEMA_signal_6430 ;
    wire new_AGEMA_signal_6431 ;
    wire new_AGEMA_signal_6432 ;
    wire new_AGEMA_signal_6433 ;
    wire new_AGEMA_signal_6434 ;
    wire new_AGEMA_signal_6435 ;
    wire new_AGEMA_signal_6436 ;
    wire new_AGEMA_signal_6437 ;
    wire new_AGEMA_signal_6438 ;
    wire new_AGEMA_signal_6439 ;
    wire new_AGEMA_signal_6440 ;
    wire new_AGEMA_signal_6441 ;
    wire new_AGEMA_signal_6442 ;
    wire new_AGEMA_signal_6443 ;
    wire new_AGEMA_signal_6444 ;
    wire new_AGEMA_signal_6445 ;
    wire new_AGEMA_signal_6446 ;
    wire new_AGEMA_signal_6447 ;
    wire new_AGEMA_signal_6448 ;
    wire new_AGEMA_signal_6449 ;
    wire new_AGEMA_signal_6450 ;
    wire new_AGEMA_signal_6451 ;
    wire new_AGEMA_signal_6452 ;
    wire new_AGEMA_signal_6453 ;
    wire new_AGEMA_signal_6454 ;
    wire new_AGEMA_signal_6455 ;
    wire new_AGEMA_signal_6456 ;
    wire new_AGEMA_signal_6457 ;
    wire new_AGEMA_signal_6458 ;
    wire new_AGEMA_signal_6459 ;
    wire new_AGEMA_signal_6460 ;
    wire new_AGEMA_signal_6461 ;
    wire new_AGEMA_signal_6462 ;
    wire new_AGEMA_signal_6463 ;
    wire new_AGEMA_signal_6464 ;
    wire new_AGEMA_signal_6465 ;
    wire new_AGEMA_signal_6466 ;
    wire new_AGEMA_signal_6467 ;
    wire new_AGEMA_signal_6468 ;
    wire new_AGEMA_signal_6469 ;
    wire new_AGEMA_signal_6470 ;
    wire new_AGEMA_signal_6471 ;
    wire new_AGEMA_signal_6472 ;
    wire new_AGEMA_signal_6473 ;
    wire new_AGEMA_signal_6474 ;
    wire new_AGEMA_signal_6475 ;
    wire new_AGEMA_signal_6476 ;
    wire new_AGEMA_signal_6477 ;
    wire new_AGEMA_signal_6478 ;
    wire new_AGEMA_signal_6479 ;
    wire new_AGEMA_signal_6480 ;
    wire new_AGEMA_signal_6481 ;
    wire new_AGEMA_signal_6482 ;
    wire new_AGEMA_signal_6483 ;
    wire new_AGEMA_signal_6484 ;
    wire new_AGEMA_signal_6485 ;
    wire new_AGEMA_signal_6486 ;
    wire new_AGEMA_signal_6487 ;
    wire new_AGEMA_signal_6488 ;
    wire new_AGEMA_signal_6489 ;
    wire new_AGEMA_signal_6490 ;
    wire new_AGEMA_signal_6491 ;
    wire new_AGEMA_signal_6492 ;
    wire new_AGEMA_signal_6493 ;
    wire new_AGEMA_signal_6494 ;
    wire new_AGEMA_signal_6495 ;
    wire new_AGEMA_signal_6496 ;
    wire new_AGEMA_signal_6497 ;
    wire new_AGEMA_signal_6498 ;
    wire new_AGEMA_signal_6499 ;
    wire new_AGEMA_signal_6500 ;
    wire new_AGEMA_signal_6501 ;
    wire new_AGEMA_signal_6502 ;
    wire new_AGEMA_signal_6503 ;
    wire new_AGEMA_signal_6504 ;
    wire new_AGEMA_signal_6505 ;
    wire new_AGEMA_signal_6506 ;
    wire new_AGEMA_signal_6507 ;
    wire new_AGEMA_signal_6508 ;
    wire new_AGEMA_signal_6509 ;
    wire new_AGEMA_signal_6510 ;
    wire new_AGEMA_signal_6511 ;
    wire new_AGEMA_signal_6512 ;
    wire new_AGEMA_signal_6513 ;
    wire new_AGEMA_signal_6514 ;
    wire new_AGEMA_signal_6515 ;
    wire new_AGEMA_signal_6516 ;
    wire new_AGEMA_signal_6517 ;
    wire new_AGEMA_signal_6518 ;
    wire new_AGEMA_signal_6519 ;
    wire new_AGEMA_signal_6520 ;
    wire new_AGEMA_signal_6521 ;
    wire new_AGEMA_signal_6522 ;
    wire new_AGEMA_signal_6523 ;
    wire new_AGEMA_signal_6524 ;
    wire new_AGEMA_signal_6525 ;
    wire new_AGEMA_signal_6526 ;
    wire new_AGEMA_signal_6527 ;
    wire new_AGEMA_signal_6528 ;
    wire new_AGEMA_signal_6529 ;
    wire new_AGEMA_signal_6530 ;
    wire new_AGEMA_signal_6531 ;
    wire new_AGEMA_signal_6532 ;
    wire new_AGEMA_signal_6533 ;
    wire new_AGEMA_signal_6534 ;
    wire new_AGEMA_signal_6535 ;
    wire new_AGEMA_signal_6536 ;
    wire new_AGEMA_signal_6537 ;
    wire new_AGEMA_signal_6538 ;
    wire new_AGEMA_signal_6539 ;
    wire new_AGEMA_signal_6540 ;
    wire new_AGEMA_signal_6541 ;
    wire new_AGEMA_signal_6542 ;
    wire new_AGEMA_signal_6543 ;
    wire new_AGEMA_signal_6544 ;
    wire new_AGEMA_signal_6545 ;
    wire new_AGEMA_signal_6546 ;
    wire new_AGEMA_signal_6547 ;
    wire new_AGEMA_signal_6548 ;
    wire new_AGEMA_signal_6549 ;
    wire new_AGEMA_signal_6550 ;
    wire new_AGEMA_signal_6551 ;
    wire new_AGEMA_signal_6552 ;
    wire new_AGEMA_signal_6553 ;
    wire new_AGEMA_signal_6554 ;
    wire new_AGEMA_signal_6555 ;
    wire new_AGEMA_signal_6556 ;
    wire new_AGEMA_signal_6557 ;
    wire new_AGEMA_signal_6558 ;
    wire new_AGEMA_signal_6559 ;
    wire new_AGEMA_signal_6560 ;
    wire new_AGEMA_signal_6561 ;
    wire new_AGEMA_signal_6562 ;
    wire new_AGEMA_signal_6563 ;
    wire new_AGEMA_signal_6564 ;
    wire new_AGEMA_signal_6565 ;
    wire new_AGEMA_signal_6566 ;
    wire new_AGEMA_signal_6567 ;
    wire new_AGEMA_signal_6568 ;
    wire new_AGEMA_signal_6569 ;
    wire new_AGEMA_signal_6570 ;
    wire new_AGEMA_signal_6571 ;
    wire new_AGEMA_signal_6572 ;
    wire new_AGEMA_signal_6573 ;
    wire new_AGEMA_signal_6574 ;
    wire new_AGEMA_signal_6575 ;
    wire new_AGEMA_signal_6576 ;
    wire new_AGEMA_signal_6577 ;
    wire new_AGEMA_signal_6578 ;
    wire new_AGEMA_signal_6579 ;
    wire new_AGEMA_signal_6580 ;
    wire new_AGEMA_signal_6581 ;
    wire new_AGEMA_signal_6582 ;
    wire new_AGEMA_signal_6583 ;
    wire new_AGEMA_signal_6584 ;
    wire new_AGEMA_signal_6585 ;
    wire new_AGEMA_signal_6586 ;
    wire new_AGEMA_signal_6587 ;
    wire new_AGEMA_signal_6588 ;
    wire new_AGEMA_signal_6589 ;
    wire new_AGEMA_signal_6590 ;
    wire new_AGEMA_signal_6591 ;
    wire new_AGEMA_signal_6592 ;
    wire new_AGEMA_signal_6593 ;
    wire new_AGEMA_signal_6594 ;
    wire new_AGEMA_signal_6595 ;
    wire new_AGEMA_signal_6596 ;
    wire new_AGEMA_signal_6597 ;
    wire new_AGEMA_signal_6598 ;
    wire new_AGEMA_signal_6599 ;
    wire new_AGEMA_signal_6600 ;
    wire new_AGEMA_signal_6601 ;
    wire new_AGEMA_signal_6602 ;
    wire new_AGEMA_signal_6603 ;
    wire new_AGEMA_signal_6604 ;
    wire new_AGEMA_signal_6605 ;
    wire new_AGEMA_signal_6606 ;
    wire new_AGEMA_signal_6607 ;
    wire new_AGEMA_signal_6608 ;
    wire new_AGEMA_signal_6609 ;
    wire new_AGEMA_signal_6610 ;
    wire new_AGEMA_signal_6611 ;
    wire new_AGEMA_signal_6612 ;
    wire new_AGEMA_signal_6613 ;
    wire new_AGEMA_signal_6614 ;
    wire new_AGEMA_signal_6615 ;
    wire new_AGEMA_signal_6616 ;
    wire new_AGEMA_signal_6617 ;
    wire new_AGEMA_signal_6618 ;
    wire new_AGEMA_signal_6619 ;
    wire new_AGEMA_signal_6620 ;
    wire new_AGEMA_signal_6621 ;
    wire new_AGEMA_signal_6622 ;
    wire new_AGEMA_signal_6623 ;
    wire new_AGEMA_signal_6624 ;
    wire new_AGEMA_signal_6625 ;
    wire new_AGEMA_signal_6626 ;
    wire new_AGEMA_signal_6627 ;
    wire new_AGEMA_signal_6628 ;
    wire new_AGEMA_signal_6629 ;
    wire new_AGEMA_signal_6630 ;
    wire new_AGEMA_signal_6631 ;
    wire new_AGEMA_signal_6632 ;
    wire new_AGEMA_signal_6633 ;
    wire new_AGEMA_signal_6634 ;
    wire new_AGEMA_signal_6635 ;
    wire new_AGEMA_signal_6636 ;
    wire new_AGEMA_signal_6637 ;
    wire new_AGEMA_signal_6638 ;
    wire new_AGEMA_signal_6639 ;
    wire new_AGEMA_signal_6640 ;
    wire new_AGEMA_signal_6641 ;
    wire new_AGEMA_signal_6642 ;
    wire new_AGEMA_signal_6643 ;
    wire new_AGEMA_signal_6644 ;
    wire new_AGEMA_signal_6645 ;
    wire new_AGEMA_signal_6646 ;
    wire new_AGEMA_signal_6647 ;
    wire new_AGEMA_signal_6648 ;
    wire new_AGEMA_signal_6649 ;
    wire new_AGEMA_signal_6650 ;
    wire new_AGEMA_signal_6651 ;
    wire new_AGEMA_signal_6652 ;
    wire new_AGEMA_signal_6653 ;
    wire new_AGEMA_signal_6654 ;
    wire new_AGEMA_signal_6655 ;
    wire new_AGEMA_signal_6656 ;
    wire new_AGEMA_signal_6657 ;
    wire new_AGEMA_signal_6658 ;
    wire new_AGEMA_signal_6659 ;
    wire new_AGEMA_signal_6660 ;
    wire new_AGEMA_signal_6661 ;
    wire new_AGEMA_signal_6662 ;
    wire new_AGEMA_signal_6663 ;
    wire new_AGEMA_signal_6664 ;
    wire new_AGEMA_signal_6665 ;
    wire new_AGEMA_signal_6666 ;
    wire new_AGEMA_signal_6667 ;
    wire new_AGEMA_signal_6668 ;
    wire new_AGEMA_signal_6669 ;
    wire new_AGEMA_signal_6670 ;
    wire new_AGEMA_signal_6671 ;
    wire new_AGEMA_signal_6672 ;
    wire new_AGEMA_signal_6673 ;
    wire new_AGEMA_signal_6674 ;
    wire new_AGEMA_signal_6675 ;
    wire new_AGEMA_signal_6676 ;
    wire new_AGEMA_signal_6677 ;
    wire new_AGEMA_signal_6678 ;
    wire new_AGEMA_signal_6679 ;
    wire new_AGEMA_signal_6680 ;
    wire new_AGEMA_signal_6681 ;
    wire new_AGEMA_signal_6682 ;
    wire new_AGEMA_signal_6683 ;
    wire new_AGEMA_signal_6684 ;
    wire new_AGEMA_signal_6685 ;
    wire new_AGEMA_signal_6686 ;
    wire new_AGEMA_signal_6687 ;
    wire new_AGEMA_signal_6688 ;
    wire new_AGEMA_signal_6689 ;
    wire new_AGEMA_signal_6690 ;
    wire new_AGEMA_signal_6691 ;
    wire new_AGEMA_signal_6692 ;
    wire new_AGEMA_signal_6693 ;
    wire new_AGEMA_signal_6694 ;
    wire new_AGEMA_signal_6695 ;
    wire new_AGEMA_signal_6696 ;
    wire new_AGEMA_signal_6697 ;
    wire new_AGEMA_signal_6698 ;
    wire new_AGEMA_signal_6699 ;
    wire new_AGEMA_signal_6700 ;
    wire new_AGEMA_signal_6701 ;
    wire new_AGEMA_signal_6702 ;
    wire new_AGEMA_signal_6703 ;
    wire new_AGEMA_signal_6704 ;
    wire new_AGEMA_signal_6705 ;
    wire new_AGEMA_signal_6706 ;
    wire new_AGEMA_signal_6707 ;
    wire new_AGEMA_signal_6708 ;
    wire new_AGEMA_signal_6709 ;
    wire new_AGEMA_signal_6710 ;
    wire new_AGEMA_signal_6711 ;
    wire new_AGEMA_signal_6712 ;
    wire new_AGEMA_signal_6713 ;
    wire new_AGEMA_signal_6714 ;
    wire new_AGEMA_signal_6715 ;
    wire new_AGEMA_signal_6716 ;
    wire new_AGEMA_signal_6717 ;
    wire new_AGEMA_signal_6718 ;
    wire new_AGEMA_signal_6719 ;
    wire new_AGEMA_signal_6720 ;
    wire new_AGEMA_signal_6721 ;
    wire new_AGEMA_signal_6722 ;
    wire new_AGEMA_signal_6723 ;
    wire new_AGEMA_signal_6724 ;
    wire new_AGEMA_signal_6725 ;
    wire new_AGEMA_signal_6726 ;
    wire new_AGEMA_signal_6727 ;
    wire new_AGEMA_signal_6728 ;
    wire new_AGEMA_signal_6729 ;
    wire new_AGEMA_signal_6730 ;
    wire new_AGEMA_signal_6731 ;
    wire new_AGEMA_signal_6732 ;
    wire new_AGEMA_signal_6733 ;
    wire new_AGEMA_signal_6734 ;
    wire new_AGEMA_signal_6735 ;
    wire new_AGEMA_signal_6736 ;
    wire new_AGEMA_signal_6737 ;
    wire new_AGEMA_signal_6738 ;
    wire new_AGEMA_signal_6739 ;
    wire new_AGEMA_signal_6740 ;
    wire new_AGEMA_signal_6741 ;
    wire new_AGEMA_signal_6742 ;
    wire new_AGEMA_signal_6743 ;
    wire new_AGEMA_signal_6744 ;
    wire new_AGEMA_signal_6745 ;
    wire new_AGEMA_signal_6746 ;
    wire new_AGEMA_signal_6747 ;
    wire new_AGEMA_signal_6748 ;
    wire new_AGEMA_signal_6749 ;
    wire new_AGEMA_signal_6750 ;
    wire new_AGEMA_signal_6751 ;
    wire new_AGEMA_signal_6752 ;
    wire new_AGEMA_signal_6753 ;
    wire new_AGEMA_signal_6754 ;
    wire new_AGEMA_signal_6755 ;
    wire new_AGEMA_signal_6756 ;
    wire new_AGEMA_signal_6757 ;
    wire new_AGEMA_signal_6758 ;
    wire new_AGEMA_signal_6759 ;
    wire new_AGEMA_signal_6760 ;
    wire new_AGEMA_signal_6761 ;
    wire new_AGEMA_signal_6762 ;
    wire new_AGEMA_signal_6763 ;
    wire new_AGEMA_signal_6764 ;
    wire new_AGEMA_signal_6765 ;
    wire new_AGEMA_signal_6766 ;
    wire new_AGEMA_signal_6767 ;
    wire new_AGEMA_signal_6768 ;
    wire new_AGEMA_signal_6769 ;
    wire new_AGEMA_signal_6770 ;
    wire new_AGEMA_signal_6771 ;
    wire new_AGEMA_signal_6772 ;
    wire new_AGEMA_signal_6773 ;
    wire new_AGEMA_signal_6774 ;
    wire new_AGEMA_signal_6775 ;
    wire new_AGEMA_signal_6776 ;
    wire new_AGEMA_signal_6777 ;
    wire new_AGEMA_signal_6778 ;
    wire new_AGEMA_signal_6779 ;
    wire new_AGEMA_signal_6780 ;
    wire new_AGEMA_signal_6781 ;
    wire new_AGEMA_signal_6782 ;
    wire new_AGEMA_signal_6783 ;
    wire new_AGEMA_signal_6784 ;
    wire new_AGEMA_signal_6785 ;
    wire new_AGEMA_signal_6786 ;
    wire new_AGEMA_signal_6787 ;
    wire new_AGEMA_signal_6788 ;
    wire new_AGEMA_signal_6789 ;
    wire new_AGEMA_signal_6790 ;
    wire new_AGEMA_signal_6791 ;
    wire new_AGEMA_signal_6792 ;
    wire new_AGEMA_signal_6793 ;
    wire new_AGEMA_signal_6794 ;
    wire new_AGEMA_signal_6795 ;
    wire new_AGEMA_signal_6796 ;
    wire new_AGEMA_signal_6797 ;
    wire new_AGEMA_signal_6798 ;
    wire new_AGEMA_signal_6799 ;
    wire new_AGEMA_signal_6800 ;
    wire new_AGEMA_signal_6801 ;
    wire new_AGEMA_signal_6802 ;
    wire new_AGEMA_signal_6803 ;
    wire new_AGEMA_signal_6804 ;
    wire new_AGEMA_signal_6805 ;
    wire new_AGEMA_signal_6806 ;
    wire new_AGEMA_signal_6807 ;
    wire new_AGEMA_signal_6808 ;
    wire new_AGEMA_signal_6809 ;
    wire new_AGEMA_signal_6810 ;
    wire new_AGEMA_signal_6811 ;
    wire new_AGEMA_signal_6812 ;
    wire new_AGEMA_signal_6813 ;
    wire new_AGEMA_signal_6814 ;
    wire new_AGEMA_signal_6815 ;
    wire new_AGEMA_signal_6816 ;
    wire new_AGEMA_signal_6817 ;
    wire new_AGEMA_signal_6818 ;
    wire new_AGEMA_signal_6819 ;
    wire new_AGEMA_signal_6820 ;
    wire new_AGEMA_signal_6821 ;
    wire new_AGEMA_signal_6822 ;
    wire new_AGEMA_signal_6823 ;
    wire new_AGEMA_signal_6824 ;
    wire new_AGEMA_signal_6825 ;
    wire new_AGEMA_signal_6826 ;
    wire new_AGEMA_signal_6827 ;
    wire new_AGEMA_signal_6828 ;
    wire new_AGEMA_signal_6829 ;
    wire new_AGEMA_signal_6830 ;
    wire new_AGEMA_signal_6831 ;
    wire new_AGEMA_signal_6832 ;
    wire new_AGEMA_signal_6833 ;
    wire new_AGEMA_signal_6834 ;
    wire new_AGEMA_signal_6835 ;
    wire new_AGEMA_signal_6836 ;
    wire new_AGEMA_signal_6837 ;
    wire new_AGEMA_signal_6838 ;
    wire new_AGEMA_signal_6839 ;
    wire new_AGEMA_signal_6840 ;
    wire new_AGEMA_signal_6841 ;
    wire new_AGEMA_signal_6842 ;
    wire new_AGEMA_signal_6843 ;
    wire new_AGEMA_signal_6844 ;
    wire new_AGEMA_signal_6845 ;
    wire new_AGEMA_signal_6846 ;
    wire new_AGEMA_signal_6847 ;
    wire new_AGEMA_signal_6848 ;
    wire new_AGEMA_signal_6849 ;
    wire new_AGEMA_signal_6850 ;
    wire new_AGEMA_signal_6851 ;
    wire new_AGEMA_signal_6852 ;
    wire new_AGEMA_signal_6853 ;
    wire new_AGEMA_signal_6854 ;
    wire new_AGEMA_signal_6855 ;
    wire new_AGEMA_signal_6856 ;
    wire new_AGEMA_signal_6857 ;
    wire new_AGEMA_signal_6858 ;
    wire new_AGEMA_signal_6859 ;
    wire new_AGEMA_signal_6860 ;
    wire new_AGEMA_signal_6861 ;
    wire new_AGEMA_signal_6862 ;
    wire new_AGEMA_signal_6863 ;
    wire new_AGEMA_signal_6864 ;
    wire new_AGEMA_signal_6865 ;
    wire new_AGEMA_signal_6866 ;
    wire new_AGEMA_signal_6867 ;
    wire new_AGEMA_signal_6868 ;
    wire new_AGEMA_signal_6869 ;
    wire new_AGEMA_signal_6870 ;
    wire new_AGEMA_signal_6871 ;
    wire new_AGEMA_signal_6872 ;
    wire new_AGEMA_signal_6873 ;
    wire new_AGEMA_signal_6874 ;
    wire new_AGEMA_signal_6875 ;
    wire new_AGEMA_signal_6876 ;
    wire new_AGEMA_signal_6877 ;
    wire new_AGEMA_signal_6878 ;
    wire new_AGEMA_signal_6879 ;
    wire new_AGEMA_signal_6880 ;
    wire new_AGEMA_signal_6881 ;
    wire new_AGEMA_signal_6882 ;
    wire new_AGEMA_signal_6883 ;
    wire new_AGEMA_signal_6884 ;
    wire new_AGEMA_signal_6885 ;
    wire new_AGEMA_signal_6886 ;
    wire new_AGEMA_signal_6887 ;
    wire new_AGEMA_signal_6888 ;
    wire new_AGEMA_signal_6889 ;
    wire new_AGEMA_signal_6890 ;
    wire new_AGEMA_signal_6891 ;
    wire new_AGEMA_signal_6892 ;
    wire new_AGEMA_signal_6893 ;
    wire new_AGEMA_signal_6894 ;
    wire new_AGEMA_signal_6895 ;
    wire new_AGEMA_signal_6896 ;
    wire new_AGEMA_signal_6897 ;
    wire new_AGEMA_signal_6898 ;
    wire new_AGEMA_signal_6899 ;
    wire new_AGEMA_signal_6900 ;
    wire new_AGEMA_signal_6901 ;
    wire new_AGEMA_signal_6902 ;
    wire new_AGEMA_signal_6903 ;
    wire new_AGEMA_signal_6904 ;
    wire new_AGEMA_signal_6905 ;
    wire new_AGEMA_signal_6906 ;
    wire new_AGEMA_signal_6907 ;
    wire new_AGEMA_signal_6908 ;
    wire new_AGEMA_signal_6909 ;
    wire new_AGEMA_signal_6910 ;
    wire new_AGEMA_signal_6911 ;
    wire new_AGEMA_signal_6912 ;
    wire new_AGEMA_signal_6913 ;
    wire new_AGEMA_signal_6914 ;
    wire new_AGEMA_signal_6915 ;
    wire new_AGEMA_signal_6916 ;
    wire new_AGEMA_signal_6917 ;
    wire new_AGEMA_signal_6918 ;
    wire new_AGEMA_signal_6919 ;
    wire new_AGEMA_signal_6920 ;
    wire new_AGEMA_signal_6921 ;
    wire new_AGEMA_signal_6922 ;
    wire new_AGEMA_signal_6923 ;
    wire new_AGEMA_signal_6924 ;
    wire new_AGEMA_signal_6925 ;
    wire new_AGEMA_signal_6926 ;
    wire new_AGEMA_signal_6927 ;
    wire new_AGEMA_signal_6928 ;
    wire new_AGEMA_signal_6929 ;
    wire new_AGEMA_signal_6930 ;
    wire new_AGEMA_signal_6931 ;
    wire new_AGEMA_signal_6932 ;
    wire new_AGEMA_signal_6933 ;
    wire new_AGEMA_signal_6934 ;
    wire new_AGEMA_signal_6935 ;
    wire new_AGEMA_signal_6936 ;
    wire new_AGEMA_signal_6937 ;
    wire new_AGEMA_signal_6938 ;
    wire new_AGEMA_signal_6939 ;
    wire new_AGEMA_signal_6940 ;
    wire new_AGEMA_signal_6941 ;
    wire new_AGEMA_signal_6942 ;
    wire new_AGEMA_signal_6943 ;
    wire new_AGEMA_signal_6944 ;
    wire new_AGEMA_signal_6945 ;
    wire new_AGEMA_signal_6946 ;
    wire new_AGEMA_signal_6947 ;
    wire new_AGEMA_signal_6948 ;
    wire new_AGEMA_signal_6949 ;
    wire new_AGEMA_signal_6950 ;
    wire new_AGEMA_signal_6951 ;
    wire new_AGEMA_signal_6952 ;
    wire new_AGEMA_signal_6953 ;
    wire new_AGEMA_signal_6954 ;
    wire new_AGEMA_signal_6955 ;
    wire new_AGEMA_signal_6956 ;
    wire new_AGEMA_signal_6957 ;
    wire new_AGEMA_signal_6958 ;
    wire new_AGEMA_signal_6959 ;
    wire new_AGEMA_signal_6960 ;
    wire new_AGEMA_signal_6961 ;
    wire new_AGEMA_signal_6962 ;
    wire new_AGEMA_signal_6963 ;
    wire new_AGEMA_signal_6964 ;
    wire new_AGEMA_signal_6965 ;
    wire new_AGEMA_signal_6966 ;
    wire new_AGEMA_signal_6967 ;
    wire new_AGEMA_signal_6968 ;
    wire new_AGEMA_signal_6969 ;
    wire new_AGEMA_signal_6970 ;
    wire new_AGEMA_signal_6971 ;
    wire new_AGEMA_signal_6972 ;
    wire new_AGEMA_signal_6973 ;
    wire new_AGEMA_signal_6974 ;
    wire new_AGEMA_signal_6975 ;
    wire new_AGEMA_signal_6976 ;
    wire new_AGEMA_signal_6977 ;
    wire new_AGEMA_signal_6978 ;
    wire new_AGEMA_signal_6979 ;
    wire new_AGEMA_signal_6980 ;
    wire new_AGEMA_signal_6981 ;
    wire new_AGEMA_signal_6982 ;
    wire new_AGEMA_signal_6983 ;
    wire new_AGEMA_signal_6984 ;
    wire new_AGEMA_signal_6985 ;
    wire new_AGEMA_signal_6986 ;
    wire new_AGEMA_signal_6987 ;
    wire new_AGEMA_signal_6988 ;
    wire new_AGEMA_signal_6989 ;
    wire new_AGEMA_signal_6990 ;
    wire new_AGEMA_signal_6991 ;
    wire new_AGEMA_signal_6992 ;
    wire new_AGEMA_signal_6993 ;
    wire new_AGEMA_signal_6994 ;
    wire new_AGEMA_signal_6995 ;
    wire new_AGEMA_signal_6996 ;
    wire new_AGEMA_signal_6997 ;
    wire new_AGEMA_signal_6998 ;
    wire new_AGEMA_signal_6999 ;
    wire new_AGEMA_signal_7000 ;
    wire new_AGEMA_signal_7001 ;
    wire new_AGEMA_signal_7002 ;
    wire new_AGEMA_signal_7003 ;
    wire new_AGEMA_signal_7004 ;
    wire new_AGEMA_signal_7005 ;
    wire new_AGEMA_signal_7006 ;
    wire new_AGEMA_signal_7007 ;
    wire new_AGEMA_signal_7008 ;
    wire new_AGEMA_signal_7009 ;
    wire new_AGEMA_signal_7010 ;
    wire new_AGEMA_signal_7011 ;
    wire new_AGEMA_signal_7012 ;
    wire new_AGEMA_signal_7013 ;
    wire new_AGEMA_signal_7014 ;
    wire new_AGEMA_signal_7015 ;
    wire new_AGEMA_signal_7016 ;
    wire new_AGEMA_signal_7017 ;
    wire new_AGEMA_signal_7018 ;
    wire new_AGEMA_signal_7019 ;
    wire new_AGEMA_signal_7020 ;
    wire new_AGEMA_signal_7021 ;
    wire new_AGEMA_signal_7022 ;
    wire new_AGEMA_signal_7023 ;
    wire new_AGEMA_signal_7024 ;
    wire new_AGEMA_signal_7025 ;
    wire new_AGEMA_signal_7026 ;
    wire new_AGEMA_signal_7027 ;
    wire new_AGEMA_signal_7028 ;
    wire new_AGEMA_signal_7029 ;
    wire new_AGEMA_signal_7030 ;
    wire new_AGEMA_signal_7031 ;
    wire new_AGEMA_signal_7032 ;
    wire new_AGEMA_signal_7033 ;
    wire new_AGEMA_signal_7034 ;
    wire new_AGEMA_signal_7035 ;
    wire new_AGEMA_signal_7036 ;
    wire new_AGEMA_signal_7037 ;
    wire new_AGEMA_signal_7038 ;
    wire new_AGEMA_signal_7039 ;
    wire new_AGEMA_signal_7040 ;
    wire new_AGEMA_signal_7041 ;
    wire new_AGEMA_signal_7042 ;
    wire new_AGEMA_signal_7043 ;
    wire new_AGEMA_signal_7044 ;
    wire new_AGEMA_signal_7045 ;
    wire new_AGEMA_signal_7046 ;
    wire new_AGEMA_signal_7047 ;
    wire new_AGEMA_signal_7048 ;
    wire new_AGEMA_signal_7049 ;
    wire new_AGEMA_signal_7050 ;
    wire new_AGEMA_signal_7051 ;
    wire new_AGEMA_signal_7052 ;
    wire new_AGEMA_signal_7053 ;
    wire new_AGEMA_signal_7054 ;
    wire new_AGEMA_signal_7055 ;
    wire new_AGEMA_signal_7056 ;
    wire new_AGEMA_signal_7057 ;
    wire new_AGEMA_signal_7058 ;
    wire new_AGEMA_signal_7059 ;
    wire new_AGEMA_signal_7060 ;
    wire new_AGEMA_signal_7061 ;
    wire new_AGEMA_signal_7062 ;
    wire new_AGEMA_signal_7063 ;
    wire new_AGEMA_signal_7064 ;
    wire new_AGEMA_signal_7065 ;
    wire new_AGEMA_signal_7066 ;
    wire new_AGEMA_signal_7067 ;
    wire new_AGEMA_signal_7068 ;
    wire new_AGEMA_signal_7069 ;
    wire new_AGEMA_signal_7070 ;
    wire new_AGEMA_signal_7071 ;
    wire new_AGEMA_signal_7072 ;
    wire new_AGEMA_signal_7073 ;
    wire new_AGEMA_signal_7074 ;
    wire new_AGEMA_signal_7075 ;
    wire new_AGEMA_signal_7076 ;
    wire new_AGEMA_signal_7077 ;
    wire new_AGEMA_signal_7078 ;
    wire new_AGEMA_signal_7079 ;
    wire new_AGEMA_signal_7080 ;
    wire new_AGEMA_signal_7081 ;
    wire new_AGEMA_signal_7082 ;
    wire new_AGEMA_signal_7083 ;
    wire new_AGEMA_signal_7084 ;
    wire new_AGEMA_signal_7085 ;
    wire new_AGEMA_signal_7086 ;
    wire new_AGEMA_signal_7087 ;
    wire new_AGEMA_signal_7088 ;
    wire new_AGEMA_signal_7089 ;
    wire new_AGEMA_signal_7090 ;
    wire new_AGEMA_signal_7091 ;
    wire new_AGEMA_signal_7092 ;
    wire new_AGEMA_signal_7093 ;
    wire new_AGEMA_signal_7094 ;
    wire new_AGEMA_signal_7095 ;
    wire new_AGEMA_signal_7096 ;
    wire new_AGEMA_signal_7097 ;
    wire new_AGEMA_signal_7098 ;
    wire new_AGEMA_signal_7099 ;
    wire new_AGEMA_signal_7100 ;
    wire new_AGEMA_signal_7101 ;
    wire new_AGEMA_signal_7102 ;
    wire new_AGEMA_signal_7103 ;
    wire new_AGEMA_signal_7104 ;
    wire new_AGEMA_signal_7105 ;
    wire new_AGEMA_signal_7106 ;
    wire new_AGEMA_signal_7107 ;
    wire new_AGEMA_signal_7108 ;
    wire new_AGEMA_signal_7109 ;
    wire new_AGEMA_signal_7110 ;
    wire new_AGEMA_signal_7111 ;
    wire new_AGEMA_signal_7112 ;
    wire new_AGEMA_signal_7113 ;
    wire new_AGEMA_signal_7114 ;
    wire new_AGEMA_signal_7115 ;
    wire new_AGEMA_signal_7116 ;
    wire new_AGEMA_signal_7117 ;
    wire new_AGEMA_signal_7118 ;
    wire new_AGEMA_signal_7119 ;
    wire new_AGEMA_signal_7120 ;
    wire new_AGEMA_signal_7121 ;
    wire new_AGEMA_signal_7122 ;
    wire new_AGEMA_signal_7123 ;
    wire new_AGEMA_signal_7124 ;
    wire new_AGEMA_signal_7125 ;
    wire new_AGEMA_signal_7126 ;
    wire new_AGEMA_signal_7127 ;
    wire new_AGEMA_signal_7128 ;
    wire new_AGEMA_signal_7129 ;
    wire new_AGEMA_signal_7130 ;
    wire new_AGEMA_signal_7131 ;
    wire new_AGEMA_signal_7132 ;
    wire new_AGEMA_signal_7133 ;
    wire new_AGEMA_signal_7134 ;
    wire new_AGEMA_signal_7135 ;
    wire new_AGEMA_signal_7136 ;
    wire new_AGEMA_signal_7137 ;
    wire new_AGEMA_signal_7138 ;
    wire new_AGEMA_signal_7139 ;
    wire new_AGEMA_signal_7140 ;
    wire new_AGEMA_signal_7141 ;
    wire new_AGEMA_signal_7142 ;
    wire new_AGEMA_signal_7143 ;
    wire new_AGEMA_signal_7144 ;
    wire new_AGEMA_signal_7145 ;
    wire new_AGEMA_signal_7146 ;
    wire new_AGEMA_signal_7147 ;
    wire new_AGEMA_signal_7148 ;
    wire new_AGEMA_signal_7149 ;
    wire new_AGEMA_signal_7150 ;
    wire new_AGEMA_signal_7151 ;
    wire new_AGEMA_signal_7152 ;
    wire new_AGEMA_signal_7153 ;
    wire new_AGEMA_signal_7154 ;
    wire new_AGEMA_signal_7155 ;
    wire new_AGEMA_signal_7156 ;
    wire new_AGEMA_signal_7157 ;
    wire new_AGEMA_signal_7158 ;
    wire new_AGEMA_signal_7159 ;
    wire new_AGEMA_signal_7160 ;
    wire new_AGEMA_signal_7161 ;
    wire new_AGEMA_signal_7162 ;
    wire new_AGEMA_signal_7163 ;
    wire new_AGEMA_signal_7164 ;
    wire new_AGEMA_signal_7165 ;
    wire new_AGEMA_signal_7166 ;
    wire new_AGEMA_signal_7167 ;
    wire new_AGEMA_signal_7168 ;
    wire new_AGEMA_signal_7169 ;
    wire new_AGEMA_signal_7170 ;
    wire new_AGEMA_signal_7171 ;
    wire new_AGEMA_signal_7172 ;
    wire new_AGEMA_signal_7173 ;
    wire new_AGEMA_signal_7174 ;
    wire new_AGEMA_signal_7175 ;
    wire new_AGEMA_signal_7176 ;
    wire new_AGEMA_signal_7177 ;
    wire new_AGEMA_signal_7178 ;
    wire new_AGEMA_signal_7179 ;
    wire new_AGEMA_signal_7180 ;
    wire new_AGEMA_signal_7181 ;
    wire new_AGEMA_signal_7182 ;
    wire new_AGEMA_signal_7183 ;
    wire new_AGEMA_signal_7184 ;
    wire new_AGEMA_signal_7185 ;
    wire new_AGEMA_signal_7186 ;
    wire new_AGEMA_signal_7187 ;
    wire new_AGEMA_signal_7188 ;
    wire new_AGEMA_signal_7189 ;
    wire new_AGEMA_signal_7190 ;
    wire new_AGEMA_signal_7191 ;
    wire new_AGEMA_signal_7192 ;
    wire new_AGEMA_signal_7193 ;
    wire new_AGEMA_signal_7194 ;
    wire new_AGEMA_signal_7195 ;
    wire new_AGEMA_signal_7196 ;
    wire new_AGEMA_signal_7197 ;
    wire new_AGEMA_signal_7198 ;
    wire new_AGEMA_signal_7199 ;
    wire new_AGEMA_signal_7200 ;
    wire new_AGEMA_signal_7201 ;
    wire new_AGEMA_signal_7202 ;
    wire new_AGEMA_signal_7203 ;
    wire new_AGEMA_signal_7204 ;
    wire new_AGEMA_signal_7205 ;
    wire new_AGEMA_signal_7206 ;
    wire new_AGEMA_signal_7207 ;
    wire new_AGEMA_signal_7208 ;
    wire new_AGEMA_signal_7209 ;
    wire new_AGEMA_signal_7210 ;
    wire new_AGEMA_signal_7211 ;
    wire new_AGEMA_signal_7212 ;
    wire new_AGEMA_signal_7213 ;
    wire new_AGEMA_signal_7214 ;
    wire new_AGEMA_signal_7215 ;
    wire new_AGEMA_signal_7216 ;
    wire new_AGEMA_signal_7217 ;
    wire new_AGEMA_signal_7218 ;
    wire new_AGEMA_signal_7219 ;
    wire new_AGEMA_signal_7220 ;
    wire new_AGEMA_signal_7221 ;
    wire new_AGEMA_signal_7222 ;
    wire new_AGEMA_signal_7223 ;
    wire new_AGEMA_signal_7224 ;
    wire new_AGEMA_signal_7225 ;
    wire new_AGEMA_signal_7226 ;
    wire new_AGEMA_signal_7227 ;
    wire new_AGEMA_signal_7228 ;
    wire new_AGEMA_signal_7229 ;
    wire new_AGEMA_signal_7230 ;
    wire new_AGEMA_signal_7231 ;
    wire new_AGEMA_signal_7232 ;
    wire new_AGEMA_signal_7233 ;
    wire new_AGEMA_signal_7234 ;
    wire new_AGEMA_signal_7235 ;
    wire new_AGEMA_signal_7236 ;
    wire new_AGEMA_signal_7237 ;
    wire new_AGEMA_signal_7238 ;
    wire new_AGEMA_signal_7239 ;
    wire new_AGEMA_signal_7240 ;
    wire new_AGEMA_signal_7241 ;
    wire new_AGEMA_signal_7242 ;
    wire new_AGEMA_signal_7243 ;
    wire new_AGEMA_signal_7244 ;
    wire new_AGEMA_signal_7245 ;
    wire new_AGEMA_signal_7246 ;
    wire new_AGEMA_signal_7247 ;
    wire new_AGEMA_signal_7248 ;
    wire new_AGEMA_signal_7249 ;
    wire new_AGEMA_signal_7250 ;
    wire new_AGEMA_signal_7251 ;
    wire new_AGEMA_signal_7252 ;
    wire new_AGEMA_signal_7253 ;
    wire new_AGEMA_signal_7254 ;
    wire new_AGEMA_signal_7255 ;
    wire new_AGEMA_signal_7256 ;
    wire new_AGEMA_signal_7257 ;
    wire new_AGEMA_signal_7258 ;
    wire new_AGEMA_signal_7259 ;
    wire new_AGEMA_signal_7260 ;
    wire new_AGEMA_signal_7261 ;
    wire new_AGEMA_signal_7262 ;
    wire new_AGEMA_signal_7263 ;
    wire new_AGEMA_signal_7264 ;
    wire new_AGEMA_signal_7265 ;
    wire new_AGEMA_signal_7266 ;
    wire new_AGEMA_signal_7267 ;
    wire new_AGEMA_signal_7268 ;
    wire new_AGEMA_signal_7269 ;
    wire new_AGEMA_signal_7270 ;
    wire new_AGEMA_signal_7271 ;
    wire new_AGEMA_signal_7272 ;
    wire new_AGEMA_signal_7273 ;
    wire new_AGEMA_signal_7274 ;
    wire new_AGEMA_signal_7275 ;
    wire new_AGEMA_signal_7276 ;
    wire new_AGEMA_signal_7277 ;
    wire new_AGEMA_signal_7278 ;
    wire new_AGEMA_signal_7279 ;
    wire new_AGEMA_signal_7280 ;
    wire new_AGEMA_signal_7281 ;
    wire new_AGEMA_signal_7282 ;
    wire new_AGEMA_signal_7283 ;
    wire new_AGEMA_signal_7284 ;
    wire new_AGEMA_signal_7285 ;
    wire new_AGEMA_signal_7286 ;
    wire new_AGEMA_signal_7287 ;
    wire new_AGEMA_signal_7288 ;
    wire new_AGEMA_signal_7289 ;
    wire new_AGEMA_signal_7290 ;
    wire new_AGEMA_signal_7291 ;
    wire new_AGEMA_signal_7292 ;
    wire new_AGEMA_signal_7293 ;
    wire new_AGEMA_signal_7294 ;
    wire new_AGEMA_signal_7295 ;
    wire new_AGEMA_signal_7296 ;
    wire new_AGEMA_signal_7297 ;
    wire new_AGEMA_signal_7298 ;
    wire new_AGEMA_signal_7299 ;
    wire new_AGEMA_signal_7300 ;
    wire new_AGEMA_signal_7301 ;
    wire new_AGEMA_signal_7302 ;
    wire new_AGEMA_signal_7303 ;
    wire new_AGEMA_signal_7304 ;
    wire new_AGEMA_signal_7305 ;
    wire new_AGEMA_signal_7306 ;
    wire new_AGEMA_signal_7307 ;
    wire new_AGEMA_signal_7308 ;
    wire new_AGEMA_signal_7309 ;
    wire new_AGEMA_signal_7310 ;
    wire new_AGEMA_signal_7311 ;
    wire new_AGEMA_signal_7312 ;
    wire new_AGEMA_signal_7313 ;
    wire new_AGEMA_signal_7314 ;
    wire new_AGEMA_signal_7315 ;
    wire new_AGEMA_signal_7316 ;
    wire new_AGEMA_signal_7317 ;
    wire new_AGEMA_signal_7318 ;
    wire new_AGEMA_signal_7319 ;
    wire new_AGEMA_signal_7320 ;
    wire new_AGEMA_signal_7321 ;
    wire new_AGEMA_signal_7322 ;
    wire new_AGEMA_signal_7323 ;
    wire new_AGEMA_signal_7324 ;
    wire new_AGEMA_signal_7325 ;
    wire new_AGEMA_signal_7326 ;
    wire new_AGEMA_signal_7327 ;
    wire new_AGEMA_signal_7328 ;
    wire new_AGEMA_signal_7329 ;
    wire new_AGEMA_signal_7330 ;
    wire new_AGEMA_signal_7331 ;
    wire new_AGEMA_signal_7332 ;
    wire new_AGEMA_signal_7333 ;
    wire new_AGEMA_signal_7334 ;
    wire new_AGEMA_signal_7335 ;
    wire new_AGEMA_signal_7336 ;
    wire new_AGEMA_signal_7337 ;
    wire new_AGEMA_signal_7338 ;
    wire new_AGEMA_signal_7339 ;
    wire new_AGEMA_signal_7340 ;
    wire new_AGEMA_signal_7341 ;
    wire new_AGEMA_signal_7342 ;
    wire new_AGEMA_signal_7343 ;
    wire new_AGEMA_signal_7344 ;
    wire new_AGEMA_signal_7345 ;
    wire new_AGEMA_signal_7346 ;
    wire new_AGEMA_signal_7347 ;
    wire new_AGEMA_signal_7348 ;
    wire new_AGEMA_signal_7349 ;
    wire new_AGEMA_signal_7350 ;
    wire new_AGEMA_signal_7351 ;
    wire new_AGEMA_signal_7352 ;
    wire new_AGEMA_signal_7353 ;
    wire new_AGEMA_signal_7354 ;
    wire new_AGEMA_signal_7355 ;
    wire new_AGEMA_signal_7356 ;
    wire new_AGEMA_signal_7357 ;
    wire new_AGEMA_signal_7358 ;
    wire new_AGEMA_signal_7359 ;
    wire new_AGEMA_signal_7360 ;
    wire new_AGEMA_signal_7361 ;
    wire new_AGEMA_signal_7362 ;
    wire new_AGEMA_signal_7363 ;
    wire new_AGEMA_signal_7364 ;
    wire new_AGEMA_signal_7365 ;
    wire new_AGEMA_signal_7366 ;
    wire new_AGEMA_signal_7367 ;
    wire new_AGEMA_signal_7368 ;
    wire new_AGEMA_signal_7369 ;
    wire new_AGEMA_signal_7370 ;
    wire new_AGEMA_signal_7371 ;
    wire new_AGEMA_signal_7372 ;
    wire new_AGEMA_signal_7373 ;
    wire new_AGEMA_signal_7374 ;
    wire new_AGEMA_signal_7375 ;
    wire new_AGEMA_signal_7376 ;
    wire new_AGEMA_signal_7377 ;
    wire new_AGEMA_signal_7378 ;
    wire new_AGEMA_signal_7379 ;
    wire new_AGEMA_signal_7380 ;
    wire new_AGEMA_signal_7381 ;
    wire new_AGEMA_signal_7382 ;
    wire new_AGEMA_signal_7383 ;
    wire new_AGEMA_signal_7384 ;
    wire new_AGEMA_signal_7385 ;
    wire new_AGEMA_signal_7386 ;
    wire new_AGEMA_signal_7387 ;
    wire new_AGEMA_signal_7388 ;
    wire new_AGEMA_signal_7389 ;
    wire new_AGEMA_signal_7390 ;
    wire new_AGEMA_signal_7391 ;
    wire new_AGEMA_signal_7392 ;
    wire new_AGEMA_signal_7393 ;
    wire new_AGEMA_signal_7394 ;
    wire new_AGEMA_signal_7395 ;
    wire new_AGEMA_signal_7396 ;
    wire new_AGEMA_signal_7397 ;
    wire new_AGEMA_signal_7398 ;
    wire new_AGEMA_signal_7399 ;
    wire new_AGEMA_signal_7400 ;
    wire new_AGEMA_signal_7401 ;
    wire new_AGEMA_signal_7402 ;
    wire new_AGEMA_signal_7403 ;
    wire new_AGEMA_signal_7404 ;
    wire new_AGEMA_signal_7405 ;
    wire new_AGEMA_signal_7406 ;
    wire new_AGEMA_signal_7407 ;
    wire new_AGEMA_signal_7408 ;
    wire new_AGEMA_signal_7409 ;
    wire new_AGEMA_signal_7410 ;
    wire new_AGEMA_signal_7411 ;
    wire new_AGEMA_signal_7412 ;
    wire new_AGEMA_signal_7413 ;
    wire new_AGEMA_signal_7414 ;
    wire new_AGEMA_signal_7415 ;
    wire new_AGEMA_signal_7416 ;
    wire new_AGEMA_signal_7417 ;
    wire new_AGEMA_signal_7418 ;
    wire new_AGEMA_signal_7419 ;
    wire new_AGEMA_signal_7420 ;
    wire new_AGEMA_signal_7421 ;
    wire new_AGEMA_signal_7422 ;
    wire new_AGEMA_signal_7423 ;
    wire new_AGEMA_signal_7424 ;
    wire new_AGEMA_signal_7425 ;
    wire new_AGEMA_signal_7426 ;
    wire new_AGEMA_signal_7427 ;
    wire new_AGEMA_signal_7428 ;
    wire new_AGEMA_signal_7429 ;
    wire new_AGEMA_signal_7430 ;
    wire new_AGEMA_signal_7431 ;
    wire new_AGEMA_signal_7432 ;
    wire new_AGEMA_signal_7433 ;
    wire new_AGEMA_signal_7434 ;
    wire new_AGEMA_signal_7435 ;
    wire new_AGEMA_signal_7436 ;
    wire new_AGEMA_signal_7437 ;
    wire new_AGEMA_signal_7438 ;
    wire new_AGEMA_signal_7439 ;
    wire new_AGEMA_signal_7440 ;
    wire new_AGEMA_signal_7441 ;
    wire new_AGEMA_signal_7442 ;
    wire new_AGEMA_signal_7443 ;
    wire new_AGEMA_signal_7444 ;
    wire new_AGEMA_signal_7445 ;
    wire new_AGEMA_signal_7446 ;
    wire new_AGEMA_signal_7447 ;
    wire new_AGEMA_signal_7448 ;
    wire new_AGEMA_signal_7449 ;
    wire new_AGEMA_signal_7450 ;
    wire new_AGEMA_signal_7451 ;
    wire new_AGEMA_signal_7452 ;
    wire new_AGEMA_signal_7453 ;
    wire new_AGEMA_signal_7454 ;
    wire new_AGEMA_signal_7455 ;
    wire new_AGEMA_signal_7456 ;
    wire new_AGEMA_signal_7457 ;
    wire new_AGEMA_signal_7458 ;
    wire new_AGEMA_signal_7459 ;
    wire new_AGEMA_signal_7460 ;
    wire new_AGEMA_signal_7461 ;
    wire new_AGEMA_signal_7462 ;
    wire new_AGEMA_signal_7463 ;
    wire new_AGEMA_signal_7464 ;
    wire new_AGEMA_signal_7465 ;
    wire new_AGEMA_signal_7466 ;
    wire new_AGEMA_signal_7467 ;
    wire new_AGEMA_signal_7468 ;
    wire new_AGEMA_signal_7469 ;
    wire new_AGEMA_signal_7470 ;
    wire new_AGEMA_signal_7471 ;
    wire new_AGEMA_signal_7472 ;
    wire new_AGEMA_signal_7473 ;
    wire new_AGEMA_signal_7474 ;
    wire new_AGEMA_signal_7475 ;
    wire new_AGEMA_signal_7476 ;
    wire new_AGEMA_signal_7477 ;
    wire new_AGEMA_signal_7478 ;
    wire new_AGEMA_signal_7479 ;
    wire new_AGEMA_signal_7480 ;
    wire new_AGEMA_signal_7481 ;
    wire new_AGEMA_signal_7482 ;
    wire new_AGEMA_signal_7483 ;
    wire new_AGEMA_signal_7484 ;
    wire new_AGEMA_signal_7485 ;
    wire new_AGEMA_signal_7486 ;
    wire new_AGEMA_signal_7487 ;
    wire new_AGEMA_signal_7488 ;
    wire new_AGEMA_signal_7489 ;
    wire new_AGEMA_signal_7490 ;
    wire new_AGEMA_signal_7491 ;
    wire new_AGEMA_signal_7492 ;
    wire new_AGEMA_signal_7493 ;
    wire new_AGEMA_signal_7494 ;
    wire new_AGEMA_signal_7495 ;
    wire new_AGEMA_signal_7496 ;
    wire new_AGEMA_signal_7497 ;
    wire new_AGEMA_signal_7498 ;
    wire new_AGEMA_signal_7499 ;
    wire new_AGEMA_signal_7500 ;
    wire new_AGEMA_signal_7501 ;
    wire new_AGEMA_signal_7502 ;
    wire new_AGEMA_signal_7503 ;
    wire new_AGEMA_signal_7504 ;
    wire new_AGEMA_signal_7505 ;
    wire new_AGEMA_signal_7506 ;
    wire new_AGEMA_signal_7507 ;
    wire new_AGEMA_signal_7508 ;
    wire new_AGEMA_signal_7509 ;
    wire new_AGEMA_signal_7510 ;
    wire new_AGEMA_signal_7511 ;
    wire new_AGEMA_signal_7512 ;
    wire new_AGEMA_signal_7513 ;
    wire new_AGEMA_signal_7514 ;
    wire new_AGEMA_signal_7515 ;
    wire new_AGEMA_signal_7516 ;
    wire new_AGEMA_signal_7517 ;
    wire new_AGEMA_signal_7518 ;
    wire new_AGEMA_signal_7519 ;
    wire new_AGEMA_signal_7520 ;
    wire new_AGEMA_signal_7521 ;
    wire new_AGEMA_signal_7522 ;
    wire new_AGEMA_signal_7523 ;
    wire new_AGEMA_signal_7524 ;
    wire new_AGEMA_signal_7525 ;
    wire new_AGEMA_signal_7526 ;
    wire new_AGEMA_signal_7527 ;
    wire new_AGEMA_signal_7528 ;
    wire new_AGEMA_signal_7529 ;
    wire new_AGEMA_signal_7530 ;
    wire new_AGEMA_signal_7531 ;
    wire new_AGEMA_signal_7532 ;
    wire new_AGEMA_signal_7533 ;
    wire new_AGEMA_signal_7534 ;
    wire new_AGEMA_signal_7535 ;
    wire new_AGEMA_signal_7536 ;
    wire new_AGEMA_signal_7537 ;
    wire new_AGEMA_signal_7538 ;
    wire new_AGEMA_signal_7539 ;
    wire new_AGEMA_signal_7540 ;
    wire new_AGEMA_signal_7541 ;
    wire new_AGEMA_signal_7542 ;
    wire new_AGEMA_signal_7543 ;
    wire new_AGEMA_signal_7544 ;
    wire new_AGEMA_signal_7545 ;
    wire new_AGEMA_signal_7546 ;
    wire new_AGEMA_signal_7547 ;
    wire new_AGEMA_signal_7548 ;
    wire new_AGEMA_signal_7549 ;
    wire new_AGEMA_signal_7550 ;
    wire new_AGEMA_signal_7551 ;
    wire new_AGEMA_signal_7552 ;
    wire new_AGEMA_signal_7553 ;
    wire new_AGEMA_signal_7554 ;
    wire new_AGEMA_signal_7555 ;
    wire new_AGEMA_signal_7556 ;
    wire new_AGEMA_signal_7557 ;
    wire new_AGEMA_signal_7558 ;
    wire new_AGEMA_signal_7559 ;
    wire new_AGEMA_signal_7560 ;
    wire new_AGEMA_signal_7561 ;
    wire new_AGEMA_signal_7562 ;
    wire new_AGEMA_signal_7563 ;
    wire new_AGEMA_signal_7564 ;
    wire new_AGEMA_signal_7565 ;
    wire new_AGEMA_signal_7566 ;
    wire new_AGEMA_signal_7567 ;
    wire new_AGEMA_signal_7568 ;
    wire new_AGEMA_signal_7569 ;
    wire new_AGEMA_signal_7570 ;
    wire new_AGEMA_signal_7571 ;
    wire new_AGEMA_signal_7572 ;
    wire new_AGEMA_signal_7573 ;
    wire new_AGEMA_signal_7574 ;
    wire new_AGEMA_signal_7575 ;
    wire new_AGEMA_signal_7576 ;
    wire new_AGEMA_signal_7577 ;
    wire new_AGEMA_signal_7578 ;
    wire new_AGEMA_signal_7579 ;
    wire new_AGEMA_signal_7580 ;
    wire new_AGEMA_signal_7581 ;
    wire new_AGEMA_signal_7582 ;
    wire new_AGEMA_signal_7583 ;
    wire new_AGEMA_signal_7584 ;
    wire new_AGEMA_signal_7585 ;
    wire new_AGEMA_signal_7586 ;
    wire new_AGEMA_signal_7587 ;
    wire new_AGEMA_signal_7588 ;
    wire new_AGEMA_signal_7589 ;
    wire new_AGEMA_signal_7590 ;
    wire new_AGEMA_signal_7591 ;
    wire new_AGEMA_signal_7592 ;
    wire new_AGEMA_signal_7593 ;
    wire new_AGEMA_signal_7594 ;
    wire new_AGEMA_signal_7595 ;
    wire new_AGEMA_signal_7596 ;
    wire new_AGEMA_signal_7597 ;
    wire new_AGEMA_signal_7598 ;
    wire new_AGEMA_signal_7599 ;
    wire new_AGEMA_signal_7600 ;
    wire new_AGEMA_signal_7601 ;
    wire new_AGEMA_signal_7602 ;
    wire new_AGEMA_signal_7603 ;
    wire new_AGEMA_signal_7604 ;
    wire new_AGEMA_signal_7605 ;
    wire new_AGEMA_signal_7606 ;
    wire new_AGEMA_signal_7607 ;
    wire new_AGEMA_signal_7608 ;
    wire new_AGEMA_signal_7609 ;
    wire new_AGEMA_signal_7610 ;
    wire new_AGEMA_signal_7611 ;
    wire new_AGEMA_signal_7612 ;
    wire new_AGEMA_signal_7613 ;
    wire new_AGEMA_signal_7614 ;
    wire new_AGEMA_signal_7615 ;
    wire new_AGEMA_signal_7616 ;
    wire new_AGEMA_signal_7617 ;
    wire new_AGEMA_signal_7618 ;
    wire new_AGEMA_signal_7619 ;
    wire new_AGEMA_signal_7620 ;
    wire new_AGEMA_signal_7621 ;
    wire new_AGEMA_signal_7622 ;
    wire new_AGEMA_signal_7623 ;
    wire new_AGEMA_signal_7624 ;
    wire new_AGEMA_signal_7625 ;
    wire new_AGEMA_signal_7626 ;
    wire new_AGEMA_signal_7627 ;
    wire new_AGEMA_signal_7628 ;
    wire new_AGEMA_signal_7629 ;
    wire new_AGEMA_signal_7630 ;
    wire new_AGEMA_signal_7631 ;
    wire new_AGEMA_signal_7632 ;
    wire new_AGEMA_signal_7633 ;
    wire new_AGEMA_signal_7634 ;
    wire new_AGEMA_signal_7635 ;
    wire new_AGEMA_signal_7636 ;
    wire new_AGEMA_signal_7637 ;
    wire new_AGEMA_signal_7638 ;
    wire new_AGEMA_signal_7639 ;
    wire new_AGEMA_signal_7640 ;
    wire new_AGEMA_signal_7641 ;
    wire new_AGEMA_signal_7642 ;
    wire new_AGEMA_signal_7643 ;
    wire new_AGEMA_signal_7644 ;
    wire new_AGEMA_signal_7645 ;
    wire new_AGEMA_signal_7646 ;
    wire new_AGEMA_signal_7647 ;
    wire new_AGEMA_signal_7648 ;
    wire new_AGEMA_signal_7649 ;
    wire new_AGEMA_signal_7650 ;
    wire new_AGEMA_signal_7651 ;
    wire new_AGEMA_signal_7652 ;
    wire new_AGEMA_signal_7653 ;
    wire new_AGEMA_signal_7654 ;
    wire new_AGEMA_signal_7655 ;
    wire new_AGEMA_signal_7656 ;
    wire new_AGEMA_signal_7657 ;
    wire new_AGEMA_signal_7658 ;
    wire new_AGEMA_signal_7659 ;
    wire new_AGEMA_signal_7660 ;
    wire new_AGEMA_signal_7661 ;
    wire new_AGEMA_signal_7662 ;
    wire new_AGEMA_signal_7663 ;
    wire new_AGEMA_signal_7664 ;
    wire new_AGEMA_signal_7665 ;
    wire new_AGEMA_signal_7666 ;
    wire new_AGEMA_signal_7667 ;
    wire new_AGEMA_signal_7668 ;
    wire new_AGEMA_signal_7669 ;
    wire new_AGEMA_signal_7670 ;
    wire new_AGEMA_signal_7671 ;
    wire new_AGEMA_signal_7672 ;
    wire new_AGEMA_signal_7673 ;
    wire new_AGEMA_signal_7674 ;
    wire new_AGEMA_signal_7675 ;
    wire new_AGEMA_signal_7676 ;
    wire new_AGEMA_signal_7677 ;
    wire new_AGEMA_signal_7678 ;
    wire new_AGEMA_signal_7679 ;
    wire new_AGEMA_signal_7680 ;
    wire new_AGEMA_signal_7681 ;
    wire new_AGEMA_signal_7682 ;
    wire new_AGEMA_signal_7683 ;
    wire new_AGEMA_signal_7684 ;
    wire new_AGEMA_signal_7685 ;
    wire new_AGEMA_signal_7686 ;
    wire new_AGEMA_signal_7687 ;
    wire new_AGEMA_signal_7688 ;
    wire new_AGEMA_signal_7689 ;
    wire new_AGEMA_signal_7690 ;
    wire new_AGEMA_signal_7691 ;
    wire new_AGEMA_signal_7692 ;
    wire new_AGEMA_signal_7693 ;
    wire new_AGEMA_signal_7694 ;
    wire new_AGEMA_signal_7695 ;
    wire new_AGEMA_signal_7696 ;
    wire new_AGEMA_signal_7697 ;
    wire new_AGEMA_signal_7698 ;
    wire new_AGEMA_signal_7699 ;
    wire new_AGEMA_signal_7700 ;
    wire new_AGEMA_signal_7701 ;
    wire new_AGEMA_signal_7702 ;
    wire new_AGEMA_signal_7703 ;
    wire new_AGEMA_signal_7704 ;
    wire new_AGEMA_signal_7705 ;
    wire new_AGEMA_signal_7706 ;
    wire new_AGEMA_signal_7707 ;
    wire new_AGEMA_signal_7708 ;
    wire new_AGEMA_signal_7709 ;
    wire new_AGEMA_signal_7710 ;
    wire new_AGEMA_signal_7711 ;
    wire new_AGEMA_signal_7712 ;
    wire new_AGEMA_signal_7713 ;
    wire new_AGEMA_signal_7714 ;
    wire new_AGEMA_signal_7715 ;
    wire new_AGEMA_signal_7716 ;
    wire new_AGEMA_signal_7717 ;
    wire new_AGEMA_signal_7718 ;
    wire new_AGEMA_signal_7719 ;
    wire new_AGEMA_signal_7720 ;
    wire new_AGEMA_signal_7721 ;
    wire new_AGEMA_signal_7722 ;
    wire new_AGEMA_signal_7723 ;
    wire new_AGEMA_signal_7724 ;
    wire new_AGEMA_signal_7725 ;
    wire new_AGEMA_signal_7726 ;
    wire new_AGEMA_signal_7727 ;
    wire new_AGEMA_signal_7728 ;
    wire new_AGEMA_signal_7729 ;
    wire new_AGEMA_signal_7730 ;
    wire new_AGEMA_signal_7731 ;
    wire new_AGEMA_signal_7732 ;
    wire new_AGEMA_signal_7733 ;
    wire new_AGEMA_signal_7734 ;
    wire new_AGEMA_signal_7735 ;
    wire new_AGEMA_signal_7736 ;
    wire new_AGEMA_signal_7737 ;
    wire new_AGEMA_signal_7738 ;
    wire new_AGEMA_signal_7739 ;
    wire new_AGEMA_signal_7740 ;
    wire new_AGEMA_signal_7741 ;
    wire new_AGEMA_signal_7742 ;
    wire new_AGEMA_signal_7743 ;
    wire new_AGEMA_signal_7744 ;
    wire new_AGEMA_signal_7745 ;
    wire new_AGEMA_signal_7746 ;
    wire new_AGEMA_signal_7747 ;
    wire new_AGEMA_signal_7748 ;
    wire new_AGEMA_signal_7749 ;
    wire new_AGEMA_signal_7750 ;
    wire new_AGEMA_signal_7751 ;
    wire new_AGEMA_signal_7752 ;
    wire new_AGEMA_signal_7753 ;
    wire new_AGEMA_signal_7754 ;
    wire new_AGEMA_signal_7755 ;
    wire new_AGEMA_signal_7756 ;
    wire new_AGEMA_signal_7757 ;
    wire new_AGEMA_signal_7758 ;
    wire new_AGEMA_signal_7759 ;
    wire new_AGEMA_signal_7760 ;
    wire new_AGEMA_signal_7761 ;
    wire new_AGEMA_signal_7762 ;
    wire new_AGEMA_signal_7763 ;
    wire new_AGEMA_signal_7764 ;
    wire new_AGEMA_signal_7765 ;
    wire new_AGEMA_signal_7766 ;
    wire new_AGEMA_signal_7767 ;
    wire new_AGEMA_signal_7768 ;
    wire new_AGEMA_signal_7769 ;
    wire new_AGEMA_signal_7770 ;
    wire new_AGEMA_signal_7771 ;
    wire new_AGEMA_signal_7772 ;
    wire new_AGEMA_signal_7773 ;
    wire new_AGEMA_signal_7774 ;
    wire new_AGEMA_signal_7775 ;
    wire new_AGEMA_signal_7776 ;
    wire new_AGEMA_signal_7777 ;
    wire new_AGEMA_signal_7778 ;
    wire new_AGEMA_signal_7779 ;
    wire new_AGEMA_signal_7780 ;
    wire new_AGEMA_signal_7781 ;
    wire new_AGEMA_signal_7782 ;
    wire new_AGEMA_signal_7783 ;
    wire new_AGEMA_signal_7784 ;
    wire new_AGEMA_signal_7785 ;
    wire new_AGEMA_signal_7786 ;
    wire new_AGEMA_signal_7787 ;
    wire new_AGEMA_signal_7788 ;
    wire new_AGEMA_signal_7789 ;
    wire new_AGEMA_signal_7790 ;
    wire new_AGEMA_signal_7791 ;
    wire new_AGEMA_signal_7792 ;
    wire new_AGEMA_signal_7796 ;
    wire new_AGEMA_signal_7797 ;
    wire new_AGEMA_signal_7798 ;
    wire new_AGEMA_signal_7799 ;
    wire new_AGEMA_signal_7800 ;
    wire new_AGEMA_signal_7801 ;
    wire new_AGEMA_signal_7802 ;
    wire new_AGEMA_signal_7803 ;
    wire new_AGEMA_signal_7804 ;
    wire new_AGEMA_signal_7805 ;
    wire new_AGEMA_signal_7806 ;
    wire new_AGEMA_signal_7807 ;
    wire new_AGEMA_signal_7808 ;
    wire new_AGEMA_signal_7809 ;
    wire new_AGEMA_signal_7810 ;
    wire new_AGEMA_signal_7811 ;
    wire new_AGEMA_signal_7812 ;
    wire new_AGEMA_signal_7813 ;
    wire new_AGEMA_signal_7814 ;
    wire new_AGEMA_signal_7815 ;
    wire new_AGEMA_signal_7816 ;
    wire new_AGEMA_signal_7817 ;
    wire new_AGEMA_signal_7818 ;
    wire new_AGEMA_signal_7819 ;
    wire new_AGEMA_signal_7820 ;
    wire new_AGEMA_signal_7821 ;
    wire new_AGEMA_signal_7822 ;
    wire new_AGEMA_signal_7826 ;
    wire new_AGEMA_signal_7827 ;
    wire new_AGEMA_signal_7828 ;
    wire new_AGEMA_signal_7832 ;
    wire new_AGEMA_signal_7833 ;
    wire new_AGEMA_signal_7834 ;
    wire new_AGEMA_signal_7838 ;
    wire new_AGEMA_signal_7839 ;
    wire new_AGEMA_signal_7840 ;
    wire new_AGEMA_signal_7844 ;
    wire new_AGEMA_signal_7845 ;
    wire new_AGEMA_signal_7846 ;
    wire new_AGEMA_signal_7850 ;
    wire new_AGEMA_signal_7851 ;
    wire new_AGEMA_signal_7852 ;
    wire new_AGEMA_signal_7856 ;
    wire new_AGEMA_signal_7857 ;
    wire new_AGEMA_signal_7858 ;
    wire new_AGEMA_signal_7862 ;
    wire new_AGEMA_signal_7863 ;
    wire new_AGEMA_signal_7864 ;
    wire new_AGEMA_signal_7865 ;
    wire new_AGEMA_signal_7866 ;
    wire new_AGEMA_signal_7867 ;
    wire new_AGEMA_signal_7868 ;
    wire new_AGEMA_signal_7869 ;
    wire new_AGEMA_signal_7870 ;
    wire new_AGEMA_signal_7871 ;
    wire new_AGEMA_signal_7872 ;
    wire new_AGEMA_signal_7873 ;
    wire new_AGEMA_signal_7874 ;
    wire new_AGEMA_signal_7875 ;
    wire new_AGEMA_signal_7876 ;
    wire new_AGEMA_signal_7877 ;
    wire new_AGEMA_signal_7878 ;
    wire new_AGEMA_signal_7879 ;
    wire new_AGEMA_signal_7880 ;
    wire new_AGEMA_signal_7881 ;
    wire new_AGEMA_signal_7882 ;
    wire new_AGEMA_signal_7883 ;
    wire new_AGEMA_signal_7884 ;
    wire new_AGEMA_signal_7885 ;
    wire new_AGEMA_signal_7886 ;
    wire new_AGEMA_signal_7887 ;
    wire new_AGEMA_signal_7888 ;
    wire new_AGEMA_signal_7889 ;
    wire new_AGEMA_signal_7890 ;
    wire new_AGEMA_signal_7891 ;
    wire new_AGEMA_signal_7892 ;
    wire new_AGEMA_signal_7893 ;
    wire new_AGEMA_signal_7894 ;
    wire new_AGEMA_signal_7895 ;
    wire new_AGEMA_signal_7896 ;
    wire new_AGEMA_signal_7897 ;
    wire new_AGEMA_signal_7898 ;
    wire new_AGEMA_signal_7899 ;
    wire new_AGEMA_signal_7900 ;
    wire new_AGEMA_signal_7901 ;
    wire new_AGEMA_signal_7902 ;
    wire new_AGEMA_signal_7903 ;
    wire new_AGEMA_signal_7904 ;
    wire new_AGEMA_signal_7905 ;
    wire new_AGEMA_signal_7906 ;
    wire new_AGEMA_signal_7907 ;
    wire new_AGEMA_signal_7908 ;
    wire new_AGEMA_signal_7909 ;
    wire new_AGEMA_signal_7910 ;
    wire new_AGEMA_signal_7911 ;
    wire new_AGEMA_signal_7912 ;
    wire new_AGEMA_signal_7913 ;
    wire new_AGEMA_signal_7914 ;
    wire new_AGEMA_signal_7915 ;
    wire new_AGEMA_signal_7916 ;
    wire new_AGEMA_signal_7917 ;
    wire new_AGEMA_signal_7918 ;
    wire new_AGEMA_signal_7919 ;
    wire new_AGEMA_signal_7920 ;
    wire new_AGEMA_signal_7921 ;
    wire new_AGEMA_signal_7922 ;
    wire new_AGEMA_signal_7923 ;
    wire new_AGEMA_signal_7924 ;
    wire new_AGEMA_signal_7925 ;
    wire new_AGEMA_signal_7926 ;
    wire new_AGEMA_signal_7927 ;
    wire new_AGEMA_signal_7928 ;
    wire new_AGEMA_signal_7929 ;
    wire new_AGEMA_signal_7930 ;
    wire new_AGEMA_signal_7931 ;
    wire new_AGEMA_signal_7932 ;
    wire new_AGEMA_signal_7933 ;
    wire new_AGEMA_signal_7934 ;
    wire new_AGEMA_signal_7935 ;
    wire new_AGEMA_signal_7936 ;
    wire new_AGEMA_signal_7937 ;
    wire new_AGEMA_signal_7938 ;
    wire new_AGEMA_signal_7939 ;
    wire new_AGEMA_signal_7940 ;
    wire new_AGEMA_signal_7941 ;
    wire new_AGEMA_signal_7942 ;
    wire new_AGEMA_signal_7943 ;
    wire new_AGEMA_signal_7944 ;
    wire new_AGEMA_signal_7945 ;
    wire new_AGEMA_signal_7946 ;
    wire new_AGEMA_signal_7947 ;
    wire new_AGEMA_signal_7948 ;
    wire new_AGEMA_signal_7949 ;
    wire new_AGEMA_signal_7950 ;
    wire new_AGEMA_signal_7951 ;
    wire new_AGEMA_signal_7952 ;
    wire new_AGEMA_signal_7953 ;
    wire new_AGEMA_signal_7954 ;
    wire new_AGEMA_signal_7955 ;
    wire new_AGEMA_signal_7956 ;
    wire new_AGEMA_signal_7957 ;

    /* cells in depth 0 */
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) U23 ( .A0_t (ctrl_n4), .A0_f (new_AGEMA_signal_5778), .B0_t (start_t), .B0_f (start_f), .Z0_t (enKS), .Z0_f (new_AGEMA_signal_5916) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U25 ( .A0_t (keyStateIn[0]), .A0_f (new_AGEMA_signal_2489), .A1_t (new_AGEMA_signal_2490), .A1_f (new_AGEMA_signal_2491), .B0_t (port_out_s0_t[0]), .B0_f (port_out_s0_f[0]), .B1_t (port_out_s1_t[0]), .B1_f (port_out_s1_f[0]), .Z0_t (StateOutXORroundKey[0]), .Z0_f (new_AGEMA_signal_2495), .Z1_t (new_AGEMA_signal_2496), .Z1_f (new_AGEMA_signal_2497) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U26 ( .A0_t (keyStateIn[1]), .A0_f (new_AGEMA_signal_2498), .A1_t (new_AGEMA_signal_2499), .A1_f (new_AGEMA_signal_2500), .B0_t (port_out_s0_t[1]), .B0_f (port_out_s0_f[1]), .B1_t (port_out_s1_t[1]), .B1_f (port_out_s1_f[1]), .Z0_t (StateOutXORroundKey[1]), .Z0_f (new_AGEMA_signal_2504), .Z1_t (new_AGEMA_signal_2505), .Z1_f (new_AGEMA_signal_2506) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U27 ( .A0_t (keyStateIn[2]), .A0_f (new_AGEMA_signal_2507), .A1_t (new_AGEMA_signal_2508), .A1_f (new_AGEMA_signal_2509), .B0_t (port_out_s0_t[2]), .B0_f (port_out_s0_f[2]), .B1_t (port_out_s1_t[2]), .B1_f (port_out_s1_f[2]), .Z0_t (StateOutXORroundKey[2]), .Z0_f (new_AGEMA_signal_2513), .Z1_t (new_AGEMA_signal_2514), .Z1_f (new_AGEMA_signal_2515) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U28 ( .A0_t (keyStateIn[3]), .A0_f (new_AGEMA_signal_2516), .A1_t (new_AGEMA_signal_2517), .A1_f (new_AGEMA_signal_2518), .B0_t (port_out_s0_t[3]), .B0_f (port_out_s0_f[3]), .B1_t (port_out_s1_t[3]), .B1_f (port_out_s1_f[3]), .Z0_t (StateOutXORroundKey[3]), .Z0_f (new_AGEMA_signal_2522), .Z1_t (new_AGEMA_signal_2523), .Z1_f (new_AGEMA_signal_2524) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U29 ( .A0_t (keyStateIn[4]), .A0_f (new_AGEMA_signal_2525), .A1_t (new_AGEMA_signal_2526), .A1_f (new_AGEMA_signal_2527), .B0_t (port_out_s0_t[4]), .B0_f (port_out_s0_f[4]), .B1_t (port_out_s1_t[4]), .B1_f (port_out_s1_f[4]), .Z0_t (StateOutXORroundKey[4]), .Z0_f (new_AGEMA_signal_2531), .Z1_t (new_AGEMA_signal_2532), .Z1_f (new_AGEMA_signal_2533) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U30 ( .A0_t (keyStateIn[5]), .A0_f (new_AGEMA_signal_2534), .A1_t (new_AGEMA_signal_2535), .A1_f (new_AGEMA_signal_2536), .B0_t (port_out_s0_t[5]), .B0_f (port_out_s0_f[5]), .B1_t (port_out_s1_t[5]), .B1_f (port_out_s1_f[5]), .Z0_t (StateOutXORroundKey[5]), .Z0_f (new_AGEMA_signal_2540), .Z1_t (new_AGEMA_signal_2541), .Z1_f (new_AGEMA_signal_2542) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U31 ( .A0_t (keyStateIn[6]), .A0_f (new_AGEMA_signal_2543), .A1_t (new_AGEMA_signal_2544), .A1_f (new_AGEMA_signal_2545), .B0_t (port_out_s0_t[6]), .B0_f (port_out_s0_f[6]), .B1_t (port_out_s1_t[6]), .B1_f (port_out_s1_f[6]), .Z0_t (StateOutXORroundKey[6]), .Z0_f (new_AGEMA_signal_2549), .Z1_t (new_AGEMA_signal_2550), .Z1_f (new_AGEMA_signal_2551) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U32 ( .A0_t (keyStateIn[7]), .A0_f (new_AGEMA_signal_2552), .A1_t (new_AGEMA_signal_2553), .A1_f (new_AGEMA_signal_2554), .B0_t (port_out_s0_t[7]), .B0_f (port_out_s0_f[7]), .B1_t (port_out_s1_t[7]), .B1_f (port_out_s1_f[7]), .Z0_t (StateOutXORroundKey[7]), .Z0_f (new_AGEMA_signal_2558), .Z1_t (new_AGEMA_signal_2559), .Z1_f (new_AGEMA_signal_2560) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) U33 ( .A0_t (notFirst), .A0_f (new_AGEMA_signal_5133), .B0_t (selXOR), .B0_f (new_AGEMA_signal_4203), .Z0_t (intselXOR), .Z0_f (new_AGEMA_signal_5158) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) ctrl_U25 ( .A0_t (ctrl_n24), .A0_f (new_AGEMA_signal_4695), .B0_t (start_t), .B0_f (start_f), .Z0_t (ctrl_nRstSeq4), .Z0_f (new_AGEMA_signal_5159) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b0)) ctrl_U24 ( .A0_t (ctrl_seq6Out_4_), .A0_f (new_AGEMA_signal_2561), .B0_t (ctrl_seq6In_1_), .B0_f (new_AGEMA_signal_2562), .Z0_t (ctrl_n22), .Z0_f (new_AGEMA_signal_2563) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1), .NL(1'b1)) ctrl_U23 ( .A0_t (ctrl_n4), .A0_f (new_AGEMA_signal_5778), .B0_t (ctrl_n19), .B0_f (new_AGEMA_signal_4694), .Z0_t (ctrl_n5), .Z0_f (new_AGEMA_signal_2571) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) ctrl_U22 ( .A0_t (selXOR), .A0_f (new_AGEMA_signal_4203), .B0_t (ctrl_n5), .B0_f (new_AGEMA_signal_2571), .Z0_t (ctrl_n19), .Z0_f (new_AGEMA_signal_4694) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) ctrl_U21 ( .A0_t (start_t), .A0_f (start_f), .B0_t (ctrl_n18), .B0_f (new_AGEMA_signal_2566), .Z0_t (selXOR), .Z0_f (new_AGEMA_signal_4203) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) ctrl_U20 ( .A0_t (ctrl_seq4Out_1_), .A0_f (new_AGEMA_signal_2564), .B0_t (ctrl_seq4In_1_), .B0_f (new_AGEMA_signal_2565), .Z0_t (ctrl_n18), .Z0_f (new_AGEMA_signal_2566) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b1), .NL(1'b1)) ctrl_U19 ( .A0_t (ctrl_n4), .A0_f (new_AGEMA_signal_5778), .B0_t (ctrl_n17), .B0_f (new_AGEMA_signal_5777), .Z0_t (enRCon), .Z0_f (new_AGEMA_signal_4178) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) ctrl_U18 ( .A0_t (enRCon), .A0_f (new_AGEMA_signal_4178), .B0_t (done_t), .B0_f (done_f), .Z0_t (ctrl_n17), .Z0_f (new_AGEMA_signal_5777) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) ctrl_U17 ( .A0_t (start_t), .A0_f (start_f), .B0_t (ctrl_n24), .B0_f (new_AGEMA_signal_4695), .Z0_t (ctrl_n14), .Z0_f (new_AGEMA_signal_5160) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) ctrl_U16 ( .A0_t (ctrl_seq4Out_1_), .A0_f (new_AGEMA_signal_2564), .B0_t (ctrl_n12), .B0_f (new_AGEMA_signal_5161), .Z0_t (ctrl_finalStep), .Z0_f (new_AGEMA_signal_5307) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) ctrl_U15 ( .A0_t (ctrl_n24), .A0_f (new_AGEMA_signal_4695), .B0_t (ctrl_seq4In_1_), .B0_f (new_AGEMA_signal_2565), .Z0_t (ctrl_n12), .Z0_f (new_AGEMA_signal_5161) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) ctrl_U14 ( .A0_t (ctrl_n10), .A0_f (new_AGEMA_signal_2570), .B0_t (ctrl_n9), .B0_f (new_AGEMA_signal_2568), .Z0_t (ctrl_n11), .Z0_f (new_AGEMA_signal_4204) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) ctrl_U13 ( .A0_t (ctrl_seq6In_3_), .A0_f (new_AGEMA_signal_2567), .B0_t (ctrl_seq6Out_4_), .B0_f (new_AGEMA_signal_2561), .Z0_t (ctrl_n9), .Z0_f (new_AGEMA_signal_2568) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) ctrl_U12 ( .A0_t (ctrl_seq6In_1_), .A0_f (new_AGEMA_signal_2562), .B0_t (ctrl_seq6In_4_), .B0_f (new_AGEMA_signal_2569), .Z0_t (ctrl_n10), .Z0_f (new_AGEMA_signal_2570) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) ctrl_U9 ( .A0_t (ctrl_seq6In_2_), .A0_f (new_AGEMA_signal_2575), .B0_t (ctrl_n11), .B0_f (new_AGEMA_signal_4204), .Z0_t (ctrl_n24), .Z0_f (new_AGEMA_signal_4695) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) ctrl_U8 ( .A0_t (start_t), .A0_f (start_f), .B0_t (ctrl_n13), .B0_f (new_AGEMA_signal_5461), .Z0_t (done_t), .Z0_f (done_f) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) ctrl_U6 ( .A0_t (ctrl_finalStep), .A0_f (new_AGEMA_signal_5307), .B0_t (intFinal), .B0_f (new_AGEMA_signal_4669), .Z0_t (ctrl_n13), .Z0_f (new_AGEMA_signal_5461) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) ctrl_U5 ( .A0_t (done_t), .A0_f (done_f), .B0_t (ctrl_n14), .B0_f (new_AGEMA_signal_5160), .Z0_t (ctrl_n4), .Z0_f (new_AGEMA_signal_5778) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) ctrl_U3 ( .A0_t (ctrl_n5), .A0_f (new_AGEMA_signal_2571), .B0_t (start_t), .B0_f (start_f), .Z0_t (selMC), .Z0_f (new_AGEMA_signal_2573) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1), .NL(1'b1)) ctrl_seq6_SFF_0_U3 ( .A0_t (ctrl_seq6_SFF_0_n2), .A0_f (new_AGEMA_signal_5780), .B0_t (ctrl_seq6_SFF_0_n1), .B0_f (new_AGEMA_signal_5779), .Z0_t (ctrl_seq6In_1_), .Z0_f (new_AGEMA_signal_2562) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) ctrl_seq6_SFF_0_U2 ( .A0_t (done_t), .A0_f (done_f), .B0_t (ctrl_seq6In_1_), .B0_f (new_AGEMA_signal_2562), .Z0_t (ctrl_seq6_SFF_0_n1), .Z0_f (new_AGEMA_signal_5779) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) ctrl_seq6_SFF_0_U1 ( .A0_t (ctrl_seq6_SFF_0_QD), .A0_f (new_AGEMA_signal_5162), .B0_t (done_t), .B0_f (done_f), .Z0_t (ctrl_seq6_SFF_0_n2), .Z0_f (new_AGEMA_signal_5780) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) ctrl_seq6_SFF_0_MUXInst_XOR1_U1 ( .A0_t (1'b1), .A0_f (1'b1), .B0_t (ctrl_n22), .B0_f (new_AGEMA_signal_2563), .Z0_t (ctrl_seq6_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_4205) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) ctrl_seq6_SFF_0_MUXInst_AND1_U1 ( .A0_t (start_t), .A0_f (start_f), .B0_t (ctrl_seq6_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_4205), .Z0_t (ctrl_seq6_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_4696) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) ctrl_seq6_SFF_0_MUXInst_XOR2_U1 ( .A0_t (ctrl_seq6_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_4696), .B0_t (1'b1), .B0_f (1'b1), .Z0_t (ctrl_seq6_SFF_0_QD), .Z0_f (new_AGEMA_signal_5162) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1), .NL(1'b1)) ctrl_seq6_SFF_1_U3 ( .A0_t (ctrl_seq6_SFF_1_n2), .A0_f (new_AGEMA_signal_5782), .B0_t (ctrl_seq6_SFF_1_n1), .B0_f (new_AGEMA_signal_5781), .Z0_t (ctrl_seq6In_2_), .Z0_f (new_AGEMA_signal_2575) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) ctrl_seq6_SFF_1_U2 ( .A0_t (done_t), .A0_f (done_f), .B0_t (ctrl_seq6In_2_), .B0_f (new_AGEMA_signal_2575), .Z0_t (ctrl_seq6_SFF_1_n1), .Z0_f (new_AGEMA_signal_5781) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) ctrl_seq6_SFF_1_U1 ( .A0_t (ctrl_seq6_SFF_1_QD), .A0_f (new_AGEMA_signal_4697), .B0_t (done_t), .B0_f (done_f), .Z0_t (ctrl_seq6_SFF_1_n2), .Z0_f (new_AGEMA_signal_5782) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) ctrl_seq6_SFF_1_MUXInst_XOR1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .B0_t (ctrl_seq6In_1_), .B0_f (new_AGEMA_signal_2562), .Z0_t (ctrl_seq6_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_2574) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) ctrl_seq6_SFF_1_MUXInst_AND1_U1 ( .A0_t (start_t), .A0_f (start_f), .B0_t (ctrl_seq6_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_2574), .Z0_t (ctrl_seq6_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_4206) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) ctrl_seq6_SFF_1_MUXInst_XOR2_U1 ( .A0_t (ctrl_seq6_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_4206), .B0_t (1'b0), .B0_f (1'b1), .Z0_t (ctrl_seq6_SFF_1_QD), .Z0_f (new_AGEMA_signal_4697) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1), .NL(1'b1)) ctrl_seq6_SFF_2_U3 ( .A0_t (ctrl_seq6_SFF_2_n2), .A0_f (new_AGEMA_signal_5784), .B0_t (ctrl_seq6_SFF_2_n1), .B0_f (new_AGEMA_signal_5783), .Z0_t (ctrl_seq6In_3_), .Z0_f (new_AGEMA_signal_2567) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) ctrl_seq6_SFF_2_U2 ( .A0_t (done_t), .A0_f (done_f), .B0_t (ctrl_seq6In_3_), .B0_f (new_AGEMA_signal_2567), .Z0_t (ctrl_seq6_SFF_2_n1), .Z0_f (new_AGEMA_signal_5783) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) ctrl_seq6_SFF_2_U1 ( .A0_t (ctrl_seq6_SFF_2_QD), .A0_f (new_AGEMA_signal_4698), .B0_t (done_t), .B0_f (done_f), .Z0_t (ctrl_seq6_SFF_2_n2), .Z0_f (new_AGEMA_signal_5784) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) ctrl_seq6_SFF_2_MUXInst_XOR1_U1 ( .A0_t (1'b1), .A0_f (1'b1), .B0_t (ctrl_seq6In_2_), .B0_f (new_AGEMA_signal_2575), .Z0_t (ctrl_seq6_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_2576) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) ctrl_seq6_SFF_2_MUXInst_AND1_U1 ( .A0_t (start_t), .A0_f (start_f), .B0_t (ctrl_seq6_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_2576), .Z0_t (ctrl_seq6_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_4207) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) ctrl_seq6_SFF_2_MUXInst_XOR2_U1 ( .A0_t (ctrl_seq6_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_4207), .B0_t (1'b1), .B0_f (1'b1), .Z0_t (ctrl_seq6_SFF_2_QD), .Z0_f (new_AGEMA_signal_4698) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1), .NL(1'b1)) ctrl_seq6_SFF_3_U3 ( .A0_t (ctrl_seq6_SFF_3_n2), .A0_f (new_AGEMA_signal_5786), .B0_t (ctrl_seq6_SFF_3_n1), .B0_f (new_AGEMA_signal_5785), .Z0_t (ctrl_seq6In_4_), .Z0_f (new_AGEMA_signal_2569) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) ctrl_seq6_SFF_3_U2 ( .A0_t (done_t), .A0_f (done_f), .B0_t (ctrl_seq6In_4_), .B0_f (new_AGEMA_signal_2569), .Z0_t (ctrl_seq6_SFF_3_n1), .Z0_f (new_AGEMA_signal_5785) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) ctrl_seq6_SFF_3_U1 ( .A0_t (ctrl_seq6_SFF_3_QD), .A0_f (new_AGEMA_signal_4699), .B0_t (done_t), .B0_f (done_f), .Z0_t (ctrl_seq6_SFF_3_n2), .Z0_f (new_AGEMA_signal_5786) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) ctrl_seq6_SFF_3_MUXInst_XOR1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .B0_t (ctrl_seq6In_3_), .B0_f (new_AGEMA_signal_2567), .Z0_t (ctrl_seq6_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_2577) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) ctrl_seq6_SFF_3_MUXInst_AND1_U1 ( .A0_t (start_t), .A0_f (start_f), .B0_t (ctrl_seq6_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_2577), .Z0_t (ctrl_seq6_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_4208) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) ctrl_seq6_SFF_3_MUXInst_XOR2_U1 ( .A0_t (ctrl_seq6_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_4208), .B0_t (1'b0), .B0_f (1'b1), .Z0_t (ctrl_seq6_SFF_3_QD), .Z0_f (new_AGEMA_signal_4699) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1), .NL(1'b1)) ctrl_seq6_SFF_4_U3 ( .A0_t (ctrl_seq6_SFF_4_n2), .A0_f (new_AGEMA_signal_5788), .B0_t (ctrl_seq6_SFF_4_n1), .B0_f (new_AGEMA_signal_5787), .Z0_t (ctrl_seq6Out_4_), .Z0_f (new_AGEMA_signal_2561) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) ctrl_seq6_SFF_4_U2 ( .A0_t (done_t), .A0_f (done_f), .B0_t (ctrl_seq6Out_4_), .B0_f (new_AGEMA_signal_2561), .Z0_t (ctrl_seq6_SFF_4_n1), .Z0_f (new_AGEMA_signal_5787) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) ctrl_seq6_SFF_4_U1 ( .A0_t (ctrl_seq6_SFF_4_QD), .A0_f (new_AGEMA_signal_4700), .B0_t (done_t), .B0_f (done_f), .Z0_t (ctrl_seq6_SFF_4_n2), .Z0_f (new_AGEMA_signal_5788) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) ctrl_seq6_SFF_4_MUXInst_XOR1_U1 ( .A0_t (1'b1), .A0_f (1'b1), .B0_t (ctrl_seq6In_4_), .B0_f (new_AGEMA_signal_2569), .Z0_t (ctrl_seq6_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_2578) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) ctrl_seq6_SFF_4_MUXInst_AND1_U1 ( .A0_t (start_t), .A0_f (start_f), .B0_t (ctrl_seq6_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_2578), .Z0_t (ctrl_seq6_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_4209) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) ctrl_seq6_SFF_4_MUXInst_XOR2_U1 ( .A0_t (ctrl_seq6_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_4209), .B0_t (1'b1), .B0_f (1'b1), .Z0_t (ctrl_seq6_SFF_4_QD), .Z0_f (new_AGEMA_signal_4700) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1), .NL(1'b1)) ctrl_seq4_SFF_0_U3 ( .A0_t (ctrl_seq4_SFF_0_n2), .A0_f (new_AGEMA_signal_5790), .B0_t (ctrl_seq4_SFF_0_n1), .B0_f (new_AGEMA_signal_5789), .Z0_t (ctrl_seq4In_1_), .Z0_f (new_AGEMA_signal_2565) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) ctrl_seq4_SFF_0_U2 ( .A0_t (done_t), .A0_f (done_f), .B0_t (ctrl_seq4In_1_), .B0_f (new_AGEMA_signal_2565), .Z0_t (ctrl_seq4_SFF_0_n1), .Z0_f (new_AGEMA_signal_5789) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) ctrl_seq4_SFF_0_U1 ( .A0_t (ctrl_seq4_SFF_0_QD), .A0_f (new_AGEMA_signal_5462), .B0_t (done_t), .B0_f (done_f), .Z0_t (ctrl_seq4_SFF_0_n2), .Z0_f (new_AGEMA_signal_5790) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) ctrl_seq4_SFF_0_MUXInst_XOR1_U1 ( .A0_t (1'b1), .A0_f (1'b1), .B0_t (ctrl_seq4Out_1_), .B0_f (new_AGEMA_signal_2564), .Z0_t (ctrl_seq4_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_2579) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) ctrl_seq4_SFF_0_MUXInst_AND1_U1 ( .A0_t (ctrl_nRstSeq4), .A0_f (new_AGEMA_signal_5159), .B0_t (ctrl_seq4_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_2579), .Z0_t (ctrl_seq4_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_5308) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) ctrl_seq4_SFF_0_MUXInst_XOR2_U1 ( .A0_t (ctrl_seq4_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_5308), .B0_t (1'b1), .B0_f (1'b1), .Z0_t (ctrl_seq4_SFF_0_QD), .Z0_f (new_AGEMA_signal_5462) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1), .NL(1'b1)) ctrl_seq4_SFF_1_U3 ( .A0_t (ctrl_seq4_SFF_1_n2), .A0_f (new_AGEMA_signal_5792), .B0_t (ctrl_seq4_SFF_1_n1), .B0_f (new_AGEMA_signal_5791), .Z0_t (ctrl_seq4Out_1_), .Z0_f (new_AGEMA_signal_2564) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) ctrl_seq4_SFF_1_U2 ( .A0_t (done_t), .A0_f (done_f), .B0_t (ctrl_seq4Out_1_), .B0_f (new_AGEMA_signal_2564), .Z0_t (ctrl_seq4_SFF_1_n1), .Z0_f (new_AGEMA_signal_5791) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) ctrl_seq4_SFF_1_U1 ( .A0_t (ctrl_seq4_SFF_1_QD), .A0_f (new_AGEMA_signal_5463), .B0_t (done_t), .B0_f (done_f), .Z0_t (ctrl_seq4_SFF_1_n2), .Z0_f (new_AGEMA_signal_5792) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) ctrl_seq4_SFF_1_MUXInst_XOR1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .B0_t (ctrl_seq4In_1_), .B0_f (new_AGEMA_signal_2565), .Z0_t (ctrl_seq4_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_2580) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) ctrl_seq4_SFF_1_MUXInst_AND1_U1 ( .A0_t (ctrl_nRstSeq4), .A0_f (new_AGEMA_signal_5159), .B0_t (ctrl_seq4_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_2580), .Z0_t (ctrl_seq4_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_5309) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) ctrl_seq4_SFF_1_MUXInst_XOR2_U1 ( .A0_t (ctrl_seq4_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_5309), .B0_t (1'b0), .B0_f (1'b1), .Z0_t (ctrl_seq4_SFF_1_QD), .Z0_f (new_AGEMA_signal_5463) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_0_XOR1_U1 ( .A0_t (SboxOut[0]), .A0_f (new_AGEMA_signal_7502), .A1_t (new_AGEMA_signal_7503), .A1_f (new_AGEMA_signal_7504), .B0_t (StateOutXORroundKey[0]), .B0_f (new_AGEMA_signal_2495), .B1_t (new_AGEMA_signal_2496), .B1_f (new_AGEMA_signal_2497), .Z0_t (MUX_StateIn_mux_inst_0_X), .Z0_f (new_AGEMA_signal_7505), .Z1_t (new_AGEMA_signal_7506), .Z1_f (new_AGEMA_signal_7507) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_0_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_4669), .B0_t (MUX_StateIn_mux_inst_0_X), .B0_f (new_AGEMA_signal_7505), .B1_t (new_AGEMA_signal_7506), .B1_f (new_AGEMA_signal_7507), .Z0_t (MUX_StateIn_mux_inst_0_Y), .Z0_f (new_AGEMA_signal_7532), .Z1_t (new_AGEMA_signal_7533), .Z1_f (new_AGEMA_signal_7534) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_0_XOR2_U1 ( .A0_t (MUX_StateIn_mux_inst_0_Y), .A0_f (new_AGEMA_signal_7532), .A1_t (new_AGEMA_signal_7533), .A1_f (new_AGEMA_signal_7534), .B0_t (SboxOut[0]), .B0_f (new_AGEMA_signal_7502), .B1_t (new_AGEMA_signal_7503), .B1_f (new_AGEMA_signal_7504), .Z0_t (StateIn[0]), .Z0_f (new_AGEMA_signal_7580), .Z1_t (new_AGEMA_signal_7581), .Z1_f (new_AGEMA_signal_7582) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_1_XOR1_U1 ( .A0_t (SboxOut[1]), .A0_f (new_AGEMA_signal_7529), .A1_t (new_AGEMA_signal_7530), .A1_f (new_AGEMA_signal_7531), .B0_t (StateOutXORroundKey[1]), .B0_f (new_AGEMA_signal_2504), .B1_t (new_AGEMA_signal_2505), .B1_f (new_AGEMA_signal_2506), .Z0_t (MUX_StateIn_mux_inst_1_X), .Z0_f (new_AGEMA_signal_7535), .Z1_t (new_AGEMA_signal_7536), .Z1_f (new_AGEMA_signal_7537) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_4669), .B0_t (MUX_StateIn_mux_inst_1_X), .B0_f (new_AGEMA_signal_7535), .B1_t (new_AGEMA_signal_7536), .B1_f (new_AGEMA_signal_7537), .Z0_t (MUX_StateIn_mux_inst_1_Y), .Z0_f (new_AGEMA_signal_7583), .Z1_t (new_AGEMA_signal_7584), .Z1_f (new_AGEMA_signal_7585) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_1_XOR2_U1 ( .A0_t (MUX_StateIn_mux_inst_1_Y), .A0_f (new_AGEMA_signal_7583), .A1_t (new_AGEMA_signal_7584), .A1_f (new_AGEMA_signal_7585), .B0_t (SboxOut[1]), .B0_f (new_AGEMA_signal_7529), .B1_t (new_AGEMA_signal_7530), .B1_f (new_AGEMA_signal_7531), .Z0_t (StateIn[1]), .Z0_f (new_AGEMA_signal_7628), .Z1_t (new_AGEMA_signal_7629), .Z1_f (new_AGEMA_signal_7630) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_2_XOR1_U1 ( .A0_t (SboxOut[2]), .A0_f (new_AGEMA_signal_7526), .A1_t (new_AGEMA_signal_7527), .A1_f (new_AGEMA_signal_7528), .B0_t (StateOutXORroundKey[2]), .B0_f (new_AGEMA_signal_2513), .B1_t (new_AGEMA_signal_2514), .B1_f (new_AGEMA_signal_2515), .Z0_t (MUX_StateIn_mux_inst_2_X), .Z0_f (new_AGEMA_signal_7538), .Z1_t (new_AGEMA_signal_7539), .Z1_f (new_AGEMA_signal_7540) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_2_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_4669), .B0_t (MUX_StateIn_mux_inst_2_X), .B0_f (new_AGEMA_signal_7538), .B1_t (new_AGEMA_signal_7539), .B1_f (new_AGEMA_signal_7540), .Z0_t (MUX_StateIn_mux_inst_2_Y), .Z0_f (new_AGEMA_signal_7586), .Z1_t (new_AGEMA_signal_7587), .Z1_f (new_AGEMA_signal_7588) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_2_XOR2_U1 ( .A0_t (MUX_StateIn_mux_inst_2_Y), .A0_f (new_AGEMA_signal_7586), .A1_t (new_AGEMA_signal_7587), .A1_f (new_AGEMA_signal_7588), .B0_t (SboxOut[2]), .B0_f (new_AGEMA_signal_7526), .B1_t (new_AGEMA_signal_7527), .B1_f (new_AGEMA_signal_7528), .Z0_t (StateIn[2]), .Z0_f (new_AGEMA_signal_7631), .Z1_t (new_AGEMA_signal_7632), .Z1_f (new_AGEMA_signal_7633) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_3_XOR1_U1 ( .A0_t (SboxOut[3]), .A0_f (new_AGEMA_signal_7523), .A1_t (new_AGEMA_signal_7524), .A1_f (new_AGEMA_signal_7525), .B0_t (StateOutXORroundKey[3]), .B0_f (new_AGEMA_signal_2522), .B1_t (new_AGEMA_signal_2523), .B1_f (new_AGEMA_signal_2524), .Z0_t (MUX_StateIn_mux_inst_3_X), .Z0_f (new_AGEMA_signal_7541), .Z1_t (new_AGEMA_signal_7542), .Z1_f (new_AGEMA_signal_7543) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_3_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_4669), .B0_t (MUX_StateIn_mux_inst_3_X), .B0_f (new_AGEMA_signal_7541), .B1_t (new_AGEMA_signal_7542), .B1_f (new_AGEMA_signal_7543), .Z0_t (MUX_StateIn_mux_inst_3_Y), .Z0_f (new_AGEMA_signal_7589), .Z1_t (new_AGEMA_signal_7590), .Z1_f (new_AGEMA_signal_7591) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_3_XOR2_U1 ( .A0_t (MUX_StateIn_mux_inst_3_Y), .A0_f (new_AGEMA_signal_7589), .A1_t (new_AGEMA_signal_7590), .A1_f (new_AGEMA_signal_7591), .B0_t (SboxOut[3]), .B0_f (new_AGEMA_signal_7523), .B1_t (new_AGEMA_signal_7524), .B1_f (new_AGEMA_signal_7525), .Z0_t (StateIn[3]), .Z0_f (new_AGEMA_signal_7634), .Z1_t (new_AGEMA_signal_7635), .Z1_f (new_AGEMA_signal_7636) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_4_XOR1_U1 ( .A0_t (SboxOut[4]), .A0_f (new_AGEMA_signal_7520), .A1_t (new_AGEMA_signal_7521), .A1_f (new_AGEMA_signal_7522), .B0_t (StateOutXORroundKey[4]), .B0_f (new_AGEMA_signal_2531), .B1_t (new_AGEMA_signal_2532), .B1_f (new_AGEMA_signal_2533), .Z0_t (MUX_StateIn_mux_inst_4_X), .Z0_f (new_AGEMA_signal_7544), .Z1_t (new_AGEMA_signal_7545), .Z1_f (new_AGEMA_signal_7546) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_4_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_4669), .B0_t (MUX_StateIn_mux_inst_4_X), .B0_f (new_AGEMA_signal_7544), .B1_t (new_AGEMA_signal_7545), .B1_f (new_AGEMA_signal_7546), .Z0_t (MUX_StateIn_mux_inst_4_Y), .Z0_f (new_AGEMA_signal_7592), .Z1_t (new_AGEMA_signal_7593), .Z1_f (new_AGEMA_signal_7594) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_4_XOR2_U1 ( .A0_t (MUX_StateIn_mux_inst_4_Y), .A0_f (new_AGEMA_signal_7592), .A1_t (new_AGEMA_signal_7593), .A1_f (new_AGEMA_signal_7594), .B0_t (SboxOut[4]), .B0_f (new_AGEMA_signal_7520), .B1_t (new_AGEMA_signal_7521), .B1_f (new_AGEMA_signal_7522), .Z0_t (StateIn[4]), .Z0_f (new_AGEMA_signal_7637), .Z1_t (new_AGEMA_signal_7638), .Z1_f (new_AGEMA_signal_7639) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_5_XOR1_U1 ( .A0_t (SboxOut[5]), .A0_f (new_AGEMA_signal_7517), .A1_t (new_AGEMA_signal_7518), .A1_f (new_AGEMA_signal_7519), .B0_t (StateOutXORroundKey[5]), .B0_f (new_AGEMA_signal_2540), .B1_t (new_AGEMA_signal_2541), .B1_f (new_AGEMA_signal_2542), .Z0_t (MUX_StateIn_mux_inst_5_X), .Z0_f (new_AGEMA_signal_7547), .Z1_t (new_AGEMA_signal_7548), .Z1_f (new_AGEMA_signal_7549) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_5_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_4669), .B0_t (MUX_StateIn_mux_inst_5_X), .B0_f (new_AGEMA_signal_7547), .B1_t (new_AGEMA_signal_7548), .B1_f (new_AGEMA_signal_7549), .Z0_t (MUX_StateIn_mux_inst_5_Y), .Z0_f (new_AGEMA_signal_7595), .Z1_t (new_AGEMA_signal_7596), .Z1_f (new_AGEMA_signal_7597) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_5_XOR2_U1 ( .A0_t (MUX_StateIn_mux_inst_5_Y), .A0_f (new_AGEMA_signal_7595), .A1_t (new_AGEMA_signal_7596), .A1_f (new_AGEMA_signal_7597), .B0_t (SboxOut[5]), .B0_f (new_AGEMA_signal_7517), .B1_t (new_AGEMA_signal_7518), .B1_f (new_AGEMA_signal_7519), .Z0_t (StateIn[5]), .Z0_f (new_AGEMA_signal_7640), .Z1_t (new_AGEMA_signal_7641), .Z1_f (new_AGEMA_signal_7642) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_6_XOR1_U1 ( .A0_t (SboxOut[6]), .A0_f (new_AGEMA_signal_7514), .A1_t (new_AGEMA_signal_7515), .A1_f (new_AGEMA_signal_7516), .B0_t (StateOutXORroundKey[6]), .B0_f (new_AGEMA_signal_2549), .B1_t (new_AGEMA_signal_2550), .B1_f (new_AGEMA_signal_2551), .Z0_t (MUX_StateIn_mux_inst_6_X), .Z0_f (new_AGEMA_signal_7550), .Z1_t (new_AGEMA_signal_7551), .Z1_f (new_AGEMA_signal_7552) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_6_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_4669), .B0_t (MUX_StateIn_mux_inst_6_X), .B0_f (new_AGEMA_signal_7550), .B1_t (new_AGEMA_signal_7551), .B1_f (new_AGEMA_signal_7552), .Z0_t (MUX_StateIn_mux_inst_6_Y), .Z0_f (new_AGEMA_signal_7598), .Z1_t (new_AGEMA_signal_7599), .Z1_f (new_AGEMA_signal_7600) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_6_XOR2_U1 ( .A0_t (MUX_StateIn_mux_inst_6_Y), .A0_f (new_AGEMA_signal_7598), .A1_t (new_AGEMA_signal_7599), .A1_f (new_AGEMA_signal_7600), .B0_t (SboxOut[6]), .B0_f (new_AGEMA_signal_7514), .B1_t (new_AGEMA_signal_7515), .B1_f (new_AGEMA_signal_7516), .Z0_t (StateIn[6]), .Z0_f (new_AGEMA_signal_7643), .Z1_t (new_AGEMA_signal_7644), .Z1_f (new_AGEMA_signal_7645) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_7_XOR1_U1 ( .A0_t (SboxOut[7]), .A0_f (new_AGEMA_signal_7511), .A1_t (new_AGEMA_signal_7512), .A1_f (new_AGEMA_signal_7513), .B0_t (StateOutXORroundKey[7]), .B0_f (new_AGEMA_signal_2558), .B1_t (new_AGEMA_signal_2559), .B1_f (new_AGEMA_signal_2560), .Z0_t (MUX_StateIn_mux_inst_7_X), .Z0_f (new_AGEMA_signal_7553), .Z1_t (new_AGEMA_signal_7554), .Z1_f (new_AGEMA_signal_7555) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_7_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_4669), .B0_t (MUX_StateIn_mux_inst_7_X), .B0_f (new_AGEMA_signal_7553), .B1_t (new_AGEMA_signal_7554), .B1_f (new_AGEMA_signal_7555), .Z0_t (MUX_StateIn_mux_inst_7_Y), .Z0_f (new_AGEMA_signal_7601), .Z1_t (new_AGEMA_signal_7602), .Z1_f (new_AGEMA_signal_7603) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateIn_mux_inst_7_XOR2_U1 ( .A0_t (MUX_StateIn_mux_inst_7_Y), .A0_f (new_AGEMA_signal_7601), .A1_t (new_AGEMA_signal_7602), .A1_f (new_AGEMA_signal_7603), .B0_t (SboxOut[7]), .B0_f (new_AGEMA_signal_7511), .B1_t (new_AGEMA_signal_7512), .B1_f (new_AGEMA_signal_7513), .Z0_t (StateIn[7]), .Z0_f (new_AGEMA_signal_7646), .Z1_t (new_AGEMA_signal_7647), .Z1_f (new_AGEMA_signal_7648) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) stateArray_U3 ( .A0_t (start_t), .A0_f (start_f), .B0_t (selMC), .B0_f (new_AGEMA_signal_2573), .Z0_t (stateArray_nReset_selMC), .Z0_f (new_AGEMA_signal_4210) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S00reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS01ser[0]), .A0_f (new_AGEMA_signal_2581), .A1_t (new_AGEMA_signal_2582), .A1_f (new_AGEMA_signal_2583), .B0_t (port_out_s0_t[0]), .B0_f (port_out_s0_f[0]), .B1_t (port_out_s1_t[0]), .B1_f (port_out_s1_f[0]), .Z0_t (stateArray_S00reg_gff_1_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_2584), .Z1_t (new_AGEMA_signal_2585), .Z1_f (new_AGEMA_signal_2586) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S00reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S00reg_gff_1_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_2584), .B1_t (new_AGEMA_signal_2585), .B1_f (new_AGEMA_signal_2586), .Z0_t (stateArray_S00reg_gff_1_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_5917), .Z1_t (new_AGEMA_signal_5918), .Z1_f (new_AGEMA_signal_5919) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S00reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (stateArray_S00reg_gff_1_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_5917), .A1_t (new_AGEMA_signal_5918), .A1_f (new_AGEMA_signal_5919), .B0_t (stateArray_outS01ser[0]), .B0_f (new_AGEMA_signal_2581), .B1_t (new_AGEMA_signal_2582), .B1_f (new_AGEMA_signal_2583), .Z0_t (port_out_s0_t[0]), .Z0_f (port_out_s0_f[0]), .Z1_t (port_out_s1_t[0]), .Z1_f (port_out_s1_f[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S00reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS01ser[1]), .A0_f (new_AGEMA_signal_2587), .A1_t (new_AGEMA_signal_2588), .A1_f (new_AGEMA_signal_2589), .B0_t (port_out_s0_t[1]), .B0_f (port_out_s0_f[1]), .B1_t (port_out_s1_t[1]), .B1_f (port_out_s1_f[1]), .Z0_t (stateArray_S00reg_gff_1_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_2590), .Z1_t (new_AGEMA_signal_2591), .Z1_f (new_AGEMA_signal_2592) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S00reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S00reg_gff_1_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_2590), .B1_t (new_AGEMA_signal_2591), .B1_f (new_AGEMA_signal_2592), .Z0_t (stateArray_S00reg_gff_1_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_5920), .Z1_t (new_AGEMA_signal_5921), .Z1_f (new_AGEMA_signal_5922) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S00reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (stateArray_S00reg_gff_1_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_5920), .A1_t (new_AGEMA_signal_5921), .A1_f (new_AGEMA_signal_5922), .B0_t (stateArray_outS01ser[1]), .B0_f (new_AGEMA_signal_2587), .B1_t (new_AGEMA_signal_2588), .B1_f (new_AGEMA_signal_2589), .Z0_t (port_out_s0_t[1]), .Z0_f (port_out_s0_f[1]), .Z1_t (port_out_s1_t[1]), .Z1_f (port_out_s1_f[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S00reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS01ser[2]), .A0_f (new_AGEMA_signal_2593), .A1_t (new_AGEMA_signal_2594), .A1_f (new_AGEMA_signal_2595), .B0_t (port_out_s0_t[2]), .B0_f (port_out_s0_f[2]), .B1_t (port_out_s1_t[2]), .B1_f (port_out_s1_f[2]), .Z0_t (stateArray_S00reg_gff_1_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_2596), .Z1_t (new_AGEMA_signal_2597), .Z1_f (new_AGEMA_signal_2598) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S00reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S00reg_gff_1_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_2596), .B1_t (new_AGEMA_signal_2597), .B1_f (new_AGEMA_signal_2598), .Z0_t (stateArray_S00reg_gff_1_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_5923), .Z1_t (new_AGEMA_signal_5924), .Z1_f (new_AGEMA_signal_5925) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S00reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (stateArray_S00reg_gff_1_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_5923), .A1_t (new_AGEMA_signal_5924), .A1_f (new_AGEMA_signal_5925), .B0_t (stateArray_outS01ser[2]), .B0_f (new_AGEMA_signal_2593), .B1_t (new_AGEMA_signal_2594), .B1_f (new_AGEMA_signal_2595), .Z0_t (port_out_s0_t[2]), .Z0_f (port_out_s0_f[2]), .Z1_t (port_out_s1_t[2]), .Z1_f (port_out_s1_f[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S00reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS01ser[3]), .A0_f (new_AGEMA_signal_2599), .A1_t (new_AGEMA_signal_2600), .A1_f (new_AGEMA_signal_2601), .B0_t (port_out_s0_t[3]), .B0_f (port_out_s0_f[3]), .B1_t (port_out_s1_t[3]), .B1_f (port_out_s1_f[3]), .Z0_t (stateArray_S00reg_gff_1_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_2602), .Z1_t (new_AGEMA_signal_2603), .Z1_f (new_AGEMA_signal_2604) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S00reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S00reg_gff_1_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_2602), .B1_t (new_AGEMA_signal_2603), .B1_f (new_AGEMA_signal_2604), .Z0_t (stateArray_S00reg_gff_1_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_5926), .Z1_t (new_AGEMA_signal_5927), .Z1_f (new_AGEMA_signal_5928) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S00reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (stateArray_S00reg_gff_1_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_5926), .A1_t (new_AGEMA_signal_5927), .A1_f (new_AGEMA_signal_5928), .B0_t (stateArray_outS01ser[3]), .B0_f (new_AGEMA_signal_2599), .B1_t (new_AGEMA_signal_2600), .B1_f (new_AGEMA_signal_2601), .Z0_t (port_out_s0_t[3]), .Z0_f (port_out_s0_f[3]), .Z1_t (port_out_s1_t[3]), .Z1_f (port_out_s1_f[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S00reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS01ser[4]), .A0_f (new_AGEMA_signal_2605), .A1_t (new_AGEMA_signal_2606), .A1_f (new_AGEMA_signal_2607), .B0_t (port_out_s0_t[4]), .B0_f (port_out_s0_f[4]), .B1_t (port_out_s1_t[4]), .B1_f (port_out_s1_f[4]), .Z0_t (stateArray_S00reg_gff_1_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_2608), .Z1_t (new_AGEMA_signal_2609), .Z1_f (new_AGEMA_signal_2610) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S00reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S00reg_gff_1_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_2608), .B1_t (new_AGEMA_signal_2609), .B1_f (new_AGEMA_signal_2610), .Z0_t (stateArray_S00reg_gff_1_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_5929), .Z1_t (new_AGEMA_signal_5930), .Z1_f (new_AGEMA_signal_5931) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S00reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (stateArray_S00reg_gff_1_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_5929), .A1_t (new_AGEMA_signal_5930), .A1_f (new_AGEMA_signal_5931), .B0_t (stateArray_outS01ser[4]), .B0_f (new_AGEMA_signal_2605), .B1_t (new_AGEMA_signal_2606), .B1_f (new_AGEMA_signal_2607), .Z0_t (port_out_s0_t[4]), .Z0_f (port_out_s0_f[4]), .Z1_t (port_out_s1_t[4]), .Z1_f (port_out_s1_f[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S00reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS01ser[5]), .A0_f (new_AGEMA_signal_2611), .A1_t (new_AGEMA_signal_2612), .A1_f (new_AGEMA_signal_2613), .B0_t (port_out_s0_t[5]), .B0_f (port_out_s0_f[5]), .B1_t (port_out_s1_t[5]), .B1_f (port_out_s1_f[5]), .Z0_t (stateArray_S00reg_gff_1_SFF_5_MUXInst_X), .Z0_f (new_AGEMA_signal_2614), .Z1_t (new_AGEMA_signal_2615), .Z1_f (new_AGEMA_signal_2616) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S00reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S00reg_gff_1_SFF_5_MUXInst_X), .B0_f (new_AGEMA_signal_2614), .B1_t (new_AGEMA_signal_2615), .B1_f (new_AGEMA_signal_2616), .Z0_t (stateArray_S00reg_gff_1_SFF_5_MUXInst_Y), .Z0_f (new_AGEMA_signal_5932), .Z1_t (new_AGEMA_signal_5933), .Z1_f (new_AGEMA_signal_5934) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S00reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (stateArray_S00reg_gff_1_SFF_5_MUXInst_Y), .A0_f (new_AGEMA_signal_5932), .A1_t (new_AGEMA_signal_5933), .A1_f (new_AGEMA_signal_5934), .B0_t (stateArray_outS01ser[5]), .B0_f (new_AGEMA_signal_2611), .B1_t (new_AGEMA_signal_2612), .B1_f (new_AGEMA_signal_2613), .Z0_t (port_out_s0_t[5]), .Z0_f (port_out_s0_f[5]), .Z1_t (port_out_s1_t[5]), .Z1_f (port_out_s1_f[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S00reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS01ser[6]), .A0_f (new_AGEMA_signal_2617), .A1_t (new_AGEMA_signal_2618), .A1_f (new_AGEMA_signal_2619), .B0_t (port_out_s0_t[6]), .B0_f (port_out_s0_f[6]), .B1_t (port_out_s1_t[6]), .B1_f (port_out_s1_f[6]), .Z0_t (stateArray_S00reg_gff_1_SFF_6_MUXInst_X), .Z0_f (new_AGEMA_signal_2620), .Z1_t (new_AGEMA_signal_2621), .Z1_f (new_AGEMA_signal_2622) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S00reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S00reg_gff_1_SFF_6_MUXInst_X), .B0_f (new_AGEMA_signal_2620), .B1_t (new_AGEMA_signal_2621), .B1_f (new_AGEMA_signal_2622), .Z0_t (stateArray_S00reg_gff_1_SFF_6_MUXInst_Y), .Z0_f (new_AGEMA_signal_5935), .Z1_t (new_AGEMA_signal_5936), .Z1_f (new_AGEMA_signal_5937) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S00reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (stateArray_S00reg_gff_1_SFF_6_MUXInst_Y), .A0_f (new_AGEMA_signal_5935), .A1_t (new_AGEMA_signal_5936), .A1_f (new_AGEMA_signal_5937), .B0_t (stateArray_outS01ser[6]), .B0_f (new_AGEMA_signal_2617), .B1_t (new_AGEMA_signal_2618), .B1_f (new_AGEMA_signal_2619), .Z0_t (port_out_s0_t[6]), .Z0_f (port_out_s0_f[6]), .Z1_t (port_out_s1_t[6]), .Z1_f (port_out_s1_f[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S00reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS01ser[7]), .A0_f (new_AGEMA_signal_2623), .A1_t (new_AGEMA_signal_2624), .A1_f (new_AGEMA_signal_2625), .B0_t (port_out_s0_t[7]), .B0_f (port_out_s0_f[7]), .B1_t (port_out_s1_t[7]), .B1_f (port_out_s1_f[7]), .Z0_t (stateArray_S00reg_gff_1_SFF_7_MUXInst_X), .Z0_f (new_AGEMA_signal_2626), .Z1_t (new_AGEMA_signal_2627), .Z1_f (new_AGEMA_signal_2628) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S00reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S00reg_gff_1_SFF_7_MUXInst_X), .B0_f (new_AGEMA_signal_2626), .B1_t (new_AGEMA_signal_2627), .B1_f (new_AGEMA_signal_2628), .Z0_t (stateArray_S00reg_gff_1_SFF_7_MUXInst_Y), .Z0_f (new_AGEMA_signal_5938), .Z1_t (new_AGEMA_signal_5939), .Z1_f (new_AGEMA_signal_5940) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S00reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (stateArray_S00reg_gff_1_SFF_7_MUXInst_Y), .A0_f (new_AGEMA_signal_5938), .A1_t (new_AGEMA_signal_5939), .A1_f (new_AGEMA_signal_5940), .B0_t (stateArray_outS01ser[7]), .B0_f (new_AGEMA_signal_2623), .B1_t (new_AGEMA_signal_2624), .B1_f (new_AGEMA_signal_2625), .Z0_t (port_out_s0_t[7]), .Z0_f (port_out_s0_f[7]), .Z1_t (port_out_s1_t[7]), .Z1_f (port_out_s1_f[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S01reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS02ser[0]), .A0_f (new_AGEMA_signal_2629), .A1_t (new_AGEMA_signal_2630), .A1_f (new_AGEMA_signal_2631), .B0_t (stateArray_outS01ser[0]), .B0_f (new_AGEMA_signal_2581), .B1_t (new_AGEMA_signal_2582), .B1_f (new_AGEMA_signal_2583), .Z0_t (stateArray_S01reg_gff_1_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_2632), .Z1_t (new_AGEMA_signal_2633), .Z1_f (new_AGEMA_signal_2634) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S01reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S01reg_gff_1_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_2632), .B1_t (new_AGEMA_signal_2633), .B1_f (new_AGEMA_signal_2634), .Z0_t (stateArray_S01reg_gff_1_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_5941), .Z1_t (new_AGEMA_signal_5942), .Z1_f (new_AGEMA_signal_5943) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S01reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (stateArray_S01reg_gff_1_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_5941), .A1_t (new_AGEMA_signal_5942), .A1_f (new_AGEMA_signal_5943), .B0_t (stateArray_outS02ser[0]), .B0_f (new_AGEMA_signal_2629), .B1_t (new_AGEMA_signal_2630), .B1_f (new_AGEMA_signal_2631), .Z0_t (stateArray_outS01ser[0]), .Z0_f (new_AGEMA_signal_2581), .Z1_t (new_AGEMA_signal_2582), .Z1_f (new_AGEMA_signal_2583) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S01reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS02ser[1]), .A0_f (new_AGEMA_signal_2635), .A1_t (new_AGEMA_signal_2636), .A1_f (new_AGEMA_signal_2637), .B0_t (stateArray_outS01ser[1]), .B0_f (new_AGEMA_signal_2587), .B1_t (new_AGEMA_signal_2588), .B1_f (new_AGEMA_signal_2589), .Z0_t (stateArray_S01reg_gff_1_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_2638), .Z1_t (new_AGEMA_signal_2639), .Z1_f (new_AGEMA_signal_2640) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S01reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S01reg_gff_1_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_2638), .B1_t (new_AGEMA_signal_2639), .B1_f (new_AGEMA_signal_2640), .Z0_t (stateArray_S01reg_gff_1_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_5944), .Z1_t (new_AGEMA_signal_5945), .Z1_f (new_AGEMA_signal_5946) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S01reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (stateArray_S01reg_gff_1_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_5944), .A1_t (new_AGEMA_signal_5945), .A1_f (new_AGEMA_signal_5946), .B0_t (stateArray_outS02ser[1]), .B0_f (new_AGEMA_signal_2635), .B1_t (new_AGEMA_signal_2636), .B1_f (new_AGEMA_signal_2637), .Z0_t (stateArray_outS01ser[1]), .Z0_f (new_AGEMA_signal_2587), .Z1_t (new_AGEMA_signal_2588), .Z1_f (new_AGEMA_signal_2589) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S01reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS02ser[2]), .A0_f (new_AGEMA_signal_2641), .A1_t (new_AGEMA_signal_2642), .A1_f (new_AGEMA_signal_2643), .B0_t (stateArray_outS01ser[2]), .B0_f (new_AGEMA_signal_2593), .B1_t (new_AGEMA_signal_2594), .B1_f (new_AGEMA_signal_2595), .Z0_t (stateArray_S01reg_gff_1_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_2644), .Z1_t (new_AGEMA_signal_2645), .Z1_f (new_AGEMA_signal_2646) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S01reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S01reg_gff_1_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_2644), .B1_t (new_AGEMA_signal_2645), .B1_f (new_AGEMA_signal_2646), .Z0_t (stateArray_S01reg_gff_1_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_5947), .Z1_t (new_AGEMA_signal_5948), .Z1_f (new_AGEMA_signal_5949) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S01reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (stateArray_S01reg_gff_1_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_5947), .A1_t (new_AGEMA_signal_5948), .A1_f (new_AGEMA_signal_5949), .B0_t (stateArray_outS02ser[2]), .B0_f (new_AGEMA_signal_2641), .B1_t (new_AGEMA_signal_2642), .B1_f (new_AGEMA_signal_2643), .Z0_t (stateArray_outS01ser[2]), .Z0_f (new_AGEMA_signal_2593), .Z1_t (new_AGEMA_signal_2594), .Z1_f (new_AGEMA_signal_2595) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S01reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS02ser[3]), .A0_f (new_AGEMA_signal_2647), .A1_t (new_AGEMA_signal_2648), .A1_f (new_AGEMA_signal_2649), .B0_t (stateArray_outS01ser[3]), .B0_f (new_AGEMA_signal_2599), .B1_t (new_AGEMA_signal_2600), .B1_f (new_AGEMA_signal_2601), .Z0_t (stateArray_S01reg_gff_1_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_2650), .Z1_t (new_AGEMA_signal_2651), .Z1_f (new_AGEMA_signal_2652) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S01reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S01reg_gff_1_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_2650), .B1_t (new_AGEMA_signal_2651), .B1_f (new_AGEMA_signal_2652), .Z0_t (stateArray_S01reg_gff_1_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_5950), .Z1_t (new_AGEMA_signal_5951), .Z1_f (new_AGEMA_signal_5952) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S01reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (stateArray_S01reg_gff_1_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_5950), .A1_t (new_AGEMA_signal_5951), .A1_f (new_AGEMA_signal_5952), .B0_t (stateArray_outS02ser[3]), .B0_f (new_AGEMA_signal_2647), .B1_t (new_AGEMA_signal_2648), .B1_f (new_AGEMA_signal_2649), .Z0_t (stateArray_outS01ser[3]), .Z0_f (new_AGEMA_signal_2599), .Z1_t (new_AGEMA_signal_2600), .Z1_f (new_AGEMA_signal_2601) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S01reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS02ser[4]), .A0_f (new_AGEMA_signal_2653), .A1_t (new_AGEMA_signal_2654), .A1_f (new_AGEMA_signal_2655), .B0_t (stateArray_outS01ser[4]), .B0_f (new_AGEMA_signal_2605), .B1_t (new_AGEMA_signal_2606), .B1_f (new_AGEMA_signal_2607), .Z0_t (stateArray_S01reg_gff_1_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_2656), .Z1_t (new_AGEMA_signal_2657), .Z1_f (new_AGEMA_signal_2658) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S01reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S01reg_gff_1_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_2656), .B1_t (new_AGEMA_signal_2657), .B1_f (new_AGEMA_signal_2658), .Z0_t (stateArray_S01reg_gff_1_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_5953), .Z1_t (new_AGEMA_signal_5954), .Z1_f (new_AGEMA_signal_5955) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S01reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (stateArray_S01reg_gff_1_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_5953), .A1_t (new_AGEMA_signal_5954), .A1_f (new_AGEMA_signal_5955), .B0_t (stateArray_outS02ser[4]), .B0_f (new_AGEMA_signal_2653), .B1_t (new_AGEMA_signal_2654), .B1_f (new_AGEMA_signal_2655), .Z0_t (stateArray_outS01ser[4]), .Z0_f (new_AGEMA_signal_2605), .Z1_t (new_AGEMA_signal_2606), .Z1_f (new_AGEMA_signal_2607) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S01reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS02ser[5]), .A0_f (new_AGEMA_signal_2659), .A1_t (new_AGEMA_signal_2660), .A1_f (new_AGEMA_signal_2661), .B0_t (stateArray_outS01ser[5]), .B0_f (new_AGEMA_signal_2611), .B1_t (new_AGEMA_signal_2612), .B1_f (new_AGEMA_signal_2613), .Z0_t (stateArray_S01reg_gff_1_SFF_5_MUXInst_X), .Z0_f (new_AGEMA_signal_2662), .Z1_t (new_AGEMA_signal_2663), .Z1_f (new_AGEMA_signal_2664) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S01reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S01reg_gff_1_SFF_5_MUXInst_X), .B0_f (new_AGEMA_signal_2662), .B1_t (new_AGEMA_signal_2663), .B1_f (new_AGEMA_signal_2664), .Z0_t (stateArray_S01reg_gff_1_SFF_5_MUXInst_Y), .Z0_f (new_AGEMA_signal_5956), .Z1_t (new_AGEMA_signal_5957), .Z1_f (new_AGEMA_signal_5958) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S01reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (stateArray_S01reg_gff_1_SFF_5_MUXInst_Y), .A0_f (new_AGEMA_signal_5956), .A1_t (new_AGEMA_signal_5957), .A1_f (new_AGEMA_signal_5958), .B0_t (stateArray_outS02ser[5]), .B0_f (new_AGEMA_signal_2659), .B1_t (new_AGEMA_signal_2660), .B1_f (new_AGEMA_signal_2661), .Z0_t (stateArray_outS01ser[5]), .Z0_f (new_AGEMA_signal_2611), .Z1_t (new_AGEMA_signal_2612), .Z1_f (new_AGEMA_signal_2613) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S01reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS02ser[6]), .A0_f (new_AGEMA_signal_2665), .A1_t (new_AGEMA_signal_2666), .A1_f (new_AGEMA_signal_2667), .B0_t (stateArray_outS01ser[6]), .B0_f (new_AGEMA_signal_2617), .B1_t (new_AGEMA_signal_2618), .B1_f (new_AGEMA_signal_2619), .Z0_t (stateArray_S01reg_gff_1_SFF_6_MUXInst_X), .Z0_f (new_AGEMA_signal_2668), .Z1_t (new_AGEMA_signal_2669), .Z1_f (new_AGEMA_signal_2670) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S01reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S01reg_gff_1_SFF_6_MUXInst_X), .B0_f (new_AGEMA_signal_2668), .B1_t (new_AGEMA_signal_2669), .B1_f (new_AGEMA_signal_2670), .Z0_t (stateArray_S01reg_gff_1_SFF_6_MUXInst_Y), .Z0_f (new_AGEMA_signal_5959), .Z1_t (new_AGEMA_signal_5960), .Z1_f (new_AGEMA_signal_5961) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S01reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (stateArray_S01reg_gff_1_SFF_6_MUXInst_Y), .A0_f (new_AGEMA_signal_5959), .A1_t (new_AGEMA_signal_5960), .A1_f (new_AGEMA_signal_5961), .B0_t (stateArray_outS02ser[6]), .B0_f (new_AGEMA_signal_2665), .B1_t (new_AGEMA_signal_2666), .B1_f (new_AGEMA_signal_2667), .Z0_t (stateArray_outS01ser[6]), .Z0_f (new_AGEMA_signal_2617), .Z1_t (new_AGEMA_signal_2618), .Z1_f (new_AGEMA_signal_2619) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S01reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS02ser[7]), .A0_f (new_AGEMA_signal_2671), .A1_t (new_AGEMA_signal_2672), .A1_f (new_AGEMA_signal_2673), .B0_t (stateArray_outS01ser[7]), .B0_f (new_AGEMA_signal_2623), .B1_t (new_AGEMA_signal_2624), .B1_f (new_AGEMA_signal_2625), .Z0_t (stateArray_S01reg_gff_1_SFF_7_MUXInst_X), .Z0_f (new_AGEMA_signal_2674), .Z1_t (new_AGEMA_signal_2675), .Z1_f (new_AGEMA_signal_2676) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S01reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S01reg_gff_1_SFF_7_MUXInst_X), .B0_f (new_AGEMA_signal_2674), .B1_t (new_AGEMA_signal_2675), .B1_f (new_AGEMA_signal_2676), .Z0_t (stateArray_S01reg_gff_1_SFF_7_MUXInst_Y), .Z0_f (new_AGEMA_signal_5962), .Z1_t (new_AGEMA_signal_5963), .Z1_f (new_AGEMA_signal_5964) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S01reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (stateArray_S01reg_gff_1_SFF_7_MUXInst_Y), .A0_f (new_AGEMA_signal_5962), .A1_t (new_AGEMA_signal_5963), .A1_f (new_AGEMA_signal_5964), .B0_t (stateArray_outS02ser[7]), .B0_f (new_AGEMA_signal_2671), .B1_t (new_AGEMA_signal_2672), .B1_f (new_AGEMA_signal_2673), .Z0_t (stateArray_outS01ser[7]), .Z0_f (new_AGEMA_signal_2623), .Z1_t (new_AGEMA_signal_2624), .Z1_f (new_AGEMA_signal_2625) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S02reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS03ser[0]), .A0_f (new_AGEMA_signal_2677), .A1_t (new_AGEMA_signal_2678), .A1_f (new_AGEMA_signal_2679), .B0_t (stateArray_outS02ser[0]), .B0_f (new_AGEMA_signal_2629), .B1_t (new_AGEMA_signal_2630), .B1_f (new_AGEMA_signal_2631), .Z0_t (stateArray_S02reg_gff_1_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_2680), .Z1_t (new_AGEMA_signal_2681), .Z1_f (new_AGEMA_signal_2682) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S02reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S02reg_gff_1_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_2680), .B1_t (new_AGEMA_signal_2681), .B1_f (new_AGEMA_signal_2682), .Z0_t (stateArray_S02reg_gff_1_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_5965), .Z1_t (new_AGEMA_signal_5966), .Z1_f (new_AGEMA_signal_5967) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S02reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (stateArray_S02reg_gff_1_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_5965), .A1_t (new_AGEMA_signal_5966), .A1_f (new_AGEMA_signal_5967), .B0_t (stateArray_outS03ser[0]), .B0_f (new_AGEMA_signal_2677), .B1_t (new_AGEMA_signal_2678), .B1_f (new_AGEMA_signal_2679), .Z0_t (stateArray_outS02ser[0]), .Z0_f (new_AGEMA_signal_2629), .Z1_t (new_AGEMA_signal_2630), .Z1_f (new_AGEMA_signal_2631) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S02reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS03ser[1]), .A0_f (new_AGEMA_signal_2683), .A1_t (new_AGEMA_signal_2684), .A1_f (new_AGEMA_signal_2685), .B0_t (stateArray_outS02ser[1]), .B0_f (new_AGEMA_signal_2635), .B1_t (new_AGEMA_signal_2636), .B1_f (new_AGEMA_signal_2637), .Z0_t (stateArray_S02reg_gff_1_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_2686), .Z1_t (new_AGEMA_signal_2687), .Z1_f (new_AGEMA_signal_2688) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S02reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S02reg_gff_1_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_2686), .B1_t (new_AGEMA_signal_2687), .B1_f (new_AGEMA_signal_2688), .Z0_t (stateArray_S02reg_gff_1_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_5968), .Z1_t (new_AGEMA_signal_5969), .Z1_f (new_AGEMA_signal_5970) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S02reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (stateArray_S02reg_gff_1_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_5968), .A1_t (new_AGEMA_signal_5969), .A1_f (new_AGEMA_signal_5970), .B0_t (stateArray_outS03ser[1]), .B0_f (new_AGEMA_signal_2683), .B1_t (new_AGEMA_signal_2684), .B1_f (new_AGEMA_signal_2685), .Z0_t (stateArray_outS02ser[1]), .Z0_f (new_AGEMA_signal_2635), .Z1_t (new_AGEMA_signal_2636), .Z1_f (new_AGEMA_signal_2637) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S02reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS03ser[2]), .A0_f (new_AGEMA_signal_2689), .A1_t (new_AGEMA_signal_2690), .A1_f (new_AGEMA_signal_2691), .B0_t (stateArray_outS02ser[2]), .B0_f (new_AGEMA_signal_2641), .B1_t (new_AGEMA_signal_2642), .B1_f (new_AGEMA_signal_2643), .Z0_t (stateArray_S02reg_gff_1_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_2692), .Z1_t (new_AGEMA_signal_2693), .Z1_f (new_AGEMA_signal_2694) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S02reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S02reg_gff_1_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_2692), .B1_t (new_AGEMA_signal_2693), .B1_f (new_AGEMA_signal_2694), .Z0_t (stateArray_S02reg_gff_1_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_5971), .Z1_t (new_AGEMA_signal_5972), .Z1_f (new_AGEMA_signal_5973) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S02reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (stateArray_S02reg_gff_1_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_5971), .A1_t (new_AGEMA_signal_5972), .A1_f (new_AGEMA_signal_5973), .B0_t (stateArray_outS03ser[2]), .B0_f (new_AGEMA_signal_2689), .B1_t (new_AGEMA_signal_2690), .B1_f (new_AGEMA_signal_2691), .Z0_t (stateArray_outS02ser[2]), .Z0_f (new_AGEMA_signal_2641), .Z1_t (new_AGEMA_signal_2642), .Z1_f (new_AGEMA_signal_2643) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S02reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS03ser[3]), .A0_f (new_AGEMA_signal_2695), .A1_t (new_AGEMA_signal_2696), .A1_f (new_AGEMA_signal_2697), .B0_t (stateArray_outS02ser[3]), .B0_f (new_AGEMA_signal_2647), .B1_t (new_AGEMA_signal_2648), .B1_f (new_AGEMA_signal_2649), .Z0_t (stateArray_S02reg_gff_1_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_2698), .Z1_t (new_AGEMA_signal_2699), .Z1_f (new_AGEMA_signal_2700) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S02reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S02reg_gff_1_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_2698), .B1_t (new_AGEMA_signal_2699), .B1_f (new_AGEMA_signal_2700), .Z0_t (stateArray_S02reg_gff_1_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_5974), .Z1_t (new_AGEMA_signal_5975), .Z1_f (new_AGEMA_signal_5976) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S02reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (stateArray_S02reg_gff_1_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_5974), .A1_t (new_AGEMA_signal_5975), .A1_f (new_AGEMA_signal_5976), .B0_t (stateArray_outS03ser[3]), .B0_f (new_AGEMA_signal_2695), .B1_t (new_AGEMA_signal_2696), .B1_f (new_AGEMA_signal_2697), .Z0_t (stateArray_outS02ser[3]), .Z0_f (new_AGEMA_signal_2647), .Z1_t (new_AGEMA_signal_2648), .Z1_f (new_AGEMA_signal_2649) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S02reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS03ser[4]), .A0_f (new_AGEMA_signal_2701), .A1_t (new_AGEMA_signal_2702), .A1_f (new_AGEMA_signal_2703), .B0_t (stateArray_outS02ser[4]), .B0_f (new_AGEMA_signal_2653), .B1_t (new_AGEMA_signal_2654), .B1_f (new_AGEMA_signal_2655), .Z0_t (stateArray_S02reg_gff_1_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_2704), .Z1_t (new_AGEMA_signal_2705), .Z1_f (new_AGEMA_signal_2706) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S02reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S02reg_gff_1_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_2704), .B1_t (new_AGEMA_signal_2705), .B1_f (new_AGEMA_signal_2706), .Z0_t (stateArray_S02reg_gff_1_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_5977), .Z1_t (new_AGEMA_signal_5978), .Z1_f (new_AGEMA_signal_5979) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S02reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (stateArray_S02reg_gff_1_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_5977), .A1_t (new_AGEMA_signal_5978), .A1_f (new_AGEMA_signal_5979), .B0_t (stateArray_outS03ser[4]), .B0_f (new_AGEMA_signal_2701), .B1_t (new_AGEMA_signal_2702), .B1_f (new_AGEMA_signal_2703), .Z0_t (stateArray_outS02ser[4]), .Z0_f (new_AGEMA_signal_2653), .Z1_t (new_AGEMA_signal_2654), .Z1_f (new_AGEMA_signal_2655) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S02reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS03ser[5]), .A0_f (new_AGEMA_signal_2707), .A1_t (new_AGEMA_signal_2708), .A1_f (new_AGEMA_signal_2709), .B0_t (stateArray_outS02ser[5]), .B0_f (new_AGEMA_signal_2659), .B1_t (new_AGEMA_signal_2660), .B1_f (new_AGEMA_signal_2661), .Z0_t (stateArray_S02reg_gff_1_SFF_5_MUXInst_X), .Z0_f (new_AGEMA_signal_2710), .Z1_t (new_AGEMA_signal_2711), .Z1_f (new_AGEMA_signal_2712) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S02reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S02reg_gff_1_SFF_5_MUXInst_X), .B0_f (new_AGEMA_signal_2710), .B1_t (new_AGEMA_signal_2711), .B1_f (new_AGEMA_signal_2712), .Z0_t (stateArray_S02reg_gff_1_SFF_5_MUXInst_Y), .Z0_f (new_AGEMA_signal_5980), .Z1_t (new_AGEMA_signal_5981), .Z1_f (new_AGEMA_signal_5982) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S02reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (stateArray_S02reg_gff_1_SFF_5_MUXInst_Y), .A0_f (new_AGEMA_signal_5980), .A1_t (new_AGEMA_signal_5981), .A1_f (new_AGEMA_signal_5982), .B0_t (stateArray_outS03ser[5]), .B0_f (new_AGEMA_signal_2707), .B1_t (new_AGEMA_signal_2708), .B1_f (new_AGEMA_signal_2709), .Z0_t (stateArray_outS02ser[5]), .Z0_f (new_AGEMA_signal_2659), .Z1_t (new_AGEMA_signal_2660), .Z1_f (new_AGEMA_signal_2661) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S02reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS03ser[6]), .A0_f (new_AGEMA_signal_2713), .A1_t (new_AGEMA_signal_2714), .A1_f (new_AGEMA_signal_2715), .B0_t (stateArray_outS02ser[6]), .B0_f (new_AGEMA_signal_2665), .B1_t (new_AGEMA_signal_2666), .B1_f (new_AGEMA_signal_2667), .Z0_t (stateArray_S02reg_gff_1_SFF_6_MUXInst_X), .Z0_f (new_AGEMA_signal_2716), .Z1_t (new_AGEMA_signal_2717), .Z1_f (new_AGEMA_signal_2718) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S02reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S02reg_gff_1_SFF_6_MUXInst_X), .B0_f (new_AGEMA_signal_2716), .B1_t (new_AGEMA_signal_2717), .B1_f (new_AGEMA_signal_2718), .Z0_t (stateArray_S02reg_gff_1_SFF_6_MUXInst_Y), .Z0_f (new_AGEMA_signal_5983), .Z1_t (new_AGEMA_signal_5984), .Z1_f (new_AGEMA_signal_5985) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S02reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (stateArray_S02reg_gff_1_SFF_6_MUXInst_Y), .A0_f (new_AGEMA_signal_5983), .A1_t (new_AGEMA_signal_5984), .A1_f (new_AGEMA_signal_5985), .B0_t (stateArray_outS03ser[6]), .B0_f (new_AGEMA_signal_2713), .B1_t (new_AGEMA_signal_2714), .B1_f (new_AGEMA_signal_2715), .Z0_t (stateArray_outS02ser[6]), .Z0_f (new_AGEMA_signal_2665), .Z1_t (new_AGEMA_signal_2666), .Z1_f (new_AGEMA_signal_2667) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S02reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS03ser[7]), .A0_f (new_AGEMA_signal_2719), .A1_t (new_AGEMA_signal_2720), .A1_f (new_AGEMA_signal_2721), .B0_t (stateArray_outS02ser[7]), .B0_f (new_AGEMA_signal_2671), .B1_t (new_AGEMA_signal_2672), .B1_f (new_AGEMA_signal_2673), .Z0_t (stateArray_S02reg_gff_1_SFF_7_MUXInst_X), .Z0_f (new_AGEMA_signal_2722), .Z1_t (new_AGEMA_signal_2723), .Z1_f (new_AGEMA_signal_2724) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S02reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S02reg_gff_1_SFF_7_MUXInst_X), .B0_f (new_AGEMA_signal_2722), .B1_t (new_AGEMA_signal_2723), .B1_f (new_AGEMA_signal_2724), .Z0_t (stateArray_S02reg_gff_1_SFF_7_MUXInst_Y), .Z0_f (new_AGEMA_signal_5986), .Z1_t (new_AGEMA_signal_5987), .Z1_f (new_AGEMA_signal_5988) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S02reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (stateArray_S02reg_gff_1_SFF_7_MUXInst_Y), .A0_f (new_AGEMA_signal_5986), .A1_t (new_AGEMA_signal_5987), .A1_f (new_AGEMA_signal_5988), .B0_t (stateArray_outS03ser[7]), .B0_f (new_AGEMA_signal_2719), .B1_t (new_AGEMA_signal_2720), .B1_f (new_AGEMA_signal_2721), .Z0_t (stateArray_outS02ser[7]), .Z0_f (new_AGEMA_signal_2671), .Z1_t (new_AGEMA_signal_2672), .Z1_f (new_AGEMA_signal_2673) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S03reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS03ser[0]), .A0_f (new_AGEMA_signal_6205), .A1_t (new_AGEMA_signal_6206), .A1_f (new_AGEMA_signal_6207), .B0_t (stateArray_outS03ser[0]), .B0_f (new_AGEMA_signal_2677), .B1_t (new_AGEMA_signal_2678), .B1_f (new_AGEMA_signal_2679), .Z0_t (stateArray_S03reg_gff_1_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_6319), .Z1_t (new_AGEMA_signal_6320), .Z1_f (new_AGEMA_signal_6321) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S03reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S03reg_gff_1_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_6319), .B1_t (new_AGEMA_signal_6320), .B1_f (new_AGEMA_signal_6321), .Z0_t (stateArray_S03reg_gff_1_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_7158), .Z1_t (new_AGEMA_signal_7159), .Z1_f (new_AGEMA_signal_7160) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S03reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (stateArray_S03reg_gff_1_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_7158), .A1_t (new_AGEMA_signal_7159), .A1_f (new_AGEMA_signal_7160), .B0_t (stateArray_inS03ser[0]), .B0_f (new_AGEMA_signal_6205), .B1_t (new_AGEMA_signal_6206), .B1_f (new_AGEMA_signal_6207), .Z0_t (stateArray_outS03ser[0]), .Z0_f (new_AGEMA_signal_2677), .Z1_t (new_AGEMA_signal_2678), .Z1_f (new_AGEMA_signal_2679) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S03reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS03ser[1]), .A0_f (new_AGEMA_signal_6364), .A1_t (new_AGEMA_signal_6365), .A1_f (new_AGEMA_signal_6366), .B0_t (stateArray_outS03ser[1]), .B0_f (new_AGEMA_signal_2683), .B1_t (new_AGEMA_signal_2684), .B1_f (new_AGEMA_signal_2685), .Z0_t (stateArray_S03reg_gff_1_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_7161), .Z1_t (new_AGEMA_signal_7162), .Z1_f (new_AGEMA_signal_7163) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S03reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S03reg_gff_1_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_7161), .B1_t (new_AGEMA_signal_7162), .B1_f (new_AGEMA_signal_7163), .Z0_t (stateArray_S03reg_gff_1_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_7274), .Z1_t (new_AGEMA_signal_7275), .Z1_f (new_AGEMA_signal_7276) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S03reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (stateArray_S03reg_gff_1_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_7274), .A1_t (new_AGEMA_signal_7275), .A1_f (new_AGEMA_signal_7276), .B0_t (stateArray_inS03ser[1]), .B0_f (new_AGEMA_signal_6364), .B1_t (new_AGEMA_signal_6365), .B1_f (new_AGEMA_signal_6366), .Z0_t (stateArray_outS03ser[1]), .Z0_f (new_AGEMA_signal_2683), .Z1_t (new_AGEMA_signal_2684), .Z1_f (new_AGEMA_signal_2685) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S03reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS03ser[2]), .A0_f (new_AGEMA_signal_6211), .A1_t (new_AGEMA_signal_6212), .A1_f (new_AGEMA_signal_6213), .B0_t (stateArray_outS03ser[2]), .B0_f (new_AGEMA_signal_2689), .B1_t (new_AGEMA_signal_2690), .B1_f (new_AGEMA_signal_2691), .Z0_t (stateArray_S03reg_gff_1_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_6322), .Z1_t (new_AGEMA_signal_6323), .Z1_f (new_AGEMA_signal_6324) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S03reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S03reg_gff_1_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_6322), .B1_t (new_AGEMA_signal_6323), .B1_f (new_AGEMA_signal_6324), .Z0_t (stateArray_S03reg_gff_1_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_7164), .Z1_t (new_AGEMA_signal_7165), .Z1_f (new_AGEMA_signal_7166) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S03reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (stateArray_S03reg_gff_1_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_7164), .A1_t (new_AGEMA_signal_7165), .A1_f (new_AGEMA_signal_7166), .B0_t (stateArray_inS03ser[2]), .B0_f (new_AGEMA_signal_6211), .B1_t (new_AGEMA_signal_6212), .B1_f (new_AGEMA_signal_6213), .Z0_t (stateArray_outS03ser[2]), .Z0_f (new_AGEMA_signal_2689), .Z1_t (new_AGEMA_signal_2690), .Z1_f (new_AGEMA_signal_2691) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S03reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS03ser[3]), .A0_f (new_AGEMA_signal_6367), .A1_t (new_AGEMA_signal_6368), .A1_f (new_AGEMA_signal_6369), .B0_t (stateArray_outS03ser[3]), .B0_f (new_AGEMA_signal_2695), .B1_t (new_AGEMA_signal_2696), .B1_f (new_AGEMA_signal_2697), .Z0_t (stateArray_S03reg_gff_1_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_7167), .Z1_t (new_AGEMA_signal_7168), .Z1_f (new_AGEMA_signal_7169) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S03reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S03reg_gff_1_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_7167), .B1_t (new_AGEMA_signal_7168), .B1_f (new_AGEMA_signal_7169), .Z0_t (stateArray_S03reg_gff_1_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_7277), .Z1_t (new_AGEMA_signal_7278), .Z1_f (new_AGEMA_signal_7279) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S03reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (stateArray_S03reg_gff_1_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_7277), .A1_t (new_AGEMA_signal_7278), .A1_f (new_AGEMA_signal_7279), .B0_t (stateArray_inS03ser[3]), .B0_f (new_AGEMA_signal_6367), .B1_t (new_AGEMA_signal_6368), .B1_f (new_AGEMA_signal_6369), .Z0_t (stateArray_outS03ser[3]), .Z0_f (new_AGEMA_signal_2695), .Z1_t (new_AGEMA_signal_2696), .Z1_f (new_AGEMA_signal_2697) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S03reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS03ser[4]), .A0_f (new_AGEMA_signal_6370), .A1_t (new_AGEMA_signal_6371), .A1_f (new_AGEMA_signal_6372), .B0_t (stateArray_outS03ser[4]), .B0_f (new_AGEMA_signal_2701), .B1_t (new_AGEMA_signal_2702), .B1_f (new_AGEMA_signal_2703), .Z0_t (stateArray_S03reg_gff_1_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_7170), .Z1_t (new_AGEMA_signal_7171), .Z1_f (new_AGEMA_signal_7172) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S03reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S03reg_gff_1_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_7170), .B1_t (new_AGEMA_signal_7171), .B1_f (new_AGEMA_signal_7172), .Z0_t (stateArray_S03reg_gff_1_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_7280), .Z1_t (new_AGEMA_signal_7281), .Z1_f (new_AGEMA_signal_7282) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S03reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (stateArray_S03reg_gff_1_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_7280), .A1_t (new_AGEMA_signal_7281), .A1_f (new_AGEMA_signal_7282), .B0_t (stateArray_inS03ser[4]), .B0_f (new_AGEMA_signal_6370), .B1_t (new_AGEMA_signal_6371), .B1_f (new_AGEMA_signal_6372), .Z0_t (stateArray_outS03ser[4]), .Z0_f (new_AGEMA_signal_2701), .Z1_t (new_AGEMA_signal_2702), .Z1_f (new_AGEMA_signal_2703) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S03reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS03ser[5]), .A0_f (new_AGEMA_signal_6220), .A1_t (new_AGEMA_signal_6221), .A1_f (new_AGEMA_signal_6222), .B0_t (stateArray_outS03ser[5]), .B0_f (new_AGEMA_signal_2707), .B1_t (new_AGEMA_signal_2708), .B1_f (new_AGEMA_signal_2709), .Z0_t (stateArray_S03reg_gff_1_SFF_5_MUXInst_X), .Z0_f (new_AGEMA_signal_6325), .Z1_t (new_AGEMA_signal_6326), .Z1_f (new_AGEMA_signal_6327) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S03reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S03reg_gff_1_SFF_5_MUXInst_X), .B0_f (new_AGEMA_signal_6325), .B1_t (new_AGEMA_signal_6326), .B1_f (new_AGEMA_signal_6327), .Z0_t (stateArray_S03reg_gff_1_SFF_5_MUXInst_Y), .Z0_f (new_AGEMA_signal_7173), .Z1_t (new_AGEMA_signal_7174), .Z1_f (new_AGEMA_signal_7175) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S03reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (stateArray_S03reg_gff_1_SFF_5_MUXInst_Y), .A0_f (new_AGEMA_signal_7173), .A1_t (new_AGEMA_signal_7174), .A1_f (new_AGEMA_signal_7175), .B0_t (stateArray_inS03ser[5]), .B0_f (new_AGEMA_signal_6220), .B1_t (new_AGEMA_signal_6221), .B1_f (new_AGEMA_signal_6222), .Z0_t (stateArray_outS03ser[5]), .Z0_f (new_AGEMA_signal_2707), .Z1_t (new_AGEMA_signal_2708), .Z1_f (new_AGEMA_signal_2709) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S03reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS03ser[6]), .A0_f (new_AGEMA_signal_6223), .A1_t (new_AGEMA_signal_6224), .A1_f (new_AGEMA_signal_6225), .B0_t (stateArray_outS03ser[6]), .B0_f (new_AGEMA_signal_2713), .B1_t (new_AGEMA_signal_2714), .B1_f (new_AGEMA_signal_2715), .Z0_t (stateArray_S03reg_gff_1_SFF_6_MUXInst_X), .Z0_f (new_AGEMA_signal_6328), .Z1_t (new_AGEMA_signal_6329), .Z1_f (new_AGEMA_signal_6330) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S03reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S03reg_gff_1_SFF_6_MUXInst_X), .B0_f (new_AGEMA_signal_6328), .B1_t (new_AGEMA_signal_6329), .B1_f (new_AGEMA_signal_6330), .Z0_t (stateArray_S03reg_gff_1_SFF_6_MUXInst_Y), .Z0_f (new_AGEMA_signal_7176), .Z1_t (new_AGEMA_signal_7177), .Z1_f (new_AGEMA_signal_7178) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S03reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (stateArray_S03reg_gff_1_SFF_6_MUXInst_Y), .A0_f (new_AGEMA_signal_7176), .A1_t (new_AGEMA_signal_7177), .A1_f (new_AGEMA_signal_7178), .B0_t (stateArray_inS03ser[6]), .B0_f (new_AGEMA_signal_6223), .B1_t (new_AGEMA_signal_6224), .B1_f (new_AGEMA_signal_6225), .Z0_t (stateArray_outS03ser[6]), .Z0_f (new_AGEMA_signal_2713), .Z1_t (new_AGEMA_signal_2714), .Z1_f (new_AGEMA_signal_2715) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S03reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS03ser[7]), .A0_f (new_AGEMA_signal_6226), .A1_t (new_AGEMA_signal_6227), .A1_f (new_AGEMA_signal_6228), .B0_t (stateArray_outS03ser[7]), .B0_f (new_AGEMA_signal_2719), .B1_t (new_AGEMA_signal_2720), .B1_f (new_AGEMA_signal_2721), .Z0_t (stateArray_S03reg_gff_1_SFF_7_MUXInst_X), .Z0_f (new_AGEMA_signal_6331), .Z1_t (new_AGEMA_signal_6332), .Z1_f (new_AGEMA_signal_6333) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S03reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S03reg_gff_1_SFF_7_MUXInst_X), .B0_f (new_AGEMA_signal_6331), .B1_t (new_AGEMA_signal_6332), .B1_f (new_AGEMA_signal_6333), .Z0_t (stateArray_S03reg_gff_1_SFF_7_MUXInst_Y), .Z0_f (new_AGEMA_signal_7179), .Z1_t (new_AGEMA_signal_7180), .Z1_f (new_AGEMA_signal_7181) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S03reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (stateArray_S03reg_gff_1_SFF_7_MUXInst_Y), .A0_f (new_AGEMA_signal_7179), .A1_t (new_AGEMA_signal_7180), .A1_f (new_AGEMA_signal_7181), .B0_t (stateArray_inS03ser[7]), .B0_f (new_AGEMA_signal_6226), .B1_t (new_AGEMA_signal_6227), .B1_f (new_AGEMA_signal_6228), .Z0_t (stateArray_outS03ser[7]), .Z0_f (new_AGEMA_signal_2719), .Z1_t (new_AGEMA_signal_2720), .Z1_f (new_AGEMA_signal_2721) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S10reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS11ser[0]), .A0_f (new_AGEMA_signal_2725), .A1_t (new_AGEMA_signal_2726), .A1_f (new_AGEMA_signal_2727), .B0_t (stateArray_outS11ser[0]), .B0_f (new_AGEMA_signal_2725), .B1_t (new_AGEMA_signal_2726), .B1_f (new_AGEMA_signal_2727), .Z0_t (stateArray_S10reg_gff_1_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_2728), .Z1_t (new_AGEMA_signal_2729), .Z1_f (new_AGEMA_signal_2730) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S10reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S10reg_gff_1_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_2728), .B1_t (new_AGEMA_signal_2729), .B1_f (new_AGEMA_signal_2730), .Z0_t (stateArray_S10reg_gff_1_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_5989), .Z1_t (new_AGEMA_signal_5990), .Z1_f (new_AGEMA_signal_5991) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S10reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (stateArray_S10reg_gff_1_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_5989), .A1_t (new_AGEMA_signal_5990), .A1_f (new_AGEMA_signal_5991), .B0_t (stateArray_outS11ser[0]), .B0_f (new_AGEMA_signal_2725), .B1_t (new_AGEMA_signal_2726), .B1_f (new_AGEMA_signal_2727), .Z0_t (MCin[16]), .Z0_f (new_AGEMA_signal_3988), .Z1_t (new_AGEMA_signal_3989), .Z1_f (new_AGEMA_signal_3990) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S10reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS11ser[1]), .A0_f (new_AGEMA_signal_2731), .A1_t (new_AGEMA_signal_2732), .A1_f (new_AGEMA_signal_2733), .B0_t (stateArray_outS11ser[1]), .B0_f (new_AGEMA_signal_2731), .B1_t (new_AGEMA_signal_2732), .B1_f (new_AGEMA_signal_2733), .Z0_t (stateArray_S10reg_gff_1_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_2734), .Z1_t (new_AGEMA_signal_2735), .Z1_f (new_AGEMA_signal_2736) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S10reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S10reg_gff_1_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_2734), .B1_t (new_AGEMA_signal_2735), .B1_f (new_AGEMA_signal_2736), .Z0_t (stateArray_S10reg_gff_1_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_5992), .Z1_t (new_AGEMA_signal_5993), .Z1_f (new_AGEMA_signal_5994) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S10reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (stateArray_S10reg_gff_1_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_5992), .A1_t (new_AGEMA_signal_5993), .A1_f (new_AGEMA_signal_5994), .B0_t (stateArray_outS11ser[1]), .B0_f (new_AGEMA_signal_2731), .B1_t (new_AGEMA_signal_2732), .B1_f (new_AGEMA_signal_2733), .Z0_t (MixColumns_line1_S02[2]), .Z0_f (new_AGEMA_signal_3982), .Z1_t (new_AGEMA_signal_3983), .Z1_f (new_AGEMA_signal_3984) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S10reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS11ser[2]), .A0_f (new_AGEMA_signal_2737), .A1_t (new_AGEMA_signal_2738), .A1_f (new_AGEMA_signal_2739), .B0_t (stateArray_outS11ser[2]), .B0_f (new_AGEMA_signal_2737), .B1_t (new_AGEMA_signal_2738), .B1_f (new_AGEMA_signal_2739), .Z0_t (stateArray_S10reg_gff_1_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_2740), .Z1_t (new_AGEMA_signal_2741), .Z1_f (new_AGEMA_signal_2742) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S10reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S10reg_gff_1_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_2740), .B1_t (new_AGEMA_signal_2741), .B1_f (new_AGEMA_signal_2742), .Z0_t (stateArray_S10reg_gff_1_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_5995), .Z1_t (new_AGEMA_signal_5996), .Z1_f (new_AGEMA_signal_5997) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S10reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (stateArray_S10reg_gff_1_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_5995), .A1_t (new_AGEMA_signal_5996), .A1_f (new_AGEMA_signal_5997), .B0_t (stateArray_outS11ser[2]), .B0_f (new_AGEMA_signal_2737), .B1_t (new_AGEMA_signal_2738), .B1_f (new_AGEMA_signal_2739), .Z0_t (MCin[18]), .Z0_f (new_AGEMA_signal_3979), .Z1_t (new_AGEMA_signal_3980), .Z1_f (new_AGEMA_signal_3981) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S10reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS11ser[3]), .A0_f (new_AGEMA_signal_2743), .A1_t (new_AGEMA_signal_2744), .A1_f (new_AGEMA_signal_2745), .B0_t (stateArray_outS11ser[3]), .B0_f (new_AGEMA_signal_2743), .B1_t (new_AGEMA_signal_2744), .B1_f (new_AGEMA_signal_2745), .Z0_t (stateArray_S10reg_gff_1_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_2746), .Z1_t (new_AGEMA_signal_2747), .Z1_f (new_AGEMA_signal_2748) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S10reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S10reg_gff_1_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_2746), .B1_t (new_AGEMA_signal_2747), .B1_f (new_AGEMA_signal_2748), .Z0_t (stateArray_S10reg_gff_1_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_5998), .Z1_t (new_AGEMA_signal_5999), .Z1_f (new_AGEMA_signal_6000) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S10reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (stateArray_S10reg_gff_1_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_5998), .A1_t (new_AGEMA_signal_5999), .A1_f (new_AGEMA_signal_6000), .B0_t (stateArray_outS11ser[3]), .B0_f (new_AGEMA_signal_2743), .B1_t (new_AGEMA_signal_2744), .B1_f (new_AGEMA_signal_2745), .Z0_t (MCin[19]), .Z0_f (new_AGEMA_signal_3994), .Z1_t (new_AGEMA_signal_3995), .Z1_f (new_AGEMA_signal_3996) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S10reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS11ser[4]), .A0_f (new_AGEMA_signal_2749), .A1_t (new_AGEMA_signal_2750), .A1_f (new_AGEMA_signal_2751), .B0_t (stateArray_outS11ser[4]), .B0_f (new_AGEMA_signal_2749), .B1_t (new_AGEMA_signal_2750), .B1_f (new_AGEMA_signal_2751), .Z0_t (stateArray_S10reg_gff_1_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_2752), .Z1_t (new_AGEMA_signal_2753), .Z1_f (new_AGEMA_signal_2754) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S10reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S10reg_gff_1_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_2752), .B1_t (new_AGEMA_signal_2753), .B1_f (new_AGEMA_signal_2754), .Z0_t (stateArray_S10reg_gff_1_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_6001), .Z1_t (new_AGEMA_signal_6002), .Z1_f (new_AGEMA_signal_6003) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S10reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (stateArray_S10reg_gff_1_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_6001), .A1_t (new_AGEMA_signal_6002), .A1_f (new_AGEMA_signal_6003), .B0_t (stateArray_outS11ser[4]), .B0_f (new_AGEMA_signal_2749), .B1_t (new_AGEMA_signal_2750), .B1_f (new_AGEMA_signal_2751), .Z0_t (MixColumns_line1_S02[5]), .Z0_f (new_AGEMA_signal_3973), .Z1_t (new_AGEMA_signal_3974), .Z1_f (new_AGEMA_signal_3975) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S10reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS11ser[5]), .A0_f (new_AGEMA_signal_2755), .A1_t (new_AGEMA_signal_2756), .A1_f (new_AGEMA_signal_2757), .B0_t (stateArray_outS11ser[5]), .B0_f (new_AGEMA_signal_2755), .B1_t (new_AGEMA_signal_2756), .B1_f (new_AGEMA_signal_2757), .Z0_t (stateArray_S10reg_gff_1_SFF_5_MUXInst_X), .Z0_f (new_AGEMA_signal_2758), .Z1_t (new_AGEMA_signal_2759), .Z1_f (new_AGEMA_signal_2760) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S10reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S10reg_gff_1_SFF_5_MUXInst_X), .B0_f (new_AGEMA_signal_2758), .B1_t (new_AGEMA_signal_2759), .B1_f (new_AGEMA_signal_2760), .Z0_t (stateArray_S10reg_gff_1_SFF_5_MUXInst_Y), .Z0_f (new_AGEMA_signal_6004), .Z1_t (new_AGEMA_signal_6005), .Z1_f (new_AGEMA_signal_6006) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S10reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (stateArray_S10reg_gff_1_SFF_5_MUXInst_Y), .A0_f (new_AGEMA_signal_6004), .A1_t (new_AGEMA_signal_6005), .A1_f (new_AGEMA_signal_6006), .B0_t (stateArray_outS11ser[5]), .B0_f (new_AGEMA_signal_2755), .B1_t (new_AGEMA_signal_2756), .B1_f (new_AGEMA_signal_2757), .Z0_t (MixColumns_line1_S02[6]), .Z0_f (new_AGEMA_signal_3967), .Z1_t (new_AGEMA_signal_3968), .Z1_f (new_AGEMA_signal_3969) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S10reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS11ser[6]), .A0_f (new_AGEMA_signal_2761), .A1_t (new_AGEMA_signal_2762), .A1_f (new_AGEMA_signal_2763), .B0_t (stateArray_outS11ser[6]), .B0_f (new_AGEMA_signal_2761), .B1_t (new_AGEMA_signal_2762), .B1_f (new_AGEMA_signal_2763), .Z0_t (stateArray_S10reg_gff_1_SFF_6_MUXInst_X), .Z0_f (new_AGEMA_signal_2764), .Z1_t (new_AGEMA_signal_2765), .Z1_f (new_AGEMA_signal_2766) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S10reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S10reg_gff_1_SFF_6_MUXInst_X), .B0_f (new_AGEMA_signal_2764), .B1_t (new_AGEMA_signal_2765), .B1_f (new_AGEMA_signal_2766), .Z0_t (stateArray_S10reg_gff_1_SFF_6_MUXInst_Y), .Z0_f (new_AGEMA_signal_6007), .Z1_t (new_AGEMA_signal_6008), .Z1_f (new_AGEMA_signal_6009) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S10reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (stateArray_S10reg_gff_1_SFF_6_MUXInst_Y), .A0_f (new_AGEMA_signal_6007), .A1_t (new_AGEMA_signal_6008), .A1_f (new_AGEMA_signal_6009), .B0_t (stateArray_outS11ser[6]), .B0_f (new_AGEMA_signal_2761), .B1_t (new_AGEMA_signal_2762), .B1_f (new_AGEMA_signal_2763), .Z0_t (MixColumns_line1_S02[7]), .Z0_f (new_AGEMA_signal_3961), .Z1_t (new_AGEMA_signal_3962), .Z1_f (new_AGEMA_signal_3963) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S10reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS11ser[7]), .A0_f (new_AGEMA_signal_2767), .A1_t (new_AGEMA_signal_2768), .A1_f (new_AGEMA_signal_2769), .B0_t (stateArray_outS11ser[7]), .B0_f (new_AGEMA_signal_2767), .B1_t (new_AGEMA_signal_2768), .B1_f (new_AGEMA_signal_2769), .Z0_t (stateArray_S10reg_gff_1_SFF_7_MUXInst_X), .Z0_f (new_AGEMA_signal_2770), .Z1_t (new_AGEMA_signal_2771), .Z1_f (new_AGEMA_signal_2772) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S10reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S10reg_gff_1_SFF_7_MUXInst_X), .B0_f (new_AGEMA_signal_2770), .B1_t (new_AGEMA_signal_2771), .B1_f (new_AGEMA_signal_2772), .Z0_t (stateArray_S10reg_gff_1_SFF_7_MUXInst_Y), .Z0_f (new_AGEMA_signal_6010), .Z1_t (new_AGEMA_signal_6011), .Z1_f (new_AGEMA_signal_6012) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S10reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (stateArray_S10reg_gff_1_SFF_7_MUXInst_Y), .A0_f (new_AGEMA_signal_6010), .A1_t (new_AGEMA_signal_6011), .A1_f (new_AGEMA_signal_6012), .B0_t (stateArray_outS11ser[7]), .B0_f (new_AGEMA_signal_2767), .B1_t (new_AGEMA_signal_2768), .B1_f (new_AGEMA_signal_2769), .Z0_t (MixColumns_line1_S02[0]), .Z0_f (new_AGEMA_signal_3958), .Z1_t (new_AGEMA_signal_3959), .Z1_f (new_AGEMA_signal_3960) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S11reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS12ser[0]), .A0_f (new_AGEMA_signal_2773), .A1_t (new_AGEMA_signal_2774), .A1_f (new_AGEMA_signal_2775), .B0_t (stateArray_outS12ser[0]), .B0_f (new_AGEMA_signal_2773), .B1_t (new_AGEMA_signal_2774), .B1_f (new_AGEMA_signal_2775), .Z0_t (stateArray_S11reg_gff_1_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_2776), .Z1_t (new_AGEMA_signal_2777), .Z1_f (new_AGEMA_signal_2778) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S11reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S11reg_gff_1_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_2776), .B1_t (new_AGEMA_signal_2777), .B1_f (new_AGEMA_signal_2778), .Z0_t (stateArray_S11reg_gff_1_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_6013), .Z1_t (new_AGEMA_signal_6014), .Z1_f (new_AGEMA_signal_6015) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S11reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (stateArray_S11reg_gff_1_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_6013), .A1_t (new_AGEMA_signal_6014), .A1_f (new_AGEMA_signal_6015), .B0_t (stateArray_outS12ser[0]), .B0_f (new_AGEMA_signal_2773), .B1_t (new_AGEMA_signal_2774), .B1_f (new_AGEMA_signal_2775), .Z0_t (stateArray_outS11ser[0]), .Z0_f (new_AGEMA_signal_2725), .Z1_t (new_AGEMA_signal_2726), .Z1_f (new_AGEMA_signal_2727) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S11reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS12ser[1]), .A0_f (new_AGEMA_signal_2779), .A1_t (new_AGEMA_signal_2780), .A1_f (new_AGEMA_signal_2781), .B0_t (stateArray_outS12ser[1]), .B0_f (new_AGEMA_signal_2779), .B1_t (new_AGEMA_signal_2780), .B1_f (new_AGEMA_signal_2781), .Z0_t (stateArray_S11reg_gff_1_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_2782), .Z1_t (new_AGEMA_signal_2783), .Z1_f (new_AGEMA_signal_2784) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S11reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S11reg_gff_1_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_2782), .B1_t (new_AGEMA_signal_2783), .B1_f (new_AGEMA_signal_2784), .Z0_t (stateArray_S11reg_gff_1_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_6016), .Z1_t (new_AGEMA_signal_6017), .Z1_f (new_AGEMA_signal_6018) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S11reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (stateArray_S11reg_gff_1_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_6016), .A1_t (new_AGEMA_signal_6017), .A1_f (new_AGEMA_signal_6018), .B0_t (stateArray_outS12ser[1]), .B0_f (new_AGEMA_signal_2779), .B1_t (new_AGEMA_signal_2780), .B1_f (new_AGEMA_signal_2781), .Z0_t (stateArray_outS11ser[1]), .Z0_f (new_AGEMA_signal_2731), .Z1_t (new_AGEMA_signal_2732), .Z1_f (new_AGEMA_signal_2733) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S11reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS12ser[2]), .A0_f (new_AGEMA_signal_2785), .A1_t (new_AGEMA_signal_2786), .A1_f (new_AGEMA_signal_2787), .B0_t (stateArray_outS12ser[2]), .B0_f (new_AGEMA_signal_2785), .B1_t (new_AGEMA_signal_2786), .B1_f (new_AGEMA_signal_2787), .Z0_t (stateArray_S11reg_gff_1_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_2788), .Z1_t (new_AGEMA_signal_2789), .Z1_f (new_AGEMA_signal_2790) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S11reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S11reg_gff_1_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_2788), .B1_t (new_AGEMA_signal_2789), .B1_f (new_AGEMA_signal_2790), .Z0_t (stateArray_S11reg_gff_1_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_6019), .Z1_t (new_AGEMA_signal_6020), .Z1_f (new_AGEMA_signal_6021) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S11reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (stateArray_S11reg_gff_1_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_6019), .A1_t (new_AGEMA_signal_6020), .A1_f (new_AGEMA_signal_6021), .B0_t (stateArray_outS12ser[2]), .B0_f (new_AGEMA_signal_2785), .B1_t (new_AGEMA_signal_2786), .B1_f (new_AGEMA_signal_2787), .Z0_t (stateArray_outS11ser[2]), .Z0_f (new_AGEMA_signal_2737), .Z1_t (new_AGEMA_signal_2738), .Z1_f (new_AGEMA_signal_2739) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S11reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS12ser[3]), .A0_f (new_AGEMA_signal_2791), .A1_t (new_AGEMA_signal_2792), .A1_f (new_AGEMA_signal_2793), .B0_t (stateArray_outS12ser[3]), .B0_f (new_AGEMA_signal_2791), .B1_t (new_AGEMA_signal_2792), .B1_f (new_AGEMA_signal_2793), .Z0_t (stateArray_S11reg_gff_1_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_2794), .Z1_t (new_AGEMA_signal_2795), .Z1_f (new_AGEMA_signal_2796) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S11reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S11reg_gff_1_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_2794), .B1_t (new_AGEMA_signal_2795), .B1_f (new_AGEMA_signal_2796), .Z0_t (stateArray_S11reg_gff_1_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_6022), .Z1_t (new_AGEMA_signal_6023), .Z1_f (new_AGEMA_signal_6024) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S11reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (stateArray_S11reg_gff_1_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_6022), .A1_t (new_AGEMA_signal_6023), .A1_f (new_AGEMA_signal_6024), .B0_t (stateArray_outS12ser[3]), .B0_f (new_AGEMA_signal_2791), .B1_t (new_AGEMA_signal_2792), .B1_f (new_AGEMA_signal_2793), .Z0_t (stateArray_outS11ser[3]), .Z0_f (new_AGEMA_signal_2743), .Z1_t (new_AGEMA_signal_2744), .Z1_f (new_AGEMA_signal_2745) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S11reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS12ser[4]), .A0_f (new_AGEMA_signal_2797), .A1_t (new_AGEMA_signal_2798), .A1_f (new_AGEMA_signal_2799), .B0_t (stateArray_outS12ser[4]), .B0_f (new_AGEMA_signal_2797), .B1_t (new_AGEMA_signal_2798), .B1_f (new_AGEMA_signal_2799), .Z0_t (stateArray_S11reg_gff_1_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_2800), .Z1_t (new_AGEMA_signal_2801), .Z1_f (new_AGEMA_signal_2802) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S11reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S11reg_gff_1_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_2800), .B1_t (new_AGEMA_signal_2801), .B1_f (new_AGEMA_signal_2802), .Z0_t (stateArray_S11reg_gff_1_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_6025), .Z1_t (new_AGEMA_signal_6026), .Z1_f (new_AGEMA_signal_6027) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S11reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (stateArray_S11reg_gff_1_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_6025), .A1_t (new_AGEMA_signal_6026), .A1_f (new_AGEMA_signal_6027), .B0_t (stateArray_outS12ser[4]), .B0_f (new_AGEMA_signal_2797), .B1_t (new_AGEMA_signal_2798), .B1_f (new_AGEMA_signal_2799), .Z0_t (stateArray_outS11ser[4]), .Z0_f (new_AGEMA_signal_2749), .Z1_t (new_AGEMA_signal_2750), .Z1_f (new_AGEMA_signal_2751) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S11reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS12ser[5]), .A0_f (new_AGEMA_signal_2803), .A1_t (new_AGEMA_signal_2804), .A1_f (new_AGEMA_signal_2805), .B0_t (stateArray_outS12ser[5]), .B0_f (new_AGEMA_signal_2803), .B1_t (new_AGEMA_signal_2804), .B1_f (new_AGEMA_signal_2805), .Z0_t (stateArray_S11reg_gff_1_SFF_5_MUXInst_X), .Z0_f (new_AGEMA_signal_2806), .Z1_t (new_AGEMA_signal_2807), .Z1_f (new_AGEMA_signal_2808) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S11reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S11reg_gff_1_SFF_5_MUXInst_X), .B0_f (new_AGEMA_signal_2806), .B1_t (new_AGEMA_signal_2807), .B1_f (new_AGEMA_signal_2808), .Z0_t (stateArray_S11reg_gff_1_SFF_5_MUXInst_Y), .Z0_f (new_AGEMA_signal_6028), .Z1_t (new_AGEMA_signal_6029), .Z1_f (new_AGEMA_signal_6030) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S11reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (stateArray_S11reg_gff_1_SFF_5_MUXInst_Y), .A0_f (new_AGEMA_signal_6028), .A1_t (new_AGEMA_signal_6029), .A1_f (new_AGEMA_signal_6030), .B0_t (stateArray_outS12ser[5]), .B0_f (new_AGEMA_signal_2803), .B1_t (new_AGEMA_signal_2804), .B1_f (new_AGEMA_signal_2805), .Z0_t (stateArray_outS11ser[5]), .Z0_f (new_AGEMA_signal_2755), .Z1_t (new_AGEMA_signal_2756), .Z1_f (new_AGEMA_signal_2757) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S11reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS12ser[6]), .A0_f (new_AGEMA_signal_2809), .A1_t (new_AGEMA_signal_2810), .A1_f (new_AGEMA_signal_2811), .B0_t (stateArray_outS12ser[6]), .B0_f (new_AGEMA_signal_2809), .B1_t (new_AGEMA_signal_2810), .B1_f (new_AGEMA_signal_2811), .Z0_t (stateArray_S11reg_gff_1_SFF_6_MUXInst_X), .Z0_f (new_AGEMA_signal_2812), .Z1_t (new_AGEMA_signal_2813), .Z1_f (new_AGEMA_signal_2814) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S11reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S11reg_gff_1_SFF_6_MUXInst_X), .B0_f (new_AGEMA_signal_2812), .B1_t (new_AGEMA_signal_2813), .B1_f (new_AGEMA_signal_2814), .Z0_t (stateArray_S11reg_gff_1_SFF_6_MUXInst_Y), .Z0_f (new_AGEMA_signal_6031), .Z1_t (new_AGEMA_signal_6032), .Z1_f (new_AGEMA_signal_6033) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S11reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (stateArray_S11reg_gff_1_SFF_6_MUXInst_Y), .A0_f (new_AGEMA_signal_6031), .A1_t (new_AGEMA_signal_6032), .A1_f (new_AGEMA_signal_6033), .B0_t (stateArray_outS12ser[6]), .B0_f (new_AGEMA_signal_2809), .B1_t (new_AGEMA_signal_2810), .B1_f (new_AGEMA_signal_2811), .Z0_t (stateArray_outS11ser[6]), .Z0_f (new_AGEMA_signal_2761), .Z1_t (new_AGEMA_signal_2762), .Z1_f (new_AGEMA_signal_2763) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S11reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS12ser[7]), .A0_f (new_AGEMA_signal_2815), .A1_t (new_AGEMA_signal_2816), .A1_f (new_AGEMA_signal_2817), .B0_t (stateArray_outS12ser[7]), .B0_f (new_AGEMA_signal_2815), .B1_t (new_AGEMA_signal_2816), .B1_f (new_AGEMA_signal_2817), .Z0_t (stateArray_S11reg_gff_1_SFF_7_MUXInst_X), .Z0_f (new_AGEMA_signal_2818), .Z1_t (new_AGEMA_signal_2819), .Z1_f (new_AGEMA_signal_2820) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S11reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S11reg_gff_1_SFF_7_MUXInst_X), .B0_f (new_AGEMA_signal_2818), .B1_t (new_AGEMA_signal_2819), .B1_f (new_AGEMA_signal_2820), .Z0_t (stateArray_S11reg_gff_1_SFF_7_MUXInst_Y), .Z0_f (new_AGEMA_signal_6034), .Z1_t (new_AGEMA_signal_6035), .Z1_f (new_AGEMA_signal_6036) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S11reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (stateArray_S11reg_gff_1_SFF_7_MUXInst_Y), .A0_f (new_AGEMA_signal_6034), .A1_t (new_AGEMA_signal_6035), .A1_f (new_AGEMA_signal_6036), .B0_t (stateArray_outS12ser[7]), .B0_f (new_AGEMA_signal_2815), .B1_t (new_AGEMA_signal_2816), .B1_f (new_AGEMA_signal_2817), .Z0_t (stateArray_outS11ser[7]), .Z0_f (new_AGEMA_signal_2767), .Z1_t (new_AGEMA_signal_2768), .Z1_f (new_AGEMA_signal_2769) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S12reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS13ser[0]), .A0_f (new_AGEMA_signal_2821), .A1_t (new_AGEMA_signal_2822), .A1_f (new_AGEMA_signal_2823), .B0_t (stateArray_outS13ser[0]), .B0_f (new_AGEMA_signal_2821), .B1_t (new_AGEMA_signal_2822), .B1_f (new_AGEMA_signal_2823), .Z0_t (stateArray_S12reg_gff_1_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_2824), .Z1_t (new_AGEMA_signal_2825), .Z1_f (new_AGEMA_signal_2826) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S12reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S12reg_gff_1_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_2824), .B1_t (new_AGEMA_signal_2825), .B1_f (new_AGEMA_signal_2826), .Z0_t (stateArray_S12reg_gff_1_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_6037), .Z1_t (new_AGEMA_signal_6038), .Z1_f (new_AGEMA_signal_6039) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S12reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (stateArray_S12reg_gff_1_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_6037), .A1_t (new_AGEMA_signal_6038), .A1_f (new_AGEMA_signal_6039), .B0_t (stateArray_outS13ser[0]), .B0_f (new_AGEMA_signal_2821), .B1_t (new_AGEMA_signal_2822), .B1_f (new_AGEMA_signal_2823), .Z0_t (stateArray_outS12ser[0]), .Z0_f (new_AGEMA_signal_2773), .Z1_t (new_AGEMA_signal_2774), .Z1_f (new_AGEMA_signal_2775) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S12reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS13ser[1]), .A0_f (new_AGEMA_signal_2827), .A1_t (new_AGEMA_signal_2828), .A1_f (new_AGEMA_signal_2829), .B0_t (stateArray_outS13ser[1]), .B0_f (new_AGEMA_signal_2827), .B1_t (new_AGEMA_signal_2828), .B1_f (new_AGEMA_signal_2829), .Z0_t (stateArray_S12reg_gff_1_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_2830), .Z1_t (new_AGEMA_signal_2831), .Z1_f (new_AGEMA_signal_2832) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S12reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S12reg_gff_1_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_2830), .B1_t (new_AGEMA_signal_2831), .B1_f (new_AGEMA_signal_2832), .Z0_t (stateArray_S12reg_gff_1_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_6040), .Z1_t (new_AGEMA_signal_6041), .Z1_f (new_AGEMA_signal_6042) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S12reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (stateArray_S12reg_gff_1_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_6040), .A1_t (new_AGEMA_signal_6041), .A1_f (new_AGEMA_signal_6042), .B0_t (stateArray_outS13ser[1]), .B0_f (new_AGEMA_signal_2827), .B1_t (new_AGEMA_signal_2828), .B1_f (new_AGEMA_signal_2829), .Z0_t (stateArray_outS12ser[1]), .Z0_f (new_AGEMA_signal_2779), .Z1_t (new_AGEMA_signal_2780), .Z1_f (new_AGEMA_signal_2781) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S12reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS13ser[2]), .A0_f (new_AGEMA_signal_2833), .A1_t (new_AGEMA_signal_2834), .A1_f (new_AGEMA_signal_2835), .B0_t (stateArray_outS13ser[2]), .B0_f (new_AGEMA_signal_2833), .B1_t (new_AGEMA_signal_2834), .B1_f (new_AGEMA_signal_2835), .Z0_t (stateArray_S12reg_gff_1_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_2836), .Z1_t (new_AGEMA_signal_2837), .Z1_f (new_AGEMA_signal_2838) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S12reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S12reg_gff_1_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_2836), .B1_t (new_AGEMA_signal_2837), .B1_f (new_AGEMA_signal_2838), .Z0_t (stateArray_S12reg_gff_1_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_6043), .Z1_t (new_AGEMA_signal_6044), .Z1_f (new_AGEMA_signal_6045) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S12reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (stateArray_S12reg_gff_1_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_6043), .A1_t (new_AGEMA_signal_6044), .A1_f (new_AGEMA_signal_6045), .B0_t (stateArray_outS13ser[2]), .B0_f (new_AGEMA_signal_2833), .B1_t (new_AGEMA_signal_2834), .B1_f (new_AGEMA_signal_2835), .Z0_t (stateArray_outS12ser[2]), .Z0_f (new_AGEMA_signal_2785), .Z1_t (new_AGEMA_signal_2786), .Z1_f (new_AGEMA_signal_2787) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S12reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS13ser[3]), .A0_f (new_AGEMA_signal_2839), .A1_t (new_AGEMA_signal_2840), .A1_f (new_AGEMA_signal_2841), .B0_t (stateArray_outS13ser[3]), .B0_f (new_AGEMA_signal_2839), .B1_t (new_AGEMA_signal_2840), .B1_f (new_AGEMA_signal_2841), .Z0_t (stateArray_S12reg_gff_1_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_2842), .Z1_t (new_AGEMA_signal_2843), .Z1_f (new_AGEMA_signal_2844) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S12reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S12reg_gff_1_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_2842), .B1_t (new_AGEMA_signal_2843), .B1_f (new_AGEMA_signal_2844), .Z0_t (stateArray_S12reg_gff_1_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_6046), .Z1_t (new_AGEMA_signal_6047), .Z1_f (new_AGEMA_signal_6048) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S12reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (stateArray_S12reg_gff_1_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_6046), .A1_t (new_AGEMA_signal_6047), .A1_f (new_AGEMA_signal_6048), .B0_t (stateArray_outS13ser[3]), .B0_f (new_AGEMA_signal_2839), .B1_t (new_AGEMA_signal_2840), .B1_f (new_AGEMA_signal_2841), .Z0_t (stateArray_outS12ser[3]), .Z0_f (new_AGEMA_signal_2791), .Z1_t (new_AGEMA_signal_2792), .Z1_f (new_AGEMA_signal_2793) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S12reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS13ser[4]), .A0_f (new_AGEMA_signal_2845), .A1_t (new_AGEMA_signal_2846), .A1_f (new_AGEMA_signal_2847), .B0_t (stateArray_outS13ser[4]), .B0_f (new_AGEMA_signal_2845), .B1_t (new_AGEMA_signal_2846), .B1_f (new_AGEMA_signal_2847), .Z0_t (stateArray_S12reg_gff_1_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_2848), .Z1_t (new_AGEMA_signal_2849), .Z1_f (new_AGEMA_signal_2850) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S12reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S12reg_gff_1_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_2848), .B1_t (new_AGEMA_signal_2849), .B1_f (new_AGEMA_signal_2850), .Z0_t (stateArray_S12reg_gff_1_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_6049), .Z1_t (new_AGEMA_signal_6050), .Z1_f (new_AGEMA_signal_6051) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S12reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (stateArray_S12reg_gff_1_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_6049), .A1_t (new_AGEMA_signal_6050), .A1_f (new_AGEMA_signal_6051), .B0_t (stateArray_outS13ser[4]), .B0_f (new_AGEMA_signal_2845), .B1_t (new_AGEMA_signal_2846), .B1_f (new_AGEMA_signal_2847), .Z0_t (stateArray_outS12ser[4]), .Z0_f (new_AGEMA_signal_2797), .Z1_t (new_AGEMA_signal_2798), .Z1_f (new_AGEMA_signal_2799) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S12reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS13ser[5]), .A0_f (new_AGEMA_signal_2851), .A1_t (new_AGEMA_signal_2852), .A1_f (new_AGEMA_signal_2853), .B0_t (stateArray_outS13ser[5]), .B0_f (new_AGEMA_signal_2851), .B1_t (new_AGEMA_signal_2852), .B1_f (new_AGEMA_signal_2853), .Z0_t (stateArray_S12reg_gff_1_SFF_5_MUXInst_X), .Z0_f (new_AGEMA_signal_2854), .Z1_t (new_AGEMA_signal_2855), .Z1_f (new_AGEMA_signal_2856) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S12reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S12reg_gff_1_SFF_5_MUXInst_X), .B0_f (new_AGEMA_signal_2854), .B1_t (new_AGEMA_signal_2855), .B1_f (new_AGEMA_signal_2856), .Z0_t (stateArray_S12reg_gff_1_SFF_5_MUXInst_Y), .Z0_f (new_AGEMA_signal_6052), .Z1_t (new_AGEMA_signal_6053), .Z1_f (new_AGEMA_signal_6054) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S12reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (stateArray_S12reg_gff_1_SFF_5_MUXInst_Y), .A0_f (new_AGEMA_signal_6052), .A1_t (new_AGEMA_signal_6053), .A1_f (new_AGEMA_signal_6054), .B0_t (stateArray_outS13ser[5]), .B0_f (new_AGEMA_signal_2851), .B1_t (new_AGEMA_signal_2852), .B1_f (new_AGEMA_signal_2853), .Z0_t (stateArray_outS12ser[5]), .Z0_f (new_AGEMA_signal_2803), .Z1_t (new_AGEMA_signal_2804), .Z1_f (new_AGEMA_signal_2805) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S12reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS13ser[6]), .A0_f (new_AGEMA_signal_2857), .A1_t (new_AGEMA_signal_2858), .A1_f (new_AGEMA_signal_2859), .B0_t (stateArray_outS13ser[6]), .B0_f (new_AGEMA_signal_2857), .B1_t (new_AGEMA_signal_2858), .B1_f (new_AGEMA_signal_2859), .Z0_t (stateArray_S12reg_gff_1_SFF_6_MUXInst_X), .Z0_f (new_AGEMA_signal_2860), .Z1_t (new_AGEMA_signal_2861), .Z1_f (new_AGEMA_signal_2862) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S12reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S12reg_gff_1_SFF_6_MUXInst_X), .B0_f (new_AGEMA_signal_2860), .B1_t (new_AGEMA_signal_2861), .B1_f (new_AGEMA_signal_2862), .Z0_t (stateArray_S12reg_gff_1_SFF_6_MUXInst_Y), .Z0_f (new_AGEMA_signal_6055), .Z1_t (new_AGEMA_signal_6056), .Z1_f (new_AGEMA_signal_6057) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S12reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (stateArray_S12reg_gff_1_SFF_6_MUXInst_Y), .A0_f (new_AGEMA_signal_6055), .A1_t (new_AGEMA_signal_6056), .A1_f (new_AGEMA_signal_6057), .B0_t (stateArray_outS13ser[6]), .B0_f (new_AGEMA_signal_2857), .B1_t (new_AGEMA_signal_2858), .B1_f (new_AGEMA_signal_2859), .Z0_t (stateArray_outS12ser[6]), .Z0_f (new_AGEMA_signal_2809), .Z1_t (new_AGEMA_signal_2810), .Z1_f (new_AGEMA_signal_2811) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S12reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS13ser[7]), .A0_f (new_AGEMA_signal_2863), .A1_t (new_AGEMA_signal_2864), .A1_f (new_AGEMA_signal_2865), .B0_t (stateArray_outS13ser[7]), .B0_f (new_AGEMA_signal_2863), .B1_t (new_AGEMA_signal_2864), .B1_f (new_AGEMA_signal_2865), .Z0_t (stateArray_S12reg_gff_1_SFF_7_MUXInst_X), .Z0_f (new_AGEMA_signal_2866), .Z1_t (new_AGEMA_signal_2867), .Z1_f (new_AGEMA_signal_2868) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S12reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S12reg_gff_1_SFF_7_MUXInst_X), .B0_f (new_AGEMA_signal_2866), .B1_t (new_AGEMA_signal_2867), .B1_f (new_AGEMA_signal_2868), .Z0_t (stateArray_S12reg_gff_1_SFF_7_MUXInst_Y), .Z0_f (new_AGEMA_signal_6058), .Z1_t (new_AGEMA_signal_6059), .Z1_f (new_AGEMA_signal_6060) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S12reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (stateArray_S12reg_gff_1_SFF_7_MUXInst_Y), .A0_f (new_AGEMA_signal_6058), .A1_t (new_AGEMA_signal_6059), .A1_f (new_AGEMA_signal_6060), .B0_t (stateArray_outS13ser[7]), .B0_f (new_AGEMA_signal_2863), .B1_t (new_AGEMA_signal_2864), .B1_f (new_AGEMA_signal_2865), .Z0_t (stateArray_outS12ser[7]), .Z0_f (new_AGEMA_signal_2815), .Z1_t (new_AGEMA_signal_2816), .Z1_f (new_AGEMA_signal_2817) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S13reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS13ser[0]), .A0_f (new_AGEMA_signal_6229), .A1_t (new_AGEMA_signal_6230), .A1_f (new_AGEMA_signal_6231), .B0_t (MCin[16]), .B0_f (new_AGEMA_signal_3988), .B1_t (new_AGEMA_signal_3989), .B1_f (new_AGEMA_signal_3990), .Z0_t (stateArray_S13reg_gff_1_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_6334), .Z1_t (new_AGEMA_signal_6335), .Z1_f (new_AGEMA_signal_6336) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S13reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S13reg_gff_1_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_6334), .B1_t (new_AGEMA_signal_6335), .B1_f (new_AGEMA_signal_6336), .Z0_t (stateArray_S13reg_gff_1_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_7182), .Z1_t (new_AGEMA_signal_7183), .Z1_f (new_AGEMA_signal_7184) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S13reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (stateArray_S13reg_gff_1_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_7182), .A1_t (new_AGEMA_signal_7183), .A1_f (new_AGEMA_signal_7184), .B0_t (stateArray_inS13ser[0]), .B0_f (new_AGEMA_signal_6229), .B1_t (new_AGEMA_signal_6230), .B1_f (new_AGEMA_signal_6231), .Z0_t (stateArray_outS13ser[0]), .Z0_f (new_AGEMA_signal_2821), .Z1_t (new_AGEMA_signal_2822), .Z1_f (new_AGEMA_signal_2823) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S13reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS13ser[1]), .A0_f (new_AGEMA_signal_6373), .A1_t (new_AGEMA_signal_6374), .A1_f (new_AGEMA_signal_6375), .B0_t (MixColumns_line1_S02[2]), .B0_f (new_AGEMA_signal_3982), .B1_t (new_AGEMA_signal_3983), .B1_f (new_AGEMA_signal_3984), .Z0_t (stateArray_S13reg_gff_1_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_7185), .Z1_t (new_AGEMA_signal_7186), .Z1_f (new_AGEMA_signal_7187) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S13reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S13reg_gff_1_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_7185), .B1_t (new_AGEMA_signal_7186), .B1_f (new_AGEMA_signal_7187), .Z0_t (stateArray_S13reg_gff_1_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_7283), .Z1_t (new_AGEMA_signal_7284), .Z1_f (new_AGEMA_signal_7285) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S13reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (stateArray_S13reg_gff_1_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_7283), .A1_t (new_AGEMA_signal_7284), .A1_f (new_AGEMA_signal_7285), .B0_t (stateArray_inS13ser[1]), .B0_f (new_AGEMA_signal_6373), .B1_t (new_AGEMA_signal_6374), .B1_f (new_AGEMA_signal_6375), .Z0_t (stateArray_outS13ser[1]), .Z0_f (new_AGEMA_signal_2827), .Z1_t (new_AGEMA_signal_2828), .Z1_f (new_AGEMA_signal_2829) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S13reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS13ser[2]), .A0_f (new_AGEMA_signal_6235), .A1_t (new_AGEMA_signal_6236), .A1_f (new_AGEMA_signal_6237), .B0_t (MCin[18]), .B0_f (new_AGEMA_signal_3979), .B1_t (new_AGEMA_signal_3980), .B1_f (new_AGEMA_signal_3981), .Z0_t (stateArray_S13reg_gff_1_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_6337), .Z1_t (new_AGEMA_signal_6338), .Z1_f (new_AGEMA_signal_6339) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S13reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S13reg_gff_1_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_6337), .B1_t (new_AGEMA_signal_6338), .B1_f (new_AGEMA_signal_6339), .Z0_t (stateArray_S13reg_gff_1_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_7188), .Z1_t (new_AGEMA_signal_7189), .Z1_f (new_AGEMA_signal_7190) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S13reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (stateArray_S13reg_gff_1_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_7188), .A1_t (new_AGEMA_signal_7189), .A1_f (new_AGEMA_signal_7190), .B0_t (stateArray_inS13ser[2]), .B0_f (new_AGEMA_signal_6235), .B1_t (new_AGEMA_signal_6236), .B1_f (new_AGEMA_signal_6237), .Z0_t (stateArray_outS13ser[2]), .Z0_f (new_AGEMA_signal_2833), .Z1_t (new_AGEMA_signal_2834), .Z1_f (new_AGEMA_signal_2835) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S13reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS13ser[3]), .A0_f (new_AGEMA_signal_6376), .A1_t (new_AGEMA_signal_6377), .A1_f (new_AGEMA_signal_6378), .B0_t (MCin[19]), .B0_f (new_AGEMA_signal_3994), .B1_t (new_AGEMA_signal_3995), .B1_f (new_AGEMA_signal_3996), .Z0_t (stateArray_S13reg_gff_1_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_7191), .Z1_t (new_AGEMA_signal_7192), .Z1_f (new_AGEMA_signal_7193) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S13reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S13reg_gff_1_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_7191), .B1_t (new_AGEMA_signal_7192), .B1_f (new_AGEMA_signal_7193), .Z0_t (stateArray_S13reg_gff_1_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_7286), .Z1_t (new_AGEMA_signal_7287), .Z1_f (new_AGEMA_signal_7288) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S13reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (stateArray_S13reg_gff_1_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_7286), .A1_t (new_AGEMA_signal_7287), .A1_f (new_AGEMA_signal_7288), .B0_t (stateArray_inS13ser[3]), .B0_f (new_AGEMA_signal_6376), .B1_t (new_AGEMA_signal_6377), .B1_f (new_AGEMA_signal_6378), .Z0_t (stateArray_outS13ser[3]), .Z0_f (new_AGEMA_signal_2839), .Z1_t (new_AGEMA_signal_2840), .Z1_f (new_AGEMA_signal_2841) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S13reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS13ser[4]), .A0_f (new_AGEMA_signal_6379), .A1_t (new_AGEMA_signal_6380), .A1_f (new_AGEMA_signal_6381), .B0_t (MixColumns_line1_S02[5]), .B0_f (new_AGEMA_signal_3973), .B1_t (new_AGEMA_signal_3974), .B1_f (new_AGEMA_signal_3975), .Z0_t (stateArray_S13reg_gff_1_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_7194), .Z1_t (new_AGEMA_signal_7195), .Z1_f (new_AGEMA_signal_7196) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S13reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S13reg_gff_1_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_7194), .B1_t (new_AGEMA_signal_7195), .B1_f (new_AGEMA_signal_7196), .Z0_t (stateArray_S13reg_gff_1_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_7289), .Z1_t (new_AGEMA_signal_7290), .Z1_f (new_AGEMA_signal_7291) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S13reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (stateArray_S13reg_gff_1_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_7289), .A1_t (new_AGEMA_signal_7290), .A1_f (new_AGEMA_signal_7291), .B0_t (stateArray_inS13ser[4]), .B0_f (new_AGEMA_signal_6379), .B1_t (new_AGEMA_signal_6380), .B1_f (new_AGEMA_signal_6381), .Z0_t (stateArray_outS13ser[4]), .Z0_f (new_AGEMA_signal_2845), .Z1_t (new_AGEMA_signal_2846), .Z1_f (new_AGEMA_signal_2847) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S13reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS13ser[5]), .A0_f (new_AGEMA_signal_6244), .A1_t (new_AGEMA_signal_6245), .A1_f (new_AGEMA_signal_6246), .B0_t (MixColumns_line1_S02[6]), .B0_f (new_AGEMA_signal_3967), .B1_t (new_AGEMA_signal_3968), .B1_f (new_AGEMA_signal_3969), .Z0_t (stateArray_S13reg_gff_1_SFF_5_MUXInst_X), .Z0_f (new_AGEMA_signal_6340), .Z1_t (new_AGEMA_signal_6341), .Z1_f (new_AGEMA_signal_6342) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S13reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S13reg_gff_1_SFF_5_MUXInst_X), .B0_f (new_AGEMA_signal_6340), .B1_t (new_AGEMA_signal_6341), .B1_f (new_AGEMA_signal_6342), .Z0_t (stateArray_S13reg_gff_1_SFF_5_MUXInst_Y), .Z0_f (new_AGEMA_signal_7197), .Z1_t (new_AGEMA_signal_7198), .Z1_f (new_AGEMA_signal_7199) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S13reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (stateArray_S13reg_gff_1_SFF_5_MUXInst_Y), .A0_f (new_AGEMA_signal_7197), .A1_t (new_AGEMA_signal_7198), .A1_f (new_AGEMA_signal_7199), .B0_t (stateArray_inS13ser[5]), .B0_f (new_AGEMA_signal_6244), .B1_t (new_AGEMA_signal_6245), .B1_f (new_AGEMA_signal_6246), .Z0_t (stateArray_outS13ser[5]), .Z0_f (new_AGEMA_signal_2851), .Z1_t (new_AGEMA_signal_2852), .Z1_f (new_AGEMA_signal_2853) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S13reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS13ser[6]), .A0_f (new_AGEMA_signal_6247), .A1_t (new_AGEMA_signal_6248), .A1_f (new_AGEMA_signal_6249), .B0_t (MixColumns_line1_S02[7]), .B0_f (new_AGEMA_signal_3961), .B1_t (new_AGEMA_signal_3962), .B1_f (new_AGEMA_signal_3963), .Z0_t (stateArray_S13reg_gff_1_SFF_6_MUXInst_X), .Z0_f (new_AGEMA_signal_6343), .Z1_t (new_AGEMA_signal_6344), .Z1_f (new_AGEMA_signal_6345) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S13reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S13reg_gff_1_SFF_6_MUXInst_X), .B0_f (new_AGEMA_signal_6343), .B1_t (new_AGEMA_signal_6344), .B1_f (new_AGEMA_signal_6345), .Z0_t (stateArray_S13reg_gff_1_SFF_6_MUXInst_Y), .Z0_f (new_AGEMA_signal_7200), .Z1_t (new_AGEMA_signal_7201), .Z1_f (new_AGEMA_signal_7202) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S13reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (stateArray_S13reg_gff_1_SFF_6_MUXInst_Y), .A0_f (new_AGEMA_signal_7200), .A1_t (new_AGEMA_signal_7201), .A1_f (new_AGEMA_signal_7202), .B0_t (stateArray_inS13ser[6]), .B0_f (new_AGEMA_signal_6247), .B1_t (new_AGEMA_signal_6248), .B1_f (new_AGEMA_signal_6249), .Z0_t (stateArray_outS13ser[6]), .Z0_f (new_AGEMA_signal_2857), .Z1_t (new_AGEMA_signal_2858), .Z1_f (new_AGEMA_signal_2859) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S13reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS13ser[7]), .A0_f (new_AGEMA_signal_6250), .A1_t (new_AGEMA_signal_6251), .A1_f (new_AGEMA_signal_6252), .B0_t (MixColumns_line1_S02[0]), .B0_f (new_AGEMA_signal_3958), .B1_t (new_AGEMA_signal_3959), .B1_f (new_AGEMA_signal_3960), .Z0_t (stateArray_S13reg_gff_1_SFF_7_MUXInst_X), .Z0_f (new_AGEMA_signal_6346), .Z1_t (new_AGEMA_signal_6347), .Z1_f (new_AGEMA_signal_6348) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S13reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S13reg_gff_1_SFF_7_MUXInst_X), .B0_f (new_AGEMA_signal_6346), .B1_t (new_AGEMA_signal_6347), .B1_f (new_AGEMA_signal_6348), .Z0_t (stateArray_S13reg_gff_1_SFF_7_MUXInst_Y), .Z0_f (new_AGEMA_signal_7203), .Z1_t (new_AGEMA_signal_7204), .Z1_f (new_AGEMA_signal_7205) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S13reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (stateArray_S13reg_gff_1_SFF_7_MUXInst_Y), .A0_f (new_AGEMA_signal_7203), .A1_t (new_AGEMA_signal_7204), .A1_f (new_AGEMA_signal_7205), .B0_t (stateArray_inS13ser[7]), .B0_f (new_AGEMA_signal_6250), .B1_t (new_AGEMA_signal_6251), .B1_f (new_AGEMA_signal_6252), .Z0_t (stateArray_outS13ser[7]), .Z0_f (new_AGEMA_signal_2863), .Z1_t (new_AGEMA_signal_2864), .Z1_f (new_AGEMA_signal_2865) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S20reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS21ser[0]), .A0_f (new_AGEMA_signal_2869), .A1_t (new_AGEMA_signal_2870), .A1_f (new_AGEMA_signal_2871), .B0_t (stateArray_outS22ser[0]), .B0_f (new_AGEMA_signal_2872), .B1_t (new_AGEMA_signal_2873), .B1_f (new_AGEMA_signal_2874), .Z0_t (stateArray_S20reg_gff_1_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_2875), .Z1_t (new_AGEMA_signal_2876), .Z1_f (new_AGEMA_signal_2877) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S20reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S20reg_gff_1_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_2875), .B1_t (new_AGEMA_signal_2876), .B1_f (new_AGEMA_signal_2877), .Z0_t (stateArray_S20reg_gff_1_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_6061), .Z1_t (new_AGEMA_signal_6062), .Z1_f (new_AGEMA_signal_6063) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S20reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (stateArray_S20reg_gff_1_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_6061), .A1_t (new_AGEMA_signal_6062), .A1_f (new_AGEMA_signal_6063), .B0_t (stateArray_outS21ser[0]), .B0_f (new_AGEMA_signal_2869), .B1_t (new_AGEMA_signal_2870), .B1_f (new_AGEMA_signal_2871), .Z0_t (MCin[8]), .Z0_f (new_AGEMA_signal_2989), .Z1_t (new_AGEMA_signal_2990), .Z1_f (new_AGEMA_signal_2991) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S20reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS21ser[1]), .A0_f (new_AGEMA_signal_2878), .A1_t (new_AGEMA_signal_2879), .A1_f (new_AGEMA_signal_2880), .B0_t (stateArray_outS22ser[1]), .B0_f (new_AGEMA_signal_2881), .B1_t (new_AGEMA_signal_2882), .B1_f (new_AGEMA_signal_2883), .Z0_t (stateArray_S20reg_gff_1_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_2884), .Z1_t (new_AGEMA_signal_2885), .Z1_f (new_AGEMA_signal_2886) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S20reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S20reg_gff_1_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_2884), .B1_t (new_AGEMA_signal_2885), .B1_f (new_AGEMA_signal_2886), .Z0_t (stateArray_S20reg_gff_1_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_6064), .Z1_t (new_AGEMA_signal_6065), .Z1_f (new_AGEMA_signal_6066) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S20reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (stateArray_S20reg_gff_1_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_6064), .A1_t (new_AGEMA_signal_6065), .A1_f (new_AGEMA_signal_6066), .B0_t (stateArray_outS21ser[1]), .B0_f (new_AGEMA_signal_2878), .B1_t (new_AGEMA_signal_2879), .B1_f (new_AGEMA_signal_2880), .Z0_t (MixColumns_line2_S02[2]), .Z0_f (new_AGEMA_signal_2995), .Z1_t (new_AGEMA_signal_2996), .Z1_f (new_AGEMA_signal_2997) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S20reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS21ser[2]), .A0_f (new_AGEMA_signal_2887), .A1_t (new_AGEMA_signal_2888), .A1_f (new_AGEMA_signal_2889), .B0_t (stateArray_outS22ser[2]), .B0_f (new_AGEMA_signal_2890), .B1_t (new_AGEMA_signal_2891), .B1_f (new_AGEMA_signal_2892), .Z0_t (stateArray_S20reg_gff_1_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_2893), .Z1_t (new_AGEMA_signal_2894), .Z1_f (new_AGEMA_signal_2895) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S20reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S20reg_gff_1_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_2893), .B1_t (new_AGEMA_signal_2894), .B1_f (new_AGEMA_signal_2895), .Z0_t (stateArray_S20reg_gff_1_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_6067), .Z1_t (new_AGEMA_signal_6068), .Z1_f (new_AGEMA_signal_6069) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S20reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (stateArray_S20reg_gff_1_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_6067), .A1_t (new_AGEMA_signal_6068), .A1_f (new_AGEMA_signal_6069), .B0_t (stateArray_outS21ser[2]), .B0_f (new_AGEMA_signal_2887), .B1_t (new_AGEMA_signal_2888), .B1_f (new_AGEMA_signal_2889), .Z0_t (MCin[10]), .Z0_f (new_AGEMA_signal_3001), .Z1_t (new_AGEMA_signal_3002), .Z1_f (new_AGEMA_signal_3003) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S20reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS21ser[3]), .A0_f (new_AGEMA_signal_2896), .A1_t (new_AGEMA_signal_2897), .A1_f (new_AGEMA_signal_2898), .B0_t (stateArray_outS22ser[3]), .B0_f (new_AGEMA_signal_2899), .B1_t (new_AGEMA_signal_2900), .B1_f (new_AGEMA_signal_2901), .Z0_t (stateArray_S20reg_gff_1_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_2902), .Z1_t (new_AGEMA_signal_2903), .Z1_f (new_AGEMA_signal_2904) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S20reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S20reg_gff_1_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_2902), .B1_t (new_AGEMA_signal_2903), .B1_f (new_AGEMA_signal_2904), .Z0_t (stateArray_S20reg_gff_1_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_6070), .Z1_t (new_AGEMA_signal_6071), .Z1_f (new_AGEMA_signal_6072) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S20reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (stateArray_S20reg_gff_1_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_6070), .A1_t (new_AGEMA_signal_6071), .A1_f (new_AGEMA_signal_6072), .B0_t (stateArray_outS21ser[3]), .B0_f (new_AGEMA_signal_2896), .B1_t (new_AGEMA_signal_2897), .B1_f (new_AGEMA_signal_2898), .Z0_t (MCin[11]), .Z0_f (new_AGEMA_signal_3007), .Z1_t (new_AGEMA_signal_3008), .Z1_f (new_AGEMA_signal_3009) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S20reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS21ser[4]), .A0_f (new_AGEMA_signal_2905), .A1_t (new_AGEMA_signal_2906), .A1_f (new_AGEMA_signal_2907), .B0_t (stateArray_outS22ser[4]), .B0_f (new_AGEMA_signal_2908), .B1_t (new_AGEMA_signal_2909), .B1_f (new_AGEMA_signal_2910), .Z0_t (stateArray_S20reg_gff_1_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_2911), .Z1_t (new_AGEMA_signal_2912), .Z1_f (new_AGEMA_signal_2913) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S20reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S20reg_gff_1_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_2911), .B1_t (new_AGEMA_signal_2912), .B1_f (new_AGEMA_signal_2913), .Z0_t (stateArray_S20reg_gff_1_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_6073), .Z1_t (new_AGEMA_signal_6074), .Z1_f (new_AGEMA_signal_6075) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S20reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (stateArray_S20reg_gff_1_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_6073), .A1_t (new_AGEMA_signal_6074), .A1_f (new_AGEMA_signal_6075), .B0_t (stateArray_outS21ser[4]), .B0_f (new_AGEMA_signal_2905), .B1_t (new_AGEMA_signal_2906), .B1_f (new_AGEMA_signal_2907), .Z0_t (MixColumns_line2_S02[5]), .Z0_f (new_AGEMA_signal_3013), .Z1_t (new_AGEMA_signal_3014), .Z1_f (new_AGEMA_signal_3015) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S20reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS21ser[5]), .A0_f (new_AGEMA_signal_2914), .A1_t (new_AGEMA_signal_2915), .A1_f (new_AGEMA_signal_2916), .B0_t (stateArray_outS22ser[5]), .B0_f (new_AGEMA_signal_2917), .B1_t (new_AGEMA_signal_2918), .B1_f (new_AGEMA_signal_2919), .Z0_t (stateArray_S20reg_gff_1_SFF_5_MUXInst_X), .Z0_f (new_AGEMA_signal_2920), .Z1_t (new_AGEMA_signal_2921), .Z1_f (new_AGEMA_signal_2922) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S20reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S20reg_gff_1_SFF_5_MUXInst_X), .B0_f (new_AGEMA_signal_2920), .B1_t (new_AGEMA_signal_2921), .B1_f (new_AGEMA_signal_2922), .Z0_t (stateArray_S20reg_gff_1_SFF_5_MUXInst_Y), .Z0_f (new_AGEMA_signal_6076), .Z1_t (new_AGEMA_signal_6077), .Z1_f (new_AGEMA_signal_6078) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S20reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (stateArray_S20reg_gff_1_SFF_5_MUXInst_Y), .A0_f (new_AGEMA_signal_6076), .A1_t (new_AGEMA_signal_6077), .A1_f (new_AGEMA_signal_6078), .B0_t (stateArray_outS21ser[5]), .B0_f (new_AGEMA_signal_2914), .B1_t (new_AGEMA_signal_2915), .B1_f (new_AGEMA_signal_2916), .Z0_t (MixColumns_line2_S02[6]), .Z0_f (new_AGEMA_signal_3019), .Z1_t (new_AGEMA_signal_3020), .Z1_f (new_AGEMA_signal_3021) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S20reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS21ser[6]), .A0_f (new_AGEMA_signal_2923), .A1_t (new_AGEMA_signal_2924), .A1_f (new_AGEMA_signal_2925), .B0_t (stateArray_outS22ser[6]), .B0_f (new_AGEMA_signal_2926), .B1_t (new_AGEMA_signal_2927), .B1_f (new_AGEMA_signal_2928), .Z0_t (stateArray_S20reg_gff_1_SFF_6_MUXInst_X), .Z0_f (new_AGEMA_signal_2929), .Z1_t (new_AGEMA_signal_2930), .Z1_f (new_AGEMA_signal_2931) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S20reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S20reg_gff_1_SFF_6_MUXInst_X), .B0_f (new_AGEMA_signal_2929), .B1_t (new_AGEMA_signal_2930), .B1_f (new_AGEMA_signal_2931), .Z0_t (stateArray_S20reg_gff_1_SFF_6_MUXInst_Y), .Z0_f (new_AGEMA_signal_6079), .Z1_t (new_AGEMA_signal_6080), .Z1_f (new_AGEMA_signal_6081) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S20reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (stateArray_S20reg_gff_1_SFF_6_MUXInst_Y), .A0_f (new_AGEMA_signal_6079), .A1_t (new_AGEMA_signal_6080), .A1_f (new_AGEMA_signal_6081), .B0_t (stateArray_outS21ser[6]), .B0_f (new_AGEMA_signal_2923), .B1_t (new_AGEMA_signal_2924), .B1_f (new_AGEMA_signal_2925), .Z0_t (MixColumns_line2_S02[7]), .Z0_f (new_AGEMA_signal_3025), .Z1_t (new_AGEMA_signal_3026), .Z1_f (new_AGEMA_signal_3027) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S20reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS21ser[7]), .A0_f (new_AGEMA_signal_2932), .A1_t (new_AGEMA_signal_2933), .A1_f (new_AGEMA_signal_2934), .B0_t (stateArray_outS22ser[7]), .B0_f (new_AGEMA_signal_2935), .B1_t (new_AGEMA_signal_2936), .B1_f (new_AGEMA_signal_2937), .Z0_t (stateArray_S20reg_gff_1_SFF_7_MUXInst_X), .Z0_f (new_AGEMA_signal_2938), .Z1_t (new_AGEMA_signal_2939), .Z1_f (new_AGEMA_signal_2940) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S20reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S20reg_gff_1_SFF_7_MUXInst_X), .B0_f (new_AGEMA_signal_2938), .B1_t (new_AGEMA_signal_2939), .B1_f (new_AGEMA_signal_2940), .Z0_t (stateArray_S20reg_gff_1_SFF_7_MUXInst_Y), .Z0_f (new_AGEMA_signal_6082), .Z1_t (new_AGEMA_signal_6083), .Z1_f (new_AGEMA_signal_6084) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S20reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (stateArray_S20reg_gff_1_SFF_7_MUXInst_Y), .A0_f (new_AGEMA_signal_6082), .A1_t (new_AGEMA_signal_6083), .A1_f (new_AGEMA_signal_6084), .B0_t (stateArray_outS21ser[7]), .B0_f (new_AGEMA_signal_2932), .B1_t (new_AGEMA_signal_2933), .B1_f (new_AGEMA_signal_2934), .Z0_t (MixColumns_line2_S02[0]), .Z0_f (new_AGEMA_signal_3031), .Z1_t (new_AGEMA_signal_3032), .Z1_f (new_AGEMA_signal_3033) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S21reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS22ser[0]), .A0_f (new_AGEMA_signal_2872), .A1_t (new_AGEMA_signal_2873), .A1_f (new_AGEMA_signal_2874), .B0_t (stateArray_outS23ser[0]), .B0_f (new_AGEMA_signal_2941), .B1_t (new_AGEMA_signal_2942), .B1_f (new_AGEMA_signal_2943), .Z0_t (stateArray_S21reg_gff_1_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_2944), .Z1_t (new_AGEMA_signal_2945), .Z1_f (new_AGEMA_signal_2946) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S21reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S21reg_gff_1_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_2944), .B1_t (new_AGEMA_signal_2945), .B1_f (new_AGEMA_signal_2946), .Z0_t (stateArray_S21reg_gff_1_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_6085), .Z1_t (new_AGEMA_signal_6086), .Z1_f (new_AGEMA_signal_6087) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S21reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (stateArray_S21reg_gff_1_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_6085), .A1_t (new_AGEMA_signal_6086), .A1_f (new_AGEMA_signal_6087), .B0_t (stateArray_outS22ser[0]), .B0_f (new_AGEMA_signal_2872), .B1_t (new_AGEMA_signal_2873), .B1_f (new_AGEMA_signal_2874), .Z0_t (stateArray_outS21ser[0]), .Z0_f (new_AGEMA_signal_2869), .Z1_t (new_AGEMA_signal_2870), .Z1_f (new_AGEMA_signal_2871) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S21reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS22ser[1]), .A0_f (new_AGEMA_signal_2881), .A1_t (new_AGEMA_signal_2882), .A1_f (new_AGEMA_signal_2883), .B0_t (stateArray_outS23ser[1]), .B0_f (new_AGEMA_signal_2947), .B1_t (new_AGEMA_signal_2948), .B1_f (new_AGEMA_signal_2949), .Z0_t (stateArray_S21reg_gff_1_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_2950), .Z1_t (new_AGEMA_signal_2951), .Z1_f (new_AGEMA_signal_2952) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S21reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S21reg_gff_1_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_2950), .B1_t (new_AGEMA_signal_2951), .B1_f (new_AGEMA_signal_2952), .Z0_t (stateArray_S21reg_gff_1_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_6088), .Z1_t (new_AGEMA_signal_6089), .Z1_f (new_AGEMA_signal_6090) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S21reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (stateArray_S21reg_gff_1_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_6088), .A1_t (new_AGEMA_signal_6089), .A1_f (new_AGEMA_signal_6090), .B0_t (stateArray_outS22ser[1]), .B0_f (new_AGEMA_signal_2881), .B1_t (new_AGEMA_signal_2882), .B1_f (new_AGEMA_signal_2883), .Z0_t (stateArray_outS21ser[1]), .Z0_f (new_AGEMA_signal_2878), .Z1_t (new_AGEMA_signal_2879), .Z1_f (new_AGEMA_signal_2880) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S21reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS22ser[2]), .A0_f (new_AGEMA_signal_2890), .A1_t (new_AGEMA_signal_2891), .A1_f (new_AGEMA_signal_2892), .B0_t (stateArray_outS23ser[2]), .B0_f (new_AGEMA_signal_2953), .B1_t (new_AGEMA_signal_2954), .B1_f (new_AGEMA_signal_2955), .Z0_t (stateArray_S21reg_gff_1_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_2956), .Z1_t (new_AGEMA_signal_2957), .Z1_f (new_AGEMA_signal_2958) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S21reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S21reg_gff_1_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_2956), .B1_t (new_AGEMA_signal_2957), .B1_f (new_AGEMA_signal_2958), .Z0_t (stateArray_S21reg_gff_1_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_6091), .Z1_t (new_AGEMA_signal_6092), .Z1_f (new_AGEMA_signal_6093) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S21reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (stateArray_S21reg_gff_1_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_6091), .A1_t (new_AGEMA_signal_6092), .A1_f (new_AGEMA_signal_6093), .B0_t (stateArray_outS22ser[2]), .B0_f (new_AGEMA_signal_2890), .B1_t (new_AGEMA_signal_2891), .B1_f (new_AGEMA_signal_2892), .Z0_t (stateArray_outS21ser[2]), .Z0_f (new_AGEMA_signal_2887), .Z1_t (new_AGEMA_signal_2888), .Z1_f (new_AGEMA_signal_2889) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S21reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS22ser[3]), .A0_f (new_AGEMA_signal_2899), .A1_t (new_AGEMA_signal_2900), .A1_f (new_AGEMA_signal_2901), .B0_t (stateArray_outS23ser[3]), .B0_f (new_AGEMA_signal_2959), .B1_t (new_AGEMA_signal_2960), .B1_f (new_AGEMA_signal_2961), .Z0_t (stateArray_S21reg_gff_1_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_2962), .Z1_t (new_AGEMA_signal_2963), .Z1_f (new_AGEMA_signal_2964) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S21reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S21reg_gff_1_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_2962), .B1_t (new_AGEMA_signal_2963), .B1_f (new_AGEMA_signal_2964), .Z0_t (stateArray_S21reg_gff_1_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_6094), .Z1_t (new_AGEMA_signal_6095), .Z1_f (new_AGEMA_signal_6096) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S21reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (stateArray_S21reg_gff_1_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_6094), .A1_t (new_AGEMA_signal_6095), .A1_f (new_AGEMA_signal_6096), .B0_t (stateArray_outS22ser[3]), .B0_f (new_AGEMA_signal_2899), .B1_t (new_AGEMA_signal_2900), .B1_f (new_AGEMA_signal_2901), .Z0_t (stateArray_outS21ser[3]), .Z0_f (new_AGEMA_signal_2896), .Z1_t (new_AGEMA_signal_2897), .Z1_f (new_AGEMA_signal_2898) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S21reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS22ser[4]), .A0_f (new_AGEMA_signal_2908), .A1_t (new_AGEMA_signal_2909), .A1_f (new_AGEMA_signal_2910), .B0_t (stateArray_outS23ser[4]), .B0_f (new_AGEMA_signal_2965), .B1_t (new_AGEMA_signal_2966), .B1_f (new_AGEMA_signal_2967), .Z0_t (stateArray_S21reg_gff_1_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_2968), .Z1_t (new_AGEMA_signal_2969), .Z1_f (new_AGEMA_signal_2970) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S21reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S21reg_gff_1_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_2968), .B1_t (new_AGEMA_signal_2969), .B1_f (new_AGEMA_signal_2970), .Z0_t (stateArray_S21reg_gff_1_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_6097), .Z1_t (new_AGEMA_signal_6098), .Z1_f (new_AGEMA_signal_6099) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S21reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (stateArray_S21reg_gff_1_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_6097), .A1_t (new_AGEMA_signal_6098), .A1_f (new_AGEMA_signal_6099), .B0_t (stateArray_outS22ser[4]), .B0_f (new_AGEMA_signal_2908), .B1_t (new_AGEMA_signal_2909), .B1_f (new_AGEMA_signal_2910), .Z0_t (stateArray_outS21ser[4]), .Z0_f (new_AGEMA_signal_2905), .Z1_t (new_AGEMA_signal_2906), .Z1_f (new_AGEMA_signal_2907) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S21reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS22ser[5]), .A0_f (new_AGEMA_signal_2917), .A1_t (new_AGEMA_signal_2918), .A1_f (new_AGEMA_signal_2919), .B0_t (stateArray_outS23ser[5]), .B0_f (new_AGEMA_signal_2971), .B1_t (new_AGEMA_signal_2972), .B1_f (new_AGEMA_signal_2973), .Z0_t (stateArray_S21reg_gff_1_SFF_5_MUXInst_X), .Z0_f (new_AGEMA_signal_2974), .Z1_t (new_AGEMA_signal_2975), .Z1_f (new_AGEMA_signal_2976) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S21reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S21reg_gff_1_SFF_5_MUXInst_X), .B0_f (new_AGEMA_signal_2974), .B1_t (new_AGEMA_signal_2975), .B1_f (new_AGEMA_signal_2976), .Z0_t (stateArray_S21reg_gff_1_SFF_5_MUXInst_Y), .Z0_f (new_AGEMA_signal_6100), .Z1_t (new_AGEMA_signal_6101), .Z1_f (new_AGEMA_signal_6102) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S21reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (stateArray_S21reg_gff_1_SFF_5_MUXInst_Y), .A0_f (new_AGEMA_signal_6100), .A1_t (new_AGEMA_signal_6101), .A1_f (new_AGEMA_signal_6102), .B0_t (stateArray_outS22ser[5]), .B0_f (new_AGEMA_signal_2917), .B1_t (new_AGEMA_signal_2918), .B1_f (new_AGEMA_signal_2919), .Z0_t (stateArray_outS21ser[5]), .Z0_f (new_AGEMA_signal_2914), .Z1_t (new_AGEMA_signal_2915), .Z1_f (new_AGEMA_signal_2916) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S21reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS22ser[6]), .A0_f (new_AGEMA_signal_2926), .A1_t (new_AGEMA_signal_2927), .A1_f (new_AGEMA_signal_2928), .B0_t (stateArray_outS23ser[6]), .B0_f (new_AGEMA_signal_2977), .B1_t (new_AGEMA_signal_2978), .B1_f (new_AGEMA_signal_2979), .Z0_t (stateArray_S21reg_gff_1_SFF_6_MUXInst_X), .Z0_f (new_AGEMA_signal_2980), .Z1_t (new_AGEMA_signal_2981), .Z1_f (new_AGEMA_signal_2982) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S21reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S21reg_gff_1_SFF_6_MUXInst_X), .B0_f (new_AGEMA_signal_2980), .B1_t (new_AGEMA_signal_2981), .B1_f (new_AGEMA_signal_2982), .Z0_t (stateArray_S21reg_gff_1_SFF_6_MUXInst_Y), .Z0_f (new_AGEMA_signal_6103), .Z1_t (new_AGEMA_signal_6104), .Z1_f (new_AGEMA_signal_6105) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S21reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (stateArray_S21reg_gff_1_SFF_6_MUXInst_Y), .A0_f (new_AGEMA_signal_6103), .A1_t (new_AGEMA_signal_6104), .A1_f (new_AGEMA_signal_6105), .B0_t (stateArray_outS22ser[6]), .B0_f (new_AGEMA_signal_2926), .B1_t (new_AGEMA_signal_2927), .B1_f (new_AGEMA_signal_2928), .Z0_t (stateArray_outS21ser[6]), .Z0_f (new_AGEMA_signal_2923), .Z1_t (new_AGEMA_signal_2924), .Z1_f (new_AGEMA_signal_2925) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S21reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS22ser[7]), .A0_f (new_AGEMA_signal_2935), .A1_t (new_AGEMA_signal_2936), .A1_f (new_AGEMA_signal_2937), .B0_t (stateArray_outS23ser[7]), .B0_f (new_AGEMA_signal_2983), .B1_t (new_AGEMA_signal_2984), .B1_f (new_AGEMA_signal_2985), .Z0_t (stateArray_S21reg_gff_1_SFF_7_MUXInst_X), .Z0_f (new_AGEMA_signal_2986), .Z1_t (new_AGEMA_signal_2987), .Z1_f (new_AGEMA_signal_2988) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S21reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S21reg_gff_1_SFF_7_MUXInst_X), .B0_f (new_AGEMA_signal_2986), .B1_t (new_AGEMA_signal_2987), .B1_f (new_AGEMA_signal_2988), .Z0_t (stateArray_S21reg_gff_1_SFF_7_MUXInst_Y), .Z0_f (new_AGEMA_signal_6106), .Z1_t (new_AGEMA_signal_6107), .Z1_f (new_AGEMA_signal_6108) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S21reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (stateArray_S21reg_gff_1_SFF_7_MUXInst_Y), .A0_f (new_AGEMA_signal_6106), .A1_t (new_AGEMA_signal_6107), .A1_f (new_AGEMA_signal_6108), .B0_t (stateArray_outS22ser[7]), .B0_f (new_AGEMA_signal_2935), .B1_t (new_AGEMA_signal_2936), .B1_f (new_AGEMA_signal_2937), .Z0_t (stateArray_outS21ser[7]), .Z0_f (new_AGEMA_signal_2932), .Z1_t (new_AGEMA_signal_2933), .Z1_f (new_AGEMA_signal_2934) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S22reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS23ser[0]), .A0_f (new_AGEMA_signal_2941), .A1_t (new_AGEMA_signal_2942), .A1_f (new_AGEMA_signal_2943), .B0_t (MCin[8]), .B0_f (new_AGEMA_signal_2989), .B1_t (new_AGEMA_signal_2990), .B1_f (new_AGEMA_signal_2991), .Z0_t (stateArray_S22reg_gff_1_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_2992), .Z1_t (new_AGEMA_signal_2993), .Z1_f (new_AGEMA_signal_2994) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S22reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S22reg_gff_1_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_2992), .B1_t (new_AGEMA_signal_2993), .B1_f (new_AGEMA_signal_2994), .Z0_t (stateArray_S22reg_gff_1_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_6109), .Z1_t (new_AGEMA_signal_6110), .Z1_f (new_AGEMA_signal_6111) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S22reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (stateArray_S22reg_gff_1_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_6109), .A1_t (new_AGEMA_signal_6110), .A1_f (new_AGEMA_signal_6111), .B0_t (stateArray_outS23ser[0]), .B0_f (new_AGEMA_signal_2941), .B1_t (new_AGEMA_signal_2942), .B1_f (new_AGEMA_signal_2943), .Z0_t (stateArray_outS22ser[0]), .Z0_f (new_AGEMA_signal_2872), .Z1_t (new_AGEMA_signal_2873), .Z1_f (new_AGEMA_signal_2874) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S22reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS23ser[1]), .A0_f (new_AGEMA_signal_2947), .A1_t (new_AGEMA_signal_2948), .A1_f (new_AGEMA_signal_2949), .B0_t (MixColumns_line2_S02[2]), .B0_f (new_AGEMA_signal_2995), .B1_t (new_AGEMA_signal_2996), .B1_f (new_AGEMA_signal_2997), .Z0_t (stateArray_S22reg_gff_1_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_2998), .Z1_t (new_AGEMA_signal_2999), .Z1_f (new_AGEMA_signal_3000) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S22reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S22reg_gff_1_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_2998), .B1_t (new_AGEMA_signal_2999), .B1_f (new_AGEMA_signal_3000), .Z0_t (stateArray_S22reg_gff_1_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_6112), .Z1_t (new_AGEMA_signal_6113), .Z1_f (new_AGEMA_signal_6114) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S22reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (stateArray_S22reg_gff_1_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_6112), .A1_t (new_AGEMA_signal_6113), .A1_f (new_AGEMA_signal_6114), .B0_t (stateArray_outS23ser[1]), .B0_f (new_AGEMA_signal_2947), .B1_t (new_AGEMA_signal_2948), .B1_f (new_AGEMA_signal_2949), .Z0_t (stateArray_outS22ser[1]), .Z0_f (new_AGEMA_signal_2881), .Z1_t (new_AGEMA_signal_2882), .Z1_f (new_AGEMA_signal_2883) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S22reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS23ser[2]), .A0_f (new_AGEMA_signal_2953), .A1_t (new_AGEMA_signal_2954), .A1_f (new_AGEMA_signal_2955), .B0_t (MCin[10]), .B0_f (new_AGEMA_signal_3001), .B1_t (new_AGEMA_signal_3002), .B1_f (new_AGEMA_signal_3003), .Z0_t (stateArray_S22reg_gff_1_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_3004), .Z1_t (new_AGEMA_signal_3005), .Z1_f (new_AGEMA_signal_3006) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S22reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S22reg_gff_1_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_3004), .B1_t (new_AGEMA_signal_3005), .B1_f (new_AGEMA_signal_3006), .Z0_t (stateArray_S22reg_gff_1_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_6115), .Z1_t (new_AGEMA_signal_6116), .Z1_f (new_AGEMA_signal_6117) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S22reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (stateArray_S22reg_gff_1_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_6115), .A1_t (new_AGEMA_signal_6116), .A1_f (new_AGEMA_signal_6117), .B0_t (stateArray_outS23ser[2]), .B0_f (new_AGEMA_signal_2953), .B1_t (new_AGEMA_signal_2954), .B1_f (new_AGEMA_signal_2955), .Z0_t (stateArray_outS22ser[2]), .Z0_f (new_AGEMA_signal_2890), .Z1_t (new_AGEMA_signal_2891), .Z1_f (new_AGEMA_signal_2892) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S22reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS23ser[3]), .A0_f (new_AGEMA_signal_2959), .A1_t (new_AGEMA_signal_2960), .A1_f (new_AGEMA_signal_2961), .B0_t (MCin[11]), .B0_f (new_AGEMA_signal_3007), .B1_t (new_AGEMA_signal_3008), .B1_f (new_AGEMA_signal_3009), .Z0_t (stateArray_S22reg_gff_1_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_3010), .Z1_t (new_AGEMA_signal_3011), .Z1_f (new_AGEMA_signal_3012) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S22reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S22reg_gff_1_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_3010), .B1_t (new_AGEMA_signal_3011), .B1_f (new_AGEMA_signal_3012), .Z0_t (stateArray_S22reg_gff_1_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_6118), .Z1_t (new_AGEMA_signal_6119), .Z1_f (new_AGEMA_signal_6120) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S22reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (stateArray_S22reg_gff_1_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_6118), .A1_t (new_AGEMA_signal_6119), .A1_f (new_AGEMA_signal_6120), .B0_t (stateArray_outS23ser[3]), .B0_f (new_AGEMA_signal_2959), .B1_t (new_AGEMA_signal_2960), .B1_f (new_AGEMA_signal_2961), .Z0_t (stateArray_outS22ser[3]), .Z0_f (new_AGEMA_signal_2899), .Z1_t (new_AGEMA_signal_2900), .Z1_f (new_AGEMA_signal_2901) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S22reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS23ser[4]), .A0_f (new_AGEMA_signal_2965), .A1_t (new_AGEMA_signal_2966), .A1_f (new_AGEMA_signal_2967), .B0_t (MixColumns_line2_S02[5]), .B0_f (new_AGEMA_signal_3013), .B1_t (new_AGEMA_signal_3014), .B1_f (new_AGEMA_signal_3015), .Z0_t (stateArray_S22reg_gff_1_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_3016), .Z1_t (new_AGEMA_signal_3017), .Z1_f (new_AGEMA_signal_3018) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S22reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S22reg_gff_1_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_3016), .B1_t (new_AGEMA_signal_3017), .B1_f (new_AGEMA_signal_3018), .Z0_t (stateArray_S22reg_gff_1_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_6121), .Z1_t (new_AGEMA_signal_6122), .Z1_f (new_AGEMA_signal_6123) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S22reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (stateArray_S22reg_gff_1_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_6121), .A1_t (new_AGEMA_signal_6122), .A1_f (new_AGEMA_signal_6123), .B0_t (stateArray_outS23ser[4]), .B0_f (new_AGEMA_signal_2965), .B1_t (new_AGEMA_signal_2966), .B1_f (new_AGEMA_signal_2967), .Z0_t (stateArray_outS22ser[4]), .Z0_f (new_AGEMA_signal_2908), .Z1_t (new_AGEMA_signal_2909), .Z1_f (new_AGEMA_signal_2910) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S22reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS23ser[5]), .A0_f (new_AGEMA_signal_2971), .A1_t (new_AGEMA_signal_2972), .A1_f (new_AGEMA_signal_2973), .B0_t (MixColumns_line2_S02[6]), .B0_f (new_AGEMA_signal_3019), .B1_t (new_AGEMA_signal_3020), .B1_f (new_AGEMA_signal_3021), .Z0_t (stateArray_S22reg_gff_1_SFF_5_MUXInst_X), .Z0_f (new_AGEMA_signal_3022), .Z1_t (new_AGEMA_signal_3023), .Z1_f (new_AGEMA_signal_3024) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S22reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S22reg_gff_1_SFF_5_MUXInst_X), .B0_f (new_AGEMA_signal_3022), .B1_t (new_AGEMA_signal_3023), .B1_f (new_AGEMA_signal_3024), .Z0_t (stateArray_S22reg_gff_1_SFF_5_MUXInst_Y), .Z0_f (new_AGEMA_signal_6124), .Z1_t (new_AGEMA_signal_6125), .Z1_f (new_AGEMA_signal_6126) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S22reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (stateArray_S22reg_gff_1_SFF_5_MUXInst_Y), .A0_f (new_AGEMA_signal_6124), .A1_t (new_AGEMA_signal_6125), .A1_f (new_AGEMA_signal_6126), .B0_t (stateArray_outS23ser[5]), .B0_f (new_AGEMA_signal_2971), .B1_t (new_AGEMA_signal_2972), .B1_f (new_AGEMA_signal_2973), .Z0_t (stateArray_outS22ser[5]), .Z0_f (new_AGEMA_signal_2917), .Z1_t (new_AGEMA_signal_2918), .Z1_f (new_AGEMA_signal_2919) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S22reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS23ser[6]), .A0_f (new_AGEMA_signal_2977), .A1_t (new_AGEMA_signal_2978), .A1_f (new_AGEMA_signal_2979), .B0_t (MixColumns_line2_S02[7]), .B0_f (new_AGEMA_signal_3025), .B1_t (new_AGEMA_signal_3026), .B1_f (new_AGEMA_signal_3027), .Z0_t (stateArray_S22reg_gff_1_SFF_6_MUXInst_X), .Z0_f (new_AGEMA_signal_3028), .Z1_t (new_AGEMA_signal_3029), .Z1_f (new_AGEMA_signal_3030) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S22reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S22reg_gff_1_SFF_6_MUXInst_X), .B0_f (new_AGEMA_signal_3028), .B1_t (new_AGEMA_signal_3029), .B1_f (new_AGEMA_signal_3030), .Z0_t (stateArray_S22reg_gff_1_SFF_6_MUXInst_Y), .Z0_f (new_AGEMA_signal_6127), .Z1_t (new_AGEMA_signal_6128), .Z1_f (new_AGEMA_signal_6129) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S22reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (stateArray_S22reg_gff_1_SFF_6_MUXInst_Y), .A0_f (new_AGEMA_signal_6127), .A1_t (new_AGEMA_signal_6128), .A1_f (new_AGEMA_signal_6129), .B0_t (stateArray_outS23ser[6]), .B0_f (new_AGEMA_signal_2977), .B1_t (new_AGEMA_signal_2978), .B1_f (new_AGEMA_signal_2979), .Z0_t (stateArray_outS22ser[6]), .Z0_f (new_AGEMA_signal_2926), .Z1_t (new_AGEMA_signal_2927), .Z1_f (new_AGEMA_signal_2928) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S22reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS23ser[7]), .A0_f (new_AGEMA_signal_2983), .A1_t (new_AGEMA_signal_2984), .A1_f (new_AGEMA_signal_2985), .B0_t (MixColumns_line2_S02[0]), .B0_f (new_AGEMA_signal_3031), .B1_t (new_AGEMA_signal_3032), .B1_f (new_AGEMA_signal_3033), .Z0_t (stateArray_S22reg_gff_1_SFF_7_MUXInst_X), .Z0_f (new_AGEMA_signal_3034), .Z1_t (new_AGEMA_signal_3035), .Z1_f (new_AGEMA_signal_3036) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S22reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S22reg_gff_1_SFF_7_MUXInst_X), .B0_f (new_AGEMA_signal_3034), .B1_t (new_AGEMA_signal_3035), .B1_f (new_AGEMA_signal_3036), .Z0_t (stateArray_S22reg_gff_1_SFF_7_MUXInst_Y), .Z0_f (new_AGEMA_signal_6130), .Z1_t (new_AGEMA_signal_6131), .Z1_f (new_AGEMA_signal_6132) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S22reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (stateArray_S22reg_gff_1_SFF_7_MUXInst_Y), .A0_f (new_AGEMA_signal_6130), .A1_t (new_AGEMA_signal_6131), .A1_f (new_AGEMA_signal_6132), .B0_t (stateArray_outS23ser[7]), .B0_f (new_AGEMA_signal_2983), .B1_t (new_AGEMA_signal_2984), .B1_f (new_AGEMA_signal_2985), .Z0_t (stateArray_outS22ser[7]), .Z0_f (new_AGEMA_signal_2935), .Z1_t (new_AGEMA_signal_2936), .Z1_f (new_AGEMA_signal_2937) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S23reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS23ser[0]), .A0_f (new_AGEMA_signal_6253), .A1_t (new_AGEMA_signal_6254), .A1_f (new_AGEMA_signal_6255), .B0_t (stateArray_outS21ser[0]), .B0_f (new_AGEMA_signal_2869), .B1_t (new_AGEMA_signal_2870), .B1_f (new_AGEMA_signal_2871), .Z0_t (stateArray_S23reg_gff_1_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_6349), .Z1_t (new_AGEMA_signal_6350), .Z1_f (new_AGEMA_signal_6351) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S23reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S23reg_gff_1_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_6349), .B1_t (new_AGEMA_signal_6350), .B1_f (new_AGEMA_signal_6351), .Z0_t (stateArray_S23reg_gff_1_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_7206), .Z1_t (new_AGEMA_signal_7207), .Z1_f (new_AGEMA_signal_7208) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S23reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (stateArray_S23reg_gff_1_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_7206), .A1_t (new_AGEMA_signal_7207), .A1_f (new_AGEMA_signal_7208), .B0_t (stateArray_inS23ser[0]), .B0_f (new_AGEMA_signal_6253), .B1_t (new_AGEMA_signal_6254), .B1_f (new_AGEMA_signal_6255), .Z0_t (stateArray_outS23ser[0]), .Z0_f (new_AGEMA_signal_2941), .Z1_t (new_AGEMA_signal_2942), .Z1_f (new_AGEMA_signal_2943) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S23reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS23ser[1]), .A0_f (new_AGEMA_signal_6382), .A1_t (new_AGEMA_signal_6383), .A1_f (new_AGEMA_signal_6384), .B0_t (stateArray_outS21ser[1]), .B0_f (new_AGEMA_signal_2878), .B1_t (new_AGEMA_signal_2879), .B1_f (new_AGEMA_signal_2880), .Z0_t (stateArray_S23reg_gff_1_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_7209), .Z1_t (new_AGEMA_signal_7210), .Z1_f (new_AGEMA_signal_7211) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S23reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S23reg_gff_1_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_7209), .B1_t (new_AGEMA_signal_7210), .B1_f (new_AGEMA_signal_7211), .Z0_t (stateArray_S23reg_gff_1_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_7292), .Z1_t (new_AGEMA_signal_7293), .Z1_f (new_AGEMA_signal_7294) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S23reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (stateArray_S23reg_gff_1_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_7292), .A1_t (new_AGEMA_signal_7293), .A1_f (new_AGEMA_signal_7294), .B0_t (stateArray_inS23ser[1]), .B0_f (new_AGEMA_signal_6382), .B1_t (new_AGEMA_signal_6383), .B1_f (new_AGEMA_signal_6384), .Z0_t (stateArray_outS23ser[1]), .Z0_f (new_AGEMA_signal_2947), .Z1_t (new_AGEMA_signal_2948), .Z1_f (new_AGEMA_signal_2949) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S23reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS23ser[2]), .A0_f (new_AGEMA_signal_6259), .A1_t (new_AGEMA_signal_6260), .A1_f (new_AGEMA_signal_6261), .B0_t (stateArray_outS21ser[2]), .B0_f (new_AGEMA_signal_2887), .B1_t (new_AGEMA_signal_2888), .B1_f (new_AGEMA_signal_2889), .Z0_t (stateArray_S23reg_gff_1_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_6352), .Z1_t (new_AGEMA_signal_6353), .Z1_f (new_AGEMA_signal_6354) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S23reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S23reg_gff_1_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_6352), .B1_t (new_AGEMA_signal_6353), .B1_f (new_AGEMA_signal_6354), .Z0_t (stateArray_S23reg_gff_1_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_7212), .Z1_t (new_AGEMA_signal_7213), .Z1_f (new_AGEMA_signal_7214) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S23reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (stateArray_S23reg_gff_1_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_7212), .A1_t (new_AGEMA_signal_7213), .A1_f (new_AGEMA_signal_7214), .B0_t (stateArray_inS23ser[2]), .B0_f (new_AGEMA_signal_6259), .B1_t (new_AGEMA_signal_6260), .B1_f (new_AGEMA_signal_6261), .Z0_t (stateArray_outS23ser[2]), .Z0_f (new_AGEMA_signal_2953), .Z1_t (new_AGEMA_signal_2954), .Z1_f (new_AGEMA_signal_2955) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S23reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS23ser[3]), .A0_f (new_AGEMA_signal_6385), .A1_t (new_AGEMA_signal_6386), .A1_f (new_AGEMA_signal_6387), .B0_t (stateArray_outS21ser[3]), .B0_f (new_AGEMA_signal_2896), .B1_t (new_AGEMA_signal_2897), .B1_f (new_AGEMA_signal_2898), .Z0_t (stateArray_S23reg_gff_1_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_7215), .Z1_t (new_AGEMA_signal_7216), .Z1_f (new_AGEMA_signal_7217) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S23reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S23reg_gff_1_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_7215), .B1_t (new_AGEMA_signal_7216), .B1_f (new_AGEMA_signal_7217), .Z0_t (stateArray_S23reg_gff_1_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_7295), .Z1_t (new_AGEMA_signal_7296), .Z1_f (new_AGEMA_signal_7297) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S23reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (stateArray_S23reg_gff_1_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_7295), .A1_t (new_AGEMA_signal_7296), .A1_f (new_AGEMA_signal_7297), .B0_t (stateArray_inS23ser[3]), .B0_f (new_AGEMA_signal_6385), .B1_t (new_AGEMA_signal_6386), .B1_f (new_AGEMA_signal_6387), .Z0_t (stateArray_outS23ser[3]), .Z0_f (new_AGEMA_signal_2959), .Z1_t (new_AGEMA_signal_2960), .Z1_f (new_AGEMA_signal_2961) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S23reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS23ser[4]), .A0_f (new_AGEMA_signal_6388), .A1_t (new_AGEMA_signal_6389), .A1_f (new_AGEMA_signal_6390), .B0_t (stateArray_outS21ser[4]), .B0_f (new_AGEMA_signal_2905), .B1_t (new_AGEMA_signal_2906), .B1_f (new_AGEMA_signal_2907), .Z0_t (stateArray_S23reg_gff_1_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_7218), .Z1_t (new_AGEMA_signal_7219), .Z1_f (new_AGEMA_signal_7220) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S23reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S23reg_gff_1_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_7218), .B1_t (new_AGEMA_signal_7219), .B1_f (new_AGEMA_signal_7220), .Z0_t (stateArray_S23reg_gff_1_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_7298), .Z1_t (new_AGEMA_signal_7299), .Z1_f (new_AGEMA_signal_7300) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S23reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (stateArray_S23reg_gff_1_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_7298), .A1_t (new_AGEMA_signal_7299), .A1_f (new_AGEMA_signal_7300), .B0_t (stateArray_inS23ser[4]), .B0_f (new_AGEMA_signal_6388), .B1_t (new_AGEMA_signal_6389), .B1_f (new_AGEMA_signal_6390), .Z0_t (stateArray_outS23ser[4]), .Z0_f (new_AGEMA_signal_2965), .Z1_t (new_AGEMA_signal_2966), .Z1_f (new_AGEMA_signal_2967) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S23reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS23ser[5]), .A0_f (new_AGEMA_signal_6268), .A1_t (new_AGEMA_signal_6269), .A1_f (new_AGEMA_signal_6270), .B0_t (stateArray_outS21ser[5]), .B0_f (new_AGEMA_signal_2914), .B1_t (new_AGEMA_signal_2915), .B1_f (new_AGEMA_signal_2916), .Z0_t (stateArray_S23reg_gff_1_SFF_5_MUXInst_X), .Z0_f (new_AGEMA_signal_6355), .Z1_t (new_AGEMA_signal_6356), .Z1_f (new_AGEMA_signal_6357) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S23reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S23reg_gff_1_SFF_5_MUXInst_X), .B0_f (new_AGEMA_signal_6355), .B1_t (new_AGEMA_signal_6356), .B1_f (new_AGEMA_signal_6357), .Z0_t (stateArray_S23reg_gff_1_SFF_5_MUXInst_Y), .Z0_f (new_AGEMA_signal_7221), .Z1_t (new_AGEMA_signal_7222), .Z1_f (new_AGEMA_signal_7223) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S23reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (stateArray_S23reg_gff_1_SFF_5_MUXInst_Y), .A0_f (new_AGEMA_signal_7221), .A1_t (new_AGEMA_signal_7222), .A1_f (new_AGEMA_signal_7223), .B0_t (stateArray_inS23ser[5]), .B0_f (new_AGEMA_signal_6268), .B1_t (new_AGEMA_signal_6269), .B1_f (new_AGEMA_signal_6270), .Z0_t (stateArray_outS23ser[5]), .Z0_f (new_AGEMA_signal_2971), .Z1_t (new_AGEMA_signal_2972), .Z1_f (new_AGEMA_signal_2973) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S23reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS23ser[6]), .A0_f (new_AGEMA_signal_6271), .A1_t (new_AGEMA_signal_6272), .A1_f (new_AGEMA_signal_6273), .B0_t (stateArray_outS21ser[6]), .B0_f (new_AGEMA_signal_2923), .B1_t (new_AGEMA_signal_2924), .B1_f (new_AGEMA_signal_2925), .Z0_t (stateArray_S23reg_gff_1_SFF_6_MUXInst_X), .Z0_f (new_AGEMA_signal_6358), .Z1_t (new_AGEMA_signal_6359), .Z1_f (new_AGEMA_signal_6360) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S23reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S23reg_gff_1_SFF_6_MUXInst_X), .B0_f (new_AGEMA_signal_6358), .B1_t (new_AGEMA_signal_6359), .B1_f (new_AGEMA_signal_6360), .Z0_t (stateArray_S23reg_gff_1_SFF_6_MUXInst_Y), .Z0_f (new_AGEMA_signal_7224), .Z1_t (new_AGEMA_signal_7225), .Z1_f (new_AGEMA_signal_7226) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S23reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (stateArray_S23reg_gff_1_SFF_6_MUXInst_Y), .A0_f (new_AGEMA_signal_7224), .A1_t (new_AGEMA_signal_7225), .A1_f (new_AGEMA_signal_7226), .B0_t (stateArray_inS23ser[6]), .B0_f (new_AGEMA_signal_6271), .B1_t (new_AGEMA_signal_6272), .B1_f (new_AGEMA_signal_6273), .Z0_t (stateArray_outS23ser[6]), .Z0_f (new_AGEMA_signal_2977), .Z1_t (new_AGEMA_signal_2978), .Z1_f (new_AGEMA_signal_2979) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S23reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS23ser[7]), .A0_f (new_AGEMA_signal_6274), .A1_t (new_AGEMA_signal_6275), .A1_f (new_AGEMA_signal_6276), .B0_t (stateArray_outS21ser[7]), .B0_f (new_AGEMA_signal_2932), .B1_t (new_AGEMA_signal_2933), .B1_f (new_AGEMA_signal_2934), .Z0_t (stateArray_S23reg_gff_1_SFF_7_MUXInst_X), .Z0_f (new_AGEMA_signal_6361), .Z1_t (new_AGEMA_signal_6362), .Z1_f (new_AGEMA_signal_6363) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S23reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S23reg_gff_1_SFF_7_MUXInst_X), .B0_f (new_AGEMA_signal_6361), .B1_t (new_AGEMA_signal_6362), .B1_f (new_AGEMA_signal_6363), .Z0_t (stateArray_S23reg_gff_1_SFF_7_MUXInst_Y), .Z0_f (new_AGEMA_signal_7227), .Z1_t (new_AGEMA_signal_7228), .Z1_f (new_AGEMA_signal_7229) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S23reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (stateArray_S23reg_gff_1_SFF_7_MUXInst_Y), .A0_f (new_AGEMA_signal_7227), .A1_t (new_AGEMA_signal_7228), .A1_f (new_AGEMA_signal_7229), .B0_t (stateArray_inS23ser[7]), .B0_f (new_AGEMA_signal_6274), .B1_t (new_AGEMA_signal_6275), .B1_f (new_AGEMA_signal_6276), .Z0_t (stateArray_outS23ser[7]), .Z0_f (new_AGEMA_signal_2983), .Z1_t (new_AGEMA_signal_2984), .Z1_f (new_AGEMA_signal_2985) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S30reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS31ser[0]), .A0_f (new_AGEMA_signal_3037), .A1_t (new_AGEMA_signal_3038), .A1_f (new_AGEMA_signal_3039), .B0_t (stateArray_outS33ser[0]), .B0_f (new_AGEMA_signal_3040), .B1_t (new_AGEMA_signal_3041), .B1_f (new_AGEMA_signal_3042), .Z0_t (stateArray_S30reg_gff_1_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_3043), .Z1_t (new_AGEMA_signal_3044), .Z1_f (new_AGEMA_signal_3045) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S30reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S30reg_gff_1_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_3043), .B1_t (new_AGEMA_signal_3044), .B1_f (new_AGEMA_signal_3045), .Z0_t (stateArray_S30reg_gff_1_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_6133), .Z1_t (new_AGEMA_signal_6134), .Z1_f (new_AGEMA_signal_6135) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S30reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (stateArray_S30reg_gff_1_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_6133), .A1_t (new_AGEMA_signal_6134), .A1_f (new_AGEMA_signal_6135), .B0_t (stateArray_outS31ser[0]), .B0_f (new_AGEMA_signal_3037), .B1_t (new_AGEMA_signal_3038), .B1_f (new_AGEMA_signal_3039), .Z0_t (MCin[0]), .Z0_f (new_AGEMA_signal_3112), .Z1_t (new_AGEMA_signal_3113), .Z1_f (new_AGEMA_signal_3114) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S30reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS31ser[1]), .A0_f (new_AGEMA_signal_3046), .A1_t (new_AGEMA_signal_3047), .A1_f (new_AGEMA_signal_3048), .B0_t (stateArray_outS33ser[1]), .B0_f (new_AGEMA_signal_3049), .B1_t (new_AGEMA_signal_3050), .B1_f (new_AGEMA_signal_3051), .Z0_t (stateArray_S30reg_gff_1_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_3052), .Z1_t (new_AGEMA_signal_3053), .Z1_f (new_AGEMA_signal_3054) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S30reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S30reg_gff_1_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_3052), .B1_t (new_AGEMA_signal_3053), .B1_f (new_AGEMA_signal_3054), .Z0_t (stateArray_S30reg_gff_1_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_6136), .Z1_t (new_AGEMA_signal_6137), .Z1_f (new_AGEMA_signal_6138) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S30reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (stateArray_S30reg_gff_1_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_6136), .A1_t (new_AGEMA_signal_6137), .A1_f (new_AGEMA_signal_6138), .B0_t (stateArray_outS31ser[1]), .B0_f (new_AGEMA_signal_3046), .B1_t (new_AGEMA_signal_3047), .B1_f (new_AGEMA_signal_3048), .Z0_t (MixColumns_line3_S02[2]), .Z0_f (new_AGEMA_signal_3121), .Z1_t (new_AGEMA_signal_3122), .Z1_f (new_AGEMA_signal_3123) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S30reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS31ser[2]), .A0_f (new_AGEMA_signal_3055), .A1_t (new_AGEMA_signal_3056), .A1_f (new_AGEMA_signal_3057), .B0_t (stateArray_outS33ser[2]), .B0_f (new_AGEMA_signal_3058), .B1_t (new_AGEMA_signal_3059), .B1_f (new_AGEMA_signal_3060), .Z0_t (stateArray_S30reg_gff_1_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_3061), .Z1_t (new_AGEMA_signal_3062), .Z1_f (new_AGEMA_signal_3063) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S30reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S30reg_gff_1_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_3061), .B1_t (new_AGEMA_signal_3062), .B1_f (new_AGEMA_signal_3063), .Z0_t (stateArray_S30reg_gff_1_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_6139), .Z1_t (new_AGEMA_signal_6140), .Z1_f (new_AGEMA_signal_6141) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S30reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (stateArray_S30reg_gff_1_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_6139), .A1_t (new_AGEMA_signal_6140), .A1_f (new_AGEMA_signal_6141), .B0_t (stateArray_outS31ser[2]), .B0_f (new_AGEMA_signal_3055), .B1_t (new_AGEMA_signal_3056), .B1_f (new_AGEMA_signal_3057), .Z0_t (MCin[2]), .Z0_f (new_AGEMA_signal_3130), .Z1_t (new_AGEMA_signal_3131), .Z1_f (new_AGEMA_signal_3132) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S30reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS31ser[3]), .A0_f (new_AGEMA_signal_3064), .A1_t (new_AGEMA_signal_3065), .A1_f (new_AGEMA_signal_3066), .B0_t (stateArray_outS33ser[3]), .B0_f (new_AGEMA_signal_3067), .B1_t (new_AGEMA_signal_3068), .B1_f (new_AGEMA_signal_3069), .Z0_t (stateArray_S30reg_gff_1_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_3070), .Z1_t (new_AGEMA_signal_3071), .Z1_f (new_AGEMA_signal_3072) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S30reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S30reg_gff_1_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_3070), .B1_t (new_AGEMA_signal_3071), .B1_f (new_AGEMA_signal_3072), .Z0_t (stateArray_S30reg_gff_1_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_6142), .Z1_t (new_AGEMA_signal_6143), .Z1_f (new_AGEMA_signal_6144) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S30reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (stateArray_S30reg_gff_1_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_6142), .A1_t (new_AGEMA_signal_6143), .A1_f (new_AGEMA_signal_6144), .B0_t (stateArray_outS31ser[3]), .B0_f (new_AGEMA_signal_3064), .B1_t (new_AGEMA_signal_3065), .B1_f (new_AGEMA_signal_3066), .Z0_t (MCin[3]), .Z0_f (new_AGEMA_signal_3139), .Z1_t (new_AGEMA_signal_3140), .Z1_f (new_AGEMA_signal_3141) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S30reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS31ser[4]), .A0_f (new_AGEMA_signal_3073), .A1_t (new_AGEMA_signal_3074), .A1_f (new_AGEMA_signal_3075), .B0_t (stateArray_outS33ser[4]), .B0_f (new_AGEMA_signal_3076), .B1_t (new_AGEMA_signal_3077), .B1_f (new_AGEMA_signal_3078), .Z0_t (stateArray_S30reg_gff_1_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_3079), .Z1_t (new_AGEMA_signal_3080), .Z1_f (new_AGEMA_signal_3081) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S30reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S30reg_gff_1_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_3079), .B1_t (new_AGEMA_signal_3080), .B1_f (new_AGEMA_signal_3081), .Z0_t (stateArray_S30reg_gff_1_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_6145), .Z1_t (new_AGEMA_signal_6146), .Z1_f (new_AGEMA_signal_6147) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S30reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (stateArray_S30reg_gff_1_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_6145), .A1_t (new_AGEMA_signal_6146), .A1_f (new_AGEMA_signal_6147), .B0_t (stateArray_outS31ser[4]), .B0_f (new_AGEMA_signal_3073), .B1_t (new_AGEMA_signal_3074), .B1_f (new_AGEMA_signal_3075), .Z0_t (MixColumns_line3_S02[5]), .Z0_f (new_AGEMA_signal_3148), .Z1_t (new_AGEMA_signal_3149), .Z1_f (new_AGEMA_signal_3150) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S30reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS31ser[5]), .A0_f (new_AGEMA_signal_3082), .A1_t (new_AGEMA_signal_3083), .A1_f (new_AGEMA_signal_3084), .B0_t (stateArray_outS33ser[5]), .B0_f (new_AGEMA_signal_3085), .B1_t (new_AGEMA_signal_3086), .B1_f (new_AGEMA_signal_3087), .Z0_t (stateArray_S30reg_gff_1_SFF_5_MUXInst_X), .Z0_f (new_AGEMA_signal_3088), .Z1_t (new_AGEMA_signal_3089), .Z1_f (new_AGEMA_signal_3090) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S30reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S30reg_gff_1_SFF_5_MUXInst_X), .B0_f (new_AGEMA_signal_3088), .B1_t (new_AGEMA_signal_3089), .B1_f (new_AGEMA_signal_3090), .Z0_t (stateArray_S30reg_gff_1_SFF_5_MUXInst_Y), .Z0_f (new_AGEMA_signal_6148), .Z1_t (new_AGEMA_signal_6149), .Z1_f (new_AGEMA_signal_6150) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S30reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (stateArray_S30reg_gff_1_SFF_5_MUXInst_Y), .A0_f (new_AGEMA_signal_6148), .A1_t (new_AGEMA_signal_6149), .A1_f (new_AGEMA_signal_6150), .B0_t (stateArray_outS31ser[5]), .B0_f (new_AGEMA_signal_3082), .B1_t (new_AGEMA_signal_3083), .B1_f (new_AGEMA_signal_3084), .Z0_t (MixColumns_line3_S02[6]), .Z0_f (new_AGEMA_signal_3157), .Z1_t (new_AGEMA_signal_3158), .Z1_f (new_AGEMA_signal_3159) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S30reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS31ser[6]), .A0_f (new_AGEMA_signal_3091), .A1_t (new_AGEMA_signal_3092), .A1_f (new_AGEMA_signal_3093), .B0_t (stateArray_outS33ser[6]), .B0_f (new_AGEMA_signal_3094), .B1_t (new_AGEMA_signal_3095), .B1_f (new_AGEMA_signal_3096), .Z0_t (stateArray_S30reg_gff_1_SFF_6_MUXInst_X), .Z0_f (new_AGEMA_signal_3097), .Z1_t (new_AGEMA_signal_3098), .Z1_f (new_AGEMA_signal_3099) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S30reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S30reg_gff_1_SFF_6_MUXInst_X), .B0_f (new_AGEMA_signal_3097), .B1_t (new_AGEMA_signal_3098), .B1_f (new_AGEMA_signal_3099), .Z0_t (stateArray_S30reg_gff_1_SFF_6_MUXInst_Y), .Z0_f (new_AGEMA_signal_6151), .Z1_t (new_AGEMA_signal_6152), .Z1_f (new_AGEMA_signal_6153) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S30reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (stateArray_S30reg_gff_1_SFF_6_MUXInst_Y), .A0_f (new_AGEMA_signal_6151), .A1_t (new_AGEMA_signal_6152), .A1_f (new_AGEMA_signal_6153), .B0_t (stateArray_outS31ser[6]), .B0_f (new_AGEMA_signal_3091), .B1_t (new_AGEMA_signal_3092), .B1_f (new_AGEMA_signal_3093), .Z0_t (MixColumns_line3_S02[7]), .Z0_f (new_AGEMA_signal_3166), .Z1_t (new_AGEMA_signal_3167), .Z1_f (new_AGEMA_signal_3168) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S30reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS31ser[7]), .A0_f (new_AGEMA_signal_3100), .A1_t (new_AGEMA_signal_3101), .A1_f (new_AGEMA_signal_3102), .B0_t (stateArray_outS33ser[7]), .B0_f (new_AGEMA_signal_3103), .B1_t (new_AGEMA_signal_3104), .B1_f (new_AGEMA_signal_3105), .Z0_t (stateArray_S30reg_gff_1_SFF_7_MUXInst_X), .Z0_f (new_AGEMA_signal_3106), .Z1_t (new_AGEMA_signal_3107), .Z1_f (new_AGEMA_signal_3108) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S30reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S30reg_gff_1_SFF_7_MUXInst_X), .B0_f (new_AGEMA_signal_3106), .B1_t (new_AGEMA_signal_3107), .B1_f (new_AGEMA_signal_3108), .Z0_t (stateArray_S30reg_gff_1_SFF_7_MUXInst_Y), .Z0_f (new_AGEMA_signal_6154), .Z1_t (new_AGEMA_signal_6155), .Z1_f (new_AGEMA_signal_6156) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S30reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (stateArray_S30reg_gff_1_SFF_7_MUXInst_Y), .A0_f (new_AGEMA_signal_6154), .A1_t (new_AGEMA_signal_6155), .A1_f (new_AGEMA_signal_6156), .B0_t (stateArray_outS31ser[7]), .B0_f (new_AGEMA_signal_3100), .B1_t (new_AGEMA_signal_3101), .B1_f (new_AGEMA_signal_3102), .Z0_t (MixColumns_line3_S02[0]), .Z0_f (new_AGEMA_signal_3175), .Z1_t (new_AGEMA_signal_3176), .Z1_f (new_AGEMA_signal_3177) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S31reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS32ser[0]), .A0_f (new_AGEMA_signal_3109), .A1_t (new_AGEMA_signal_3110), .A1_f (new_AGEMA_signal_3111), .B0_t (MCin[0]), .B0_f (new_AGEMA_signal_3112), .B1_t (new_AGEMA_signal_3113), .B1_f (new_AGEMA_signal_3114), .Z0_t (stateArray_S31reg_gff_1_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_3115), .Z1_t (new_AGEMA_signal_3116), .Z1_f (new_AGEMA_signal_3117) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S31reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S31reg_gff_1_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_3115), .B1_t (new_AGEMA_signal_3116), .B1_f (new_AGEMA_signal_3117), .Z0_t (stateArray_S31reg_gff_1_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_6157), .Z1_t (new_AGEMA_signal_6158), .Z1_f (new_AGEMA_signal_6159) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S31reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (stateArray_S31reg_gff_1_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_6157), .A1_t (new_AGEMA_signal_6158), .A1_f (new_AGEMA_signal_6159), .B0_t (stateArray_outS32ser[0]), .B0_f (new_AGEMA_signal_3109), .B1_t (new_AGEMA_signal_3110), .B1_f (new_AGEMA_signal_3111), .Z0_t (stateArray_outS31ser[0]), .Z0_f (new_AGEMA_signal_3037), .Z1_t (new_AGEMA_signal_3038), .Z1_f (new_AGEMA_signal_3039) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S31reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS32ser[1]), .A0_f (new_AGEMA_signal_3118), .A1_t (new_AGEMA_signal_3119), .A1_f (new_AGEMA_signal_3120), .B0_t (MixColumns_line3_S02[2]), .B0_f (new_AGEMA_signal_3121), .B1_t (new_AGEMA_signal_3122), .B1_f (new_AGEMA_signal_3123), .Z0_t (stateArray_S31reg_gff_1_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_3124), .Z1_t (new_AGEMA_signal_3125), .Z1_f (new_AGEMA_signal_3126) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S31reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S31reg_gff_1_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_3124), .B1_t (new_AGEMA_signal_3125), .B1_f (new_AGEMA_signal_3126), .Z0_t (stateArray_S31reg_gff_1_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_6160), .Z1_t (new_AGEMA_signal_6161), .Z1_f (new_AGEMA_signal_6162) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S31reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (stateArray_S31reg_gff_1_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_6160), .A1_t (new_AGEMA_signal_6161), .A1_f (new_AGEMA_signal_6162), .B0_t (stateArray_outS32ser[1]), .B0_f (new_AGEMA_signal_3118), .B1_t (new_AGEMA_signal_3119), .B1_f (new_AGEMA_signal_3120), .Z0_t (stateArray_outS31ser[1]), .Z0_f (new_AGEMA_signal_3046), .Z1_t (new_AGEMA_signal_3047), .Z1_f (new_AGEMA_signal_3048) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S31reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS32ser[2]), .A0_f (new_AGEMA_signal_3127), .A1_t (new_AGEMA_signal_3128), .A1_f (new_AGEMA_signal_3129), .B0_t (MCin[2]), .B0_f (new_AGEMA_signal_3130), .B1_t (new_AGEMA_signal_3131), .B1_f (new_AGEMA_signal_3132), .Z0_t (stateArray_S31reg_gff_1_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_3133), .Z1_t (new_AGEMA_signal_3134), .Z1_f (new_AGEMA_signal_3135) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S31reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S31reg_gff_1_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_3133), .B1_t (new_AGEMA_signal_3134), .B1_f (new_AGEMA_signal_3135), .Z0_t (stateArray_S31reg_gff_1_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_6163), .Z1_t (new_AGEMA_signal_6164), .Z1_f (new_AGEMA_signal_6165) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S31reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (stateArray_S31reg_gff_1_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_6163), .A1_t (new_AGEMA_signal_6164), .A1_f (new_AGEMA_signal_6165), .B0_t (stateArray_outS32ser[2]), .B0_f (new_AGEMA_signal_3127), .B1_t (new_AGEMA_signal_3128), .B1_f (new_AGEMA_signal_3129), .Z0_t (stateArray_outS31ser[2]), .Z0_f (new_AGEMA_signal_3055), .Z1_t (new_AGEMA_signal_3056), .Z1_f (new_AGEMA_signal_3057) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S31reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS32ser[3]), .A0_f (new_AGEMA_signal_3136), .A1_t (new_AGEMA_signal_3137), .A1_f (new_AGEMA_signal_3138), .B0_t (MCin[3]), .B0_f (new_AGEMA_signal_3139), .B1_t (new_AGEMA_signal_3140), .B1_f (new_AGEMA_signal_3141), .Z0_t (stateArray_S31reg_gff_1_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_3142), .Z1_t (new_AGEMA_signal_3143), .Z1_f (new_AGEMA_signal_3144) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S31reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S31reg_gff_1_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_3142), .B1_t (new_AGEMA_signal_3143), .B1_f (new_AGEMA_signal_3144), .Z0_t (stateArray_S31reg_gff_1_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_6166), .Z1_t (new_AGEMA_signal_6167), .Z1_f (new_AGEMA_signal_6168) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S31reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (stateArray_S31reg_gff_1_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_6166), .A1_t (new_AGEMA_signal_6167), .A1_f (new_AGEMA_signal_6168), .B0_t (stateArray_outS32ser[3]), .B0_f (new_AGEMA_signal_3136), .B1_t (new_AGEMA_signal_3137), .B1_f (new_AGEMA_signal_3138), .Z0_t (stateArray_outS31ser[3]), .Z0_f (new_AGEMA_signal_3064), .Z1_t (new_AGEMA_signal_3065), .Z1_f (new_AGEMA_signal_3066) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S31reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS32ser[4]), .A0_f (new_AGEMA_signal_3145), .A1_t (new_AGEMA_signal_3146), .A1_f (new_AGEMA_signal_3147), .B0_t (MixColumns_line3_S02[5]), .B0_f (new_AGEMA_signal_3148), .B1_t (new_AGEMA_signal_3149), .B1_f (new_AGEMA_signal_3150), .Z0_t (stateArray_S31reg_gff_1_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_3151), .Z1_t (new_AGEMA_signal_3152), .Z1_f (new_AGEMA_signal_3153) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S31reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S31reg_gff_1_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_3151), .B1_t (new_AGEMA_signal_3152), .B1_f (new_AGEMA_signal_3153), .Z0_t (stateArray_S31reg_gff_1_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_6169), .Z1_t (new_AGEMA_signal_6170), .Z1_f (new_AGEMA_signal_6171) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S31reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (stateArray_S31reg_gff_1_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_6169), .A1_t (new_AGEMA_signal_6170), .A1_f (new_AGEMA_signal_6171), .B0_t (stateArray_outS32ser[4]), .B0_f (new_AGEMA_signal_3145), .B1_t (new_AGEMA_signal_3146), .B1_f (new_AGEMA_signal_3147), .Z0_t (stateArray_outS31ser[4]), .Z0_f (new_AGEMA_signal_3073), .Z1_t (new_AGEMA_signal_3074), .Z1_f (new_AGEMA_signal_3075) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S31reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS32ser[5]), .A0_f (new_AGEMA_signal_3154), .A1_t (new_AGEMA_signal_3155), .A1_f (new_AGEMA_signal_3156), .B0_t (MixColumns_line3_S02[6]), .B0_f (new_AGEMA_signal_3157), .B1_t (new_AGEMA_signal_3158), .B1_f (new_AGEMA_signal_3159), .Z0_t (stateArray_S31reg_gff_1_SFF_5_MUXInst_X), .Z0_f (new_AGEMA_signal_3160), .Z1_t (new_AGEMA_signal_3161), .Z1_f (new_AGEMA_signal_3162) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S31reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S31reg_gff_1_SFF_5_MUXInst_X), .B0_f (new_AGEMA_signal_3160), .B1_t (new_AGEMA_signal_3161), .B1_f (new_AGEMA_signal_3162), .Z0_t (stateArray_S31reg_gff_1_SFF_5_MUXInst_Y), .Z0_f (new_AGEMA_signal_6172), .Z1_t (new_AGEMA_signal_6173), .Z1_f (new_AGEMA_signal_6174) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S31reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (stateArray_S31reg_gff_1_SFF_5_MUXInst_Y), .A0_f (new_AGEMA_signal_6172), .A1_t (new_AGEMA_signal_6173), .A1_f (new_AGEMA_signal_6174), .B0_t (stateArray_outS32ser[5]), .B0_f (new_AGEMA_signal_3154), .B1_t (new_AGEMA_signal_3155), .B1_f (new_AGEMA_signal_3156), .Z0_t (stateArray_outS31ser[5]), .Z0_f (new_AGEMA_signal_3082), .Z1_t (new_AGEMA_signal_3083), .Z1_f (new_AGEMA_signal_3084) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S31reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS32ser[6]), .A0_f (new_AGEMA_signal_3163), .A1_t (new_AGEMA_signal_3164), .A1_f (new_AGEMA_signal_3165), .B0_t (MixColumns_line3_S02[7]), .B0_f (new_AGEMA_signal_3166), .B1_t (new_AGEMA_signal_3167), .B1_f (new_AGEMA_signal_3168), .Z0_t (stateArray_S31reg_gff_1_SFF_6_MUXInst_X), .Z0_f (new_AGEMA_signal_3169), .Z1_t (new_AGEMA_signal_3170), .Z1_f (new_AGEMA_signal_3171) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S31reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S31reg_gff_1_SFF_6_MUXInst_X), .B0_f (new_AGEMA_signal_3169), .B1_t (new_AGEMA_signal_3170), .B1_f (new_AGEMA_signal_3171), .Z0_t (stateArray_S31reg_gff_1_SFF_6_MUXInst_Y), .Z0_f (new_AGEMA_signal_6175), .Z1_t (new_AGEMA_signal_6176), .Z1_f (new_AGEMA_signal_6177) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S31reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (stateArray_S31reg_gff_1_SFF_6_MUXInst_Y), .A0_f (new_AGEMA_signal_6175), .A1_t (new_AGEMA_signal_6176), .A1_f (new_AGEMA_signal_6177), .B0_t (stateArray_outS32ser[6]), .B0_f (new_AGEMA_signal_3163), .B1_t (new_AGEMA_signal_3164), .B1_f (new_AGEMA_signal_3165), .Z0_t (stateArray_outS31ser[6]), .Z0_f (new_AGEMA_signal_3091), .Z1_t (new_AGEMA_signal_3092), .Z1_f (new_AGEMA_signal_3093) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S31reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS32ser[7]), .A0_f (new_AGEMA_signal_3172), .A1_t (new_AGEMA_signal_3173), .A1_f (new_AGEMA_signal_3174), .B0_t (MixColumns_line3_S02[0]), .B0_f (new_AGEMA_signal_3175), .B1_t (new_AGEMA_signal_3176), .B1_f (new_AGEMA_signal_3177), .Z0_t (stateArray_S31reg_gff_1_SFF_7_MUXInst_X), .Z0_f (new_AGEMA_signal_3178), .Z1_t (new_AGEMA_signal_3179), .Z1_f (new_AGEMA_signal_3180) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S31reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S31reg_gff_1_SFF_7_MUXInst_X), .B0_f (new_AGEMA_signal_3178), .B1_t (new_AGEMA_signal_3179), .B1_f (new_AGEMA_signal_3180), .Z0_t (stateArray_S31reg_gff_1_SFF_7_MUXInst_Y), .Z0_f (new_AGEMA_signal_6178), .Z1_t (new_AGEMA_signal_6179), .Z1_f (new_AGEMA_signal_6180) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S31reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (stateArray_S31reg_gff_1_SFF_7_MUXInst_Y), .A0_f (new_AGEMA_signal_6178), .A1_t (new_AGEMA_signal_6179), .A1_f (new_AGEMA_signal_6180), .B0_t (stateArray_outS32ser[7]), .B0_f (new_AGEMA_signal_3172), .B1_t (new_AGEMA_signal_3173), .B1_f (new_AGEMA_signal_3174), .Z0_t (stateArray_outS31ser[7]), .Z0_f (new_AGEMA_signal_3100), .Z1_t (new_AGEMA_signal_3101), .Z1_f (new_AGEMA_signal_3102) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S32reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS33ser[0]), .A0_f (new_AGEMA_signal_3040), .A1_t (new_AGEMA_signal_3041), .A1_f (new_AGEMA_signal_3042), .B0_t (stateArray_outS31ser[0]), .B0_f (new_AGEMA_signal_3037), .B1_t (new_AGEMA_signal_3038), .B1_f (new_AGEMA_signal_3039), .Z0_t (stateArray_S32reg_gff_1_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_3181), .Z1_t (new_AGEMA_signal_3182), .Z1_f (new_AGEMA_signal_3183) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S32reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S32reg_gff_1_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_3181), .B1_t (new_AGEMA_signal_3182), .B1_f (new_AGEMA_signal_3183), .Z0_t (stateArray_S32reg_gff_1_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_6181), .Z1_t (new_AGEMA_signal_6182), .Z1_f (new_AGEMA_signal_6183) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S32reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (stateArray_S32reg_gff_1_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_6181), .A1_t (new_AGEMA_signal_6182), .A1_f (new_AGEMA_signal_6183), .B0_t (stateArray_outS33ser[0]), .B0_f (new_AGEMA_signal_3040), .B1_t (new_AGEMA_signal_3041), .B1_f (new_AGEMA_signal_3042), .Z0_t (stateArray_outS32ser[0]), .Z0_f (new_AGEMA_signal_3109), .Z1_t (new_AGEMA_signal_3110), .Z1_f (new_AGEMA_signal_3111) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S32reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS33ser[1]), .A0_f (new_AGEMA_signal_3049), .A1_t (new_AGEMA_signal_3050), .A1_f (new_AGEMA_signal_3051), .B0_t (stateArray_outS31ser[1]), .B0_f (new_AGEMA_signal_3046), .B1_t (new_AGEMA_signal_3047), .B1_f (new_AGEMA_signal_3048), .Z0_t (stateArray_S32reg_gff_1_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_3184), .Z1_t (new_AGEMA_signal_3185), .Z1_f (new_AGEMA_signal_3186) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S32reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S32reg_gff_1_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_3184), .B1_t (new_AGEMA_signal_3185), .B1_f (new_AGEMA_signal_3186), .Z0_t (stateArray_S32reg_gff_1_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_6184), .Z1_t (new_AGEMA_signal_6185), .Z1_f (new_AGEMA_signal_6186) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S32reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (stateArray_S32reg_gff_1_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_6184), .A1_t (new_AGEMA_signal_6185), .A1_f (new_AGEMA_signal_6186), .B0_t (stateArray_outS33ser[1]), .B0_f (new_AGEMA_signal_3049), .B1_t (new_AGEMA_signal_3050), .B1_f (new_AGEMA_signal_3051), .Z0_t (stateArray_outS32ser[1]), .Z0_f (new_AGEMA_signal_3118), .Z1_t (new_AGEMA_signal_3119), .Z1_f (new_AGEMA_signal_3120) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S32reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS33ser[2]), .A0_f (new_AGEMA_signal_3058), .A1_t (new_AGEMA_signal_3059), .A1_f (new_AGEMA_signal_3060), .B0_t (stateArray_outS31ser[2]), .B0_f (new_AGEMA_signal_3055), .B1_t (new_AGEMA_signal_3056), .B1_f (new_AGEMA_signal_3057), .Z0_t (stateArray_S32reg_gff_1_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_3187), .Z1_t (new_AGEMA_signal_3188), .Z1_f (new_AGEMA_signal_3189) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S32reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S32reg_gff_1_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_3187), .B1_t (new_AGEMA_signal_3188), .B1_f (new_AGEMA_signal_3189), .Z0_t (stateArray_S32reg_gff_1_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_6187), .Z1_t (new_AGEMA_signal_6188), .Z1_f (new_AGEMA_signal_6189) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S32reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (stateArray_S32reg_gff_1_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_6187), .A1_t (new_AGEMA_signal_6188), .A1_f (new_AGEMA_signal_6189), .B0_t (stateArray_outS33ser[2]), .B0_f (new_AGEMA_signal_3058), .B1_t (new_AGEMA_signal_3059), .B1_f (new_AGEMA_signal_3060), .Z0_t (stateArray_outS32ser[2]), .Z0_f (new_AGEMA_signal_3127), .Z1_t (new_AGEMA_signal_3128), .Z1_f (new_AGEMA_signal_3129) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S32reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS33ser[3]), .A0_f (new_AGEMA_signal_3067), .A1_t (new_AGEMA_signal_3068), .A1_f (new_AGEMA_signal_3069), .B0_t (stateArray_outS31ser[3]), .B0_f (new_AGEMA_signal_3064), .B1_t (new_AGEMA_signal_3065), .B1_f (new_AGEMA_signal_3066), .Z0_t (stateArray_S32reg_gff_1_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_3190), .Z1_t (new_AGEMA_signal_3191), .Z1_f (new_AGEMA_signal_3192) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S32reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S32reg_gff_1_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_3190), .B1_t (new_AGEMA_signal_3191), .B1_f (new_AGEMA_signal_3192), .Z0_t (stateArray_S32reg_gff_1_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_6190), .Z1_t (new_AGEMA_signal_6191), .Z1_f (new_AGEMA_signal_6192) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S32reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (stateArray_S32reg_gff_1_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_6190), .A1_t (new_AGEMA_signal_6191), .A1_f (new_AGEMA_signal_6192), .B0_t (stateArray_outS33ser[3]), .B0_f (new_AGEMA_signal_3067), .B1_t (new_AGEMA_signal_3068), .B1_f (new_AGEMA_signal_3069), .Z0_t (stateArray_outS32ser[3]), .Z0_f (new_AGEMA_signal_3136), .Z1_t (new_AGEMA_signal_3137), .Z1_f (new_AGEMA_signal_3138) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S32reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS33ser[4]), .A0_f (new_AGEMA_signal_3076), .A1_t (new_AGEMA_signal_3077), .A1_f (new_AGEMA_signal_3078), .B0_t (stateArray_outS31ser[4]), .B0_f (new_AGEMA_signal_3073), .B1_t (new_AGEMA_signal_3074), .B1_f (new_AGEMA_signal_3075), .Z0_t (stateArray_S32reg_gff_1_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_3193), .Z1_t (new_AGEMA_signal_3194), .Z1_f (new_AGEMA_signal_3195) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S32reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S32reg_gff_1_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_3193), .B1_t (new_AGEMA_signal_3194), .B1_f (new_AGEMA_signal_3195), .Z0_t (stateArray_S32reg_gff_1_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_6193), .Z1_t (new_AGEMA_signal_6194), .Z1_f (new_AGEMA_signal_6195) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S32reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (stateArray_S32reg_gff_1_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_6193), .A1_t (new_AGEMA_signal_6194), .A1_f (new_AGEMA_signal_6195), .B0_t (stateArray_outS33ser[4]), .B0_f (new_AGEMA_signal_3076), .B1_t (new_AGEMA_signal_3077), .B1_f (new_AGEMA_signal_3078), .Z0_t (stateArray_outS32ser[4]), .Z0_f (new_AGEMA_signal_3145), .Z1_t (new_AGEMA_signal_3146), .Z1_f (new_AGEMA_signal_3147) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S32reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS33ser[5]), .A0_f (new_AGEMA_signal_3085), .A1_t (new_AGEMA_signal_3086), .A1_f (new_AGEMA_signal_3087), .B0_t (stateArray_outS31ser[5]), .B0_f (new_AGEMA_signal_3082), .B1_t (new_AGEMA_signal_3083), .B1_f (new_AGEMA_signal_3084), .Z0_t (stateArray_S32reg_gff_1_SFF_5_MUXInst_X), .Z0_f (new_AGEMA_signal_3196), .Z1_t (new_AGEMA_signal_3197), .Z1_f (new_AGEMA_signal_3198) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S32reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S32reg_gff_1_SFF_5_MUXInst_X), .B0_f (new_AGEMA_signal_3196), .B1_t (new_AGEMA_signal_3197), .B1_f (new_AGEMA_signal_3198), .Z0_t (stateArray_S32reg_gff_1_SFF_5_MUXInst_Y), .Z0_f (new_AGEMA_signal_6196), .Z1_t (new_AGEMA_signal_6197), .Z1_f (new_AGEMA_signal_6198) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S32reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (stateArray_S32reg_gff_1_SFF_5_MUXInst_Y), .A0_f (new_AGEMA_signal_6196), .A1_t (new_AGEMA_signal_6197), .A1_f (new_AGEMA_signal_6198), .B0_t (stateArray_outS33ser[5]), .B0_f (new_AGEMA_signal_3085), .B1_t (new_AGEMA_signal_3086), .B1_f (new_AGEMA_signal_3087), .Z0_t (stateArray_outS32ser[5]), .Z0_f (new_AGEMA_signal_3154), .Z1_t (new_AGEMA_signal_3155), .Z1_f (new_AGEMA_signal_3156) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S32reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS33ser[6]), .A0_f (new_AGEMA_signal_3094), .A1_t (new_AGEMA_signal_3095), .A1_f (new_AGEMA_signal_3096), .B0_t (stateArray_outS31ser[6]), .B0_f (new_AGEMA_signal_3091), .B1_t (new_AGEMA_signal_3092), .B1_f (new_AGEMA_signal_3093), .Z0_t (stateArray_S32reg_gff_1_SFF_6_MUXInst_X), .Z0_f (new_AGEMA_signal_3199), .Z1_t (new_AGEMA_signal_3200), .Z1_f (new_AGEMA_signal_3201) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S32reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S32reg_gff_1_SFF_6_MUXInst_X), .B0_f (new_AGEMA_signal_3199), .B1_t (new_AGEMA_signal_3200), .B1_f (new_AGEMA_signal_3201), .Z0_t (stateArray_S32reg_gff_1_SFF_6_MUXInst_Y), .Z0_f (new_AGEMA_signal_6199), .Z1_t (new_AGEMA_signal_6200), .Z1_f (new_AGEMA_signal_6201) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S32reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (stateArray_S32reg_gff_1_SFF_6_MUXInst_Y), .A0_f (new_AGEMA_signal_6199), .A1_t (new_AGEMA_signal_6200), .A1_f (new_AGEMA_signal_6201), .B0_t (stateArray_outS33ser[6]), .B0_f (new_AGEMA_signal_3094), .B1_t (new_AGEMA_signal_3095), .B1_f (new_AGEMA_signal_3096), .Z0_t (stateArray_outS32ser[6]), .Z0_f (new_AGEMA_signal_3163), .Z1_t (new_AGEMA_signal_3164), .Z1_f (new_AGEMA_signal_3165) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S32reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (stateArray_outS33ser[7]), .A0_f (new_AGEMA_signal_3103), .A1_t (new_AGEMA_signal_3104), .A1_f (new_AGEMA_signal_3105), .B0_t (stateArray_outS31ser[7]), .B0_f (new_AGEMA_signal_3100), .B1_t (new_AGEMA_signal_3101), .B1_f (new_AGEMA_signal_3102), .Z0_t (stateArray_S32reg_gff_1_SFF_7_MUXInst_X), .Z0_f (new_AGEMA_signal_3202), .Z1_t (new_AGEMA_signal_3203), .Z1_f (new_AGEMA_signal_3204) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S32reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S32reg_gff_1_SFF_7_MUXInst_X), .B0_f (new_AGEMA_signal_3202), .B1_t (new_AGEMA_signal_3203), .B1_f (new_AGEMA_signal_3204), .Z0_t (stateArray_S32reg_gff_1_SFF_7_MUXInst_Y), .Z0_f (new_AGEMA_signal_6202), .Z1_t (new_AGEMA_signal_6203), .Z1_f (new_AGEMA_signal_6204) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S32reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (stateArray_S32reg_gff_1_SFF_7_MUXInst_Y), .A0_f (new_AGEMA_signal_6202), .A1_t (new_AGEMA_signal_6203), .A1_f (new_AGEMA_signal_6204), .B0_t (stateArray_outS33ser[7]), .B0_f (new_AGEMA_signal_3103), .B1_t (new_AGEMA_signal_3104), .B1_f (new_AGEMA_signal_3105), .Z0_t (stateArray_outS32ser[7]), .Z0_f (new_AGEMA_signal_3172), .Z1_t (new_AGEMA_signal_3173), .Z1_f (new_AGEMA_signal_3174) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S33reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS33ser[0]), .A0_f (new_AGEMA_signal_7865), .A1_t (new_AGEMA_signal_7866), .A1_f (new_AGEMA_signal_7867), .B0_t (stateArray_outS32ser[0]), .B0_f (new_AGEMA_signal_3109), .B1_t (new_AGEMA_signal_3110), .B1_f (new_AGEMA_signal_3111), .Z0_t (stateArray_S33reg_gff_1_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_7889), .Z1_t (new_AGEMA_signal_7890), .Z1_f (new_AGEMA_signal_7891) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S33reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S33reg_gff_1_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_7889), .B1_t (new_AGEMA_signal_7890), .B1_f (new_AGEMA_signal_7891), .Z0_t (stateArray_S33reg_gff_1_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_7913), .Z1_t (new_AGEMA_signal_7914), .Z1_f (new_AGEMA_signal_7915) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S33reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (stateArray_S33reg_gff_1_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_7913), .A1_t (new_AGEMA_signal_7914), .A1_f (new_AGEMA_signal_7915), .B0_t (stateArray_inS33ser[0]), .B0_f (new_AGEMA_signal_7865), .B1_t (new_AGEMA_signal_7866), .B1_f (new_AGEMA_signal_7867), .Z0_t (stateArray_outS33ser[0]), .Z0_f (new_AGEMA_signal_3040), .Z1_t (new_AGEMA_signal_3041), .Z1_f (new_AGEMA_signal_3042) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S33reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS33ser[1]), .A0_f (new_AGEMA_signal_7892), .A1_t (new_AGEMA_signal_7893), .A1_f (new_AGEMA_signal_7894), .B0_t (stateArray_outS32ser[1]), .B0_f (new_AGEMA_signal_3118), .B1_t (new_AGEMA_signal_3119), .B1_f (new_AGEMA_signal_3120), .Z0_t (stateArray_S33reg_gff_1_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_7916), .Z1_t (new_AGEMA_signal_7917), .Z1_f (new_AGEMA_signal_7918) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S33reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S33reg_gff_1_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_7916), .B1_t (new_AGEMA_signal_7917), .B1_f (new_AGEMA_signal_7918), .Z0_t (stateArray_S33reg_gff_1_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_7937), .Z1_t (new_AGEMA_signal_7938), .Z1_f (new_AGEMA_signal_7939) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S33reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (stateArray_S33reg_gff_1_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_7937), .A1_t (new_AGEMA_signal_7938), .A1_f (new_AGEMA_signal_7939), .B0_t (stateArray_inS33ser[1]), .B0_f (new_AGEMA_signal_7892), .B1_t (new_AGEMA_signal_7893), .B1_f (new_AGEMA_signal_7894), .Z0_t (stateArray_outS33ser[1]), .Z0_f (new_AGEMA_signal_3049), .Z1_t (new_AGEMA_signal_3050), .Z1_f (new_AGEMA_signal_3051) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S33reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS33ser[2]), .A0_f (new_AGEMA_signal_7895), .A1_t (new_AGEMA_signal_7896), .A1_f (new_AGEMA_signal_7897), .B0_t (stateArray_outS32ser[2]), .B0_f (new_AGEMA_signal_3127), .B1_t (new_AGEMA_signal_3128), .B1_f (new_AGEMA_signal_3129), .Z0_t (stateArray_S33reg_gff_1_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_7919), .Z1_t (new_AGEMA_signal_7920), .Z1_f (new_AGEMA_signal_7921) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S33reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S33reg_gff_1_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_7919), .B1_t (new_AGEMA_signal_7920), .B1_f (new_AGEMA_signal_7921), .Z0_t (stateArray_S33reg_gff_1_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_7940), .Z1_t (new_AGEMA_signal_7941), .Z1_f (new_AGEMA_signal_7942) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S33reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (stateArray_S33reg_gff_1_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_7940), .A1_t (new_AGEMA_signal_7941), .A1_f (new_AGEMA_signal_7942), .B0_t (stateArray_inS33ser[2]), .B0_f (new_AGEMA_signal_7895), .B1_t (new_AGEMA_signal_7896), .B1_f (new_AGEMA_signal_7897), .Z0_t (stateArray_outS33ser[2]), .Z0_f (new_AGEMA_signal_3058), .Z1_t (new_AGEMA_signal_3059), .Z1_f (new_AGEMA_signal_3060) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S33reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS33ser[3]), .A0_f (new_AGEMA_signal_7898), .A1_t (new_AGEMA_signal_7899), .A1_f (new_AGEMA_signal_7900), .B0_t (stateArray_outS32ser[3]), .B0_f (new_AGEMA_signal_3136), .B1_t (new_AGEMA_signal_3137), .B1_f (new_AGEMA_signal_3138), .Z0_t (stateArray_S33reg_gff_1_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_7922), .Z1_t (new_AGEMA_signal_7923), .Z1_f (new_AGEMA_signal_7924) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S33reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S33reg_gff_1_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_7922), .B1_t (new_AGEMA_signal_7923), .B1_f (new_AGEMA_signal_7924), .Z0_t (stateArray_S33reg_gff_1_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_7943), .Z1_t (new_AGEMA_signal_7944), .Z1_f (new_AGEMA_signal_7945) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S33reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (stateArray_S33reg_gff_1_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_7943), .A1_t (new_AGEMA_signal_7944), .A1_f (new_AGEMA_signal_7945), .B0_t (stateArray_inS33ser[3]), .B0_f (new_AGEMA_signal_7898), .B1_t (new_AGEMA_signal_7899), .B1_f (new_AGEMA_signal_7900), .Z0_t (stateArray_outS33ser[3]), .Z0_f (new_AGEMA_signal_3067), .Z1_t (new_AGEMA_signal_3068), .Z1_f (new_AGEMA_signal_3069) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S33reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS33ser[4]), .A0_f (new_AGEMA_signal_7901), .A1_t (new_AGEMA_signal_7902), .A1_f (new_AGEMA_signal_7903), .B0_t (stateArray_outS32ser[4]), .B0_f (new_AGEMA_signal_3145), .B1_t (new_AGEMA_signal_3146), .B1_f (new_AGEMA_signal_3147), .Z0_t (stateArray_S33reg_gff_1_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_7925), .Z1_t (new_AGEMA_signal_7926), .Z1_f (new_AGEMA_signal_7927) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S33reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S33reg_gff_1_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_7925), .B1_t (new_AGEMA_signal_7926), .B1_f (new_AGEMA_signal_7927), .Z0_t (stateArray_S33reg_gff_1_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_7946), .Z1_t (new_AGEMA_signal_7947), .Z1_f (new_AGEMA_signal_7948) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S33reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (stateArray_S33reg_gff_1_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_7946), .A1_t (new_AGEMA_signal_7947), .A1_f (new_AGEMA_signal_7948), .B0_t (stateArray_inS33ser[4]), .B0_f (new_AGEMA_signal_7901), .B1_t (new_AGEMA_signal_7902), .B1_f (new_AGEMA_signal_7903), .Z0_t (stateArray_outS33ser[4]), .Z0_f (new_AGEMA_signal_3076), .Z1_t (new_AGEMA_signal_3077), .Z1_f (new_AGEMA_signal_3078) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S33reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS33ser[5]), .A0_f (new_AGEMA_signal_7904), .A1_t (new_AGEMA_signal_7905), .A1_f (new_AGEMA_signal_7906), .B0_t (stateArray_outS32ser[5]), .B0_f (new_AGEMA_signal_3154), .B1_t (new_AGEMA_signal_3155), .B1_f (new_AGEMA_signal_3156), .Z0_t (stateArray_S33reg_gff_1_SFF_5_MUXInst_X), .Z0_f (new_AGEMA_signal_7928), .Z1_t (new_AGEMA_signal_7929), .Z1_f (new_AGEMA_signal_7930) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S33reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S33reg_gff_1_SFF_5_MUXInst_X), .B0_f (new_AGEMA_signal_7928), .B1_t (new_AGEMA_signal_7929), .B1_f (new_AGEMA_signal_7930), .Z0_t (stateArray_S33reg_gff_1_SFF_5_MUXInst_Y), .Z0_f (new_AGEMA_signal_7949), .Z1_t (new_AGEMA_signal_7950), .Z1_f (new_AGEMA_signal_7951) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S33reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (stateArray_S33reg_gff_1_SFF_5_MUXInst_Y), .A0_f (new_AGEMA_signal_7949), .A1_t (new_AGEMA_signal_7950), .A1_f (new_AGEMA_signal_7951), .B0_t (stateArray_inS33ser[5]), .B0_f (new_AGEMA_signal_7904), .B1_t (new_AGEMA_signal_7905), .B1_f (new_AGEMA_signal_7906), .Z0_t (stateArray_outS33ser[5]), .Z0_f (new_AGEMA_signal_3085), .Z1_t (new_AGEMA_signal_3086), .Z1_f (new_AGEMA_signal_3087) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S33reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS33ser[6]), .A0_f (new_AGEMA_signal_7907), .A1_t (new_AGEMA_signal_7908), .A1_f (new_AGEMA_signal_7909), .B0_t (stateArray_outS32ser[6]), .B0_f (new_AGEMA_signal_3163), .B1_t (new_AGEMA_signal_3164), .B1_f (new_AGEMA_signal_3165), .Z0_t (stateArray_S33reg_gff_1_SFF_6_MUXInst_X), .Z0_f (new_AGEMA_signal_7931), .Z1_t (new_AGEMA_signal_7932), .Z1_f (new_AGEMA_signal_7933) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S33reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S33reg_gff_1_SFF_6_MUXInst_X), .B0_f (new_AGEMA_signal_7931), .B1_t (new_AGEMA_signal_7932), .B1_f (new_AGEMA_signal_7933), .Z0_t (stateArray_S33reg_gff_1_SFF_6_MUXInst_Y), .Z0_f (new_AGEMA_signal_7952), .Z1_t (new_AGEMA_signal_7953), .Z1_f (new_AGEMA_signal_7954) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S33reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (stateArray_S33reg_gff_1_SFF_6_MUXInst_Y), .A0_f (new_AGEMA_signal_7952), .A1_t (new_AGEMA_signal_7953), .A1_f (new_AGEMA_signal_7954), .B0_t (stateArray_inS33ser[6]), .B0_f (new_AGEMA_signal_7907), .B1_t (new_AGEMA_signal_7908), .B1_f (new_AGEMA_signal_7909), .Z0_t (stateArray_outS33ser[6]), .Z0_f (new_AGEMA_signal_3094), .Z1_t (new_AGEMA_signal_3095), .Z1_f (new_AGEMA_signal_3096) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S33reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (stateArray_inS33ser[7]), .A0_f (new_AGEMA_signal_7910), .A1_t (new_AGEMA_signal_7911), .A1_f (new_AGEMA_signal_7912), .B0_t (stateArray_outS32ser[7]), .B0_f (new_AGEMA_signal_3172), .B1_t (new_AGEMA_signal_3173), .B1_f (new_AGEMA_signal_3174), .Z0_t (stateArray_S33reg_gff_1_SFF_7_MUXInst_X), .Z0_f (new_AGEMA_signal_7934), .Z1_t (new_AGEMA_signal_7935), .Z1_f (new_AGEMA_signal_7936) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_S33reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (ctrl_n4), .A1_f (new_AGEMA_signal_5778), .B0_t (stateArray_S33reg_gff_1_SFF_7_MUXInst_X), .B0_f (new_AGEMA_signal_7934), .B1_t (new_AGEMA_signal_7935), .B1_f (new_AGEMA_signal_7936), .Z0_t (stateArray_S33reg_gff_1_SFF_7_MUXInst_Y), .Z0_f (new_AGEMA_signal_7955), .Z1_t (new_AGEMA_signal_7956), .Z1_f (new_AGEMA_signal_7957) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateArray_S33reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (stateArray_S33reg_gff_1_SFF_7_MUXInst_Y), .A0_f (new_AGEMA_signal_7955), .A1_t (new_AGEMA_signal_7956), .A1_f (new_AGEMA_signal_7957), .B0_t (stateArray_inS33ser[7]), .B0_f (new_AGEMA_signal_7910), .B1_t (new_AGEMA_signal_7911), .B1_f (new_AGEMA_signal_7912), .Z0_t (stateArray_outS33ser[7]), .Z0_f (new_AGEMA_signal_3103), .Z1_t (new_AGEMA_signal_3104), .Z1_f (new_AGEMA_signal_3105) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_0_XOR1_U1 ( .A0_t (MCin[16]), .A0_f (new_AGEMA_signal_3988), .A1_t (new_AGEMA_signal_3989), .A1_f (new_AGEMA_signal_3990), .B0_t (StateInMC[24]), .B0_f (new_AGEMA_signal_5536), .B1_t (new_AGEMA_signal_5537), .B1_f (new_AGEMA_signal_5538), .Z0_t (stateArray_MUX_inS03ser_mux_inst_0_X), .Z0_f (new_AGEMA_signal_5633), .Z1_t (new_AGEMA_signal_5634), .Z1_f (new_AGEMA_signal_5635) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_0_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (stateArray_nReset_selMC), .A1_f (new_AGEMA_signal_4210), .B0_t (stateArray_MUX_inS03ser_mux_inst_0_X), .B0_f (new_AGEMA_signal_5633), .B1_t (new_AGEMA_signal_5634), .B1_f (new_AGEMA_signal_5635), .Z0_t (stateArray_MUX_inS03ser_mux_inst_0_Y), .Z0_f (new_AGEMA_signal_5793), .Z1_t (new_AGEMA_signal_5794), .Z1_f (new_AGEMA_signal_5795) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_0_XOR2_U1 ( .A0_t (stateArray_MUX_inS03ser_mux_inst_0_Y), .A0_f (new_AGEMA_signal_5793), .A1_t (new_AGEMA_signal_5794), .A1_f (new_AGEMA_signal_5795), .B0_t (MCin[16]), .B0_f (new_AGEMA_signal_3988), .B1_t (new_AGEMA_signal_3989), .B1_f (new_AGEMA_signal_3990), .Z0_t (stateArray_inS03ser[0]), .Z0_f (new_AGEMA_signal_6205), .Z1_t (new_AGEMA_signal_6206), .Z1_f (new_AGEMA_signal_6207) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_1_XOR1_U1 ( .A0_t (MixColumns_line1_S02[2]), .A0_f (new_AGEMA_signal_3982), .A1_t (new_AGEMA_signal_3983), .A1_f (new_AGEMA_signal_3984), .B0_t (StateInMC[25]), .B0_f (new_AGEMA_signal_5705), .B1_t (new_AGEMA_signal_5706), .B1_f (new_AGEMA_signal_5707), .Z0_t (stateArray_MUX_inS03ser_mux_inst_1_X), .Z0_f (new_AGEMA_signal_5796), .Z1_t (new_AGEMA_signal_5797), .Z1_f (new_AGEMA_signal_5798) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (stateArray_nReset_selMC), .A1_f (new_AGEMA_signal_4210), .B0_t (stateArray_MUX_inS03ser_mux_inst_1_X), .B0_f (new_AGEMA_signal_5796), .B1_t (new_AGEMA_signal_5797), .B1_f (new_AGEMA_signal_5798), .Z0_t (stateArray_MUX_inS03ser_mux_inst_1_Y), .Z0_f (new_AGEMA_signal_6208), .Z1_t (new_AGEMA_signal_6209), .Z1_f (new_AGEMA_signal_6210) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_1_XOR2_U1 ( .A0_t (stateArray_MUX_inS03ser_mux_inst_1_Y), .A0_f (new_AGEMA_signal_6208), .A1_t (new_AGEMA_signal_6209), .A1_f (new_AGEMA_signal_6210), .B0_t (MixColumns_line1_S02[2]), .B0_f (new_AGEMA_signal_3982), .B1_t (new_AGEMA_signal_3983), .B1_f (new_AGEMA_signal_3984), .Z0_t (stateArray_inS03ser[1]), .Z0_f (new_AGEMA_signal_6364), .Z1_t (new_AGEMA_signal_6365), .Z1_f (new_AGEMA_signal_6366) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_2_XOR1_U1 ( .A0_t (MCin[18]), .A0_f (new_AGEMA_signal_3979), .A1_t (new_AGEMA_signal_3980), .A1_f (new_AGEMA_signal_3981), .B0_t (StateInMC[26]), .B0_f (new_AGEMA_signal_5542), .B1_t (new_AGEMA_signal_5543), .B1_f (new_AGEMA_signal_5544), .Z0_t (stateArray_MUX_inS03ser_mux_inst_2_X), .Z0_f (new_AGEMA_signal_5636), .Z1_t (new_AGEMA_signal_5637), .Z1_f (new_AGEMA_signal_5638) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_2_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (stateArray_nReset_selMC), .A1_f (new_AGEMA_signal_4210), .B0_t (stateArray_MUX_inS03ser_mux_inst_2_X), .B0_f (new_AGEMA_signal_5636), .B1_t (new_AGEMA_signal_5637), .B1_f (new_AGEMA_signal_5638), .Z0_t (stateArray_MUX_inS03ser_mux_inst_2_Y), .Z0_f (new_AGEMA_signal_5799), .Z1_t (new_AGEMA_signal_5800), .Z1_f (new_AGEMA_signal_5801) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_2_XOR2_U1 ( .A0_t (stateArray_MUX_inS03ser_mux_inst_2_Y), .A0_f (new_AGEMA_signal_5799), .A1_t (new_AGEMA_signal_5800), .A1_f (new_AGEMA_signal_5801), .B0_t (MCin[18]), .B0_f (new_AGEMA_signal_3979), .B1_t (new_AGEMA_signal_3980), .B1_f (new_AGEMA_signal_3981), .Z0_t (stateArray_inS03ser[2]), .Z0_f (new_AGEMA_signal_6211), .Z1_t (new_AGEMA_signal_6212), .Z1_f (new_AGEMA_signal_6213) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_3_XOR1_U1 ( .A0_t (MCin[19]), .A0_f (new_AGEMA_signal_3994), .A1_t (new_AGEMA_signal_3995), .A1_f (new_AGEMA_signal_3996), .B0_t (StateInMC[27]), .B0_f (new_AGEMA_signal_5708), .B1_t (new_AGEMA_signal_5709), .B1_f (new_AGEMA_signal_5710), .Z0_t (stateArray_MUX_inS03ser_mux_inst_3_X), .Z0_f (new_AGEMA_signal_5802), .Z1_t (new_AGEMA_signal_5803), .Z1_f (new_AGEMA_signal_5804) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_3_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (stateArray_nReset_selMC), .A1_f (new_AGEMA_signal_4210), .B0_t (stateArray_MUX_inS03ser_mux_inst_3_X), .B0_f (new_AGEMA_signal_5802), .B1_t (new_AGEMA_signal_5803), .B1_f (new_AGEMA_signal_5804), .Z0_t (stateArray_MUX_inS03ser_mux_inst_3_Y), .Z0_f (new_AGEMA_signal_6214), .Z1_t (new_AGEMA_signal_6215), .Z1_f (new_AGEMA_signal_6216) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_3_XOR2_U1 ( .A0_t (stateArray_MUX_inS03ser_mux_inst_3_Y), .A0_f (new_AGEMA_signal_6214), .A1_t (new_AGEMA_signal_6215), .A1_f (new_AGEMA_signal_6216), .B0_t (MCin[19]), .B0_f (new_AGEMA_signal_3994), .B1_t (new_AGEMA_signal_3995), .B1_f (new_AGEMA_signal_3996), .Z0_t (stateArray_inS03ser[3]), .Z0_f (new_AGEMA_signal_6367), .Z1_t (new_AGEMA_signal_6368), .Z1_f (new_AGEMA_signal_6369) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_4_XOR1_U1 ( .A0_t (MixColumns_line1_S02[5]), .A0_f (new_AGEMA_signal_3973), .A1_t (new_AGEMA_signal_3974), .A1_f (new_AGEMA_signal_3975), .B0_t (StateInMC[28]), .B0_f (new_AGEMA_signal_5711), .B1_t (new_AGEMA_signal_5712), .B1_f (new_AGEMA_signal_5713), .Z0_t (stateArray_MUX_inS03ser_mux_inst_4_X), .Z0_f (new_AGEMA_signal_5805), .Z1_t (new_AGEMA_signal_5806), .Z1_f (new_AGEMA_signal_5807) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_4_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (stateArray_nReset_selMC), .A1_f (new_AGEMA_signal_4210), .B0_t (stateArray_MUX_inS03ser_mux_inst_4_X), .B0_f (new_AGEMA_signal_5805), .B1_t (new_AGEMA_signal_5806), .B1_f (new_AGEMA_signal_5807), .Z0_t (stateArray_MUX_inS03ser_mux_inst_4_Y), .Z0_f (new_AGEMA_signal_6217), .Z1_t (new_AGEMA_signal_6218), .Z1_f (new_AGEMA_signal_6219) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_4_XOR2_U1 ( .A0_t (stateArray_MUX_inS03ser_mux_inst_4_Y), .A0_f (new_AGEMA_signal_6217), .A1_t (new_AGEMA_signal_6218), .A1_f (new_AGEMA_signal_6219), .B0_t (MixColumns_line1_S02[5]), .B0_f (new_AGEMA_signal_3973), .B1_t (new_AGEMA_signal_3974), .B1_f (new_AGEMA_signal_3975), .Z0_t (stateArray_inS03ser[4]), .Z0_f (new_AGEMA_signal_6370), .Z1_t (new_AGEMA_signal_6371), .Z1_f (new_AGEMA_signal_6372) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_5_XOR1_U1 ( .A0_t (MixColumns_line1_S02[6]), .A0_f (new_AGEMA_signal_3967), .A1_t (new_AGEMA_signal_3968), .A1_f (new_AGEMA_signal_3969), .B0_t (StateInMC[29]), .B0_f (new_AGEMA_signal_5551), .B1_t (new_AGEMA_signal_5552), .B1_f (new_AGEMA_signal_5553), .Z0_t (stateArray_MUX_inS03ser_mux_inst_5_X), .Z0_f (new_AGEMA_signal_5639), .Z1_t (new_AGEMA_signal_5640), .Z1_f (new_AGEMA_signal_5641) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_5_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (stateArray_nReset_selMC), .A1_f (new_AGEMA_signal_4210), .B0_t (stateArray_MUX_inS03ser_mux_inst_5_X), .B0_f (new_AGEMA_signal_5639), .B1_t (new_AGEMA_signal_5640), .B1_f (new_AGEMA_signal_5641), .Z0_t (stateArray_MUX_inS03ser_mux_inst_5_Y), .Z0_f (new_AGEMA_signal_5808), .Z1_t (new_AGEMA_signal_5809), .Z1_f (new_AGEMA_signal_5810) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_5_XOR2_U1 ( .A0_t (stateArray_MUX_inS03ser_mux_inst_5_Y), .A0_f (new_AGEMA_signal_5808), .A1_t (new_AGEMA_signal_5809), .A1_f (new_AGEMA_signal_5810), .B0_t (MixColumns_line1_S02[6]), .B0_f (new_AGEMA_signal_3967), .B1_t (new_AGEMA_signal_3968), .B1_f (new_AGEMA_signal_3969), .Z0_t (stateArray_inS03ser[5]), .Z0_f (new_AGEMA_signal_6220), .Z1_t (new_AGEMA_signal_6221), .Z1_f (new_AGEMA_signal_6222) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_6_XOR1_U1 ( .A0_t (MixColumns_line1_S02[7]), .A0_f (new_AGEMA_signal_3961), .A1_t (new_AGEMA_signal_3962), .A1_f (new_AGEMA_signal_3963), .B0_t (StateInMC[30]), .B0_f (new_AGEMA_signal_5554), .B1_t (new_AGEMA_signal_5555), .B1_f (new_AGEMA_signal_5556), .Z0_t (stateArray_MUX_inS03ser_mux_inst_6_X), .Z0_f (new_AGEMA_signal_5642), .Z1_t (new_AGEMA_signal_5643), .Z1_f (new_AGEMA_signal_5644) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_6_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (stateArray_nReset_selMC), .A1_f (new_AGEMA_signal_4210), .B0_t (stateArray_MUX_inS03ser_mux_inst_6_X), .B0_f (new_AGEMA_signal_5642), .B1_t (new_AGEMA_signal_5643), .B1_f (new_AGEMA_signal_5644), .Z0_t (stateArray_MUX_inS03ser_mux_inst_6_Y), .Z0_f (new_AGEMA_signal_5811), .Z1_t (new_AGEMA_signal_5812), .Z1_f (new_AGEMA_signal_5813) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_6_XOR2_U1 ( .A0_t (stateArray_MUX_inS03ser_mux_inst_6_Y), .A0_f (new_AGEMA_signal_5811), .A1_t (new_AGEMA_signal_5812), .A1_f (new_AGEMA_signal_5813), .B0_t (MixColumns_line1_S02[7]), .B0_f (new_AGEMA_signal_3961), .B1_t (new_AGEMA_signal_3962), .B1_f (new_AGEMA_signal_3963), .Z0_t (stateArray_inS03ser[6]), .Z0_f (new_AGEMA_signal_6223), .Z1_t (new_AGEMA_signal_6224), .Z1_f (new_AGEMA_signal_6225) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_7_XOR1_U1 ( .A0_t (MixColumns_line1_S02[0]), .A0_f (new_AGEMA_signal_3958), .A1_t (new_AGEMA_signal_3959), .A1_f (new_AGEMA_signal_3960), .B0_t (StateInMC[31]), .B0_f (new_AGEMA_signal_5557), .B1_t (new_AGEMA_signal_5558), .B1_f (new_AGEMA_signal_5559), .Z0_t (stateArray_MUX_inS03ser_mux_inst_7_X), .Z0_f (new_AGEMA_signal_5645), .Z1_t (new_AGEMA_signal_5646), .Z1_f (new_AGEMA_signal_5647) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_7_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (stateArray_nReset_selMC), .A1_f (new_AGEMA_signal_4210), .B0_t (stateArray_MUX_inS03ser_mux_inst_7_X), .B0_f (new_AGEMA_signal_5645), .B1_t (new_AGEMA_signal_5646), .B1_f (new_AGEMA_signal_5647), .Z0_t (stateArray_MUX_inS03ser_mux_inst_7_Y), .Z0_f (new_AGEMA_signal_5814), .Z1_t (new_AGEMA_signal_5815), .Z1_f (new_AGEMA_signal_5816) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS03ser_mux_inst_7_XOR2_U1 ( .A0_t (stateArray_MUX_inS03ser_mux_inst_7_Y), .A0_f (new_AGEMA_signal_5814), .A1_t (new_AGEMA_signal_5815), .A1_f (new_AGEMA_signal_5816), .B0_t (MixColumns_line1_S02[0]), .B0_f (new_AGEMA_signal_3958), .B1_t (new_AGEMA_signal_3959), .B1_f (new_AGEMA_signal_3960), .Z0_t (stateArray_inS03ser[7]), .Z0_f (new_AGEMA_signal_6226), .Z1_t (new_AGEMA_signal_6227), .Z1_f (new_AGEMA_signal_6228) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_0_XOR1_U1 ( .A0_t (MCin[8]), .A0_f (new_AGEMA_signal_2989), .A1_t (new_AGEMA_signal_2990), .A1_f (new_AGEMA_signal_2991), .B0_t (StateInMC[16]), .B0_f (new_AGEMA_signal_5512), .B1_t (new_AGEMA_signal_5513), .B1_f (new_AGEMA_signal_5514), .Z0_t (stateArray_MUX_inS13ser_mux_inst_0_X), .Z0_f (new_AGEMA_signal_5648), .Z1_t (new_AGEMA_signal_5649), .Z1_f (new_AGEMA_signal_5650) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_0_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (stateArray_nReset_selMC), .A1_f (new_AGEMA_signal_4210), .B0_t (stateArray_MUX_inS13ser_mux_inst_0_X), .B0_f (new_AGEMA_signal_5648), .B1_t (new_AGEMA_signal_5649), .B1_f (new_AGEMA_signal_5650), .Z0_t (stateArray_MUX_inS13ser_mux_inst_0_Y), .Z0_f (new_AGEMA_signal_5817), .Z1_t (new_AGEMA_signal_5818), .Z1_f (new_AGEMA_signal_5819) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_0_XOR2_U1 ( .A0_t (stateArray_MUX_inS13ser_mux_inst_0_Y), .A0_f (new_AGEMA_signal_5817), .A1_t (new_AGEMA_signal_5818), .A1_f (new_AGEMA_signal_5819), .B0_t (MCin[8]), .B0_f (new_AGEMA_signal_2989), .B1_t (new_AGEMA_signal_2990), .B1_f (new_AGEMA_signal_2991), .Z0_t (stateArray_inS13ser[0]), .Z0_f (new_AGEMA_signal_6229), .Z1_t (new_AGEMA_signal_6230), .Z1_f (new_AGEMA_signal_6231) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_1_XOR1_U1 ( .A0_t (MixColumns_line2_S02[2]), .A0_f (new_AGEMA_signal_2995), .A1_t (new_AGEMA_signal_2996), .A1_f (new_AGEMA_signal_2997), .B0_t (StateInMC[17]), .B0_f (new_AGEMA_signal_5696), .B1_t (new_AGEMA_signal_5697), .B1_f (new_AGEMA_signal_5698), .Z0_t (stateArray_MUX_inS13ser_mux_inst_1_X), .Z0_f (new_AGEMA_signal_5820), .Z1_t (new_AGEMA_signal_5821), .Z1_f (new_AGEMA_signal_5822) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (stateArray_nReset_selMC), .A1_f (new_AGEMA_signal_4210), .B0_t (stateArray_MUX_inS13ser_mux_inst_1_X), .B0_f (new_AGEMA_signal_5820), .B1_t (new_AGEMA_signal_5821), .B1_f (new_AGEMA_signal_5822), .Z0_t (stateArray_MUX_inS13ser_mux_inst_1_Y), .Z0_f (new_AGEMA_signal_6232), .Z1_t (new_AGEMA_signal_6233), .Z1_f (new_AGEMA_signal_6234) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_1_XOR2_U1 ( .A0_t (stateArray_MUX_inS13ser_mux_inst_1_Y), .A0_f (new_AGEMA_signal_6232), .A1_t (new_AGEMA_signal_6233), .A1_f (new_AGEMA_signal_6234), .B0_t (MixColumns_line2_S02[2]), .B0_f (new_AGEMA_signal_2995), .B1_t (new_AGEMA_signal_2996), .B1_f (new_AGEMA_signal_2997), .Z0_t (stateArray_inS13ser[1]), .Z0_f (new_AGEMA_signal_6373), .Z1_t (new_AGEMA_signal_6374), .Z1_f (new_AGEMA_signal_6375) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_2_XOR1_U1 ( .A0_t (MCin[10]), .A0_f (new_AGEMA_signal_3001), .A1_t (new_AGEMA_signal_3002), .A1_f (new_AGEMA_signal_3003), .B0_t (StateInMC[18]), .B0_f (new_AGEMA_signal_5518), .B1_t (new_AGEMA_signal_5519), .B1_f (new_AGEMA_signal_5520), .Z0_t (stateArray_MUX_inS13ser_mux_inst_2_X), .Z0_f (new_AGEMA_signal_5651), .Z1_t (new_AGEMA_signal_5652), .Z1_f (new_AGEMA_signal_5653) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_2_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (stateArray_nReset_selMC), .A1_f (new_AGEMA_signal_4210), .B0_t (stateArray_MUX_inS13ser_mux_inst_2_X), .B0_f (new_AGEMA_signal_5651), .B1_t (new_AGEMA_signal_5652), .B1_f (new_AGEMA_signal_5653), .Z0_t (stateArray_MUX_inS13ser_mux_inst_2_Y), .Z0_f (new_AGEMA_signal_5823), .Z1_t (new_AGEMA_signal_5824), .Z1_f (new_AGEMA_signal_5825) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_2_XOR2_U1 ( .A0_t (stateArray_MUX_inS13ser_mux_inst_2_Y), .A0_f (new_AGEMA_signal_5823), .A1_t (new_AGEMA_signal_5824), .A1_f (new_AGEMA_signal_5825), .B0_t (MCin[10]), .B0_f (new_AGEMA_signal_3001), .B1_t (new_AGEMA_signal_3002), .B1_f (new_AGEMA_signal_3003), .Z0_t (stateArray_inS13ser[2]), .Z0_f (new_AGEMA_signal_6235), .Z1_t (new_AGEMA_signal_6236), .Z1_f (new_AGEMA_signal_6237) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_3_XOR1_U1 ( .A0_t (MCin[11]), .A0_f (new_AGEMA_signal_3007), .A1_t (new_AGEMA_signal_3008), .A1_f (new_AGEMA_signal_3009), .B0_t (StateInMC[19]), .B0_f (new_AGEMA_signal_5699), .B1_t (new_AGEMA_signal_5700), .B1_f (new_AGEMA_signal_5701), .Z0_t (stateArray_MUX_inS13ser_mux_inst_3_X), .Z0_f (new_AGEMA_signal_5826), .Z1_t (new_AGEMA_signal_5827), .Z1_f (new_AGEMA_signal_5828) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_3_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (stateArray_nReset_selMC), .A1_f (new_AGEMA_signal_4210), .B0_t (stateArray_MUX_inS13ser_mux_inst_3_X), .B0_f (new_AGEMA_signal_5826), .B1_t (new_AGEMA_signal_5827), .B1_f (new_AGEMA_signal_5828), .Z0_t (stateArray_MUX_inS13ser_mux_inst_3_Y), .Z0_f (new_AGEMA_signal_6238), .Z1_t (new_AGEMA_signal_6239), .Z1_f (new_AGEMA_signal_6240) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_3_XOR2_U1 ( .A0_t (stateArray_MUX_inS13ser_mux_inst_3_Y), .A0_f (new_AGEMA_signal_6238), .A1_t (new_AGEMA_signal_6239), .A1_f (new_AGEMA_signal_6240), .B0_t (MCin[11]), .B0_f (new_AGEMA_signal_3007), .B1_t (new_AGEMA_signal_3008), .B1_f (new_AGEMA_signal_3009), .Z0_t (stateArray_inS13ser[3]), .Z0_f (new_AGEMA_signal_6376), .Z1_t (new_AGEMA_signal_6377), .Z1_f (new_AGEMA_signal_6378) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_4_XOR1_U1 ( .A0_t (MixColumns_line2_S02[5]), .A0_f (new_AGEMA_signal_3013), .A1_t (new_AGEMA_signal_3014), .A1_f (new_AGEMA_signal_3015), .B0_t (StateInMC[20]), .B0_f (new_AGEMA_signal_5702), .B1_t (new_AGEMA_signal_5703), .B1_f (new_AGEMA_signal_5704), .Z0_t (stateArray_MUX_inS13ser_mux_inst_4_X), .Z0_f (new_AGEMA_signal_5829), .Z1_t (new_AGEMA_signal_5830), .Z1_f (new_AGEMA_signal_5831) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_4_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (stateArray_nReset_selMC), .A1_f (new_AGEMA_signal_4210), .B0_t (stateArray_MUX_inS13ser_mux_inst_4_X), .B0_f (new_AGEMA_signal_5829), .B1_t (new_AGEMA_signal_5830), .B1_f (new_AGEMA_signal_5831), .Z0_t (stateArray_MUX_inS13ser_mux_inst_4_Y), .Z0_f (new_AGEMA_signal_6241), .Z1_t (new_AGEMA_signal_6242), .Z1_f (new_AGEMA_signal_6243) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_4_XOR2_U1 ( .A0_t (stateArray_MUX_inS13ser_mux_inst_4_Y), .A0_f (new_AGEMA_signal_6241), .A1_t (new_AGEMA_signal_6242), .A1_f (new_AGEMA_signal_6243), .B0_t (MixColumns_line2_S02[5]), .B0_f (new_AGEMA_signal_3013), .B1_t (new_AGEMA_signal_3014), .B1_f (new_AGEMA_signal_3015), .Z0_t (stateArray_inS13ser[4]), .Z0_f (new_AGEMA_signal_6379), .Z1_t (new_AGEMA_signal_6380), .Z1_f (new_AGEMA_signal_6381) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_5_XOR1_U1 ( .A0_t (MixColumns_line2_S02[6]), .A0_f (new_AGEMA_signal_3019), .A1_t (new_AGEMA_signal_3020), .A1_f (new_AGEMA_signal_3021), .B0_t (StateInMC[21]), .B0_f (new_AGEMA_signal_5527), .B1_t (new_AGEMA_signal_5528), .B1_f (new_AGEMA_signal_5529), .Z0_t (stateArray_MUX_inS13ser_mux_inst_5_X), .Z0_f (new_AGEMA_signal_5654), .Z1_t (new_AGEMA_signal_5655), .Z1_f (new_AGEMA_signal_5656) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_5_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (stateArray_nReset_selMC), .A1_f (new_AGEMA_signal_4210), .B0_t (stateArray_MUX_inS13ser_mux_inst_5_X), .B0_f (new_AGEMA_signal_5654), .B1_t (new_AGEMA_signal_5655), .B1_f (new_AGEMA_signal_5656), .Z0_t (stateArray_MUX_inS13ser_mux_inst_5_Y), .Z0_f (new_AGEMA_signal_5832), .Z1_t (new_AGEMA_signal_5833), .Z1_f (new_AGEMA_signal_5834) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_5_XOR2_U1 ( .A0_t (stateArray_MUX_inS13ser_mux_inst_5_Y), .A0_f (new_AGEMA_signal_5832), .A1_t (new_AGEMA_signal_5833), .A1_f (new_AGEMA_signal_5834), .B0_t (MixColumns_line2_S02[6]), .B0_f (new_AGEMA_signal_3019), .B1_t (new_AGEMA_signal_3020), .B1_f (new_AGEMA_signal_3021), .Z0_t (stateArray_inS13ser[5]), .Z0_f (new_AGEMA_signal_6244), .Z1_t (new_AGEMA_signal_6245), .Z1_f (new_AGEMA_signal_6246) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_6_XOR1_U1 ( .A0_t (MixColumns_line2_S02[7]), .A0_f (new_AGEMA_signal_3025), .A1_t (new_AGEMA_signal_3026), .A1_f (new_AGEMA_signal_3027), .B0_t (StateInMC[22]), .B0_f (new_AGEMA_signal_5530), .B1_t (new_AGEMA_signal_5531), .B1_f (new_AGEMA_signal_5532), .Z0_t (stateArray_MUX_inS13ser_mux_inst_6_X), .Z0_f (new_AGEMA_signal_5657), .Z1_t (new_AGEMA_signal_5658), .Z1_f (new_AGEMA_signal_5659) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_6_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (stateArray_nReset_selMC), .A1_f (new_AGEMA_signal_4210), .B0_t (stateArray_MUX_inS13ser_mux_inst_6_X), .B0_f (new_AGEMA_signal_5657), .B1_t (new_AGEMA_signal_5658), .B1_f (new_AGEMA_signal_5659), .Z0_t (stateArray_MUX_inS13ser_mux_inst_6_Y), .Z0_f (new_AGEMA_signal_5835), .Z1_t (new_AGEMA_signal_5836), .Z1_f (new_AGEMA_signal_5837) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_6_XOR2_U1 ( .A0_t (stateArray_MUX_inS13ser_mux_inst_6_Y), .A0_f (new_AGEMA_signal_5835), .A1_t (new_AGEMA_signal_5836), .A1_f (new_AGEMA_signal_5837), .B0_t (MixColumns_line2_S02[7]), .B0_f (new_AGEMA_signal_3025), .B1_t (new_AGEMA_signal_3026), .B1_f (new_AGEMA_signal_3027), .Z0_t (stateArray_inS13ser[6]), .Z0_f (new_AGEMA_signal_6247), .Z1_t (new_AGEMA_signal_6248), .Z1_f (new_AGEMA_signal_6249) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_7_XOR1_U1 ( .A0_t (MixColumns_line2_S02[0]), .A0_f (new_AGEMA_signal_3031), .A1_t (new_AGEMA_signal_3032), .A1_f (new_AGEMA_signal_3033), .B0_t (StateInMC[23]), .B0_f (new_AGEMA_signal_5533), .B1_t (new_AGEMA_signal_5534), .B1_f (new_AGEMA_signal_5535), .Z0_t (stateArray_MUX_inS13ser_mux_inst_7_X), .Z0_f (new_AGEMA_signal_5660), .Z1_t (new_AGEMA_signal_5661), .Z1_f (new_AGEMA_signal_5662) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_7_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (stateArray_nReset_selMC), .A1_f (new_AGEMA_signal_4210), .B0_t (stateArray_MUX_inS13ser_mux_inst_7_X), .B0_f (new_AGEMA_signal_5660), .B1_t (new_AGEMA_signal_5661), .B1_f (new_AGEMA_signal_5662), .Z0_t (stateArray_MUX_inS13ser_mux_inst_7_Y), .Z0_f (new_AGEMA_signal_5838), .Z1_t (new_AGEMA_signal_5839), .Z1_f (new_AGEMA_signal_5840) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS13ser_mux_inst_7_XOR2_U1 ( .A0_t (stateArray_MUX_inS13ser_mux_inst_7_Y), .A0_f (new_AGEMA_signal_5838), .A1_t (new_AGEMA_signal_5839), .A1_f (new_AGEMA_signal_5840), .B0_t (MixColumns_line2_S02[0]), .B0_f (new_AGEMA_signal_3031), .B1_t (new_AGEMA_signal_3032), .B1_f (new_AGEMA_signal_3033), .Z0_t (stateArray_inS13ser[7]), .Z0_f (new_AGEMA_signal_6250), .Z1_t (new_AGEMA_signal_6251), .Z1_f (new_AGEMA_signal_6252) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_0_XOR1_U1 ( .A0_t (MCin[0]), .A0_f (new_AGEMA_signal_3112), .A1_t (new_AGEMA_signal_3113), .A1_f (new_AGEMA_signal_3114), .B0_t (StateInMC[8]), .B0_f (new_AGEMA_signal_5488), .B1_t (new_AGEMA_signal_5489), .B1_f (new_AGEMA_signal_5490), .Z0_t (stateArray_MUX_inS23ser_mux_inst_0_X), .Z0_f (new_AGEMA_signal_5663), .Z1_t (new_AGEMA_signal_5664), .Z1_f (new_AGEMA_signal_5665) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_0_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (stateArray_nReset_selMC), .A1_f (new_AGEMA_signal_4210), .B0_t (stateArray_MUX_inS23ser_mux_inst_0_X), .B0_f (new_AGEMA_signal_5663), .B1_t (new_AGEMA_signal_5664), .B1_f (new_AGEMA_signal_5665), .Z0_t (stateArray_MUX_inS23ser_mux_inst_0_Y), .Z0_f (new_AGEMA_signal_5841), .Z1_t (new_AGEMA_signal_5842), .Z1_f (new_AGEMA_signal_5843) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_0_XOR2_U1 ( .A0_t (stateArray_MUX_inS23ser_mux_inst_0_Y), .A0_f (new_AGEMA_signal_5841), .A1_t (new_AGEMA_signal_5842), .A1_f (new_AGEMA_signal_5843), .B0_t (MCin[0]), .B0_f (new_AGEMA_signal_3112), .B1_t (new_AGEMA_signal_3113), .B1_f (new_AGEMA_signal_3114), .Z0_t (stateArray_inS23ser[0]), .Z0_f (new_AGEMA_signal_6253), .Z1_t (new_AGEMA_signal_6254), .Z1_f (new_AGEMA_signal_6255) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_1_XOR1_U1 ( .A0_t (MixColumns_line3_S02[2]), .A0_f (new_AGEMA_signal_3121), .A1_t (new_AGEMA_signal_3122), .A1_f (new_AGEMA_signal_3123), .B0_t (StateInMC[9]), .B0_f (new_AGEMA_signal_5687), .B1_t (new_AGEMA_signal_5688), .B1_f (new_AGEMA_signal_5689), .Z0_t (stateArray_MUX_inS23ser_mux_inst_1_X), .Z0_f (new_AGEMA_signal_5844), .Z1_t (new_AGEMA_signal_5845), .Z1_f (new_AGEMA_signal_5846) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (stateArray_nReset_selMC), .A1_f (new_AGEMA_signal_4210), .B0_t (stateArray_MUX_inS23ser_mux_inst_1_X), .B0_f (new_AGEMA_signal_5844), .B1_t (new_AGEMA_signal_5845), .B1_f (new_AGEMA_signal_5846), .Z0_t (stateArray_MUX_inS23ser_mux_inst_1_Y), .Z0_f (new_AGEMA_signal_6256), .Z1_t (new_AGEMA_signal_6257), .Z1_f (new_AGEMA_signal_6258) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_1_XOR2_U1 ( .A0_t (stateArray_MUX_inS23ser_mux_inst_1_Y), .A0_f (new_AGEMA_signal_6256), .A1_t (new_AGEMA_signal_6257), .A1_f (new_AGEMA_signal_6258), .B0_t (MixColumns_line3_S02[2]), .B0_f (new_AGEMA_signal_3121), .B1_t (new_AGEMA_signal_3122), .B1_f (new_AGEMA_signal_3123), .Z0_t (stateArray_inS23ser[1]), .Z0_f (new_AGEMA_signal_6382), .Z1_t (new_AGEMA_signal_6383), .Z1_f (new_AGEMA_signal_6384) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_2_XOR1_U1 ( .A0_t (MCin[2]), .A0_f (new_AGEMA_signal_3130), .A1_t (new_AGEMA_signal_3131), .A1_f (new_AGEMA_signal_3132), .B0_t (StateInMC[10]), .B0_f (new_AGEMA_signal_5494), .B1_t (new_AGEMA_signal_5495), .B1_f (new_AGEMA_signal_5496), .Z0_t (stateArray_MUX_inS23ser_mux_inst_2_X), .Z0_f (new_AGEMA_signal_5666), .Z1_t (new_AGEMA_signal_5667), .Z1_f (new_AGEMA_signal_5668) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_2_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (stateArray_nReset_selMC), .A1_f (new_AGEMA_signal_4210), .B0_t (stateArray_MUX_inS23ser_mux_inst_2_X), .B0_f (new_AGEMA_signal_5666), .B1_t (new_AGEMA_signal_5667), .B1_f (new_AGEMA_signal_5668), .Z0_t (stateArray_MUX_inS23ser_mux_inst_2_Y), .Z0_f (new_AGEMA_signal_5847), .Z1_t (new_AGEMA_signal_5848), .Z1_f (new_AGEMA_signal_5849) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_2_XOR2_U1 ( .A0_t (stateArray_MUX_inS23ser_mux_inst_2_Y), .A0_f (new_AGEMA_signal_5847), .A1_t (new_AGEMA_signal_5848), .A1_f (new_AGEMA_signal_5849), .B0_t (MCin[2]), .B0_f (new_AGEMA_signal_3130), .B1_t (new_AGEMA_signal_3131), .B1_f (new_AGEMA_signal_3132), .Z0_t (stateArray_inS23ser[2]), .Z0_f (new_AGEMA_signal_6259), .Z1_t (new_AGEMA_signal_6260), .Z1_f (new_AGEMA_signal_6261) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_3_XOR1_U1 ( .A0_t (MCin[3]), .A0_f (new_AGEMA_signal_3139), .A1_t (new_AGEMA_signal_3140), .A1_f (new_AGEMA_signal_3141), .B0_t (StateInMC[11]), .B0_f (new_AGEMA_signal_5690), .B1_t (new_AGEMA_signal_5691), .B1_f (new_AGEMA_signal_5692), .Z0_t (stateArray_MUX_inS23ser_mux_inst_3_X), .Z0_f (new_AGEMA_signal_5850), .Z1_t (new_AGEMA_signal_5851), .Z1_f (new_AGEMA_signal_5852) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_3_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (stateArray_nReset_selMC), .A1_f (new_AGEMA_signal_4210), .B0_t (stateArray_MUX_inS23ser_mux_inst_3_X), .B0_f (new_AGEMA_signal_5850), .B1_t (new_AGEMA_signal_5851), .B1_f (new_AGEMA_signal_5852), .Z0_t (stateArray_MUX_inS23ser_mux_inst_3_Y), .Z0_f (new_AGEMA_signal_6262), .Z1_t (new_AGEMA_signal_6263), .Z1_f (new_AGEMA_signal_6264) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_3_XOR2_U1 ( .A0_t (stateArray_MUX_inS23ser_mux_inst_3_Y), .A0_f (new_AGEMA_signal_6262), .A1_t (new_AGEMA_signal_6263), .A1_f (new_AGEMA_signal_6264), .B0_t (MCin[3]), .B0_f (new_AGEMA_signal_3139), .B1_t (new_AGEMA_signal_3140), .B1_f (new_AGEMA_signal_3141), .Z0_t (stateArray_inS23ser[3]), .Z0_f (new_AGEMA_signal_6385), .Z1_t (new_AGEMA_signal_6386), .Z1_f (new_AGEMA_signal_6387) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_4_XOR1_U1 ( .A0_t (MixColumns_line3_S02[5]), .A0_f (new_AGEMA_signal_3148), .A1_t (new_AGEMA_signal_3149), .A1_f (new_AGEMA_signal_3150), .B0_t (StateInMC[12]), .B0_f (new_AGEMA_signal_5693), .B1_t (new_AGEMA_signal_5694), .B1_f (new_AGEMA_signal_5695), .Z0_t (stateArray_MUX_inS23ser_mux_inst_4_X), .Z0_f (new_AGEMA_signal_5853), .Z1_t (new_AGEMA_signal_5854), .Z1_f (new_AGEMA_signal_5855) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_4_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (stateArray_nReset_selMC), .A1_f (new_AGEMA_signal_4210), .B0_t (stateArray_MUX_inS23ser_mux_inst_4_X), .B0_f (new_AGEMA_signal_5853), .B1_t (new_AGEMA_signal_5854), .B1_f (new_AGEMA_signal_5855), .Z0_t (stateArray_MUX_inS23ser_mux_inst_4_Y), .Z0_f (new_AGEMA_signal_6265), .Z1_t (new_AGEMA_signal_6266), .Z1_f (new_AGEMA_signal_6267) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_4_XOR2_U1 ( .A0_t (stateArray_MUX_inS23ser_mux_inst_4_Y), .A0_f (new_AGEMA_signal_6265), .A1_t (new_AGEMA_signal_6266), .A1_f (new_AGEMA_signal_6267), .B0_t (MixColumns_line3_S02[5]), .B0_f (new_AGEMA_signal_3148), .B1_t (new_AGEMA_signal_3149), .B1_f (new_AGEMA_signal_3150), .Z0_t (stateArray_inS23ser[4]), .Z0_f (new_AGEMA_signal_6388), .Z1_t (new_AGEMA_signal_6389), .Z1_f (new_AGEMA_signal_6390) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_5_XOR1_U1 ( .A0_t (MixColumns_line3_S02[6]), .A0_f (new_AGEMA_signal_3157), .A1_t (new_AGEMA_signal_3158), .A1_f (new_AGEMA_signal_3159), .B0_t (StateInMC[13]), .B0_f (new_AGEMA_signal_5503), .B1_t (new_AGEMA_signal_5504), .B1_f (new_AGEMA_signal_5505), .Z0_t (stateArray_MUX_inS23ser_mux_inst_5_X), .Z0_f (new_AGEMA_signal_5669), .Z1_t (new_AGEMA_signal_5670), .Z1_f (new_AGEMA_signal_5671) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_5_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (stateArray_nReset_selMC), .A1_f (new_AGEMA_signal_4210), .B0_t (stateArray_MUX_inS23ser_mux_inst_5_X), .B0_f (new_AGEMA_signal_5669), .B1_t (new_AGEMA_signal_5670), .B1_f (new_AGEMA_signal_5671), .Z0_t (stateArray_MUX_inS23ser_mux_inst_5_Y), .Z0_f (new_AGEMA_signal_5856), .Z1_t (new_AGEMA_signal_5857), .Z1_f (new_AGEMA_signal_5858) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_5_XOR2_U1 ( .A0_t (stateArray_MUX_inS23ser_mux_inst_5_Y), .A0_f (new_AGEMA_signal_5856), .A1_t (new_AGEMA_signal_5857), .A1_f (new_AGEMA_signal_5858), .B0_t (MixColumns_line3_S02[6]), .B0_f (new_AGEMA_signal_3157), .B1_t (new_AGEMA_signal_3158), .B1_f (new_AGEMA_signal_3159), .Z0_t (stateArray_inS23ser[5]), .Z0_f (new_AGEMA_signal_6268), .Z1_t (new_AGEMA_signal_6269), .Z1_f (new_AGEMA_signal_6270) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_6_XOR1_U1 ( .A0_t (MixColumns_line3_S02[7]), .A0_f (new_AGEMA_signal_3166), .A1_t (new_AGEMA_signal_3167), .A1_f (new_AGEMA_signal_3168), .B0_t (StateInMC[14]), .B0_f (new_AGEMA_signal_5506), .B1_t (new_AGEMA_signal_5507), .B1_f (new_AGEMA_signal_5508), .Z0_t (stateArray_MUX_inS23ser_mux_inst_6_X), .Z0_f (new_AGEMA_signal_5672), .Z1_t (new_AGEMA_signal_5673), .Z1_f (new_AGEMA_signal_5674) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_6_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (stateArray_nReset_selMC), .A1_f (new_AGEMA_signal_4210), .B0_t (stateArray_MUX_inS23ser_mux_inst_6_X), .B0_f (new_AGEMA_signal_5672), .B1_t (new_AGEMA_signal_5673), .B1_f (new_AGEMA_signal_5674), .Z0_t (stateArray_MUX_inS23ser_mux_inst_6_Y), .Z0_f (new_AGEMA_signal_5859), .Z1_t (new_AGEMA_signal_5860), .Z1_f (new_AGEMA_signal_5861) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_6_XOR2_U1 ( .A0_t (stateArray_MUX_inS23ser_mux_inst_6_Y), .A0_f (new_AGEMA_signal_5859), .A1_t (new_AGEMA_signal_5860), .A1_f (new_AGEMA_signal_5861), .B0_t (MixColumns_line3_S02[7]), .B0_f (new_AGEMA_signal_3166), .B1_t (new_AGEMA_signal_3167), .B1_f (new_AGEMA_signal_3168), .Z0_t (stateArray_inS23ser[6]), .Z0_f (new_AGEMA_signal_6271), .Z1_t (new_AGEMA_signal_6272), .Z1_f (new_AGEMA_signal_6273) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_7_XOR1_U1 ( .A0_t (MixColumns_line3_S02[0]), .A0_f (new_AGEMA_signal_3175), .A1_t (new_AGEMA_signal_3176), .A1_f (new_AGEMA_signal_3177), .B0_t (StateInMC[15]), .B0_f (new_AGEMA_signal_5509), .B1_t (new_AGEMA_signal_5510), .B1_f (new_AGEMA_signal_5511), .Z0_t (stateArray_MUX_inS23ser_mux_inst_7_X), .Z0_f (new_AGEMA_signal_5675), .Z1_t (new_AGEMA_signal_5676), .Z1_f (new_AGEMA_signal_5677) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_7_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (stateArray_nReset_selMC), .A1_f (new_AGEMA_signal_4210), .B0_t (stateArray_MUX_inS23ser_mux_inst_7_X), .B0_f (new_AGEMA_signal_5675), .B1_t (new_AGEMA_signal_5676), .B1_f (new_AGEMA_signal_5677), .Z0_t (stateArray_MUX_inS23ser_mux_inst_7_Y), .Z0_f (new_AGEMA_signal_5862), .Z1_t (new_AGEMA_signal_5863), .Z1_f (new_AGEMA_signal_5864) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS23ser_mux_inst_7_XOR2_U1 ( .A0_t (stateArray_MUX_inS23ser_mux_inst_7_Y), .A0_f (new_AGEMA_signal_5862), .A1_t (new_AGEMA_signal_5863), .A1_f (new_AGEMA_signal_5864), .B0_t (MixColumns_line3_S02[0]), .B0_f (new_AGEMA_signal_3175), .B1_t (new_AGEMA_signal_3176), .B1_f (new_AGEMA_signal_3177), .Z0_t (stateArray_inS23ser[7]), .Z0_f (new_AGEMA_signal_6274), .Z1_t (new_AGEMA_signal_6275), .Z1_f (new_AGEMA_signal_6276) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_0_XOR1_U1 ( .A0_t (StateIn[0]), .A0_f (new_AGEMA_signal_7580), .A1_t (new_AGEMA_signal_7581), .A1_f (new_AGEMA_signal_7582), .B0_t (StateInMC[0]), .B0_f (new_AGEMA_signal_5464), .B1_t (new_AGEMA_signal_5465), .B1_f (new_AGEMA_signal_5466), .Z0_t (stateArray_MUX_input_MC_mux_inst_0_X), .Z0_f (new_AGEMA_signal_7649), .Z1_t (new_AGEMA_signal_7650), .Z1_f (new_AGEMA_signal_7651) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_0_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (stateArray_MUX_input_MC_mux_inst_0_X), .B0_f (new_AGEMA_signal_7649), .B1_t (new_AGEMA_signal_7650), .B1_f (new_AGEMA_signal_7651), .Z0_t (stateArray_MUX_input_MC_mux_inst_0_Y), .Z0_f (new_AGEMA_signal_7676), .Z1_t (new_AGEMA_signal_7677), .Z1_f (new_AGEMA_signal_7678) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_0_XOR2_U1 ( .A0_t (stateArray_MUX_input_MC_mux_inst_0_Y), .A0_f (new_AGEMA_signal_7676), .A1_t (new_AGEMA_signal_7677), .A1_f (new_AGEMA_signal_7678), .B0_t (StateIn[0]), .B0_f (new_AGEMA_signal_7580), .B1_t (new_AGEMA_signal_7581), .B1_f (new_AGEMA_signal_7582), .Z0_t (stateArray_input_MC[0]), .Z0_f (new_AGEMA_signal_7724), .Z1_t (new_AGEMA_signal_7725), .Z1_f (new_AGEMA_signal_7726) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_1_XOR1_U1 ( .A0_t (StateIn[1]), .A0_f (new_AGEMA_signal_7628), .A1_t (new_AGEMA_signal_7629), .A1_f (new_AGEMA_signal_7630), .B0_t (StateInMC[1]), .B0_f (new_AGEMA_signal_5678), .B1_t (new_AGEMA_signal_5679), .B1_f (new_AGEMA_signal_5680), .Z0_t (stateArray_MUX_input_MC_mux_inst_1_X), .Z0_f (new_AGEMA_signal_7679), .Z1_t (new_AGEMA_signal_7680), .Z1_f (new_AGEMA_signal_7681) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (stateArray_MUX_input_MC_mux_inst_1_X), .B0_f (new_AGEMA_signal_7679), .B1_t (new_AGEMA_signal_7680), .B1_f (new_AGEMA_signal_7681), .Z0_t (stateArray_MUX_input_MC_mux_inst_1_Y), .Z0_f (new_AGEMA_signal_7727), .Z1_t (new_AGEMA_signal_7728), .Z1_f (new_AGEMA_signal_7729) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_1_XOR2_U1 ( .A0_t (stateArray_MUX_input_MC_mux_inst_1_Y), .A0_f (new_AGEMA_signal_7727), .A1_t (new_AGEMA_signal_7728), .A1_f (new_AGEMA_signal_7729), .B0_t (StateIn[1]), .B0_f (new_AGEMA_signal_7628), .B1_t (new_AGEMA_signal_7629), .B1_f (new_AGEMA_signal_7630), .Z0_t (stateArray_input_MC[1]), .Z0_f (new_AGEMA_signal_7772), .Z1_t (new_AGEMA_signal_7773), .Z1_f (new_AGEMA_signal_7774) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_2_XOR1_U1 ( .A0_t (StateIn[2]), .A0_f (new_AGEMA_signal_7631), .A1_t (new_AGEMA_signal_7632), .A1_f (new_AGEMA_signal_7633), .B0_t (StateInMC[2]), .B0_f (new_AGEMA_signal_5470), .B1_t (new_AGEMA_signal_5471), .B1_f (new_AGEMA_signal_5472), .Z0_t (stateArray_MUX_input_MC_mux_inst_2_X), .Z0_f (new_AGEMA_signal_7682), .Z1_t (new_AGEMA_signal_7683), .Z1_f (new_AGEMA_signal_7684) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_2_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (stateArray_MUX_input_MC_mux_inst_2_X), .B0_f (new_AGEMA_signal_7682), .B1_t (new_AGEMA_signal_7683), .B1_f (new_AGEMA_signal_7684), .Z0_t (stateArray_MUX_input_MC_mux_inst_2_Y), .Z0_f (new_AGEMA_signal_7730), .Z1_t (new_AGEMA_signal_7731), .Z1_f (new_AGEMA_signal_7732) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_2_XOR2_U1 ( .A0_t (stateArray_MUX_input_MC_mux_inst_2_Y), .A0_f (new_AGEMA_signal_7730), .A1_t (new_AGEMA_signal_7731), .A1_f (new_AGEMA_signal_7732), .B0_t (StateIn[2]), .B0_f (new_AGEMA_signal_7631), .B1_t (new_AGEMA_signal_7632), .B1_f (new_AGEMA_signal_7633), .Z0_t (stateArray_input_MC[2]), .Z0_f (new_AGEMA_signal_7775), .Z1_t (new_AGEMA_signal_7776), .Z1_f (new_AGEMA_signal_7777) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_3_XOR1_U1 ( .A0_t (StateIn[3]), .A0_f (new_AGEMA_signal_7634), .A1_t (new_AGEMA_signal_7635), .A1_f (new_AGEMA_signal_7636), .B0_t (StateInMC[3]), .B0_f (new_AGEMA_signal_5681), .B1_t (new_AGEMA_signal_5682), .B1_f (new_AGEMA_signal_5683), .Z0_t (stateArray_MUX_input_MC_mux_inst_3_X), .Z0_f (new_AGEMA_signal_7685), .Z1_t (new_AGEMA_signal_7686), .Z1_f (new_AGEMA_signal_7687) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_3_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (stateArray_MUX_input_MC_mux_inst_3_X), .B0_f (new_AGEMA_signal_7685), .B1_t (new_AGEMA_signal_7686), .B1_f (new_AGEMA_signal_7687), .Z0_t (stateArray_MUX_input_MC_mux_inst_3_Y), .Z0_f (new_AGEMA_signal_7733), .Z1_t (new_AGEMA_signal_7734), .Z1_f (new_AGEMA_signal_7735) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_3_XOR2_U1 ( .A0_t (stateArray_MUX_input_MC_mux_inst_3_Y), .A0_f (new_AGEMA_signal_7733), .A1_t (new_AGEMA_signal_7734), .A1_f (new_AGEMA_signal_7735), .B0_t (StateIn[3]), .B0_f (new_AGEMA_signal_7634), .B1_t (new_AGEMA_signal_7635), .B1_f (new_AGEMA_signal_7636), .Z0_t (stateArray_input_MC[3]), .Z0_f (new_AGEMA_signal_7778), .Z1_t (new_AGEMA_signal_7779), .Z1_f (new_AGEMA_signal_7780) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_4_XOR1_U1 ( .A0_t (StateIn[4]), .A0_f (new_AGEMA_signal_7637), .A1_t (new_AGEMA_signal_7638), .A1_f (new_AGEMA_signal_7639), .B0_t (StateInMC[4]), .B0_f (new_AGEMA_signal_5684), .B1_t (new_AGEMA_signal_5685), .B1_f (new_AGEMA_signal_5686), .Z0_t (stateArray_MUX_input_MC_mux_inst_4_X), .Z0_f (new_AGEMA_signal_7688), .Z1_t (new_AGEMA_signal_7689), .Z1_f (new_AGEMA_signal_7690) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_4_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (stateArray_MUX_input_MC_mux_inst_4_X), .B0_f (new_AGEMA_signal_7688), .B1_t (new_AGEMA_signal_7689), .B1_f (new_AGEMA_signal_7690), .Z0_t (stateArray_MUX_input_MC_mux_inst_4_Y), .Z0_f (new_AGEMA_signal_7736), .Z1_t (new_AGEMA_signal_7737), .Z1_f (new_AGEMA_signal_7738) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_4_XOR2_U1 ( .A0_t (stateArray_MUX_input_MC_mux_inst_4_Y), .A0_f (new_AGEMA_signal_7736), .A1_t (new_AGEMA_signal_7737), .A1_f (new_AGEMA_signal_7738), .B0_t (StateIn[4]), .B0_f (new_AGEMA_signal_7637), .B1_t (new_AGEMA_signal_7638), .B1_f (new_AGEMA_signal_7639), .Z0_t (stateArray_input_MC[4]), .Z0_f (new_AGEMA_signal_7781), .Z1_t (new_AGEMA_signal_7782), .Z1_f (new_AGEMA_signal_7783) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_5_XOR1_U1 ( .A0_t (StateIn[5]), .A0_f (new_AGEMA_signal_7640), .A1_t (new_AGEMA_signal_7641), .A1_f (new_AGEMA_signal_7642), .B0_t (StateInMC[5]), .B0_f (new_AGEMA_signal_5479), .B1_t (new_AGEMA_signal_5480), .B1_f (new_AGEMA_signal_5481), .Z0_t (stateArray_MUX_input_MC_mux_inst_5_X), .Z0_f (new_AGEMA_signal_7691), .Z1_t (new_AGEMA_signal_7692), .Z1_f (new_AGEMA_signal_7693) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_5_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (stateArray_MUX_input_MC_mux_inst_5_X), .B0_f (new_AGEMA_signal_7691), .B1_t (new_AGEMA_signal_7692), .B1_f (new_AGEMA_signal_7693), .Z0_t (stateArray_MUX_input_MC_mux_inst_5_Y), .Z0_f (new_AGEMA_signal_7739), .Z1_t (new_AGEMA_signal_7740), .Z1_f (new_AGEMA_signal_7741) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_5_XOR2_U1 ( .A0_t (stateArray_MUX_input_MC_mux_inst_5_Y), .A0_f (new_AGEMA_signal_7739), .A1_t (new_AGEMA_signal_7740), .A1_f (new_AGEMA_signal_7741), .B0_t (StateIn[5]), .B0_f (new_AGEMA_signal_7640), .B1_t (new_AGEMA_signal_7641), .B1_f (new_AGEMA_signal_7642), .Z0_t (stateArray_input_MC[5]), .Z0_f (new_AGEMA_signal_7784), .Z1_t (new_AGEMA_signal_7785), .Z1_f (new_AGEMA_signal_7786) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_6_XOR1_U1 ( .A0_t (StateIn[6]), .A0_f (new_AGEMA_signal_7643), .A1_t (new_AGEMA_signal_7644), .A1_f (new_AGEMA_signal_7645), .B0_t (StateInMC[6]), .B0_f (new_AGEMA_signal_5482), .B1_t (new_AGEMA_signal_5483), .B1_f (new_AGEMA_signal_5484), .Z0_t (stateArray_MUX_input_MC_mux_inst_6_X), .Z0_f (new_AGEMA_signal_7694), .Z1_t (new_AGEMA_signal_7695), .Z1_f (new_AGEMA_signal_7696) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_6_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (stateArray_MUX_input_MC_mux_inst_6_X), .B0_f (new_AGEMA_signal_7694), .B1_t (new_AGEMA_signal_7695), .B1_f (new_AGEMA_signal_7696), .Z0_t (stateArray_MUX_input_MC_mux_inst_6_Y), .Z0_f (new_AGEMA_signal_7742), .Z1_t (new_AGEMA_signal_7743), .Z1_f (new_AGEMA_signal_7744) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_6_XOR2_U1 ( .A0_t (stateArray_MUX_input_MC_mux_inst_6_Y), .A0_f (new_AGEMA_signal_7742), .A1_t (new_AGEMA_signal_7743), .A1_f (new_AGEMA_signal_7744), .B0_t (StateIn[6]), .B0_f (new_AGEMA_signal_7643), .B1_t (new_AGEMA_signal_7644), .B1_f (new_AGEMA_signal_7645), .Z0_t (stateArray_input_MC[6]), .Z0_f (new_AGEMA_signal_7787), .Z1_t (new_AGEMA_signal_7788), .Z1_f (new_AGEMA_signal_7789) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_7_XOR1_U1 ( .A0_t (StateIn[7]), .A0_f (new_AGEMA_signal_7646), .A1_t (new_AGEMA_signal_7647), .A1_f (new_AGEMA_signal_7648), .B0_t (StateInMC[7]), .B0_f (new_AGEMA_signal_5485), .B1_t (new_AGEMA_signal_5486), .B1_f (new_AGEMA_signal_5487), .Z0_t (stateArray_MUX_input_MC_mux_inst_7_X), .Z0_f (new_AGEMA_signal_7697), .Z1_t (new_AGEMA_signal_7698), .Z1_f (new_AGEMA_signal_7699) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_7_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (stateArray_MUX_input_MC_mux_inst_7_X), .B0_f (new_AGEMA_signal_7697), .B1_t (new_AGEMA_signal_7698), .B1_f (new_AGEMA_signal_7699), .Z0_t (stateArray_MUX_input_MC_mux_inst_7_Y), .Z0_f (new_AGEMA_signal_7745), .Z1_t (new_AGEMA_signal_7746), .Z1_f (new_AGEMA_signal_7747) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_input_MC_mux_inst_7_XOR2_U1 ( .A0_t (stateArray_MUX_input_MC_mux_inst_7_Y), .A0_f (new_AGEMA_signal_7745), .A1_t (new_AGEMA_signal_7746), .A1_f (new_AGEMA_signal_7747), .B0_t (StateIn[7]), .B0_f (new_AGEMA_signal_7646), .B1_t (new_AGEMA_signal_7647), .B1_f (new_AGEMA_signal_7648), .Z0_t (stateArray_input_MC[7]), .Z0_f (new_AGEMA_signal_7790), .Z1_t (new_AGEMA_signal_7791), .Z1_f (new_AGEMA_signal_7792) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_0_XOR1_U1 ( .A0_t (port_in_s0_t[0]), .A0_f (port_in_s0_f[0]), .A1_t (port_in_s1_t[0]), .A1_f (port_in_s1_f[0]), .B0_t (stateArray_input_MC[0]), .B0_f (new_AGEMA_signal_7724), .B1_t (new_AGEMA_signal_7725), .B1_f (new_AGEMA_signal_7726), .Z0_t (stateArray_MUX_inS33ser_mux_inst_0_X), .Z0_f (new_AGEMA_signal_7796), .Z1_t (new_AGEMA_signal_7797), .Z1_f (new_AGEMA_signal_7798) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_0_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (stateArray_MUX_inS33ser_mux_inst_0_X), .B0_f (new_AGEMA_signal_7796), .B1_t (new_AGEMA_signal_7797), .B1_f (new_AGEMA_signal_7798), .Z0_t (stateArray_MUX_inS33ser_mux_inst_0_Y), .Z0_f (new_AGEMA_signal_7820), .Z1_t (new_AGEMA_signal_7821), .Z1_f (new_AGEMA_signal_7822) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_0_XOR2_U1 ( .A0_t (stateArray_MUX_inS33ser_mux_inst_0_Y), .A0_f (new_AGEMA_signal_7820), .A1_t (new_AGEMA_signal_7821), .A1_f (new_AGEMA_signal_7822), .B0_t (port_in_s0_t[0]), .B0_f (port_in_s0_f[0]), .B1_t (port_in_s1_t[0]), .B1_f (port_in_s1_f[0]), .Z0_t (stateArray_inS33ser[0]), .Z0_f (new_AGEMA_signal_7865), .Z1_t (new_AGEMA_signal_7866), .Z1_f (new_AGEMA_signal_7867) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_1_XOR1_U1 ( .A0_t (port_in_s0_t[1]), .A0_f (port_in_s0_f[1]), .A1_t (port_in_s1_t[1]), .A1_f (port_in_s1_f[1]), .B0_t (stateArray_input_MC[1]), .B0_f (new_AGEMA_signal_7772), .B1_t (new_AGEMA_signal_7773), .B1_f (new_AGEMA_signal_7774), .Z0_t (stateArray_MUX_inS33ser_mux_inst_1_X), .Z0_f (new_AGEMA_signal_7826), .Z1_t (new_AGEMA_signal_7827), .Z1_f (new_AGEMA_signal_7828) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (stateArray_MUX_inS33ser_mux_inst_1_X), .B0_f (new_AGEMA_signal_7826), .B1_t (new_AGEMA_signal_7827), .B1_f (new_AGEMA_signal_7828), .Z0_t (stateArray_MUX_inS33ser_mux_inst_1_Y), .Z0_f (new_AGEMA_signal_7868), .Z1_t (new_AGEMA_signal_7869), .Z1_f (new_AGEMA_signal_7870) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_1_XOR2_U1 ( .A0_t (stateArray_MUX_inS33ser_mux_inst_1_Y), .A0_f (new_AGEMA_signal_7868), .A1_t (new_AGEMA_signal_7869), .A1_f (new_AGEMA_signal_7870), .B0_t (port_in_s0_t[1]), .B0_f (port_in_s0_f[1]), .B1_t (port_in_s1_t[1]), .B1_f (port_in_s1_f[1]), .Z0_t (stateArray_inS33ser[1]), .Z0_f (new_AGEMA_signal_7892), .Z1_t (new_AGEMA_signal_7893), .Z1_f (new_AGEMA_signal_7894) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_2_XOR1_U1 ( .A0_t (port_in_s0_t[2]), .A0_f (port_in_s0_f[2]), .A1_t (port_in_s1_t[2]), .A1_f (port_in_s1_f[2]), .B0_t (stateArray_input_MC[2]), .B0_f (new_AGEMA_signal_7775), .B1_t (new_AGEMA_signal_7776), .B1_f (new_AGEMA_signal_7777), .Z0_t (stateArray_MUX_inS33ser_mux_inst_2_X), .Z0_f (new_AGEMA_signal_7832), .Z1_t (new_AGEMA_signal_7833), .Z1_f (new_AGEMA_signal_7834) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_2_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (stateArray_MUX_inS33ser_mux_inst_2_X), .B0_f (new_AGEMA_signal_7832), .B1_t (new_AGEMA_signal_7833), .B1_f (new_AGEMA_signal_7834), .Z0_t (stateArray_MUX_inS33ser_mux_inst_2_Y), .Z0_f (new_AGEMA_signal_7871), .Z1_t (new_AGEMA_signal_7872), .Z1_f (new_AGEMA_signal_7873) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_2_XOR2_U1 ( .A0_t (stateArray_MUX_inS33ser_mux_inst_2_Y), .A0_f (new_AGEMA_signal_7871), .A1_t (new_AGEMA_signal_7872), .A1_f (new_AGEMA_signal_7873), .B0_t (port_in_s0_t[2]), .B0_f (port_in_s0_f[2]), .B1_t (port_in_s1_t[2]), .B1_f (port_in_s1_f[2]), .Z0_t (stateArray_inS33ser[2]), .Z0_f (new_AGEMA_signal_7895), .Z1_t (new_AGEMA_signal_7896), .Z1_f (new_AGEMA_signal_7897) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_3_XOR1_U1 ( .A0_t (port_in_s0_t[3]), .A0_f (port_in_s0_f[3]), .A1_t (port_in_s1_t[3]), .A1_f (port_in_s1_f[3]), .B0_t (stateArray_input_MC[3]), .B0_f (new_AGEMA_signal_7778), .B1_t (new_AGEMA_signal_7779), .B1_f (new_AGEMA_signal_7780), .Z0_t (stateArray_MUX_inS33ser_mux_inst_3_X), .Z0_f (new_AGEMA_signal_7838), .Z1_t (new_AGEMA_signal_7839), .Z1_f (new_AGEMA_signal_7840) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_3_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (stateArray_MUX_inS33ser_mux_inst_3_X), .B0_f (new_AGEMA_signal_7838), .B1_t (new_AGEMA_signal_7839), .B1_f (new_AGEMA_signal_7840), .Z0_t (stateArray_MUX_inS33ser_mux_inst_3_Y), .Z0_f (new_AGEMA_signal_7874), .Z1_t (new_AGEMA_signal_7875), .Z1_f (new_AGEMA_signal_7876) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_3_XOR2_U1 ( .A0_t (stateArray_MUX_inS33ser_mux_inst_3_Y), .A0_f (new_AGEMA_signal_7874), .A1_t (new_AGEMA_signal_7875), .A1_f (new_AGEMA_signal_7876), .B0_t (port_in_s0_t[3]), .B0_f (port_in_s0_f[3]), .B1_t (port_in_s1_t[3]), .B1_f (port_in_s1_f[3]), .Z0_t (stateArray_inS33ser[3]), .Z0_f (new_AGEMA_signal_7898), .Z1_t (new_AGEMA_signal_7899), .Z1_f (new_AGEMA_signal_7900) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_4_XOR1_U1 ( .A0_t (port_in_s0_t[4]), .A0_f (port_in_s0_f[4]), .A1_t (port_in_s1_t[4]), .A1_f (port_in_s1_f[4]), .B0_t (stateArray_input_MC[4]), .B0_f (new_AGEMA_signal_7781), .B1_t (new_AGEMA_signal_7782), .B1_f (new_AGEMA_signal_7783), .Z0_t (stateArray_MUX_inS33ser_mux_inst_4_X), .Z0_f (new_AGEMA_signal_7844), .Z1_t (new_AGEMA_signal_7845), .Z1_f (new_AGEMA_signal_7846) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_4_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (stateArray_MUX_inS33ser_mux_inst_4_X), .B0_f (new_AGEMA_signal_7844), .B1_t (new_AGEMA_signal_7845), .B1_f (new_AGEMA_signal_7846), .Z0_t (stateArray_MUX_inS33ser_mux_inst_4_Y), .Z0_f (new_AGEMA_signal_7877), .Z1_t (new_AGEMA_signal_7878), .Z1_f (new_AGEMA_signal_7879) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_4_XOR2_U1 ( .A0_t (stateArray_MUX_inS33ser_mux_inst_4_Y), .A0_f (new_AGEMA_signal_7877), .A1_t (new_AGEMA_signal_7878), .A1_f (new_AGEMA_signal_7879), .B0_t (port_in_s0_t[4]), .B0_f (port_in_s0_f[4]), .B1_t (port_in_s1_t[4]), .B1_f (port_in_s1_f[4]), .Z0_t (stateArray_inS33ser[4]), .Z0_f (new_AGEMA_signal_7901), .Z1_t (new_AGEMA_signal_7902), .Z1_f (new_AGEMA_signal_7903) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_5_XOR1_U1 ( .A0_t (port_in_s0_t[5]), .A0_f (port_in_s0_f[5]), .A1_t (port_in_s1_t[5]), .A1_f (port_in_s1_f[5]), .B0_t (stateArray_input_MC[5]), .B0_f (new_AGEMA_signal_7784), .B1_t (new_AGEMA_signal_7785), .B1_f (new_AGEMA_signal_7786), .Z0_t (stateArray_MUX_inS33ser_mux_inst_5_X), .Z0_f (new_AGEMA_signal_7850), .Z1_t (new_AGEMA_signal_7851), .Z1_f (new_AGEMA_signal_7852) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_5_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (stateArray_MUX_inS33ser_mux_inst_5_X), .B0_f (new_AGEMA_signal_7850), .B1_t (new_AGEMA_signal_7851), .B1_f (new_AGEMA_signal_7852), .Z0_t (stateArray_MUX_inS33ser_mux_inst_5_Y), .Z0_f (new_AGEMA_signal_7880), .Z1_t (new_AGEMA_signal_7881), .Z1_f (new_AGEMA_signal_7882) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_5_XOR2_U1 ( .A0_t (stateArray_MUX_inS33ser_mux_inst_5_Y), .A0_f (new_AGEMA_signal_7880), .A1_t (new_AGEMA_signal_7881), .A1_f (new_AGEMA_signal_7882), .B0_t (port_in_s0_t[5]), .B0_f (port_in_s0_f[5]), .B1_t (port_in_s1_t[5]), .B1_f (port_in_s1_f[5]), .Z0_t (stateArray_inS33ser[5]), .Z0_f (new_AGEMA_signal_7904), .Z1_t (new_AGEMA_signal_7905), .Z1_f (new_AGEMA_signal_7906) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_6_XOR1_U1 ( .A0_t (port_in_s0_t[6]), .A0_f (port_in_s0_f[6]), .A1_t (port_in_s1_t[6]), .A1_f (port_in_s1_f[6]), .B0_t (stateArray_input_MC[6]), .B0_f (new_AGEMA_signal_7787), .B1_t (new_AGEMA_signal_7788), .B1_f (new_AGEMA_signal_7789), .Z0_t (stateArray_MUX_inS33ser_mux_inst_6_X), .Z0_f (new_AGEMA_signal_7856), .Z1_t (new_AGEMA_signal_7857), .Z1_f (new_AGEMA_signal_7858) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_6_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (stateArray_MUX_inS33ser_mux_inst_6_X), .B0_f (new_AGEMA_signal_7856), .B1_t (new_AGEMA_signal_7857), .B1_f (new_AGEMA_signal_7858), .Z0_t (stateArray_MUX_inS33ser_mux_inst_6_Y), .Z0_f (new_AGEMA_signal_7883), .Z1_t (new_AGEMA_signal_7884), .Z1_f (new_AGEMA_signal_7885) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_6_XOR2_U1 ( .A0_t (stateArray_MUX_inS33ser_mux_inst_6_Y), .A0_f (new_AGEMA_signal_7883), .A1_t (new_AGEMA_signal_7884), .A1_f (new_AGEMA_signal_7885), .B0_t (port_in_s0_t[6]), .B0_f (port_in_s0_f[6]), .B1_t (port_in_s1_t[6]), .B1_f (port_in_s1_f[6]), .Z0_t (stateArray_inS33ser[6]), .Z0_f (new_AGEMA_signal_7907), .Z1_t (new_AGEMA_signal_7908), .Z1_f (new_AGEMA_signal_7909) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_7_XOR1_U1 ( .A0_t (port_in_s0_t[7]), .A0_f (port_in_s0_f[7]), .A1_t (port_in_s1_t[7]), .A1_f (port_in_s1_f[7]), .B0_t (stateArray_input_MC[7]), .B0_f (new_AGEMA_signal_7790), .B1_t (new_AGEMA_signal_7791), .B1_f (new_AGEMA_signal_7792), .Z0_t (stateArray_MUX_inS33ser_mux_inst_7_X), .Z0_f (new_AGEMA_signal_7862), .Z1_t (new_AGEMA_signal_7863), .Z1_f (new_AGEMA_signal_7864) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_7_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (stateArray_MUX_inS33ser_mux_inst_7_X), .B0_f (new_AGEMA_signal_7862), .B1_t (new_AGEMA_signal_7863), .B1_f (new_AGEMA_signal_7864), .Z0_t (stateArray_MUX_inS33ser_mux_inst_7_Y), .Z0_f (new_AGEMA_signal_7886), .Z1_t (new_AGEMA_signal_7887), .Z1_f (new_AGEMA_signal_7888) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateArray_MUX_inS33ser_mux_inst_7_XOR2_U1 ( .A0_t (stateArray_MUX_inS33ser_mux_inst_7_Y), .A0_f (new_AGEMA_signal_7886), .A1_t (new_AGEMA_signal_7887), .A1_f (new_AGEMA_signal_7888), .B0_t (port_in_s0_t[7]), .B0_f (port_in_s0_f[7]), .B1_t (port_in_s1_t[7]), .B1_f (port_in_s1_f[7]), .Z0_t (stateArray_inS33ser[7]), .Z0_f (new_AGEMA_signal_7910), .Z1_t (new_AGEMA_signal_7911), .Z1_f (new_AGEMA_signal_7912) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_0_XOR1_U1 ( .A0_t (MCout[0]), .A0_f (new_AGEMA_signal_5130), .A1_t (new_AGEMA_signal_5131), .A1_f (new_AGEMA_signal_5132), .B0_t (MCin[0]), .B0_f (new_AGEMA_signal_3112), .B1_t (new_AGEMA_signal_3113), .B1_f (new_AGEMA_signal_3114), .Z0_t (MUX_StateInMC_mux_inst_0_X), .Z0_f (new_AGEMA_signal_5163), .Z1_t (new_AGEMA_signal_5164), .Z1_f (new_AGEMA_signal_5165) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_0_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_4669), .B0_t (MUX_StateInMC_mux_inst_0_X), .B0_f (new_AGEMA_signal_5163), .B1_t (new_AGEMA_signal_5164), .B1_f (new_AGEMA_signal_5165), .Z0_t (MUX_StateInMC_mux_inst_0_Y), .Z0_f (new_AGEMA_signal_5310), .Z1_t (new_AGEMA_signal_5311), .Z1_f (new_AGEMA_signal_5312) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_0_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_0_Y), .A0_f (new_AGEMA_signal_5310), .A1_t (new_AGEMA_signal_5311), .A1_f (new_AGEMA_signal_5312), .B0_t (MCout[0]), .B0_f (new_AGEMA_signal_5130), .B1_t (new_AGEMA_signal_5131), .B1_f (new_AGEMA_signal_5132), .Z0_t (StateInMC[0]), .Z0_f (new_AGEMA_signal_5464), .Z1_t (new_AGEMA_signal_5465), .Z1_f (new_AGEMA_signal_5466) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_1_XOR1_U1 ( .A0_t (MCout[1]), .A0_f (new_AGEMA_signal_5280), .A1_t (new_AGEMA_signal_5281), .A1_f (new_AGEMA_signal_5282), .B0_t (MixColumns_line3_S02[2]), .B0_f (new_AGEMA_signal_3121), .B1_t (new_AGEMA_signal_3122), .B1_f (new_AGEMA_signal_3123), .Z0_t (MUX_StateInMC_mux_inst_1_X), .Z0_f (new_AGEMA_signal_5313), .Z1_t (new_AGEMA_signal_5314), .Z1_f (new_AGEMA_signal_5315) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_4669), .B0_t (MUX_StateInMC_mux_inst_1_X), .B0_f (new_AGEMA_signal_5313), .B1_t (new_AGEMA_signal_5314), .B1_f (new_AGEMA_signal_5315), .Z0_t (MUX_StateInMC_mux_inst_1_Y), .Z0_f (new_AGEMA_signal_5467), .Z1_t (new_AGEMA_signal_5468), .Z1_f (new_AGEMA_signal_5469) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_1_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_1_Y), .A0_f (new_AGEMA_signal_5467), .A1_t (new_AGEMA_signal_5468), .A1_f (new_AGEMA_signal_5469), .B0_t (MCout[1]), .B0_f (new_AGEMA_signal_5280), .B1_t (new_AGEMA_signal_5281), .B1_f (new_AGEMA_signal_5282), .Z0_t (StateInMC[1]), .Z0_f (new_AGEMA_signal_5678), .Z1_t (new_AGEMA_signal_5679), .Z1_f (new_AGEMA_signal_5680) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_2_XOR1_U1 ( .A0_t (MCout[2]), .A0_f (new_AGEMA_signal_5124), .A1_t (new_AGEMA_signal_5125), .A1_f (new_AGEMA_signal_5126), .B0_t (MCin[2]), .B0_f (new_AGEMA_signal_3130), .B1_t (new_AGEMA_signal_3131), .B1_f (new_AGEMA_signal_3132), .Z0_t (MUX_StateInMC_mux_inst_2_X), .Z0_f (new_AGEMA_signal_5166), .Z1_t (new_AGEMA_signal_5167), .Z1_f (new_AGEMA_signal_5168) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_2_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_4669), .B0_t (MUX_StateInMC_mux_inst_2_X), .B0_f (new_AGEMA_signal_5166), .B1_t (new_AGEMA_signal_5167), .B1_f (new_AGEMA_signal_5168), .Z0_t (MUX_StateInMC_mux_inst_2_Y), .Z0_f (new_AGEMA_signal_5316), .Z1_t (new_AGEMA_signal_5317), .Z1_f (new_AGEMA_signal_5318) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_2_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_2_Y), .A0_f (new_AGEMA_signal_5316), .A1_t (new_AGEMA_signal_5317), .A1_f (new_AGEMA_signal_5318), .B0_t (MCout[2]), .B0_f (new_AGEMA_signal_5124), .B1_t (new_AGEMA_signal_5125), .B1_f (new_AGEMA_signal_5126), .Z0_t (StateInMC[2]), .Z0_f (new_AGEMA_signal_5470), .Z1_t (new_AGEMA_signal_5471), .Z1_f (new_AGEMA_signal_5472) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_3_XOR1_U1 ( .A0_t (MCout[3]), .A0_f (new_AGEMA_signal_5277), .A1_t (new_AGEMA_signal_5278), .A1_f (new_AGEMA_signal_5279), .B0_t (MCin[3]), .B0_f (new_AGEMA_signal_3139), .B1_t (new_AGEMA_signal_3140), .B1_f (new_AGEMA_signal_3141), .Z0_t (MUX_StateInMC_mux_inst_3_X), .Z0_f (new_AGEMA_signal_5319), .Z1_t (new_AGEMA_signal_5320), .Z1_f (new_AGEMA_signal_5321) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_3_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_4669), .B0_t (MUX_StateInMC_mux_inst_3_X), .B0_f (new_AGEMA_signal_5319), .B1_t (new_AGEMA_signal_5320), .B1_f (new_AGEMA_signal_5321), .Z0_t (MUX_StateInMC_mux_inst_3_Y), .Z0_f (new_AGEMA_signal_5473), .Z1_t (new_AGEMA_signal_5474), .Z1_f (new_AGEMA_signal_5475) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_3_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_3_Y), .A0_f (new_AGEMA_signal_5473), .A1_t (new_AGEMA_signal_5474), .A1_f (new_AGEMA_signal_5475), .B0_t (MCout[3]), .B0_f (new_AGEMA_signal_5277), .B1_t (new_AGEMA_signal_5278), .B1_f (new_AGEMA_signal_5279), .Z0_t (StateInMC[3]), .Z0_f (new_AGEMA_signal_5681), .Z1_t (new_AGEMA_signal_5682), .Z1_f (new_AGEMA_signal_5683) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_4_XOR1_U1 ( .A0_t (MCout[4]), .A0_f (new_AGEMA_signal_5274), .A1_t (new_AGEMA_signal_5275), .A1_f (new_AGEMA_signal_5276), .B0_t (MixColumns_line3_S02[5]), .B0_f (new_AGEMA_signal_3148), .B1_t (new_AGEMA_signal_3149), .B1_f (new_AGEMA_signal_3150), .Z0_t (MUX_StateInMC_mux_inst_4_X), .Z0_f (new_AGEMA_signal_5322), .Z1_t (new_AGEMA_signal_5323), .Z1_f (new_AGEMA_signal_5324) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_4_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_4669), .B0_t (MUX_StateInMC_mux_inst_4_X), .B0_f (new_AGEMA_signal_5322), .B1_t (new_AGEMA_signal_5323), .B1_f (new_AGEMA_signal_5324), .Z0_t (MUX_StateInMC_mux_inst_4_Y), .Z0_f (new_AGEMA_signal_5476), .Z1_t (new_AGEMA_signal_5477), .Z1_f (new_AGEMA_signal_5478) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_4_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_4_Y), .A0_f (new_AGEMA_signal_5476), .A1_t (new_AGEMA_signal_5477), .A1_f (new_AGEMA_signal_5478), .B0_t (MCout[4]), .B0_f (new_AGEMA_signal_5274), .B1_t (new_AGEMA_signal_5275), .B1_f (new_AGEMA_signal_5276), .Z0_t (StateInMC[4]), .Z0_f (new_AGEMA_signal_5684), .Z1_t (new_AGEMA_signal_5685), .Z1_f (new_AGEMA_signal_5686) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_5_XOR1_U1 ( .A0_t (MCout[5]), .A0_f (new_AGEMA_signal_5115), .A1_t (new_AGEMA_signal_5116), .A1_f (new_AGEMA_signal_5117), .B0_t (MixColumns_line3_S02[6]), .B0_f (new_AGEMA_signal_3157), .B1_t (new_AGEMA_signal_3158), .B1_f (new_AGEMA_signal_3159), .Z0_t (MUX_StateInMC_mux_inst_5_X), .Z0_f (new_AGEMA_signal_5169), .Z1_t (new_AGEMA_signal_5170), .Z1_f (new_AGEMA_signal_5171) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_5_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_4669), .B0_t (MUX_StateInMC_mux_inst_5_X), .B0_f (new_AGEMA_signal_5169), .B1_t (new_AGEMA_signal_5170), .B1_f (new_AGEMA_signal_5171), .Z0_t (MUX_StateInMC_mux_inst_5_Y), .Z0_f (new_AGEMA_signal_5325), .Z1_t (new_AGEMA_signal_5326), .Z1_f (new_AGEMA_signal_5327) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_5_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_5_Y), .A0_f (new_AGEMA_signal_5325), .A1_t (new_AGEMA_signal_5326), .A1_f (new_AGEMA_signal_5327), .B0_t (MCout[5]), .B0_f (new_AGEMA_signal_5115), .B1_t (new_AGEMA_signal_5116), .B1_f (new_AGEMA_signal_5117), .Z0_t (StateInMC[5]), .Z0_f (new_AGEMA_signal_5479), .Z1_t (new_AGEMA_signal_5480), .Z1_f (new_AGEMA_signal_5481) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_6_XOR1_U1 ( .A0_t (MCout[6]), .A0_f (new_AGEMA_signal_5112), .A1_t (new_AGEMA_signal_5113), .A1_f (new_AGEMA_signal_5114), .B0_t (MixColumns_line3_S02[7]), .B0_f (new_AGEMA_signal_3166), .B1_t (new_AGEMA_signal_3167), .B1_f (new_AGEMA_signal_3168), .Z0_t (MUX_StateInMC_mux_inst_6_X), .Z0_f (new_AGEMA_signal_5172), .Z1_t (new_AGEMA_signal_5173), .Z1_f (new_AGEMA_signal_5174) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_6_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_4669), .B0_t (MUX_StateInMC_mux_inst_6_X), .B0_f (new_AGEMA_signal_5172), .B1_t (new_AGEMA_signal_5173), .B1_f (new_AGEMA_signal_5174), .Z0_t (MUX_StateInMC_mux_inst_6_Y), .Z0_f (new_AGEMA_signal_5328), .Z1_t (new_AGEMA_signal_5329), .Z1_f (new_AGEMA_signal_5330) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_6_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_6_Y), .A0_f (new_AGEMA_signal_5328), .A1_t (new_AGEMA_signal_5329), .A1_f (new_AGEMA_signal_5330), .B0_t (MCout[6]), .B0_f (new_AGEMA_signal_5112), .B1_t (new_AGEMA_signal_5113), .B1_f (new_AGEMA_signal_5114), .Z0_t (StateInMC[6]), .Z0_f (new_AGEMA_signal_5482), .Z1_t (new_AGEMA_signal_5483), .Z1_f (new_AGEMA_signal_5484) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_7_XOR1_U1 ( .A0_t (MCout[7]), .A0_f (new_AGEMA_signal_5109), .A1_t (new_AGEMA_signal_5110), .A1_f (new_AGEMA_signal_5111), .B0_t (MixColumns_line3_S02[0]), .B0_f (new_AGEMA_signal_3175), .B1_t (new_AGEMA_signal_3176), .B1_f (new_AGEMA_signal_3177), .Z0_t (MUX_StateInMC_mux_inst_7_X), .Z0_f (new_AGEMA_signal_5175), .Z1_t (new_AGEMA_signal_5176), .Z1_f (new_AGEMA_signal_5177) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_7_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_4669), .B0_t (MUX_StateInMC_mux_inst_7_X), .B0_f (new_AGEMA_signal_5175), .B1_t (new_AGEMA_signal_5176), .B1_f (new_AGEMA_signal_5177), .Z0_t (MUX_StateInMC_mux_inst_7_Y), .Z0_f (new_AGEMA_signal_5331), .Z1_t (new_AGEMA_signal_5332), .Z1_f (new_AGEMA_signal_5333) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_7_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_7_Y), .A0_f (new_AGEMA_signal_5331), .A1_t (new_AGEMA_signal_5332), .A1_f (new_AGEMA_signal_5333), .B0_t (MCout[7]), .B0_f (new_AGEMA_signal_5109), .B1_t (new_AGEMA_signal_5110), .B1_f (new_AGEMA_signal_5111), .Z0_t (StateInMC[7]), .Z0_f (new_AGEMA_signal_5485), .Z1_t (new_AGEMA_signal_5486), .Z1_f (new_AGEMA_signal_5487) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_8_XOR1_U1 ( .A0_t (MCout[8]), .A0_f (new_AGEMA_signal_5106), .A1_t (new_AGEMA_signal_5107), .A1_f (new_AGEMA_signal_5108), .B0_t (MCin[8]), .B0_f (new_AGEMA_signal_2989), .B1_t (new_AGEMA_signal_2990), .B1_f (new_AGEMA_signal_2991), .Z0_t (MUX_StateInMC_mux_inst_8_X), .Z0_f (new_AGEMA_signal_5178), .Z1_t (new_AGEMA_signal_5179), .Z1_f (new_AGEMA_signal_5180) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_8_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_4669), .B0_t (MUX_StateInMC_mux_inst_8_X), .B0_f (new_AGEMA_signal_5178), .B1_t (new_AGEMA_signal_5179), .B1_f (new_AGEMA_signal_5180), .Z0_t (MUX_StateInMC_mux_inst_8_Y), .Z0_f (new_AGEMA_signal_5334), .Z1_t (new_AGEMA_signal_5335), .Z1_f (new_AGEMA_signal_5336) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_8_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_8_Y), .A0_f (new_AGEMA_signal_5334), .A1_t (new_AGEMA_signal_5335), .A1_f (new_AGEMA_signal_5336), .B0_t (MCout[8]), .B0_f (new_AGEMA_signal_5106), .B1_t (new_AGEMA_signal_5107), .B1_f (new_AGEMA_signal_5108), .Z0_t (StateInMC[8]), .Z0_f (new_AGEMA_signal_5488), .Z1_t (new_AGEMA_signal_5489), .Z1_f (new_AGEMA_signal_5490) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_9_XOR1_U1 ( .A0_t (MCout[9]), .A0_f (new_AGEMA_signal_5271), .A1_t (new_AGEMA_signal_5272), .A1_f (new_AGEMA_signal_5273), .B0_t (MixColumns_line2_S02[2]), .B0_f (new_AGEMA_signal_2995), .B1_t (new_AGEMA_signal_2996), .B1_f (new_AGEMA_signal_2997), .Z0_t (MUX_StateInMC_mux_inst_9_X), .Z0_f (new_AGEMA_signal_5337), .Z1_t (new_AGEMA_signal_5338), .Z1_f (new_AGEMA_signal_5339) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_9_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_4669), .B0_t (MUX_StateInMC_mux_inst_9_X), .B0_f (new_AGEMA_signal_5337), .B1_t (new_AGEMA_signal_5338), .B1_f (new_AGEMA_signal_5339), .Z0_t (MUX_StateInMC_mux_inst_9_Y), .Z0_f (new_AGEMA_signal_5491), .Z1_t (new_AGEMA_signal_5492), .Z1_f (new_AGEMA_signal_5493) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_9_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_9_Y), .A0_f (new_AGEMA_signal_5491), .A1_t (new_AGEMA_signal_5492), .A1_f (new_AGEMA_signal_5493), .B0_t (MCout[9]), .B0_f (new_AGEMA_signal_5271), .B1_t (new_AGEMA_signal_5272), .B1_f (new_AGEMA_signal_5273), .Z0_t (StateInMC[9]), .Z0_f (new_AGEMA_signal_5687), .Z1_t (new_AGEMA_signal_5688), .Z1_f (new_AGEMA_signal_5689) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_10_XOR1_U1 ( .A0_t (MCout[10]), .A0_f (new_AGEMA_signal_5100), .A1_t (new_AGEMA_signal_5101), .A1_f (new_AGEMA_signal_5102), .B0_t (MCin[10]), .B0_f (new_AGEMA_signal_3001), .B1_t (new_AGEMA_signal_3002), .B1_f (new_AGEMA_signal_3003), .Z0_t (MUX_StateInMC_mux_inst_10_X), .Z0_f (new_AGEMA_signal_5181), .Z1_t (new_AGEMA_signal_5182), .Z1_f (new_AGEMA_signal_5183) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_10_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_4669), .B0_t (MUX_StateInMC_mux_inst_10_X), .B0_f (new_AGEMA_signal_5181), .B1_t (new_AGEMA_signal_5182), .B1_f (new_AGEMA_signal_5183), .Z0_t (MUX_StateInMC_mux_inst_10_Y), .Z0_f (new_AGEMA_signal_5340), .Z1_t (new_AGEMA_signal_5341), .Z1_f (new_AGEMA_signal_5342) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_10_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_10_Y), .A0_f (new_AGEMA_signal_5340), .A1_t (new_AGEMA_signal_5341), .A1_f (new_AGEMA_signal_5342), .B0_t (MCout[10]), .B0_f (new_AGEMA_signal_5100), .B1_t (new_AGEMA_signal_5101), .B1_f (new_AGEMA_signal_5102), .Z0_t (StateInMC[10]), .Z0_f (new_AGEMA_signal_5494), .Z1_t (new_AGEMA_signal_5495), .Z1_f (new_AGEMA_signal_5496) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_11_XOR1_U1 ( .A0_t (MCout[11]), .A0_f (new_AGEMA_signal_5268), .A1_t (new_AGEMA_signal_5269), .A1_f (new_AGEMA_signal_5270), .B0_t (MCin[11]), .B0_f (new_AGEMA_signal_3007), .B1_t (new_AGEMA_signal_3008), .B1_f (new_AGEMA_signal_3009), .Z0_t (MUX_StateInMC_mux_inst_11_X), .Z0_f (new_AGEMA_signal_5343), .Z1_t (new_AGEMA_signal_5344), .Z1_f (new_AGEMA_signal_5345) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_11_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_4669), .B0_t (MUX_StateInMC_mux_inst_11_X), .B0_f (new_AGEMA_signal_5343), .B1_t (new_AGEMA_signal_5344), .B1_f (new_AGEMA_signal_5345), .Z0_t (MUX_StateInMC_mux_inst_11_Y), .Z0_f (new_AGEMA_signal_5497), .Z1_t (new_AGEMA_signal_5498), .Z1_f (new_AGEMA_signal_5499) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_11_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_11_Y), .A0_f (new_AGEMA_signal_5497), .A1_t (new_AGEMA_signal_5498), .A1_f (new_AGEMA_signal_5499), .B0_t (MCout[11]), .B0_f (new_AGEMA_signal_5268), .B1_t (new_AGEMA_signal_5269), .B1_f (new_AGEMA_signal_5270), .Z0_t (StateInMC[11]), .Z0_f (new_AGEMA_signal_5690), .Z1_t (new_AGEMA_signal_5691), .Z1_f (new_AGEMA_signal_5692) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_12_XOR1_U1 ( .A0_t (MCout[12]), .A0_f (new_AGEMA_signal_5265), .A1_t (new_AGEMA_signal_5266), .A1_f (new_AGEMA_signal_5267), .B0_t (MixColumns_line2_S02[5]), .B0_f (new_AGEMA_signal_3013), .B1_t (new_AGEMA_signal_3014), .B1_f (new_AGEMA_signal_3015), .Z0_t (MUX_StateInMC_mux_inst_12_X), .Z0_f (new_AGEMA_signal_5346), .Z1_t (new_AGEMA_signal_5347), .Z1_f (new_AGEMA_signal_5348) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_12_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_4669), .B0_t (MUX_StateInMC_mux_inst_12_X), .B0_f (new_AGEMA_signal_5346), .B1_t (new_AGEMA_signal_5347), .B1_f (new_AGEMA_signal_5348), .Z0_t (MUX_StateInMC_mux_inst_12_Y), .Z0_f (new_AGEMA_signal_5500), .Z1_t (new_AGEMA_signal_5501), .Z1_f (new_AGEMA_signal_5502) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_12_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_12_Y), .A0_f (new_AGEMA_signal_5500), .A1_t (new_AGEMA_signal_5501), .A1_f (new_AGEMA_signal_5502), .B0_t (MCout[12]), .B0_f (new_AGEMA_signal_5265), .B1_t (new_AGEMA_signal_5266), .B1_f (new_AGEMA_signal_5267), .Z0_t (StateInMC[12]), .Z0_f (new_AGEMA_signal_5693), .Z1_t (new_AGEMA_signal_5694), .Z1_f (new_AGEMA_signal_5695) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_13_XOR1_U1 ( .A0_t (MCout[13]), .A0_f (new_AGEMA_signal_5091), .A1_t (new_AGEMA_signal_5092), .A1_f (new_AGEMA_signal_5093), .B0_t (MixColumns_line2_S02[6]), .B0_f (new_AGEMA_signal_3019), .B1_t (new_AGEMA_signal_3020), .B1_f (new_AGEMA_signal_3021), .Z0_t (MUX_StateInMC_mux_inst_13_X), .Z0_f (new_AGEMA_signal_5184), .Z1_t (new_AGEMA_signal_5185), .Z1_f (new_AGEMA_signal_5186) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_13_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_4669), .B0_t (MUX_StateInMC_mux_inst_13_X), .B0_f (new_AGEMA_signal_5184), .B1_t (new_AGEMA_signal_5185), .B1_f (new_AGEMA_signal_5186), .Z0_t (MUX_StateInMC_mux_inst_13_Y), .Z0_f (new_AGEMA_signal_5349), .Z1_t (new_AGEMA_signal_5350), .Z1_f (new_AGEMA_signal_5351) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_13_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_13_Y), .A0_f (new_AGEMA_signal_5349), .A1_t (new_AGEMA_signal_5350), .A1_f (new_AGEMA_signal_5351), .B0_t (MCout[13]), .B0_f (new_AGEMA_signal_5091), .B1_t (new_AGEMA_signal_5092), .B1_f (new_AGEMA_signal_5093), .Z0_t (StateInMC[13]), .Z0_f (new_AGEMA_signal_5503), .Z1_t (new_AGEMA_signal_5504), .Z1_f (new_AGEMA_signal_5505) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_14_XOR1_U1 ( .A0_t (MCout[14]), .A0_f (new_AGEMA_signal_5088), .A1_t (new_AGEMA_signal_5089), .A1_f (new_AGEMA_signal_5090), .B0_t (MixColumns_line2_S02[7]), .B0_f (new_AGEMA_signal_3025), .B1_t (new_AGEMA_signal_3026), .B1_f (new_AGEMA_signal_3027), .Z0_t (MUX_StateInMC_mux_inst_14_X), .Z0_f (new_AGEMA_signal_5187), .Z1_t (new_AGEMA_signal_5188), .Z1_f (new_AGEMA_signal_5189) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_14_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_4669), .B0_t (MUX_StateInMC_mux_inst_14_X), .B0_f (new_AGEMA_signal_5187), .B1_t (new_AGEMA_signal_5188), .B1_f (new_AGEMA_signal_5189), .Z0_t (MUX_StateInMC_mux_inst_14_Y), .Z0_f (new_AGEMA_signal_5352), .Z1_t (new_AGEMA_signal_5353), .Z1_f (new_AGEMA_signal_5354) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_14_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_14_Y), .A0_f (new_AGEMA_signal_5352), .A1_t (new_AGEMA_signal_5353), .A1_f (new_AGEMA_signal_5354), .B0_t (MCout[14]), .B0_f (new_AGEMA_signal_5088), .B1_t (new_AGEMA_signal_5089), .B1_f (new_AGEMA_signal_5090), .Z0_t (StateInMC[14]), .Z0_f (new_AGEMA_signal_5506), .Z1_t (new_AGEMA_signal_5507), .Z1_f (new_AGEMA_signal_5508) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_15_XOR1_U1 ( .A0_t (MCout[15]), .A0_f (new_AGEMA_signal_5085), .A1_t (new_AGEMA_signal_5086), .A1_f (new_AGEMA_signal_5087), .B0_t (MixColumns_line2_S02[0]), .B0_f (new_AGEMA_signal_3031), .B1_t (new_AGEMA_signal_3032), .B1_f (new_AGEMA_signal_3033), .Z0_t (MUX_StateInMC_mux_inst_15_X), .Z0_f (new_AGEMA_signal_5190), .Z1_t (new_AGEMA_signal_5191), .Z1_f (new_AGEMA_signal_5192) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_15_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_4669), .B0_t (MUX_StateInMC_mux_inst_15_X), .B0_f (new_AGEMA_signal_5190), .B1_t (new_AGEMA_signal_5191), .B1_f (new_AGEMA_signal_5192), .Z0_t (MUX_StateInMC_mux_inst_15_Y), .Z0_f (new_AGEMA_signal_5355), .Z1_t (new_AGEMA_signal_5356), .Z1_f (new_AGEMA_signal_5357) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_15_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_15_Y), .A0_f (new_AGEMA_signal_5355), .A1_t (new_AGEMA_signal_5356), .A1_f (new_AGEMA_signal_5357), .B0_t (MCout[15]), .B0_f (new_AGEMA_signal_5085), .B1_t (new_AGEMA_signal_5086), .B1_f (new_AGEMA_signal_5087), .Z0_t (StateInMC[15]), .Z0_f (new_AGEMA_signal_5509), .Z1_t (new_AGEMA_signal_5510), .Z1_f (new_AGEMA_signal_5511) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_16_XOR1_U1 ( .A0_t (MCout[16]), .A0_f (new_AGEMA_signal_5082), .A1_t (new_AGEMA_signal_5083), .A1_f (new_AGEMA_signal_5084), .B0_t (MCin[16]), .B0_f (new_AGEMA_signal_3988), .B1_t (new_AGEMA_signal_3989), .B1_f (new_AGEMA_signal_3990), .Z0_t (MUX_StateInMC_mux_inst_16_X), .Z0_f (new_AGEMA_signal_5193), .Z1_t (new_AGEMA_signal_5194), .Z1_f (new_AGEMA_signal_5195) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_16_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_4669), .B0_t (MUX_StateInMC_mux_inst_16_X), .B0_f (new_AGEMA_signal_5193), .B1_t (new_AGEMA_signal_5194), .B1_f (new_AGEMA_signal_5195), .Z0_t (MUX_StateInMC_mux_inst_16_Y), .Z0_f (new_AGEMA_signal_5358), .Z1_t (new_AGEMA_signal_5359), .Z1_f (new_AGEMA_signal_5360) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_16_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_16_Y), .A0_f (new_AGEMA_signal_5358), .A1_t (new_AGEMA_signal_5359), .A1_f (new_AGEMA_signal_5360), .B0_t (MCout[16]), .B0_f (new_AGEMA_signal_5082), .B1_t (new_AGEMA_signal_5083), .B1_f (new_AGEMA_signal_5084), .Z0_t (StateInMC[16]), .Z0_f (new_AGEMA_signal_5512), .Z1_t (new_AGEMA_signal_5513), .Z1_f (new_AGEMA_signal_5514) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_17_XOR1_U1 ( .A0_t (MCout[17]), .A0_f (new_AGEMA_signal_5262), .A1_t (new_AGEMA_signal_5263), .A1_f (new_AGEMA_signal_5264), .B0_t (MixColumns_line1_S02[2]), .B0_f (new_AGEMA_signal_3982), .B1_t (new_AGEMA_signal_3983), .B1_f (new_AGEMA_signal_3984), .Z0_t (MUX_StateInMC_mux_inst_17_X), .Z0_f (new_AGEMA_signal_5361), .Z1_t (new_AGEMA_signal_5362), .Z1_f (new_AGEMA_signal_5363) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_17_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_4669), .B0_t (MUX_StateInMC_mux_inst_17_X), .B0_f (new_AGEMA_signal_5361), .B1_t (new_AGEMA_signal_5362), .B1_f (new_AGEMA_signal_5363), .Z0_t (MUX_StateInMC_mux_inst_17_Y), .Z0_f (new_AGEMA_signal_5515), .Z1_t (new_AGEMA_signal_5516), .Z1_f (new_AGEMA_signal_5517) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_17_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_17_Y), .A0_f (new_AGEMA_signal_5515), .A1_t (new_AGEMA_signal_5516), .A1_f (new_AGEMA_signal_5517), .B0_t (MCout[17]), .B0_f (new_AGEMA_signal_5262), .B1_t (new_AGEMA_signal_5263), .B1_f (new_AGEMA_signal_5264), .Z0_t (StateInMC[17]), .Z0_f (new_AGEMA_signal_5696), .Z1_t (new_AGEMA_signal_5697), .Z1_f (new_AGEMA_signal_5698) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_18_XOR1_U1 ( .A0_t (MCout[18]), .A0_f (new_AGEMA_signal_5076), .A1_t (new_AGEMA_signal_5077), .A1_f (new_AGEMA_signal_5078), .B0_t (MCin[18]), .B0_f (new_AGEMA_signal_3979), .B1_t (new_AGEMA_signal_3980), .B1_f (new_AGEMA_signal_3981), .Z0_t (MUX_StateInMC_mux_inst_18_X), .Z0_f (new_AGEMA_signal_5196), .Z1_t (new_AGEMA_signal_5197), .Z1_f (new_AGEMA_signal_5198) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_18_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_4669), .B0_t (MUX_StateInMC_mux_inst_18_X), .B0_f (new_AGEMA_signal_5196), .B1_t (new_AGEMA_signal_5197), .B1_f (new_AGEMA_signal_5198), .Z0_t (MUX_StateInMC_mux_inst_18_Y), .Z0_f (new_AGEMA_signal_5364), .Z1_t (new_AGEMA_signal_5365), .Z1_f (new_AGEMA_signal_5366) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_18_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_18_Y), .A0_f (new_AGEMA_signal_5364), .A1_t (new_AGEMA_signal_5365), .A1_f (new_AGEMA_signal_5366), .B0_t (MCout[18]), .B0_f (new_AGEMA_signal_5076), .B1_t (new_AGEMA_signal_5077), .B1_f (new_AGEMA_signal_5078), .Z0_t (StateInMC[18]), .Z0_f (new_AGEMA_signal_5518), .Z1_t (new_AGEMA_signal_5519), .Z1_f (new_AGEMA_signal_5520) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_19_XOR1_U1 ( .A0_t (MCout[19]), .A0_f (new_AGEMA_signal_5259), .A1_t (new_AGEMA_signal_5260), .A1_f (new_AGEMA_signal_5261), .B0_t (MCin[19]), .B0_f (new_AGEMA_signal_3994), .B1_t (new_AGEMA_signal_3995), .B1_f (new_AGEMA_signal_3996), .Z0_t (MUX_StateInMC_mux_inst_19_X), .Z0_f (new_AGEMA_signal_5367), .Z1_t (new_AGEMA_signal_5368), .Z1_f (new_AGEMA_signal_5369) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_19_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_4669), .B0_t (MUX_StateInMC_mux_inst_19_X), .B0_f (new_AGEMA_signal_5367), .B1_t (new_AGEMA_signal_5368), .B1_f (new_AGEMA_signal_5369), .Z0_t (MUX_StateInMC_mux_inst_19_Y), .Z0_f (new_AGEMA_signal_5521), .Z1_t (new_AGEMA_signal_5522), .Z1_f (new_AGEMA_signal_5523) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_19_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_19_Y), .A0_f (new_AGEMA_signal_5521), .A1_t (new_AGEMA_signal_5522), .A1_f (new_AGEMA_signal_5523), .B0_t (MCout[19]), .B0_f (new_AGEMA_signal_5259), .B1_t (new_AGEMA_signal_5260), .B1_f (new_AGEMA_signal_5261), .Z0_t (StateInMC[19]), .Z0_f (new_AGEMA_signal_5699), .Z1_t (new_AGEMA_signal_5700), .Z1_f (new_AGEMA_signal_5701) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_20_XOR1_U1 ( .A0_t (MCout[20]), .A0_f (new_AGEMA_signal_5256), .A1_t (new_AGEMA_signal_5257), .A1_f (new_AGEMA_signal_5258), .B0_t (MixColumns_line1_S02[5]), .B0_f (new_AGEMA_signal_3973), .B1_t (new_AGEMA_signal_3974), .B1_f (new_AGEMA_signal_3975), .Z0_t (MUX_StateInMC_mux_inst_20_X), .Z0_f (new_AGEMA_signal_5370), .Z1_t (new_AGEMA_signal_5371), .Z1_f (new_AGEMA_signal_5372) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_20_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_4669), .B0_t (MUX_StateInMC_mux_inst_20_X), .B0_f (new_AGEMA_signal_5370), .B1_t (new_AGEMA_signal_5371), .B1_f (new_AGEMA_signal_5372), .Z0_t (MUX_StateInMC_mux_inst_20_Y), .Z0_f (new_AGEMA_signal_5524), .Z1_t (new_AGEMA_signal_5525), .Z1_f (new_AGEMA_signal_5526) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_20_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_20_Y), .A0_f (new_AGEMA_signal_5524), .A1_t (new_AGEMA_signal_5525), .A1_f (new_AGEMA_signal_5526), .B0_t (MCout[20]), .B0_f (new_AGEMA_signal_5256), .B1_t (new_AGEMA_signal_5257), .B1_f (new_AGEMA_signal_5258), .Z0_t (StateInMC[20]), .Z0_f (new_AGEMA_signal_5702), .Z1_t (new_AGEMA_signal_5703), .Z1_f (new_AGEMA_signal_5704) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_21_XOR1_U1 ( .A0_t (MCout[21]), .A0_f (new_AGEMA_signal_5067), .A1_t (new_AGEMA_signal_5068), .A1_f (new_AGEMA_signal_5069), .B0_t (MixColumns_line1_S02[6]), .B0_f (new_AGEMA_signal_3967), .B1_t (new_AGEMA_signal_3968), .B1_f (new_AGEMA_signal_3969), .Z0_t (MUX_StateInMC_mux_inst_21_X), .Z0_f (new_AGEMA_signal_5199), .Z1_t (new_AGEMA_signal_5200), .Z1_f (new_AGEMA_signal_5201) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_21_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_4669), .B0_t (MUX_StateInMC_mux_inst_21_X), .B0_f (new_AGEMA_signal_5199), .B1_t (new_AGEMA_signal_5200), .B1_f (new_AGEMA_signal_5201), .Z0_t (MUX_StateInMC_mux_inst_21_Y), .Z0_f (new_AGEMA_signal_5373), .Z1_t (new_AGEMA_signal_5374), .Z1_f (new_AGEMA_signal_5375) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_21_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_21_Y), .A0_f (new_AGEMA_signal_5373), .A1_t (new_AGEMA_signal_5374), .A1_f (new_AGEMA_signal_5375), .B0_t (MCout[21]), .B0_f (new_AGEMA_signal_5067), .B1_t (new_AGEMA_signal_5068), .B1_f (new_AGEMA_signal_5069), .Z0_t (StateInMC[21]), .Z0_f (new_AGEMA_signal_5527), .Z1_t (new_AGEMA_signal_5528), .Z1_f (new_AGEMA_signal_5529) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_22_XOR1_U1 ( .A0_t (MCout[22]), .A0_f (new_AGEMA_signal_5064), .A1_t (new_AGEMA_signal_5065), .A1_f (new_AGEMA_signal_5066), .B0_t (MixColumns_line1_S02[7]), .B0_f (new_AGEMA_signal_3961), .B1_t (new_AGEMA_signal_3962), .B1_f (new_AGEMA_signal_3963), .Z0_t (MUX_StateInMC_mux_inst_22_X), .Z0_f (new_AGEMA_signal_5202), .Z1_t (new_AGEMA_signal_5203), .Z1_f (new_AGEMA_signal_5204) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_22_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_4669), .B0_t (MUX_StateInMC_mux_inst_22_X), .B0_f (new_AGEMA_signal_5202), .B1_t (new_AGEMA_signal_5203), .B1_f (new_AGEMA_signal_5204), .Z0_t (MUX_StateInMC_mux_inst_22_Y), .Z0_f (new_AGEMA_signal_5376), .Z1_t (new_AGEMA_signal_5377), .Z1_f (new_AGEMA_signal_5378) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_22_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_22_Y), .A0_f (new_AGEMA_signal_5376), .A1_t (new_AGEMA_signal_5377), .A1_f (new_AGEMA_signal_5378), .B0_t (MCout[22]), .B0_f (new_AGEMA_signal_5064), .B1_t (new_AGEMA_signal_5065), .B1_f (new_AGEMA_signal_5066), .Z0_t (StateInMC[22]), .Z0_f (new_AGEMA_signal_5530), .Z1_t (new_AGEMA_signal_5531), .Z1_f (new_AGEMA_signal_5532) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_23_XOR1_U1 ( .A0_t (MCout[23]), .A0_f (new_AGEMA_signal_5061), .A1_t (new_AGEMA_signal_5062), .A1_f (new_AGEMA_signal_5063), .B0_t (MixColumns_line1_S02[0]), .B0_f (new_AGEMA_signal_3958), .B1_t (new_AGEMA_signal_3959), .B1_f (new_AGEMA_signal_3960), .Z0_t (MUX_StateInMC_mux_inst_23_X), .Z0_f (new_AGEMA_signal_5205), .Z1_t (new_AGEMA_signal_5206), .Z1_f (new_AGEMA_signal_5207) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_23_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_4669), .B0_t (MUX_StateInMC_mux_inst_23_X), .B0_f (new_AGEMA_signal_5205), .B1_t (new_AGEMA_signal_5206), .B1_f (new_AGEMA_signal_5207), .Z0_t (MUX_StateInMC_mux_inst_23_Y), .Z0_f (new_AGEMA_signal_5379), .Z1_t (new_AGEMA_signal_5380), .Z1_f (new_AGEMA_signal_5381) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_23_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_23_Y), .A0_f (new_AGEMA_signal_5379), .A1_t (new_AGEMA_signal_5380), .A1_f (new_AGEMA_signal_5381), .B0_t (MCout[23]), .B0_f (new_AGEMA_signal_5061), .B1_t (new_AGEMA_signal_5062), .B1_f (new_AGEMA_signal_5063), .Z0_t (StateInMC[23]), .Z0_f (new_AGEMA_signal_5533), .Z1_t (new_AGEMA_signal_5534), .Z1_f (new_AGEMA_signal_5535) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_24_XOR1_U1 ( .A0_t (MCout[24]), .A0_f (new_AGEMA_signal_5058), .A1_t (new_AGEMA_signal_5059), .A1_f (new_AGEMA_signal_5060), .B0_t (port_out_s0_t[0]), .B0_f (port_out_s0_f[0]), .B1_t (port_out_s1_t[0]), .B1_f (port_out_s1_f[0]), .Z0_t (MUX_StateInMC_mux_inst_24_X), .Z0_f (new_AGEMA_signal_5208), .Z1_t (new_AGEMA_signal_5209), .Z1_f (new_AGEMA_signal_5210) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_24_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_4669), .B0_t (MUX_StateInMC_mux_inst_24_X), .B0_f (new_AGEMA_signal_5208), .B1_t (new_AGEMA_signal_5209), .B1_f (new_AGEMA_signal_5210), .Z0_t (MUX_StateInMC_mux_inst_24_Y), .Z0_f (new_AGEMA_signal_5382), .Z1_t (new_AGEMA_signal_5383), .Z1_f (new_AGEMA_signal_5384) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_24_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_24_Y), .A0_f (new_AGEMA_signal_5382), .A1_t (new_AGEMA_signal_5383), .A1_f (new_AGEMA_signal_5384), .B0_t (MCout[24]), .B0_f (new_AGEMA_signal_5058), .B1_t (new_AGEMA_signal_5059), .B1_f (new_AGEMA_signal_5060), .Z0_t (StateInMC[24]), .Z0_f (new_AGEMA_signal_5536), .Z1_t (new_AGEMA_signal_5537), .Z1_f (new_AGEMA_signal_5538) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_25_XOR1_U1 ( .A0_t (MCout[25]), .A0_f (new_AGEMA_signal_5253), .A1_t (new_AGEMA_signal_5254), .A1_f (new_AGEMA_signal_5255), .B0_t (port_out_s0_t[1]), .B0_f (port_out_s0_f[1]), .B1_t (port_out_s1_t[1]), .B1_f (port_out_s1_f[1]), .Z0_t (MUX_StateInMC_mux_inst_25_X), .Z0_f (new_AGEMA_signal_5385), .Z1_t (new_AGEMA_signal_5386), .Z1_f (new_AGEMA_signal_5387) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_25_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_4669), .B0_t (MUX_StateInMC_mux_inst_25_X), .B0_f (new_AGEMA_signal_5385), .B1_t (new_AGEMA_signal_5386), .B1_f (new_AGEMA_signal_5387), .Z0_t (MUX_StateInMC_mux_inst_25_Y), .Z0_f (new_AGEMA_signal_5539), .Z1_t (new_AGEMA_signal_5540), .Z1_f (new_AGEMA_signal_5541) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_25_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_25_Y), .A0_f (new_AGEMA_signal_5539), .A1_t (new_AGEMA_signal_5540), .A1_f (new_AGEMA_signal_5541), .B0_t (MCout[25]), .B0_f (new_AGEMA_signal_5253), .B1_t (new_AGEMA_signal_5254), .B1_f (new_AGEMA_signal_5255), .Z0_t (StateInMC[25]), .Z0_f (new_AGEMA_signal_5705), .Z1_t (new_AGEMA_signal_5706), .Z1_f (new_AGEMA_signal_5707) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_26_XOR1_U1 ( .A0_t (MCout[26]), .A0_f (new_AGEMA_signal_5052), .A1_t (new_AGEMA_signal_5053), .A1_f (new_AGEMA_signal_5054), .B0_t (port_out_s0_t[2]), .B0_f (port_out_s0_f[2]), .B1_t (port_out_s1_t[2]), .B1_f (port_out_s1_f[2]), .Z0_t (MUX_StateInMC_mux_inst_26_X), .Z0_f (new_AGEMA_signal_5211), .Z1_t (new_AGEMA_signal_5212), .Z1_f (new_AGEMA_signal_5213) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_26_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_4669), .B0_t (MUX_StateInMC_mux_inst_26_X), .B0_f (new_AGEMA_signal_5211), .B1_t (new_AGEMA_signal_5212), .B1_f (new_AGEMA_signal_5213), .Z0_t (MUX_StateInMC_mux_inst_26_Y), .Z0_f (new_AGEMA_signal_5388), .Z1_t (new_AGEMA_signal_5389), .Z1_f (new_AGEMA_signal_5390) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_26_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_26_Y), .A0_f (new_AGEMA_signal_5388), .A1_t (new_AGEMA_signal_5389), .A1_f (new_AGEMA_signal_5390), .B0_t (MCout[26]), .B0_f (new_AGEMA_signal_5052), .B1_t (new_AGEMA_signal_5053), .B1_f (new_AGEMA_signal_5054), .Z0_t (StateInMC[26]), .Z0_f (new_AGEMA_signal_5542), .Z1_t (new_AGEMA_signal_5543), .Z1_f (new_AGEMA_signal_5544) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_27_XOR1_U1 ( .A0_t (MCout[27]), .A0_f (new_AGEMA_signal_5250), .A1_t (new_AGEMA_signal_5251), .A1_f (new_AGEMA_signal_5252), .B0_t (port_out_s0_t[3]), .B0_f (port_out_s0_f[3]), .B1_t (port_out_s1_t[3]), .B1_f (port_out_s1_f[3]), .Z0_t (MUX_StateInMC_mux_inst_27_X), .Z0_f (new_AGEMA_signal_5391), .Z1_t (new_AGEMA_signal_5392), .Z1_f (new_AGEMA_signal_5393) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_27_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_4669), .B0_t (MUX_StateInMC_mux_inst_27_X), .B0_f (new_AGEMA_signal_5391), .B1_t (new_AGEMA_signal_5392), .B1_f (new_AGEMA_signal_5393), .Z0_t (MUX_StateInMC_mux_inst_27_Y), .Z0_f (new_AGEMA_signal_5545), .Z1_t (new_AGEMA_signal_5546), .Z1_f (new_AGEMA_signal_5547) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_27_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_27_Y), .A0_f (new_AGEMA_signal_5545), .A1_t (new_AGEMA_signal_5546), .A1_f (new_AGEMA_signal_5547), .B0_t (MCout[27]), .B0_f (new_AGEMA_signal_5250), .B1_t (new_AGEMA_signal_5251), .B1_f (new_AGEMA_signal_5252), .Z0_t (StateInMC[27]), .Z0_f (new_AGEMA_signal_5708), .Z1_t (new_AGEMA_signal_5709), .Z1_f (new_AGEMA_signal_5710) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_28_XOR1_U1 ( .A0_t (MCout[28]), .A0_f (new_AGEMA_signal_5247), .A1_t (new_AGEMA_signal_5248), .A1_f (new_AGEMA_signal_5249), .B0_t (port_out_s0_t[4]), .B0_f (port_out_s0_f[4]), .B1_t (port_out_s1_t[4]), .B1_f (port_out_s1_f[4]), .Z0_t (MUX_StateInMC_mux_inst_28_X), .Z0_f (new_AGEMA_signal_5394), .Z1_t (new_AGEMA_signal_5395), .Z1_f (new_AGEMA_signal_5396) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_28_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_4669), .B0_t (MUX_StateInMC_mux_inst_28_X), .B0_f (new_AGEMA_signal_5394), .B1_t (new_AGEMA_signal_5395), .B1_f (new_AGEMA_signal_5396), .Z0_t (MUX_StateInMC_mux_inst_28_Y), .Z0_f (new_AGEMA_signal_5548), .Z1_t (new_AGEMA_signal_5549), .Z1_f (new_AGEMA_signal_5550) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_28_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_28_Y), .A0_f (new_AGEMA_signal_5548), .A1_t (new_AGEMA_signal_5549), .A1_f (new_AGEMA_signal_5550), .B0_t (MCout[28]), .B0_f (new_AGEMA_signal_5247), .B1_t (new_AGEMA_signal_5248), .B1_f (new_AGEMA_signal_5249), .Z0_t (StateInMC[28]), .Z0_f (new_AGEMA_signal_5711), .Z1_t (new_AGEMA_signal_5712), .Z1_f (new_AGEMA_signal_5713) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_29_XOR1_U1 ( .A0_t (MCout[29]), .A0_f (new_AGEMA_signal_5043), .A1_t (new_AGEMA_signal_5044), .A1_f (new_AGEMA_signal_5045), .B0_t (port_out_s0_t[5]), .B0_f (port_out_s0_f[5]), .B1_t (port_out_s1_t[5]), .B1_f (port_out_s1_f[5]), .Z0_t (MUX_StateInMC_mux_inst_29_X), .Z0_f (new_AGEMA_signal_5214), .Z1_t (new_AGEMA_signal_5215), .Z1_f (new_AGEMA_signal_5216) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_29_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_4669), .B0_t (MUX_StateInMC_mux_inst_29_X), .B0_f (new_AGEMA_signal_5214), .B1_t (new_AGEMA_signal_5215), .B1_f (new_AGEMA_signal_5216), .Z0_t (MUX_StateInMC_mux_inst_29_Y), .Z0_f (new_AGEMA_signal_5397), .Z1_t (new_AGEMA_signal_5398), .Z1_f (new_AGEMA_signal_5399) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_29_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_29_Y), .A0_f (new_AGEMA_signal_5397), .A1_t (new_AGEMA_signal_5398), .A1_f (new_AGEMA_signal_5399), .B0_t (MCout[29]), .B0_f (new_AGEMA_signal_5043), .B1_t (new_AGEMA_signal_5044), .B1_f (new_AGEMA_signal_5045), .Z0_t (StateInMC[29]), .Z0_f (new_AGEMA_signal_5551), .Z1_t (new_AGEMA_signal_5552), .Z1_f (new_AGEMA_signal_5553) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_30_XOR1_U1 ( .A0_t (MCout[30]), .A0_f (new_AGEMA_signal_5040), .A1_t (new_AGEMA_signal_5041), .A1_f (new_AGEMA_signal_5042), .B0_t (port_out_s0_t[6]), .B0_f (port_out_s0_f[6]), .B1_t (port_out_s1_t[6]), .B1_f (port_out_s1_f[6]), .Z0_t (MUX_StateInMC_mux_inst_30_X), .Z0_f (new_AGEMA_signal_5217), .Z1_t (new_AGEMA_signal_5218), .Z1_f (new_AGEMA_signal_5219) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_30_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_4669), .B0_t (MUX_StateInMC_mux_inst_30_X), .B0_f (new_AGEMA_signal_5217), .B1_t (new_AGEMA_signal_5218), .B1_f (new_AGEMA_signal_5219), .Z0_t (MUX_StateInMC_mux_inst_30_Y), .Z0_f (new_AGEMA_signal_5400), .Z1_t (new_AGEMA_signal_5401), .Z1_f (new_AGEMA_signal_5402) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_30_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_30_Y), .A0_f (new_AGEMA_signal_5400), .A1_t (new_AGEMA_signal_5401), .A1_f (new_AGEMA_signal_5402), .B0_t (MCout[30]), .B0_f (new_AGEMA_signal_5040), .B1_t (new_AGEMA_signal_5041), .B1_f (new_AGEMA_signal_5042), .Z0_t (StateInMC[30]), .Z0_f (new_AGEMA_signal_5554), .Z1_t (new_AGEMA_signal_5555), .Z1_f (new_AGEMA_signal_5556) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_31_XOR1_U1 ( .A0_t (MCout[31]), .A0_f (new_AGEMA_signal_5037), .A1_t (new_AGEMA_signal_5038), .A1_f (new_AGEMA_signal_5039), .B0_t (port_out_s0_t[7]), .B0_f (port_out_s0_f[7]), .B1_t (port_out_s1_t[7]), .B1_f (port_out_s1_f[7]), .Z0_t (MUX_StateInMC_mux_inst_31_X), .Z0_f (new_AGEMA_signal_5220), .Z1_t (new_AGEMA_signal_5221), .Z1_f (new_AGEMA_signal_5222) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_31_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intFinal), .A1_f (new_AGEMA_signal_4669), .B0_t (MUX_StateInMC_mux_inst_31_X), .B0_f (new_AGEMA_signal_5220), .B1_t (new_AGEMA_signal_5221), .B1_f (new_AGEMA_signal_5222), .Z0_t (MUX_StateInMC_mux_inst_31_Y), .Z0_f (new_AGEMA_signal_5403), .Z1_t (new_AGEMA_signal_5404), .Z1_f (new_AGEMA_signal_5405) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_StateInMC_mux_inst_31_XOR2_U1 ( .A0_t (MUX_StateInMC_mux_inst_31_Y), .A0_f (new_AGEMA_signal_5403), .A1_t (new_AGEMA_signal_5404), .A1_f (new_AGEMA_signal_5405), .B0_t (MCout[31]), .B0_f (new_AGEMA_signal_5037), .B1_t (new_AGEMA_signal_5038), .B1_f (new_AGEMA_signal_5039), .Z0_t (StateInMC[31]), .Z0_f (new_AGEMA_signal_5557), .Z1_t (new_AGEMA_signal_5558), .Z1_f (new_AGEMA_signal_5559) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_U32 ( .A0_t (KeyArray_outS01ser_7_), .A0_f (new_AGEMA_signal_3205), .A1_t (new_AGEMA_signal_3206), .A1_f (new_AGEMA_signal_3207), .B0_t (keyStateIn[7]), .B0_f (new_AGEMA_signal_2552), .B1_t (new_AGEMA_signal_2553), .B1_f (new_AGEMA_signal_2554), .Z0_t (KeyArray_outS01ser_XOR_00[7]), .Z0_f (new_AGEMA_signal_3208), .Z1_t (new_AGEMA_signal_3209), .Z1_f (new_AGEMA_signal_3210) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_U31 ( .A0_t (KeyArray_outS01ser_6_), .A0_f (new_AGEMA_signal_3211), .A1_t (new_AGEMA_signal_3212), .A1_f (new_AGEMA_signal_3213), .B0_t (keyStateIn[6]), .B0_f (new_AGEMA_signal_2543), .B1_t (new_AGEMA_signal_2544), .B1_f (new_AGEMA_signal_2545), .Z0_t (KeyArray_outS01ser_XOR_00[6]), .Z0_f (new_AGEMA_signal_3214), .Z1_t (new_AGEMA_signal_3215), .Z1_f (new_AGEMA_signal_3216) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_U30 ( .A0_t (KeyArray_outS01ser_5_), .A0_f (new_AGEMA_signal_3217), .A1_t (new_AGEMA_signal_3218), .A1_f (new_AGEMA_signal_3219), .B0_t (keyStateIn[5]), .B0_f (new_AGEMA_signal_2534), .B1_t (new_AGEMA_signal_2535), .B1_f (new_AGEMA_signal_2536), .Z0_t (KeyArray_outS01ser_XOR_00[5]), .Z0_f (new_AGEMA_signal_3220), .Z1_t (new_AGEMA_signal_3221), .Z1_f (new_AGEMA_signal_3222) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_U29 ( .A0_t (KeyArray_outS01ser_4_), .A0_f (new_AGEMA_signal_3223), .A1_t (new_AGEMA_signal_3224), .A1_f (new_AGEMA_signal_3225), .B0_t (keyStateIn[4]), .B0_f (new_AGEMA_signal_2525), .B1_t (new_AGEMA_signal_2526), .B1_f (new_AGEMA_signal_2527), .Z0_t (KeyArray_outS01ser_XOR_00[4]), .Z0_f (new_AGEMA_signal_3226), .Z1_t (new_AGEMA_signal_3227), .Z1_f (new_AGEMA_signal_3228) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_U28 ( .A0_t (KeyArray_outS01ser_3_), .A0_f (new_AGEMA_signal_3229), .A1_t (new_AGEMA_signal_3230), .A1_f (new_AGEMA_signal_3231), .B0_t (keyStateIn[3]), .B0_f (new_AGEMA_signal_2516), .B1_t (new_AGEMA_signal_2517), .B1_f (new_AGEMA_signal_2518), .Z0_t (KeyArray_outS01ser_XOR_00[3]), .Z0_f (new_AGEMA_signal_3232), .Z1_t (new_AGEMA_signal_3233), .Z1_f (new_AGEMA_signal_3234) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_U27 ( .A0_t (KeyArray_outS01ser_2_), .A0_f (new_AGEMA_signal_3235), .A1_t (new_AGEMA_signal_3236), .A1_f (new_AGEMA_signal_3237), .B0_t (keyStateIn[2]), .B0_f (new_AGEMA_signal_2507), .B1_t (new_AGEMA_signal_2508), .B1_f (new_AGEMA_signal_2509), .Z0_t (KeyArray_outS01ser_XOR_00[2]), .Z0_f (new_AGEMA_signal_3238), .Z1_t (new_AGEMA_signal_3239), .Z1_f (new_AGEMA_signal_3240) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_U26 ( .A0_t (KeyArray_outS01ser_1_), .A0_f (new_AGEMA_signal_3241), .A1_t (new_AGEMA_signal_3242), .A1_f (new_AGEMA_signal_3243), .B0_t (keyStateIn[1]), .B0_f (new_AGEMA_signal_2498), .B1_t (new_AGEMA_signal_2499), .B1_f (new_AGEMA_signal_2500), .Z0_t (KeyArray_outS01ser_XOR_00[1]), .Z0_f (new_AGEMA_signal_3244), .Z1_t (new_AGEMA_signal_3245), .Z1_f (new_AGEMA_signal_3246) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_U25 ( .A0_t (KeyArray_outS01ser_0_), .A0_f (new_AGEMA_signal_3247), .A1_t (new_AGEMA_signal_3248), .A1_f (new_AGEMA_signal_3249), .B0_t (keyStateIn[0]), .B0_f (new_AGEMA_signal_2489), .B1_t (new_AGEMA_signal_2490), .B1_f (new_AGEMA_signal_2491), .Z0_t (KeyArray_outS01ser_XOR_00[0]), .Z0_f (new_AGEMA_signal_3250), .Z1_t (new_AGEMA_signal_3251), .Z1_f (new_AGEMA_signal_3252) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) KeyArray_U24 ( .A0_t (start_t), .A0_f (start_f), .B0_t (intselXOR), .B0_f (new_AGEMA_signal_5158), .Z0_t (KeyArray_nReset_selXOR), .Z0_f (new_AGEMA_signal_5406) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_U23 ( .A0_t (KeyArray_n32), .A0_f (new_AGEMA_signal_7556), .A1_t (new_AGEMA_signal_7557), .A1_f (new_AGEMA_signal_7558), .B0_t (keyStateIn[7]), .B0_f (new_AGEMA_signal_2552), .B1_t (new_AGEMA_signal_2553), .B1_f (new_AGEMA_signal_2554), .Z0_t (KeyArray_inS30par[7]), .Z0_f (new_AGEMA_signal_7604), .Z1_t (new_AGEMA_signal_7605), .Z1_f (new_AGEMA_signal_7606) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_U22 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (roundConstant[7]), .A1_f (new_AGEMA_signal_4179), .B0_t (SboxOut[7]), .B0_f (new_AGEMA_signal_7511), .B1_t (new_AGEMA_signal_7512), .B1_f (new_AGEMA_signal_7513), .Z0_t (KeyArray_n32), .Z0_f (new_AGEMA_signal_7556), .Z1_t (new_AGEMA_signal_7557), .Z1_f (new_AGEMA_signal_7558) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_U21 ( .A0_t (KeyArray_n31), .A0_f (new_AGEMA_signal_7559), .A1_t (new_AGEMA_signal_7560), .A1_f (new_AGEMA_signal_7561), .B0_t (keyStateIn[6]), .B0_f (new_AGEMA_signal_2543), .B1_t (new_AGEMA_signal_2544), .B1_f (new_AGEMA_signal_2545), .Z0_t (KeyArray_inS30par[6]), .Z0_f (new_AGEMA_signal_7607), .Z1_t (new_AGEMA_signal_7608), .Z1_f (new_AGEMA_signal_7609) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_U20 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (roundConstant[6]), .A1_f (new_AGEMA_signal_4181), .B0_t (SboxOut[6]), .B0_f (new_AGEMA_signal_7514), .B1_t (new_AGEMA_signal_7515), .B1_f (new_AGEMA_signal_7516), .Z0_t (KeyArray_n31), .Z0_f (new_AGEMA_signal_7559), .Z1_t (new_AGEMA_signal_7560), .Z1_f (new_AGEMA_signal_7561) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_U19 ( .A0_t (KeyArray_n30), .A0_f (new_AGEMA_signal_7562), .A1_t (new_AGEMA_signal_7563), .A1_f (new_AGEMA_signal_7564), .B0_t (keyStateIn[5]), .B0_f (new_AGEMA_signal_2534), .B1_t (new_AGEMA_signal_2535), .B1_f (new_AGEMA_signal_2536), .Z0_t (KeyArray_inS30par[5]), .Z0_f (new_AGEMA_signal_7610), .Z1_t (new_AGEMA_signal_7611), .Z1_f (new_AGEMA_signal_7612) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_U18 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (roundConstant[5]), .A1_f (new_AGEMA_signal_4183), .B0_t (SboxOut[5]), .B0_f (new_AGEMA_signal_7517), .B1_t (new_AGEMA_signal_7518), .B1_f (new_AGEMA_signal_7519), .Z0_t (KeyArray_n30), .Z0_f (new_AGEMA_signal_7562), .Z1_t (new_AGEMA_signal_7563), .Z1_f (new_AGEMA_signal_7564) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_U17 ( .A0_t (KeyArray_n29), .A0_f (new_AGEMA_signal_7565), .A1_t (new_AGEMA_signal_7566), .A1_f (new_AGEMA_signal_7567), .B0_t (keyStateIn[4]), .B0_f (new_AGEMA_signal_2525), .B1_t (new_AGEMA_signal_2526), .B1_f (new_AGEMA_signal_2527), .Z0_t (KeyArray_inS30par[4]), .Z0_f (new_AGEMA_signal_7613), .Z1_t (new_AGEMA_signal_7614), .Z1_f (new_AGEMA_signal_7615) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_U16 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (roundConstant[4]), .A1_f (new_AGEMA_signal_4185), .B0_t (SboxOut[4]), .B0_f (new_AGEMA_signal_7520), .B1_t (new_AGEMA_signal_7521), .B1_f (new_AGEMA_signal_7522), .Z0_t (KeyArray_n29), .Z0_f (new_AGEMA_signal_7565), .Z1_t (new_AGEMA_signal_7566), .Z1_f (new_AGEMA_signal_7567) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_U15 ( .A0_t (KeyArray_n28), .A0_f (new_AGEMA_signal_7568), .A1_t (new_AGEMA_signal_7569), .A1_f (new_AGEMA_signal_7570), .B0_t (keyStateIn[3]), .B0_f (new_AGEMA_signal_2516), .B1_t (new_AGEMA_signal_2517), .B1_f (new_AGEMA_signal_2518), .Z0_t (KeyArray_inS30par[3]), .Z0_f (new_AGEMA_signal_7616), .Z1_t (new_AGEMA_signal_7617), .Z1_f (new_AGEMA_signal_7618) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_U14 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (roundConstant[3]), .A1_f (new_AGEMA_signal_4187), .B0_t (SboxOut[3]), .B0_f (new_AGEMA_signal_7523), .B1_t (new_AGEMA_signal_7524), .B1_f (new_AGEMA_signal_7525), .Z0_t (KeyArray_n28), .Z0_f (new_AGEMA_signal_7568), .Z1_t (new_AGEMA_signal_7569), .Z1_f (new_AGEMA_signal_7570) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_U13 ( .A0_t (KeyArray_n27), .A0_f (new_AGEMA_signal_7571), .A1_t (new_AGEMA_signal_7572), .A1_f (new_AGEMA_signal_7573), .B0_t (keyStateIn[2]), .B0_f (new_AGEMA_signal_2507), .B1_t (new_AGEMA_signal_2508), .B1_f (new_AGEMA_signal_2509), .Z0_t (KeyArray_inS30par[2]), .Z0_f (new_AGEMA_signal_7619), .Z1_t (new_AGEMA_signal_7620), .Z1_f (new_AGEMA_signal_7621) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_U12 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (roundConstant[2]), .A1_f (new_AGEMA_signal_4189), .B0_t (SboxOut[2]), .B0_f (new_AGEMA_signal_7526), .B1_t (new_AGEMA_signal_7527), .B1_f (new_AGEMA_signal_7528), .Z0_t (KeyArray_n27), .Z0_f (new_AGEMA_signal_7571), .Z1_t (new_AGEMA_signal_7572), .Z1_f (new_AGEMA_signal_7573) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_U11 ( .A0_t (KeyArray_n26), .A0_f (new_AGEMA_signal_7574), .A1_t (new_AGEMA_signal_7575), .A1_f (new_AGEMA_signal_7576), .B0_t (keyStateIn[1]), .B0_f (new_AGEMA_signal_2498), .B1_t (new_AGEMA_signal_2499), .B1_f (new_AGEMA_signal_2500), .Z0_t (KeyArray_inS30par[1]), .Z0_f (new_AGEMA_signal_7622), .Z1_t (new_AGEMA_signal_7623), .Z1_f (new_AGEMA_signal_7624) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_U10 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (roundConstant[1]), .A1_f (new_AGEMA_signal_4191), .B0_t (SboxOut[1]), .B0_f (new_AGEMA_signal_7529), .B1_t (new_AGEMA_signal_7530), .B1_f (new_AGEMA_signal_7531), .Z0_t (KeyArray_n26), .Z0_f (new_AGEMA_signal_7574), .Z1_t (new_AGEMA_signal_7575), .Z1_f (new_AGEMA_signal_7576) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_U9 ( .A0_t (KeyArray_n25), .A0_f (new_AGEMA_signal_7508), .A1_t (new_AGEMA_signal_7509), .A1_f (new_AGEMA_signal_7510), .B0_t (keyStateIn[0]), .B0_f (new_AGEMA_signal_2489), .B1_t (new_AGEMA_signal_2490), .B1_f (new_AGEMA_signal_2491), .Z0_t (KeyArray_inS30par[0]), .Z0_f (new_AGEMA_signal_7577), .Z1_t (new_AGEMA_signal_7578), .Z1_f (new_AGEMA_signal_7579) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_U8 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (roundConstant[0]), .A1_f (new_AGEMA_signal_4193), .B0_t (SboxOut[0]), .B0_f (new_AGEMA_signal_7502), .B1_t (new_AGEMA_signal_7503), .B1_f (new_AGEMA_signal_7504), .Z0_t (KeyArray_n25), .Z0_f (new_AGEMA_signal_7508), .Z1_t (new_AGEMA_signal_7509), .Z1_f (new_AGEMA_signal_7510) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S00reg_gff_1_SFF_0_U3 ( .A0_t (KeyArray_S00reg_gff_1_SFF_0_n2), .A0_f (new_AGEMA_signal_7230), .A1_t (new_AGEMA_signal_7231), .A1_f (new_AGEMA_signal_7232), .B0_t (KeyArray_S00reg_gff_1_SFF_0_n1), .B0_f (new_AGEMA_signal_6391), .B1_t (new_AGEMA_signal_6392), .B1_f (new_AGEMA_signal_6393), .Z0_t (keyStateIn[0]), .Z0_f (new_AGEMA_signal_2489), .Z1_t (new_AGEMA_signal_2490), .Z1_f (new_AGEMA_signal_2491) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_0_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (keyStateIn[0]), .B0_f (new_AGEMA_signal_2489), .B1_t (new_AGEMA_signal_2490), .B1_f (new_AGEMA_signal_2491), .Z0_t (KeyArray_S00reg_gff_1_SFF_0_n1), .Z0_f (new_AGEMA_signal_6391), .Z1_t (new_AGEMA_signal_6392), .Z1_f (new_AGEMA_signal_6393) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_0_U1 ( .A0_t (KeyArray_S00reg_gff_1_SFF_0_QD), .A0_f (new_AGEMA_signal_6394), .A1_t (new_AGEMA_signal_6395), .A1_f (new_AGEMA_signal_6396), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S00reg_gff_1_SFF_0_n2), .Z0_f (new_AGEMA_signal_7230), .Z1_t (new_AGEMA_signal_7231), .Z1_f (new_AGEMA_signal_7232) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS00ser[0]), .A0_f (new_AGEMA_signal_5714), .A1_t (new_AGEMA_signal_5715), .A1_f (new_AGEMA_signal_5716), .B0_t (KeyArray_outS10ser[0]), .B0_f (new_AGEMA_signal_3397), .B1_t (new_AGEMA_signal_3398), .B1_f (new_AGEMA_signal_3399), .Z0_t (KeyArray_S00reg_gff_1_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_5865), .Z1_t (new_AGEMA_signal_5866), .Z1_f (new_AGEMA_signal_5867) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S00reg_gff_1_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_5865), .B1_t (new_AGEMA_signal_5866), .B1_f (new_AGEMA_signal_5867), .Z0_t (KeyArray_S00reg_gff_1_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_6277), .Z1_t (new_AGEMA_signal_6278), .Z1_f (new_AGEMA_signal_6279) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S00reg_gff_1_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_6277), .A1_t (new_AGEMA_signal_6278), .A1_f (new_AGEMA_signal_6279), .B0_t (KeyArray_inS00ser[0]), .B0_f (new_AGEMA_signal_5714), .B1_t (new_AGEMA_signal_5715), .B1_f (new_AGEMA_signal_5716), .Z0_t (KeyArray_S00reg_gff_1_SFF_0_QD), .Z0_f (new_AGEMA_signal_6394), .Z1_t (new_AGEMA_signal_6395), .Z1_f (new_AGEMA_signal_6396) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S00reg_gff_1_SFF_1_U3 ( .A0_t (KeyArray_S00reg_gff_1_SFF_1_n2), .A0_f (new_AGEMA_signal_7233), .A1_t (new_AGEMA_signal_7234), .A1_f (new_AGEMA_signal_7235), .B0_t (KeyArray_S00reg_gff_1_SFF_1_n1), .B0_f (new_AGEMA_signal_6397), .B1_t (new_AGEMA_signal_6398), .B1_f (new_AGEMA_signal_6399), .Z0_t (keyStateIn[1]), .Z0_f (new_AGEMA_signal_2498), .Z1_t (new_AGEMA_signal_2499), .Z1_f (new_AGEMA_signal_2500) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_1_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (keyStateIn[1]), .B0_f (new_AGEMA_signal_2498), .B1_t (new_AGEMA_signal_2499), .B1_f (new_AGEMA_signal_2500), .Z0_t (KeyArray_S00reg_gff_1_SFF_1_n1), .Z0_f (new_AGEMA_signal_6397), .Z1_t (new_AGEMA_signal_6398), .Z1_f (new_AGEMA_signal_6399) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_1_U1 ( .A0_t (KeyArray_S00reg_gff_1_SFF_1_QD), .A0_f (new_AGEMA_signal_6400), .A1_t (new_AGEMA_signal_6401), .A1_f (new_AGEMA_signal_6402), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S00reg_gff_1_SFF_1_n2), .Z0_f (new_AGEMA_signal_7233), .Z1_t (new_AGEMA_signal_7234), .Z1_f (new_AGEMA_signal_7235) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS00ser[1]), .A0_f (new_AGEMA_signal_5717), .A1_t (new_AGEMA_signal_5718), .A1_f (new_AGEMA_signal_5719), .B0_t (KeyArray_outS10ser[1]), .B0_f (new_AGEMA_signal_3406), .B1_t (new_AGEMA_signal_3407), .B1_f (new_AGEMA_signal_3408), .Z0_t (KeyArray_S00reg_gff_1_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_5868), .Z1_t (new_AGEMA_signal_5869), .Z1_f (new_AGEMA_signal_5870) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S00reg_gff_1_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_5868), .B1_t (new_AGEMA_signal_5869), .B1_f (new_AGEMA_signal_5870), .Z0_t (KeyArray_S00reg_gff_1_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_6280), .Z1_t (new_AGEMA_signal_6281), .Z1_f (new_AGEMA_signal_6282) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S00reg_gff_1_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_6280), .A1_t (new_AGEMA_signal_6281), .A1_f (new_AGEMA_signal_6282), .B0_t (KeyArray_inS00ser[1]), .B0_f (new_AGEMA_signal_5717), .B1_t (new_AGEMA_signal_5718), .B1_f (new_AGEMA_signal_5719), .Z0_t (KeyArray_S00reg_gff_1_SFF_1_QD), .Z0_f (new_AGEMA_signal_6400), .Z1_t (new_AGEMA_signal_6401), .Z1_f (new_AGEMA_signal_6402) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S00reg_gff_1_SFF_2_U3 ( .A0_t (KeyArray_S00reg_gff_1_SFF_2_n2), .A0_f (new_AGEMA_signal_7236), .A1_t (new_AGEMA_signal_7237), .A1_f (new_AGEMA_signal_7238), .B0_t (KeyArray_S00reg_gff_1_SFF_2_n1), .B0_f (new_AGEMA_signal_6403), .B1_t (new_AGEMA_signal_6404), .B1_f (new_AGEMA_signal_6405), .Z0_t (keyStateIn[2]), .Z0_f (new_AGEMA_signal_2507), .Z1_t (new_AGEMA_signal_2508), .Z1_f (new_AGEMA_signal_2509) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_2_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (keyStateIn[2]), .B0_f (new_AGEMA_signal_2507), .B1_t (new_AGEMA_signal_2508), .B1_f (new_AGEMA_signal_2509), .Z0_t (KeyArray_S00reg_gff_1_SFF_2_n1), .Z0_f (new_AGEMA_signal_6403), .Z1_t (new_AGEMA_signal_6404), .Z1_f (new_AGEMA_signal_6405) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_2_U1 ( .A0_t (KeyArray_S00reg_gff_1_SFF_2_QD), .A0_f (new_AGEMA_signal_6406), .A1_t (new_AGEMA_signal_6407), .A1_f (new_AGEMA_signal_6408), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S00reg_gff_1_SFF_2_n2), .Z0_f (new_AGEMA_signal_7236), .Z1_t (new_AGEMA_signal_7237), .Z1_f (new_AGEMA_signal_7238) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS00ser[2]), .A0_f (new_AGEMA_signal_5720), .A1_t (new_AGEMA_signal_5721), .A1_f (new_AGEMA_signal_5722), .B0_t (KeyArray_outS10ser[2]), .B0_f (new_AGEMA_signal_3415), .B1_t (new_AGEMA_signal_3416), .B1_f (new_AGEMA_signal_3417), .Z0_t (KeyArray_S00reg_gff_1_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_5871), .Z1_t (new_AGEMA_signal_5872), .Z1_f (new_AGEMA_signal_5873) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S00reg_gff_1_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_5871), .B1_t (new_AGEMA_signal_5872), .B1_f (new_AGEMA_signal_5873), .Z0_t (KeyArray_S00reg_gff_1_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_6283), .Z1_t (new_AGEMA_signal_6284), .Z1_f (new_AGEMA_signal_6285) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S00reg_gff_1_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_6283), .A1_t (new_AGEMA_signal_6284), .A1_f (new_AGEMA_signal_6285), .B0_t (KeyArray_inS00ser[2]), .B0_f (new_AGEMA_signal_5720), .B1_t (new_AGEMA_signal_5721), .B1_f (new_AGEMA_signal_5722), .Z0_t (KeyArray_S00reg_gff_1_SFF_2_QD), .Z0_f (new_AGEMA_signal_6406), .Z1_t (new_AGEMA_signal_6407), .Z1_f (new_AGEMA_signal_6408) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S00reg_gff_1_SFF_3_U3 ( .A0_t (KeyArray_S00reg_gff_1_SFF_3_n2), .A0_f (new_AGEMA_signal_7239), .A1_t (new_AGEMA_signal_7240), .A1_f (new_AGEMA_signal_7241), .B0_t (KeyArray_S00reg_gff_1_SFF_3_n1), .B0_f (new_AGEMA_signal_6409), .B1_t (new_AGEMA_signal_6410), .B1_f (new_AGEMA_signal_6411), .Z0_t (keyStateIn[3]), .Z0_f (new_AGEMA_signal_2516), .Z1_t (new_AGEMA_signal_2517), .Z1_f (new_AGEMA_signal_2518) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_3_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (keyStateIn[3]), .B0_f (new_AGEMA_signal_2516), .B1_t (new_AGEMA_signal_2517), .B1_f (new_AGEMA_signal_2518), .Z0_t (KeyArray_S00reg_gff_1_SFF_3_n1), .Z0_f (new_AGEMA_signal_6409), .Z1_t (new_AGEMA_signal_6410), .Z1_f (new_AGEMA_signal_6411) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_3_U1 ( .A0_t (KeyArray_S00reg_gff_1_SFF_3_QD), .A0_f (new_AGEMA_signal_6412), .A1_t (new_AGEMA_signal_6413), .A1_f (new_AGEMA_signal_6414), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S00reg_gff_1_SFF_3_n2), .Z0_f (new_AGEMA_signal_7239), .Z1_t (new_AGEMA_signal_7240), .Z1_f (new_AGEMA_signal_7241) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS00ser[3]), .A0_f (new_AGEMA_signal_5723), .A1_t (new_AGEMA_signal_5724), .A1_f (new_AGEMA_signal_5725), .B0_t (KeyArray_outS10ser[3]), .B0_f (new_AGEMA_signal_3424), .B1_t (new_AGEMA_signal_3425), .B1_f (new_AGEMA_signal_3426), .Z0_t (KeyArray_S00reg_gff_1_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_5874), .Z1_t (new_AGEMA_signal_5875), .Z1_f (new_AGEMA_signal_5876) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S00reg_gff_1_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_5874), .B1_t (new_AGEMA_signal_5875), .B1_f (new_AGEMA_signal_5876), .Z0_t (KeyArray_S00reg_gff_1_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_6286), .Z1_t (new_AGEMA_signal_6287), .Z1_f (new_AGEMA_signal_6288) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S00reg_gff_1_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_6286), .A1_t (new_AGEMA_signal_6287), .A1_f (new_AGEMA_signal_6288), .B0_t (KeyArray_inS00ser[3]), .B0_f (new_AGEMA_signal_5723), .B1_t (new_AGEMA_signal_5724), .B1_f (new_AGEMA_signal_5725), .Z0_t (KeyArray_S00reg_gff_1_SFF_3_QD), .Z0_f (new_AGEMA_signal_6412), .Z1_t (new_AGEMA_signal_6413), .Z1_f (new_AGEMA_signal_6414) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S00reg_gff_1_SFF_4_U3 ( .A0_t (KeyArray_S00reg_gff_1_SFF_4_n2), .A0_f (new_AGEMA_signal_7242), .A1_t (new_AGEMA_signal_7243), .A1_f (new_AGEMA_signal_7244), .B0_t (KeyArray_S00reg_gff_1_SFF_4_n1), .B0_f (new_AGEMA_signal_6415), .B1_t (new_AGEMA_signal_6416), .B1_f (new_AGEMA_signal_6417), .Z0_t (keyStateIn[4]), .Z0_f (new_AGEMA_signal_2525), .Z1_t (new_AGEMA_signal_2526), .Z1_f (new_AGEMA_signal_2527) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_4_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (keyStateIn[4]), .B0_f (new_AGEMA_signal_2525), .B1_t (new_AGEMA_signal_2526), .B1_f (new_AGEMA_signal_2527), .Z0_t (KeyArray_S00reg_gff_1_SFF_4_n1), .Z0_f (new_AGEMA_signal_6415), .Z1_t (new_AGEMA_signal_6416), .Z1_f (new_AGEMA_signal_6417) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_4_U1 ( .A0_t (KeyArray_S00reg_gff_1_SFF_4_QD), .A0_f (new_AGEMA_signal_6418), .A1_t (new_AGEMA_signal_6419), .A1_f (new_AGEMA_signal_6420), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S00reg_gff_1_SFF_4_n2), .Z0_f (new_AGEMA_signal_7242), .Z1_t (new_AGEMA_signal_7243), .Z1_f (new_AGEMA_signal_7244) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS00ser[4]), .A0_f (new_AGEMA_signal_5726), .A1_t (new_AGEMA_signal_5727), .A1_f (new_AGEMA_signal_5728), .B0_t (KeyArray_outS10ser[4]), .B0_f (new_AGEMA_signal_3433), .B1_t (new_AGEMA_signal_3434), .B1_f (new_AGEMA_signal_3435), .Z0_t (KeyArray_S00reg_gff_1_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_5877), .Z1_t (new_AGEMA_signal_5878), .Z1_f (new_AGEMA_signal_5879) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S00reg_gff_1_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_5877), .B1_t (new_AGEMA_signal_5878), .B1_f (new_AGEMA_signal_5879), .Z0_t (KeyArray_S00reg_gff_1_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_6289), .Z1_t (new_AGEMA_signal_6290), .Z1_f (new_AGEMA_signal_6291) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S00reg_gff_1_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_6289), .A1_t (new_AGEMA_signal_6290), .A1_f (new_AGEMA_signal_6291), .B0_t (KeyArray_inS00ser[4]), .B0_f (new_AGEMA_signal_5726), .B1_t (new_AGEMA_signal_5727), .B1_f (new_AGEMA_signal_5728), .Z0_t (KeyArray_S00reg_gff_1_SFF_4_QD), .Z0_f (new_AGEMA_signal_6418), .Z1_t (new_AGEMA_signal_6419), .Z1_f (new_AGEMA_signal_6420) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S00reg_gff_1_SFF_5_U3 ( .A0_t (KeyArray_S00reg_gff_1_SFF_5_n2), .A0_f (new_AGEMA_signal_7245), .A1_t (new_AGEMA_signal_7246), .A1_f (new_AGEMA_signal_7247), .B0_t (KeyArray_S00reg_gff_1_SFF_5_n1), .B0_f (new_AGEMA_signal_6421), .B1_t (new_AGEMA_signal_6422), .B1_f (new_AGEMA_signal_6423), .Z0_t (keyStateIn[5]), .Z0_f (new_AGEMA_signal_2534), .Z1_t (new_AGEMA_signal_2535), .Z1_f (new_AGEMA_signal_2536) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_5_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (keyStateIn[5]), .B0_f (new_AGEMA_signal_2534), .B1_t (new_AGEMA_signal_2535), .B1_f (new_AGEMA_signal_2536), .Z0_t (KeyArray_S00reg_gff_1_SFF_5_n1), .Z0_f (new_AGEMA_signal_6421), .Z1_t (new_AGEMA_signal_6422), .Z1_f (new_AGEMA_signal_6423) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_5_U1 ( .A0_t (KeyArray_S00reg_gff_1_SFF_5_QD), .A0_f (new_AGEMA_signal_6424), .A1_t (new_AGEMA_signal_6425), .A1_f (new_AGEMA_signal_6426), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S00reg_gff_1_SFF_5_n2), .Z0_f (new_AGEMA_signal_7245), .Z1_t (new_AGEMA_signal_7246), .Z1_f (new_AGEMA_signal_7247) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS00ser[5]), .A0_f (new_AGEMA_signal_5729), .A1_t (new_AGEMA_signal_5730), .A1_f (new_AGEMA_signal_5731), .B0_t (KeyArray_outS10ser[5]), .B0_f (new_AGEMA_signal_3442), .B1_t (new_AGEMA_signal_3443), .B1_f (new_AGEMA_signal_3444), .Z0_t (KeyArray_S00reg_gff_1_SFF_5_MUXInst_X), .Z0_f (new_AGEMA_signal_5880), .Z1_t (new_AGEMA_signal_5881), .Z1_f (new_AGEMA_signal_5882) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S00reg_gff_1_SFF_5_MUXInst_X), .B0_f (new_AGEMA_signal_5880), .B1_t (new_AGEMA_signal_5881), .B1_f (new_AGEMA_signal_5882), .Z0_t (KeyArray_S00reg_gff_1_SFF_5_MUXInst_Y), .Z0_f (new_AGEMA_signal_6292), .Z1_t (new_AGEMA_signal_6293), .Z1_f (new_AGEMA_signal_6294) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S00reg_gff_1_SFF_5_MUXInst_Y), .A0_f (new_AGEMA_signal_6292), .A1_t (new_AGEMA_signal_6293), .A1_f (new_AGEMA_signal_6294), .B0_t (KeyArray_inS00ser[5]), .B0_f (new_AGEMA_signal_5729), .B1_t (new_AGEMA_signal_5730), .B1_f (new_AGEMA_signal_5731), .Z0_t (KeyArray_S00reg_gff_1_SFF_5_QD), .Z0_f (new_AGEMA_signal_6424), .Z1_t (new_AGEMA_signal_6425), .Z1_f (new_AGEMA_signal_6426) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S00reg_gff_1_SFF_6_U3 ( .A0_t (KeyArray_S00reg_gff_1_SFF_6_n2), .A0_f (new_AGEMA_signal_7248), .A1_t (new_AGEMA_signal_7249), .A1_f (new_AGEMA_signal_7250), .B0_t (KeyArray_S00reg_gff_1_SFF_6_n1), .B0_f (new_AGEMA_signal_6427), .B1_t (new_AGEMA_signal_6428), .B1_f (new_AGEMA_signal_6429), .Z0_t (keyStateIn[6]), .Z0_f (new_AGEMA_signal_2543), .Z1_t (new_AGEMA_signal_2544), .Z1_f (new_AGEMA_signal_2545) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_6_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (keyStateIn[6]), .B0_f (new_AGEMA_signal_2543), .B1_t (new_AGEMA_signal_2544), .B1_f (new_AGEMA_signal_2545), .Z0_t (KeyArray_S00reg_gff_1_SFF_6_n1), .Z0_f (new_AGEMA_signal_6427), .Z1_t (new_AGEMA_signal_6428), .Z1_f (new_AGEMA_signal_6429) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_6_U1 ( .A0_t (KeyArray_S00reg_gff_1_SFF_6_QD), .A0_f (new_AGEMA_signal_6430), .A1_t (new_AGEMA_signal_6431), .A1_f (new_AGEMA_signal_6432), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S00reg_gff_1_SFF_6_n2), .Z0_f (new_AGEMA_signal_7248), .Z1_t (new_AGEMA_signal_7249), .Z1_f (new_AGEMA_signal_7250) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS00ser[6]), .A0_f (new_AGEMA_signal_5732), .A1_t (new_AGEMA_signal_5733), .A1_f (new_AGEMA_signal_5734), .B0_t (KeyArray_outS10ser[6]), .B0_f (new_AGEMA_signal_3451), .B1_t (new_AGEMA_signal_3452), .B1_f (new_AGEMA_signal_3453), .Z0_t (KeyArray_S00reg_gff_1_SFF_6_MUXInst_X), .Z0_f (new_AGEMA_signal_5883), .Z1_t (new_AGEMA_signal_5884), .Z1_f (new_AGEMA_signal_5885) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S00reg_gff_1_SFF_6_MUXInst_X), .B0_f (new_AGEMA_signal_5883), .B1_t (new_AGEMA_signal_5884), .B1_f (new_AGEMA_signal_5885), .Z0_t (KeyArray_S00reg_gff_1_SFF_6_MUXInst_Y), .Z0_f (new_AGEMA_signal_6295), .Z1_t (new_AGEMA_signal_6296), .Z1_f (new_AGEMA_signal_6297) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S00reg_gff_1_SFF_6_MUXInst_Y), .A0_f (new_AGEMA_signal_6295), .A1_t (new_AGEMA_signal_6296), .A1_f (new_AGEMA_signal_6297), .B0_t (KeyArray_inS00ser[6]), .B0_f (new_AGEMA_signal_5732), .B1_t (new_AGEMA_signal_5733), .B1_f (new_AGEMA_signal_5734), .Z0_t (KeyArray_S00reg_gff_1_SFF_6_QD), .Z0_f (new_AGEMA_signal_6430), .Z1_t (new_AGEMA_signal_6431), .Z1_f (new_AGEMA_signal_6432) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S00reg_gff_1_SFF_7_U3 ( .A0_t (KeyArray_S00reg_gff_1_SFF_7_n2), .A0_f (new_AGEMA_signal_7251), .A1_t (new_AGEMA_signal_7252), .A1_f (new_AGEMA_signal_7253), .B0_t (KeyArray_S00reg_gff_1_SFF_7_n1), .B0_f (new_AGEMA_signal_6433), .B1_t (new_AGEMA_signal_6434), .B1_f (new_AGEMA_signal_6435), .Z0_t (keyStateIn[7]), .Z0_f (new_AGEMA_signal_2552), .Z1_t (new_AGEMA_signal_2553), .Z1_f (new_AGEMA_signal_2554) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_7_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (keyStateIn[7]), .B0_f (new_AGEMA_signal_2552), .B1_t (new_AGEMA_signal_2553), .B1_f (new_AGEMA_signal_2554), .Z0_t (KeyArray_S00reg_gff_1_SFF_7_n1), .Z0_f (new_AGEMA_signal_6433), .Z1_t (new_AGEMA_signal_6434), .Z1_f (new_AGEMA_signal_6435) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_7_U1 ( .A0_t (KeyArray_S00reg_gff_1_SFF_7_QD), .A0_f (new_AGEMA_signal_6436), .A1_t (new_AGEMA_signal_6437), .A1_f (new_AGEMA_signal_6438), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S00reg_gff_1_SFF_7_n2), .Z0_f (new_AGEMA_signal_7251), .Z1_t (new_AGEMA_signal_7252), .Z1_f (new_AGEMA_signal_7253) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS00ser[7]), .A0_f (new_AGEMA_signal_5735), .A1_t (new_AGEMA_signal_5736), .A1_f (new_AGEMA_signal_5737), .B0_t (KeyArray_outS10ser[7]), .B0_f (new_AGEMA_signal_3460), .B1_t (new_AGEMA_signal_3461), .B1_f (new_AGEMA_signal_3462), .Z0_t (KeyArray_S00reg_gff_1_SFF_7_MUXInst_X), .Z0_f (new_AGEMA_signal_5886), .Z1_t (new_AGEMA_signal_5887), .Z1_f (new_AGEMA_signal_5888) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S00reg_gff_1_SFF_7_MUXInst_X), .B0_f (new_AGEMA_signal_5886), .B1_t (new_AGEMA_signal_5887), .B1_f (new_AGEMA_signal_5888), .Z0_t (KeyArray_S00reg_gff_1_SFF_7_MUXInst_Y), .Z0_f (new_AGEMA_signal_6298), .Z1_t (new_AGEMA_signal_6299), .Z1_f (new_AGEMA_signal_6300) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S00reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S00reg_gff_1_SFF_7_MUXInst_Y), .A0_f (new_AGEMA_signal_6298), .A1_t (new_AGEMA_signal_6299), .A1_f (new_AGEMA_signal_6300), .B0_t (KeyArray_inS00ser[7]), .B0_f (new_AGEMA_signal_5735), .B1_t (new_AGEMA_signal_5736), .B1_f (new_AGEMA_signal_5737), .Z0_t (KeyArray_S00reg_gff_1_SFF_7_QD), .Z0_f (new_AGEMA_signal_6436), .Z1_t (new_AGEMA_signal_6437), .Z1_f (new_AGEMA_signal_6438) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S01reg_gff_1_SFF_0_U3 ( .A0_t (KeyArray_S01reg_gff_1_SFF_0_n2), .A0_f (new_AGEMA_signal_6442), .A1_t (new_AGEMA_signal_6443), .A1_f (new_AGEMA_signal_6444), .B0_t (KeyArray_S01reg_gff_1_SFF_0_n1), .B0_f (new_AGEMA_signal_6439), .B1_t (new_AGEMA_signal_6440), .B1_f (new_AGEMA_signal_6441), .Z0_t (KeyArray_outS01ser_0_), .Z0_f (new_AGEMA_signal_3247), .Z1_t (new_AGEMA_signal_3248), .Z1_f (new_AGEMA_signal_3249) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_0_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS01ser_0_), .B0_f (new_AGEMA_signal_3247), .B1_t (new_AGEMA_signal_3248), .B1_f (new_AGEMA_signal_3249), .Z0_t (KeyArray_S01reg_gff_1_SFF_0_n1), .Z0_f (new_AGEMA_signal_6439), .Z1_t (new_AGEMA_signal_6440), .Z1_f (new_AGEMA_signal_6441) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_0_U1 ( .A0_t (KeyArray_S01reg_gff_1_SFF_0_QD), .A0_f (new_AGEMA_signal_4701), .A1_t (new_AGEMA_signal_4702), .A1_f (new_AGEMA_signal_4703), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S01reg_gff_1_SFF_0_n2), .Z0_f (new_AGEMA_signal_6442), .Z1_t (new_AGEMA_signal_6443), .Z1_f (new_AGEMA_signal_6444) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS02ser[0]), .A0_f (new_AGEMA_signal_3253), .A1_t (new_AGEMA_signal_3254), .A1_f (new_AGEMA_signal_3255), .B0_t (KeyArray_outS11ser[0]), .B0_f (new_AGEMA_signal_3256), .B1_t (new_AGEMA_signal_3257), .B1_f (new_AGEMA_signal_3258), .Z0_t (KeyArray_S01reg_gff_1_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_3259), .Z1_t (new_AGEMA_signal_3260), .Z1_f (new_AGEMA_signal_3261) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S01reg_gff_1_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_3259), .B1_t (new_AGEMA_signal_3260), .B1_f (new_AGEMA_signal_3261), .Z0_t (KeyArray_S01reg_gff_1_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_4211), .Z1_t (new_AGEMA_signal_4212), .Z1_f (new_AGEMA_signal_4213) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S01reg_gff_1_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_4211), .A1_t (new_AGEMA_signal_4212), .A1_f (new_AGEMA_signal_4213), .B0_t (KeyArray_outS02ser[0]), .B0_f (new_AGEMA_signal_3253), .B1_t (new_AGEMA_signal_3254), .B1_f (new_AGEMA_signal_3255), .Z0_t (KeyArray_S01reg_gff_1_SFF_0_QD), .Z0_f (new_AGEMA_signal_4701), .Z1_t (new_AGEMA_signal_4702), .Z1_f (new_AGEMA_signal_4703) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S01reg_gff_1_SFF_1_U3 ( .A0_t (KeyArray_S01reg_gff_1_SFF_1_n2), .A0_f (new_AGEMA_signal_6448), .A1_t (new_AGEMA_signal_6449), .A1_f (new_AGEMA_signal_6450), .B0_t (KeyArray_S01reg_gff_1_SFF_1_n1), .B0_f (new_AGEMA_signal_6445), .B1_t (new_AGEMA_signal_6446), .B1_f (new_AGEMA_signal_6447), .Z0_t (KeyArray_outS01ser_1_), .Z0_f (new_AGEMA_signal_3241), .Z1_t (new_AGEMA_signal_3242), .Z1_f (new_AGEMA_signal_3243) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_1_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS01ser_1_), .B0_f (new_AGEMA_signal_3241), .B1_t (new_AGEMA_signal_3242), .B1_f (new_AGEMA_signal_3243), .Z0_t (KeyArray_S01reg_gff_1_SFF_1_n1), .Z0_f (new_AGEMA_signal_6445), .Z1_t (new_AGEMA_signal_6446), .Z1_f (new_AGEMA_signal_6447) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_1_U1 ( .A0_t (KeyArray_S01reg_gff_1_SFF_1_QD), .A0_f (new_AGEMA_signal_4704), .A1_t (new_AGEMA_signal_4705), .A1_f (new_AGEMA_signal_4706), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S01reg_gff_1_SFF_1_n2), .Z0_f (new_AGEMA_signal_6448), .Z1_t (new_AGEMA_signal_6449), .Z1_f (new_AGEMA_signal_6450) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS02ser[1]), .A0_f (new_AGEMA_signal_3262), .A1_t (new_AGEMA_signal_3263), .A1_f (new_AGEMA_signal_3264), .B0_t (KeyArray_outS11ser[1]), .B0_f (new_AGEMA_signal_3265), .B1_t (new_AGEMA_signal_3266), .B1_f (new_AGEMA_signal_3267), .Z0_t (KeyArray_S01reg_gff_1_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_3268), .Z1_t (new_AGEMA_signal_3269), .Z1_f (new_AGEMA_signal_3270) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S01reg_gff_1_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_3268), .B1_t (new_AGEMA_signal_3269), .B1_f (new_AGEMA_signal_3270), .Z0_t (KeyArray_S01reg_gff_1_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_4214), .Z1_t (new_AGEMA_signal_4215), .Z1_f (new_AGEMA_signal_4216) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S01reg_gff_1_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_4214), .A1_t (new_AGEMA_signal_4215), .A1_f (new_AGEMA_signal_4216), .B0_t (KeyArray_outS02ser[1]), .B0_f (new_AGEMA_signal_3262), .B1_t (new_AGEMA_signal_3263), .B1_f (new_AGEMA_signal_3264), .Z0_t (KeyArray_S01reg_gff_1_SFF_1_QD), .Z0_f (new_AGEMA_signal_4704), .Z1_t (new_AGEMA_signal_4705), .Z1_f (new_AGEMA_signal_4706) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S01reg_gff_1_SFF_2_U3 ( .A0_t (KeyArray_S01reg_gff_1_SFF_2_n2), .A0_f (new_AGEMA_signal_6454), .A1_t (new_AGEMA_signal_6455), .A1_f (new_AGEMA_signal_6456), .B0_t (KeyArray_S01reg_gff_1_SFF_2_n1), .B0_f (new_AGEMA_signal_6451), .B1_t (new_AGEMA_signal_6452), .B1_f (new_AGEMA_signal_6453), .Z0_t (KeyArray_outS01ser_2_), .Z0_f (new_AGEMA_signal_3235), .Z1_t (new_AGEMA_signal_3236), .Z1_f (new_AGEMA_signal_3237) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_2_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS01ser_2_), .B0_f (new_AGEMA_signal_3235), .B1_t (new_AGEMA_signal_3236), .B1_f (new_AGEMA_signal_3237), .Z0_t (KeyArray_S01reg_gff_1_SFF_2_n1), .Z0_f (new_AGEMA_signal_6451), .Z1_t (new_AGEMA_signal_6452), .Z1_f (new_AGEMA_signal_6453) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_2_U1 ( .A0_t (KeyArray_S01reg_gff_1_SFF_2_QD), .A0_f (new_AGEMA_signal_4707), .A1_t (new_AGEMA_signal_4708), .A1_f (new_AGEMA_signal_4709), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S01reg_gff_1_SFF_2_n2), .Z0_f (new_AGEMA_signal_6454), .Z1_t (new_AGEMA_signal_6455), .Z1_f (new_AGEMA_signal_6456) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS02ser[2]), .A0_f (new_AGEMA_signal_3271), .A1_t (new_AGEMA_signal_3272), .A1_f (new_AGEMA_signal_3273), .B0_t (KeyArray_outS11ser[2]), .B0_f (new_AGEMA_signal_3274), .B1_t (new_AGEMA_signal_3275), .B1_f (new_AGEMA_signal_3276), .Z0_t (KeyArray_S01reg_gff_1_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_3277), .Z1_t (new_AGEMA_signal_3278), .Z1_f (new_AGEMA_signal_3279) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S01reg_gff_1_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_3277), .B1_t (new_AGEMA_signal_3278), .B1_f (new_AGEMA_signal_3279), .Z0_t (KeyArray_S01reg_gff_1_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_4217), .Z1_t (new_AGEMA_signal_4218), .Z1_f (new_AGEMA_signal_4219) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S01reg_gff_1_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_4217), .A1_t (new_AGEMA_signal_4218), .A1_f (new_AGEMA_signal_4219), .B0_t (KeyArray_outS02ser[2]), .B0_f (new_AGEMA_signal_3271), .B1_t (new_AGEMA_signal_3272), .B1_f (new_AGEMA_signal_3273), .Z0_t (KeyArray_S01reg_gff_1_SFF_2_QD), .Z0_f (new_AGEMA_signal_4707), .Z1_t (new_AGEMA_signal_4708), .Z1_f (new_AGEMA_signal_4709) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S01reg_gff_1_SFF_3_U3 ( .A0_t (KeyArray_S01reg_gff_1_SFF_3_n2), .A0_f (new_AGEMA_signal_6460), .A1_t (new_AGEMA_signal_6461), .A1_f (new_AGEMA_signal_6462), .B0_t (KeyArray_S01reg_gff_1_SFF_3_n1), .B0_f (new_AGEMA_signal_6457), .B1_t (new_AGEMA_signal_6458), .B1_f (new_AGEMA_signal_6459), .Z0_t (KeyArray_outS01ser_3_), .Z0_f (new_AGEMA_signal_3229), .Z1_t (new_AGEMA_signal_3230), .Z1_f (new_AGEMA_signal_3231) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_3_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS01ser_3_), .B0_f (new_AGEMA_signal_3229), .B1_t (new_AGEMA_signal_3230), .B1_f (new_AGEMA_signal_3231), .Z0_t (KeyArray_S01reg_gff_1_SFF_3_n1), .Z0_f (new_AGEMA_signal_6457), .Z1_t (new_AGEMA_signal_6458), .Z1_f (new_AGEMA_signal_6459) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_3_U1 ( .A0_t (KeyArray_S01reg_gff_1_SFF_3_QD), .A0_f (new_AGEMA_signal_4710), .A1_t (new_AGEMA_signal_4711), .A1_f (new_AGEMA_signal_4712), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S01reg_gff_1_SFF_3_n2), .Z0_f (new_AGEMA_signal_6460), .Z1_t (new_AGEMA_signal_6461), .Z1_f (new_AGEMA_signal_6462) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS02ser[3]), .A0_f (new_AGEMA_signal_3280), .A1_t (new_AGEMA_signal_3281), .A1_f (new_AGEMA_signal_3282), .B0_t (KeyArray_outS11ser[3]), .B0_f (new_AGEMA_signal_3283), .B1_t (new_AGEMA_signal_3284), .B1_f (new_AGEMA_signal_3285), .Z0_t (KeyArray_S01reg_gff_1_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_3286), .Z1_t (new_AGEMA_signal_3287), .Z1_f (new_AGEMA_signal_3288) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S01reg_gff_1_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_3286), .B1_t (new_AGEMA_signal_3287), .B1_f (new_AGEMA_signal_3288), .Z0_t (KeyArray_S01reg_gff_1_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_4220), .Z1_t (new_AGEMA_signal_4221), .Z1_f (new_AGEMA_signal_4222) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S01reg_gff_1_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_4220), .A1_t (new_AGEMA_signal_4221), .A1_f (new_AGEMA_signal_4222), .B0_t (KeyArray_outS02ser[3]), .B0_f (new_AGEMA_signal_3280), .B1_t (new_AGEMA_signal_3281), .B1_f (new_AGEMA_signal_3282), .Z0_t (KeyArray_S01reg_gff_1_SFF_3_QD), .Z0_f (new_AGEMA_signal_4710), .Z1_t (new_AGEMA_signal_4711), .Z1_f (new_AGEMA_signal_4712) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S01reg_gff_1_SFF_4_U3 ( .A0_t (KeyArray_S01reg_gff_1_SFF_4_n2), .A0_f (new_AGEMA_signal_6466), .A1_t (new_AGEMA_signal_6467), .A1_f (new_AGEMA_signal_6468), .B0_t (KeyArray_S01reg_gff_1_SFF_4_n1), .B0_f (new_AGEMA_signal_6463), .B1_t (new_AGEMA_signal_6464), .B1_f (new_AGEMA_signal_6465), .Z0_t (KeyArray_outS01ser_4_), .Z0_f (new_AGEMA_signal_3223), .Z1_t (new_AGEMA_signal_3224), .Z1_f (new_AGEMA_signal_3225) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_4_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS01ser_4_), .B0_f (new_AGEMA_signal_3223), .B1_t (new_AGEMA_signal_3224), .B1_f (new_AGEMA_signal_3225), .Z0_t (KeyArray_S01reg_gff_1_SFF_4_n1), .Z0_f (new_AGEMA_signal_6463), .Z1_t (new_AGEMA_signal_6464), .Z1_f (new_AGEMA_signal_6465) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_4_U1 ( .A0_t (KeyArray_S01reg_gff_1_SFF_4_QD), .A0_f (new_AGEMA_signal_4713), .A1_t (new_AGEMA_signal_4714), .A1_f (new_AGEMA_signal_4715), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S01reg_gff_1_SFF_4_n2), .Z0_f (new_AGEMA_signal_6466), .Z1_t (new_AGEMA_signal_6467), .Z1_f (new_AGEMA_signal_6468) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS02ser[4]), .A0_f (new_AGEMA_signal_3289), .A1_t (new_AGEMA_signal_3290), .A1_f (new_AGEMA_signal_3291), .B0_t (KeyArray_outS11ser[4]), .B0_f (new_AGEMA_signal_3292), .B1_t (new_AGEMA_signal_3293), .B1_f (new_AGEMA_signal_3294), .Z0_t (KeyArray_S01reg_gff_1_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_3295), .Z1_t (new_AGEMA_signal_3296), .Z1_f (new_AGEMA_signal_3297) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S01reg_gff_1_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_3295), .B1_t (new_AGEMA_signal_3296), .B1_f (new_AGEMA_signal_3297), .Z0_t (KeyArray_S01reg_gff_1_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_4223), .Z1_t (new_AGEMA_signal_4224), .Z1_f (new_AGEMA_signal_4225) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S01reg_gff_1_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_4223), .A1_t (new_AGEMA_signal_4224), .A1_f (new_AGEMA_signal_4225), .B0_t (KeyArray_outS02ser[4]), .B0_f (new_AGEMA_signal_3289), .B1_t (new_AGEMA_signal_3290), .B1_f (new_AGEMA_signal_3291), .Z0_t (KeyArray_S01reg_gff_1_SFF_4_QD), .Z0_f (new_AGEMA_signal_4713), .Z1_t (new_AGEMA_signal_4714), .Z1_f (new_AGEMA_signal_4715) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S01reg_gff_1_SFF_5_U3 ( .A0_t (KeyArray_S01reg_gff_1_SFF_5_n2), .A0_f (new_AGEMA_signal_6472), .A1_t (new_AGEMA_signal_6473), .A1_f (new_AGEMA_signal_6474), .B0_t (KeyArray_S01reg_gff_1_SFF_5_n1), .B0_f (new_AGEMA_signal_6469), .B1_t (new_AGEMA_signal_6470), .B1_f (new_AGEMA_signal_6471), .Z0_t (KeyArray_outS01ser_5_), .Z0_f (new_AGEMA_signal_3217), .Z1_t (new_AGEMA_signal_3218), .Z1_f (new_AGEMA_signal_3219) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_5_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS01ser_5_), .B0_f (new_AGEMA_signal_3217), .B1_t (new_AGEMA_signal_3218), .B1_f (new_AGEMA_signal_3219), .Z0_t (KeyArray_S01reg_gff_1_SFF_5_n1), .Z0_f (new_AGEMA_signal_6469), .Z1_t (new_AGEMA_signal_6470), .Z1_f (new_AGEMA_signal_6471) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_5_U1 ( .A0_t (KeyArray_S01reg_gff_1_SFF_5_QD), .A0_f (new_AGEMA_signal_4716), .A1_t (new_AGEMA_signal_4717), .A1_f (new_AGEMA_signal_4718), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S01reg_gff_1_SFF_5_n2), .Z0_f (new_AGEMA_signal_6472), .Z1_t (new_AGEMA_signal_6473), .Z1_f (new_AGEMA_signal_6474) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS02ser[5]), .A0_f (new_AGEMA_signal_3298), .A1_t (new_AGEMA_signal_3299), .A1_f (new_AGEMA_signal_3300), .B0_t (KeyArray_outS11ser[5]), .B0_f (new_AGEMA_signal_3301), .B1_t (new_AGEMA_signal_3302), .B1_f (new_AGEMA_signal_3303), .Z0_t (KeyArray_S01reg_gff_1_SFF_5_MUXInst_X), .Z0_f (new_AGEMA_signal_3304), .Z1_t (new_AGEMA_signal_3305), .Z1_f (new_AGEMA_signal_3306) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S01reg_gff_1_SFF_5_MUXInst_X), .B0_f (new_AGEMA_signal_3304), .B1_t (new_AGEMA_signal_3305), .B1_f (new_AGEMA_signal_3306), .Z0_t (KeyArray_S01reg_gff_1_SFF_5_MUXInst_Y), .Z0_f (new_AGEMA_signal_4226), .Z1_t (new_AGEMA_signal_4227), .Z1_f (new_AGEMA_signal_4228) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S01reg_gff_1_SFF_5_MUXInst_Y), .A0_f (new_AGEMA_signal_4226), .A1_t (new_AGEMA_signal_4227), .A1_f (new_AGEMA_signal_4228), .B0_t (KeyArray_outS02ser[5]), .B0_f (new_AGEMA_signal_3298), .B1_t (new_AGEMA_signal_3299), .B1_f (new_AGEMA_signal_3300), .Z0_t (KeyArray_S01reg_gff_1_SFF_5_QD), .Z0_f (new_AGEMA_signal_4716), .Z1_t (new_AGEMA_signal_4717), .Z1_f (new_AGEMA_signal_4718) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S01reg_gff_1_SFF_6_U3 ( .A0_t (KeyArray_S01reg_gff_1_SFF_6_n2), .A0_f (new_AGEMA_signal_6478), .A1_t (new_AGEMA_signal_6479), .A1_f (new_AGEMA_signal_6480), .B0_t (KeyArray_S01reg_gff_1_SFF_6_n1), .B0_f (new_AGEMA_signal_6475), .B1_t (new_AGEMA_signal_6476), .B1_f (new_AGEMA_signal_6477), .Z0_t (KeyArray_outS01ser_6_), .Z0_f (new_AGEMA_signal_3211), .Z1_t (new_AGEMA_signal_3212), .Z1_f (new_AGEMA_signal_3213) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_6_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS01ser_6_), .B0_f (new_AGEMA_signal_3211), .B1_t (new_AGEMA_signal_3212), .B1_f (new_AGEMA_signal_3213), .Z0_t (KeyArray_S01reg_gff_1_SFF_6_n1), .Z0_f (new_AGEMA_signal_6475), .Z1_t (new_AGEMA_signal_6476), .Z1_f (new_AGEMA_signal_6477) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_6_U1 ( .A0_t (KeyArray_S01reg_gff_1_SFF_6_QD), .A0_f (new_AGEMA_signal_4719), .A1_t (new_AGEMA_signal_4720), .A1_f (new_AGEMA_signal_4721), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S01reg_gff_1_SFF_6_n2), .Z0_f (new_AGEMA_signal_6478), .Z1_t (new_AGEMA_signal_6479), .Z1_f (new_AGEMA_signal_6480) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS02ser[6]), .A0_f (new_AGEMA_signal_3307), .A1_t (new_AGEMA_signal_3308), .A1_f (new_AGEMA_signal_3309), .B0_t (KeyArray_outS11ser[6]), .B0_f (new_AGEMA_signal_3310), .B1_t (new_AGEMA_signal_3311), .B1_f (new_AGEMA_signal_3312), .Z0_t (KeyArray_S01reg_gff_1_SFF_6_MUXInst_X), .Z0_f (new_AGEMA_signal_3313), .Z1_t (new_AGEMA_signal_3314), .Z1_f (new_AGEMA_signal_3315) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S01reg_gff_1_SFF_6_MUXInst_X), .B0_f (new_AGEMA_signal_3313), .B1_t (new_AGEMA_signal_3314), .B1_f (new_AGEMA_signal_3315), .Z0_t (KeyArray_S01reg_gff_1_SFF_6_MUXInst_Y), .Z0_f (new_AGEMA_signal_4229), .Z1_t (new_AGEMA_signal_4230), .Z1_f (new_AGEMA_signal_4231) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S01reg_gff_1_SFF_6_MUXInst_Y), .A0_f (new_AGEMA_signal_4229), .A1_t (new_AGEMA_signal_4230), .A1_f (new_AGEMA_signal_4231), .B0_t (KeyArray_outS02ser[6]), .B0_f (new_AGEMA_signal_3307), .B1_t (new_AGEMA_signal_3308), .B1_f (new_AGEMA_signal_3309), .Z0_t (KeyArray_S01reg_gff_1_SFF_6_QD), .Z0_f (new_AGEMA_signal_4719), .Z1_t (new_AGEMA_signal_4720), .Z1_f (new_AGEMA_signal_4721) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S01reg_gff_1_SFF_7_U3 ( .A0_t (KeyArray_S01reg_gff_1_SFF_7_n2), .A0_f (new_AGEMA_signal_6484), .A1_t (new_AGEMA_signal_6485), .A1_f (new_AGEMA_signal_6486), .B0_t (KeyArray_S01reg_gff_1_SFF_7_n1), .B0_f (new_AGEMA_signal_6481), .B1_t (new_AGEMA_signal_6482), .B1_f (new_AGEMA_signal_6483), .Z0_t (KeyArray_outS01ser_7_), .Z0_f (new_AGEMA_signal_3205), .Z1_t (new_AGEMA_signal_3206), .Z1_f (new_AGEMA_signal_3207) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_7_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS01ser_7_), .B0_f (new_AGEMA_signal_3205), .B1_t (new_AGEMA_signal_3206), .B1_f (new_AGEMA_signal_3207), .Z0_t (KeyArray_S01reg_gff_1_SFF_7_n1), .Z0_f (new_AGEMA_signal_6481), .Z1_t (new_AGEMA_signal_6482), .Z1_f (new_AGEMA_signal_6483) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_7_U1 ( .A0_t (KeyArray_S01reg_gff_1_SFF_7_QD), .A0_f (new_AGEMA_signal_4722), .A1_t (new_AGEMA_signal_4723), .A1_f (new_AGEMA_signal_4724), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S01reg_gff_1_SFF_7_n2), .Z0_f (new_AGEMA_signal_6484), .Z1_t (new_AGEMA_signal_6485), .Z1_f (new_AGEMA_signal_6486) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS02ser[7]), .A0_f (new_AGEMA_signal_3316), .A1_t (new_AGEMA_signal_3317), .A1_f (new_AGEMA_signal_3318), .B0_t (KeyArray_outS11ser[7]), .B0_f (new_AGEMA_signal_3319), .B1_t (new_AGEMA_signal_3320), .B1_f (new_AGEMA_signal_3321), .Z0_t (KeyArray_S01reg_gff_1_SFF_7_MUXInst_X), .Z0_f (new_AGEMA_signal_3322), .Z1_t (new_AGEMA_signal_3323), .Z1_f (new_AGEMA_signal_3324) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S01reg_gff_1_SFF_7_MUXInst_X), .B0_f (new_AGEMA_signal_3322), .B1_t (new_AGEMA_signal_3323), .B1_f (new_AGEMA_signal_3324), .Z0_t (KeyArray_S01reg_gff_1_SFF_7_MUXInst_Y), .Z0_f (new_AGEMA_signal_4232), .Z1_t (new_AGEMA_signal_4233), .Z1_f (new_AGEMA_signal_4234) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S01reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S01reg_gff_1_SFF_7_MUXInst_Y), .A0_f (new_AGEMA_signal_4232), .A1_t (new_AGEMA_signal_4233), .A1_f (new_AGEMA_signal_4234), .B0_t (KeyArray_outS02ser[7]), .B0_f (new_AGEMA_signal_3316), .B1_t (new_AGEMA_signal_3317), .B1_f (new_AGEMA_signal_3318), .Z0_t (KeyArray_S01reg_gff_1_SFF_7_QD), .Z0_f (new_AGEMA_signal_4722), .Z1_t (new_AGEMA_signal_4723), .Z1_f (new_AGEMA_signal_4724) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S02reg_gff_1_SFF_0_U3 ( .A0_t (KeyArray_S02reg_gff_1_SFF_0_n2), .A0_f (new_AGEMA_signal_6490), .A1_t (new_AGEMA_signal_6491), .A1_f (new_AGEMA_signal_6492), .B0_t (KeyArray_S02reg_gff_1_SFF_0_n1), .B0_f (new_AGEMA_signal_6487), .B1_t (new_AGEMA_signal_6488), .B1_f (new_AGEMA_signal_6489), .Z0_t (KeyArray_outS02ser[0]), .Z0_f (new_AGEMA_signal_3253), .Z1_t (new_AGEMA_signal_3254), .Z1_f (new_AGEMA_signal_3255) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_0_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS02ser[0]), .B0_f (new_AGEMA_signal_3253), .B1_t (new_AGEMA_signal_3254), .B1_f (new_AGEMA_signal_3255), .Z0_t (KeyArray_S02reg_gff_1_SFF_0_n1), .Z0_f (new_AGEMA_signal_6487), .Z1_t (new_AGEMA_signal_6488), .Z1_f (new_AGEMA_signal_6489) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_0_U1 ( .A0_t (KeyArray_S02reg_gff_1_SFF_0_QD), .A0_f (new_AGEMA_signal_4725), .A1_t (new_AGEMA_signal_4726), .A1_f (new_AGEMA_signal_4727), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S02reg_gff_1_SFF_0_n2), .Z0_f (new_AGEMA_signal_6490), .Z1_t (new_AGEMA_signal_6491), .Z1_f (new_AGEMA_signal_6492) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS03ser[0]), .A0_f (new_AGEMA_signal_3325), .A1_t (new_AGEMA_signal_3326), .A1_f (new_AGEMA_signal_3327), .B0_t (KeyArray_outS12ser[0]), .B0_f (new_AGEMA_signal_3328), .B1_t (new_AGEMA_signal_3329), .B1_f (new_AGEMA_signal_3330), .Z0_t (KeyArray_S02reg_gff_1_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_3331), .Z1_t (new_AGEMA_signal_3332), .Z1_f (new_AGEMA_signal_3333) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S02reg_gff_1_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_3331), .B1_t (new_AGEMA_signal_3332), .B1_f (new_AGEMA_signal_3333), .Z0_t (KeyArray_S02reg_gff_1_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_4235), .Z1_t (new_AGEMA_signal_4236), .Z1_f (new_AGEMA_signal_4237) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S02reg_gff_1_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_4235), .A1_t (new_AGEMA_signal_4236), .A1_f (new_AGEMA_signal_4237), .B0_t (KeyArray_outS03ser[0]), .B0_f (new_AGEMA_signal_3325), .B1_t (new_AGEMA_signal_3326), .B1_f (new_AGEMA_signal_3327), .Z0_t (KeyArray_S02reg_gff_1_SFF_0_QD), .Z0_f (new_AGEMA_signal_4725), .Z1_t (new_AGEMA_signal_4726), .Z1_f (new_AGEMA_signal_4727) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S02reg_gff_1_SFF_1_U3 ( .A0_t (KeyArray_S02reg_gff_1_SFF_1_n2), .A0_f (new_AGEMA_signal_6496), .A1_t (new_AGEMA_signal_6497), .A1_f (new_AGEMA_signal_6498), .B0_t (KeyArray_S02reg_gff_1_SFF_1_n1), .B0_f (new_AGEMA_signal_6493), .B1_t (new_AGEMA_signal_6494), .B1_f (new_AGEMA_signal_6495), .Z0_t (KeyArray_outS02ser[1]), .Z0_f (new_AGEMA_signal_3262), .Z1_t (new_AGEMA_signal_3263), .Z1_f (new_AGEMA_signal_3264) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_1_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS02ser[1]), .B0_f (new_AGEMA_signal_3262), .B1_t (new_AGEMA_signal_3263), .B1_f (new_AGEMA_signal_3264), .Z0_t (KeyArray_S02reg_gff_1_SFF_1_n1), .Z0_f (new_AGEMA_signal_6493), .Z1_t (new_AGEMA_signal_6494), .Z1_f (new_AGEMA_signal_6495) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_1_U1 ( .A0_t (KeyArray_S02reg_gff_1_SFF_1_QD), .A0_f (new_AGEMA_signal_4728), .A1_t (new_AGEMA_signal_4729), .A1_f (new_AGEMA_signal_4730), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S02reg_gff_1_SFF_1_n2), .Z0_f (new_AGEMA_signal_6496), .Z1_t (new_AGEMA_signal_6497), .Z1_f (new_AGEMA_signal_6498) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS03ser[1]), .A0_f (new_AGEMA_signal_3334), .A1_t (new_AGEMA_signal_3335), .A1_f (new_AGEMA_signal_3336), .B0_t (KeyArray_outS12ser[1]), .B0_f (new_AGEMA_signal_3337), .B1_t (new_AGEMA_signal_3338), .B1_f (new_AGEMA_signal_3339), .Z0_t (KeyArray_S02reg_gff_1_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_3340), .Z1_t (new_AGEMA_signal_3341), .Z1_f (new_AGEMA_signal_3342) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S02reg_gff_1_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_3340), .B1_t (new_AGEMA_signal_3341), .B1_f (new_AGEMA_signal_3342), .Z0_t (KeyArray_S02reg_gff_1_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_4238), .Z1_t (new_AGEMA_signal_4239), .Z1_f (new_AGEMA_signal_4240) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S02reg_gff_1_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_4238), .A1_t (new_AGEMA_signal_4239), .A1_f (new_AGEMA_signal_4240), .B0_t (KeyArray_outS03ser[1]), .B0_f (new_AGEMA_signal_3334), .B1_t (new_AGEMA_signal_3335), .B1_f (new_AGEMA_signal_3336), .Z0_t (KeyArray_S02reg_gff_1_SFF_1_QD), .Z0_f (new_AGEMA_signal_4728), .Z1_t (new_AGEMA_signal_4729), .Z1_f (new_AGEMA_signal_4730) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S02reg_gff_1_SFF_2_U3 ( .A0_t (KeyArray_S02reg_gff_1_SFF_2_n2), .A0_f (new_AGEMA_signal_6502), .A1_t (new_AGEMA_signal_6503), .A1_f (new_AGEMA_signal_6504), .B0_t (KeyArray_S02reg_gff_1_SFF_2_n1), .B0_f (new_AGEMA_signal_6499), .B1_t (new_AGEMA_signal_6500), .B1_f (new_AGEMA_signal_6501), .Z0_t (KeyArray_outS02ser[2]), .Z0_f (new_AGEMA_signal_3271), .Z1_t (new_AGEMA_signal_3272), .Z1_f (new_AGEMA_signal_3273) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_2_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS02ser[2]), .B0_f (new_AGEMA_signal_3271), .B1_t (new_AGEMA_signal_3272), .B1_f (new_AGEMA_signal_3273), .Z0_t (KeyArray_S02reg_gff_1_SFF_2_n1), .Z0_f (new_AGEMA_signal_6499), .Z1_t (new_AGEMA_signal_6500), .Z1_f (new_AGEMA_signal_6501) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_2_U1 ( .A0_t (KeyArray_S02reg_gff_1_SFF_2_QD), .A0_f (new_AGEMA_signal_4731), .A1_t (new_AGEMA_signal_4732), .A1_f (new_AGEMA_signal_4733), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S02reg_gff_1_SFF_2_n2), .Z0_f (new_AGEMA_signal_6502), .Z1_t (new_AGEMA_signal_6503), .Z1_f (new_AGEMA_signal_6504) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS03ser[2]), .A0_f (new_AGEMA_signal_3343), .A1_t (new_AGEMA_signal_3344), .A1_f (new_AGEMA_signal_3345), .B0_t (KeyArray_outS12ser[2]), .B0_f (new_AGEMA_signal_3346), .B1_t (new_AGEMA_signal_3347), .B1_f (new_AGEMA_signal_3348), .Z0_t (KeyArray_S02reg_gff_1_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_3349), .Z1_t (new_AGEMA_signal_3350), .Z1_f (new_AGEMA_signal_3351) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S02reg_gff_1_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_3349), .B1_t (new_AGEMA_signal_3350), .B1_f (new_AGEMA_signal_3351), .Z0_t (KeyArray_S02reg_gff_1_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_4241), .Z1_t (new_AGEMA_signal_4242), .Z1_f (new_AGEMA_signal_4243) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S02reg_gff_1_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_4241), .A1_t (new_AGEMA_signal_4242), .A1_f (new_AGEMA_signal_4243), .B0_t (KeyArray_outS03ser[2]), .B0_f (new_AGEMA_signal_3343), .B1_t (new_AGEMA_signal_3344), .B1_f (new_AGEMA_signal_3345), .Z0_t (KeyArray_S02reg_gff_1_SFF_2_QD), .Z0_f (new_AGEMA_signal_4731), .Z1_t (new_AGEMA_signal_4732), .Z1_f (new_AGEMA_signal_4733) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S02reg_gff_1_SFF_3_U3 ( .A0_t (KeyArray_S02reg_gff_1_SFF_3_n2), .A0_f (new_AGEMA_signal_6508), .A1_t (new_AGEMA_signal_6509), .A1_f (new_AGEMA_signal_6510), .B0_t (KeyArray_S02reg_gff_1_SFF_3_n1), .B0_f (new_AGEMA_signal_6505), .B1_t (new_AGEMA_signal_6506), .B1_f (new_AGEMA_signal_6507), .Z0_t (KeyArray_outS02ser[3]), .Z0_f (new_AGEMA_signal_3280), .Z1_t (new_AGEMA_signal_3281), .Z1_f (new_AGEMA_signal_3282) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_3_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS02ser[3]), .B0_f (new_AGEMA_signal_3280), .B1_t (new_AGEMA_signal_3281), .B1_f (new_AGEMA_signal_3282), .Z0_t (KeyArray_S02reg_gff_1_SFF_3_n1), .Z0_f (new_AGEMA_signal_6505), .Z1_t (new_AGEMA_signal_6506), .Z1_f (new_AGEMA_signal_6507) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_3_U1 ( .A0_t (KeyArray_S02reg_gff_1_SFF_3_QD), .A0_f (new_AGEMA_signal_4734), .A1_t (new_AGEMA_signal_4735), .A1_f (new_AGEMA_signal_4736), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S02reg_gff_1_SFF_3_n2), .Z0_f (new_AGEMA_signal_6508), .Z1_t (new_AGEMA_signal_6509), .Z1_f (new_AGEMA_signal_6510) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS03ser[3]), .A0_f (new_AGEMA_signal_3352), .A1_t (new_AGEMA_signal_3353), .A1_f (new_AGEMA_signal_3354), .B0_t (KeyArray_outS12ser[3]), .B0_f (new_AGEMA_signal_3355), .B1_t (new_AGEMA_signal_3356), .B1_f (new_AGEMA_signal_3357), .Z0_t (KeyArray_S02reg_gff_1_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_3358), .Z1_t (new_AGEMA_signal_3359), .Z1_f (new_AGEMA_signal_3360) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S02reg_gff_1_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_3358), .B1_t (new_AGEMA_signal_3359), .B1_f (new_AGEMA_signal_3360), .Z0_t (KeyArray_S02reg_gff_1_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_4244), .Z1_t (new_AGEMA_signal_4245), .Z1_f (new_AGEMA_signal_4246) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S02reg_gff_1_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_4244), .A1_t (new_AGEMA_signal_4245), .A1_f (new_AGEMA_signal_4246), .B0_t (KeyArray_outS03ser[3]), .B0_f (new_AGEMA_signal_3352), .B1_t (new_AGEMA_signal_3353), .B1_f (new_AGEMA_signal_3354), .Z0_t (KeyArray_S02reg_gff_1_SFF_3_QD), .Z0_f (new_AGEMA_signal_4734), .Z1_t (new_AGEMA_signal_4735), .Z1_f (new_AGEMA_signal_4736) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S02reg_gff_1_SFF_4_U3 ( .A0_t (KeyArray_S02reg_gff_1_SFF_4_n2), .A0_f (new_AGEMA_signal_6514), .A1_t (new_AGEMA_signal_6515), .A1_f (new_AGEMA_signal_6516), .B0_t (KeyArray_S02reg_gff_1_SFF_4_n1), .B0_f (new_AGEMA_signal_6511), .B1_t (new_AGEMA_signal_6512), .B1_f (new_AGEMA_signal_6513), .Z0_t (KeyArray_outS02ser[4]), .Z0_f (new_AGEMA_signal_3289), .Z1_t (new_AGEMA_signal_3290), .Z1_f (new_AGEMA_signal_3291) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_4_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS02ser[4]), .B0_f (new_AGEMA_signal_3289), .B1_t (new_AGEMA_signal_3290), .B1_f (new_AGEMA_signal_3291), .Z0_t (KeyArray_S02reg_gff_1_SFF_4_n1), .Z0_f (new_AGEMA_signal_6511), .Z1_t (new_AGEMA_signal_6512), .Z1_f (new_AGEMA_signal_6513) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_4_U1 ( .A0_t (KeyArray_S02reg_gff_1_SFF_4_QD), .A0_f (new_AGEMA_signal_4737), .A1_t (new_AGEMA_signal_4738), .A1_f (new_AGEMA_signal_4739), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S02reg_gff_1_SFF_4_n2), .Z0_f (new_AGEMA_signal_6514), .Z1_t (new_AGEMA_signal_6515), .Z1_f (new_AGEMA_signal_6516) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS03ser[4]), .A0_f (new_AGEMA_signal_3361), .A1_t (new_AGEMA_signal_3362), .A1_f (new_AGEMA_signal_3363), .B0_t (KeyArray_outS12ser[4]), .B0_f (new_AGEMA_signal_3364), .B1_t (new_AGEMA_signal_3365), .B1_f (new_AGEMA_signal_3366), .Z0_t (KeyArray_S02reg_gff_1_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_3367), .Z1_t (new_AGEMA_signal_3368), .Z1_f (new_AGEMA_signal_3369) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S02reg_gff_1_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_3367), .B1_t (new_AGEMA_signal_3368), .B1_f (new_AGEMA_signal_3369), .Z0_t (KeyArray_S02reg_gff_1_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_4247), .Z1_t (new_AGEMA_signal_4248), .Z1_f (new_AGEMA_signal_4249) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S02reg_gff_1_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_4247), .A1_t (new_AGEMA_signal_4248), .A1_f (new_AGEMA_signal_4249), .B0_t (KeyArray_outS03ser[4]), .B0_f (new_AGEMA_signal_3361), .B1_t (new_AGEMA_signal_3362), .B1_f (new_AGEMA_signal_3363), .Z0_t (KeyArray_S02reg_gff_1_SFF_4_QD), .Z0_f (new_AGEMA_signal_4737), .Z1_t (new_AGEMA_signal_4738), .Z1_f (new_AGEMA_signal_4739) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S02reg_gff_1_SFF_5_U3 ( .A0_t (KeyArray_S02reg_gff_1_SFF_5_n2), .A0_f (new_AGEMA_signal_6520), .A1_t (new_AGEMA_signal_6521), .A1_f (new_AGEMA_signal_6522), .B0_t (KeyArray_S02reg_gff_1_SFF_5_n1), .B0_f (new_AGEMA_signal_6517), .B1_t (new_AGEMA_signal_6518), .B1_f (new_AGEMA_signal_6519), .Z0_t (KeyArray_outS02ser[5]), .Z0_f (new_AGEMA_signal_3298), .Z1_t (new_AGEMA_signal_3299), .Z1_f (new_AGEMA_signal_3300) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_5_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS02ser[5]), .B0_f (new_AGEMA_signal_3298), .B1_t (new_AGEMA_signal_3299), .B1_f (new_AGEMA_signal_3300), .Z0_t (KeyArray_S02reg_gff_1_SFF_5_n1), .Z0_f (new_AGEMA_signal_6517), .Z1_t (new_AGEMA_signal_6518), .Z1_f (new_AGEMA_signal_6519) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_5_U1 ( .A0_t (KeyArray_S02reg_gff_1_SFF_5_QD), .A0_f (new_AGEMA_signal_4740), .A1_t (new_AGEMA_signal_4741), .A1_f (new_AGEMA_signal_4742), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S02reg_gff_1_SFF_5_n2), .Z0_f (new_AGEMA_signal_6520), .Z1_t (new_AGEMA_signal_6521), .Z1_f (new_AGEMA_signal_6522) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS03ser[5]), .A0_f (new_AGEMA_signal_3370), .A1_t (new_AGEMA_signal_3371), .A1_f (new_AGEMA_signal_3372), .B0_t (KeyArray_outS12ser[5]), .B0_f (new_AGEMA_signal_3373), .B1_t (new_AGEMA_signal_3374), .B1_f (new_AGEMA_signal_3375), .Z0_t (KeyArray_S02reg_gff_1_SFF_5_MUXInst_X), .Z0_f (new_AGEMA_signal_3376), .Z1_t (new_AGEMA_signal_3377), .Z1_f (new_AGEMA_signal_3378) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S02reg_gff_1_SFF_5_MUXInst_X), .B0_f (new_AGEMA_signal_3376), .B1_t (new_AGEMA_signal_3377), .B1_f (new_AGEMA_signal_3378), .Z0_t (KeyArray_S02reg_gff_1_SFF_5_MUXInst_Y), .Z0_f (new_AGEMA_signal_4250), .Z1_t (new_AGEMA_signal_4251), .Z1_f (new_AGEMA_signal_4252) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S02reg_gff_1_SFF_5_MUXInst_Y), .A0_f (new_AGEMA_signal_4250), .A1_t (new_AGEMA_signal_4251), .A1_f (new_AGEMA_signal_4252), .B0_t (KeyArray_outS03ser[5]), .B0_f (new_AGEMA_signal_3370), .B1_t (new_AGEMA_signal_3371), .B1_f (new_AGEMA_signal_3372), .Z0_t (KeyArray_S02reg_gff_1_SFF_5_QD), .Z0_f (new_AGEMA_signal_4740), .Z1_t (new_AGEMA_signal_4741), .Z1_f (new_AGEMA_signal_4742) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S02reg_gff_1_SFF_6_U3 ( .A0_t (KeyArray_S02reg_gff_1_SFF_6_n2), .A0_f (new_AGEMA_signal_6526), .A1_t (new_AGEMA_signal_6527), .A1_f (new_AGEMA_signal_6528), .B0_t (KeyArray_S02reg_gff_1_SFF_6_n1), .B0_f (new_AGEMA_signal_6523), .B1_t (new_AGEMA_signal_6524), .B1_f (new_AGEMA_signal_6525), .Z0_t (KeyArray_outS02ser[6]), .Z0_f (new_AGEMA_signal_3307), .Z1_t (new_AGEMA_signal_3308), .Z1_f (new_AGEMA_signal_3309) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_6_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS02ser[6]), .B0_f (new_AGEMA_signal_3307), .B1_t (new_AGEMA_signal_3308), .B1_f (new_AGEMA_signal_3309), .Z0_t (KeyArray_S02reg_gff_1_SFF_6_n1), .Z0_f (new_AGEMA_signal_6523), .Z1_t (new_AGEMA_signal_6524), .Z1_f (new_AGEMA_signal_6525) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_6_U1 ( .A0_t (KeyArray_S02reg_gff_1_SFF_6_QD), .A0_f (new_AGEMA_signal_4743), .A1_t (new_AGEMA_signal_4744), .A1_f (new_AGEMA_signal_4745), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S02reg_gff_1_SFF_6_n2), .Z0_f (new_AGEMA_signal_6526), .Z1_t (new_AGEMA_signal_6527), .Z1_f (new_AGEMA_signal_6528) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS03ser[6]), .A0_f (new_AGEMA_signal_3379), .A1_t (new_AGEMA_signal_3380), .A1_f (new_AGEMA_signal_3381), .B0_t (KeyArray_outS12ser[6]), .B0_f (new_AGEMA_signal_3382), .B1_t (new_AGEMA_signal_3383), .B1_f (new_AGEMA_signal_3384), .Z0_t (KeyArray_S02reg_gff_1_SFF_6_MUXInst_X), .Z0_f (new_AGEMA_signal_3385), .Z1_t (new_AGEMA_signal_3386), .Z1_f (new_AGEMA_signal_3387) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S02reg_gff_1_SFF_6_MUXInst_X), .B0_f (new_AGEMA_signal_3385), .B1_t (new_AGEMA_signal_3386), .B1_f (new_AGEMA_signal_3387), .Z0_t (KeyArray_S02reg_gff_1_SFF_6_MUXInst_Y), .Z0_f (new_AGEMA_signal_4253), .Z1_t (new_AGEMA_signal_4254), .Z1_f (new_AGEMA_signal_4255) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S02reg_gff_1_SFF_6_MUXInst_Y), .A0_f (new_AGEMA_signal_4253), .A1_t (new_AGEMA_signal_4254), .A1_f (new_AGEMA_signal_4255), .B0_t (KeyArray_outS03ser[6]), .B0_f (new_AGEMA_signal_3379), .B1_t (new_AGEMA_signal_3380), .B1_f (new_AGEMA_signal_3381), .Z0_t (KeyArray_S02reg_gff_1_SFF_6_QD), .Z0_f (new_AGEMA_signal_4743), .Z1_t (new_AGEMA_signal_4744), .Z1_f (new_AGEMA_signal_4745) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S02reg_gff_1_SFF_7_U3 ( .A0_t (KeyArray_S02reg_gff_1_SFF_7_n2), .A0_f (new_AGEMA_signal_6532), .A1_t (new_AGEMA_signal_6533), .A1_f (new_AGEMA_signal_6534), .B0_t (KeyArray_S02reg_gff_1_SFF_7_n1), .B0_f (new_AGEMA_signal_6529), .B1_t (new_AGEMA_signal_6530), .B1_f (new_AGEMA_signal_6531), .Z0_t (KeyArray_outS02ser[7]), .Z0_f (new_AGEMA_signal_3316), .Z1_t (new_AGEMA_signal_3317), .Z1_f (new_AGEMA_signal_3318) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_7_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS02ser[7]), .B0_f (new_AGEMA_signal_3316), .B1_t (new_AGEMA_signal_3317), .B1_f (new_AGEMA_signal_3318), .Z0_t (KeyArray_S02reg_gff_1_SFF_7_n1), .Z0_f (new_AGEMA_signal_6529), .Z1_t (new_AGEMA_signal_6530), .Z1_f (new_AGEMA_signal_6531) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_7_U1 ( .A0_t (KeyArray_S02reg_gff_1_SFF_7_QD), .A0_f (new_AGEMA_signal_4746), .A1_t (new_AGEMA_signal_4747), .A1_f (new_AGEMA_signal_4748), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S02reg_gff_1_SFF_7_n2), .Z0_f (new_AGEMA_signal_6532), .Z1_t (new_AGEMA_signal_6533), .Z1_f (new_AGEMA_signal_6534) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS03ser[7]), .A0_f (new_AGEMA_signal_3388), .A1_t (new_AGEMA_signal_3389), .A1_f (new_AGEMA_signal_3390), .B0_t (KeyArray_outS12ser[7]), .B0_f (new_AGEMA_signal_3391), .B1_t (new_AGEMA_signal_3392), .B1_f (new_AGEMA_signal_3393), .Z0_t (KeyArray_S02reg_gff_1_SFF_7_MUXInst_X), .Z0_f (new_AGEMA_signal_3394), .Z1_t (new_AGEMA_signal_3395), .Z1_f (new_AGEMA_signal_3396) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S02reg_gff_1_SFF_7_MUXInst_X), .B0_f (new_AGEMA_signal_3394), .B1_t (new_AGEMA_signal_3395), .B1_f (new_AGEMA_signal_3396), .Z0_t (KeyArray_S02reg_gff_1_SFF_7_MUXInst_Y), .Z0_f (new_AGEMA_signal_4256), .Z1_t (new_AGEMA_signal_4257), .Z1_f (new_AGEMA_signal_4258) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S02reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S02reg_gff_1_SFF_7_MUXInst_Y), .A0_f (new_AGEMA_signal_4256), .A1_t (new_AGEMA_signal_4257), .A1_f (new_AGEMA_signal_4258), .B0_t (KeyArray_outS03ser[7]), .B0_f (new_AGEMA_signal_3388), .B1_t (new_AGEMA_signal_3389), .B1_f (new_AGEMA_signal_3390), .Z0_t (KeyArray_S02reg_gff_1_SFF_7_QD), .Z0_f (new_AGEMA_signal_4746), .Z1_t (new_AGEMA_signal_4747), .Z1_f (new_AGEMA_signal_4748) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S03reg_gff_1_SFF_0_U3 ( .A0_t (KeyArray_S03reg_gff_1_SFF_0_n2), .A0_f (new_AGEMA_signal_6538), .A1_t (new_AGEMA_signal_6539), .A1_f (new_AGEMA_signal_6540), .B0_t (KeyArray_S03reg_gff_1_SFF_0_n1), .B0_f (new_AGEMA_signal_6535), .B1_t (new_AGEMA_signal_6536), .B1_f (new_AGEMA_signal_6537), .Z0_t (KeyArray_outS03ser[0]), .Z0_f (new_AGEMA_signal_3325), .Z1_t (new_AGEMA_signal_3326), .Z1_f (new_AGEMA_signal_3327) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_0_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS03ser[0]), .B0_f (new_AGEMA_signal_3325), .B1_t (new_AGEMA_signal_3326), .B1_f (new_AGEMA_signal_3327), .Z0_t (KeyArray_S03reg_gff_1_SFF_0_n1), .Z0_f (new_AGEMA_signal_6535), .Z1_t (new_AGEMA_signal_6536), .Z1_f (new_AGEMA_signal_6537) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_0_U1 ( .A0_t (KeyArray_S03reg_gff_1_SFF_0_QD), .A0_f (new_AGEMA_signal_4749), .A1_t (new_AGEMA_signal_4750), .A1_f (new_AGEMA_signal_4751), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S03reg_gff_1_SFF_0_n2), .Z0_f (new_AGEMA_signal_6538), .Z1_t (new_AGEMA_signal_6539), .Z1_f (new_AGEMA_signal_6540) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS10ser[0]), .A0_f (new_AGEMA_signal_3397), .A1_t (new_AGEMA_signal_3398), .A1_f (new_AGEMA_signal_3399), .B0_t (keySBIn[0]), .B0_f (new_AGEMA_signal_3400), .B1_t (new_AGEMA_signal_3401), .B1_f (new_AGEMA_signal_3402), .Z0_t (KeyArray_S03reg_gff_1_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_3403), .Z1_t (new_AGEMA_signal_3404), .Z1_f (new_AGEMA_signal_3405) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S03reg_gff_1_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_3403), .B1_t (new_AGEMA_signal_3404), .B1_f (new_AGEMA_signal_3405), .Z0_t (KeyArray_S03reg_gff_1_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_4259), .Z1_t (new_AGEMA_signal_4260), .Z1_f (new_AGEMA_signal_4261) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S03reg_gff_1_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_4259), .A1_t (new_AGEMA_signal_4260), .A1_f (new_AGEMA_signal_4261), .B0_t (KeyArray_outS10ser[0]), .B0_f (new_AGEMA_signal_3397), .B1_t (new_AGEMA_signal_3398), .B1_f (new_AGEMA_signal_3399), .Z0_t (KeyArray_S03reg_gff_1_SFF_0_QD), .Z0_f (new_AGEMA_signal_4749), .Z1_t (new_AGEMA_signal_4750), .Z1_f (new_AGEMA_signal_4751) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S03reg_gff_1_SFF_1_U3 ( .A0_t (KeyArray_S03reg_gff_1_SFF_1_n2), .A0_f (new_AGEMA_signal_6544), .A1_t (new_AGEMA_signal_6545), .A1_f (new_AGEMA_signal_6546), .B0_t (KeyArray_S03reg_gff_1_SFF_1_n1), .B0_f (new_AGEMA_signal_6541), .B1_t (new_AGEMA_signal_6542), .B1_f (new_AGEMA_signal_6543), .Z0_t (KeyArray_outS03ser[1]), .Z0_f (new_AGEMA_signal_3334), .Z1_t (new_AGEMA_signal_3335), .Z1_f (new_AGEMA_signal_3336) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_1_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS03ser[1]), .B0_f (new_AGEMA_signal_3334), .B1_t (new_AGEMA_signal_3335), .B1_f (new_AGEMA_signal_3336), .Z0_t (KeyArray_S03reg_gff_1_SFF_1_n1), .Z0_f (new_AGEMA_signal_6541), .Z1_t (new_AGEMA_signal_6542), .Z1_f (new_AGEMA_signal_6543) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_1_U1 ( .A0_t (KeyArray_S03reg_gff_1_SFF_1_QD), .A0_f (new_AGEMA_signal_4752), .A1_t (new_AGEMA_signal_4753), .A1_f (new_AGEMA_signal_4754), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S03reg_gff_1_SFF_1_n2), .Z0_f (new_AGEMA_signal_6544), .Z1_t (new_AGEMA_signal_6545), .Z1_f (new_AGEMA_signal_6546) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS10ser[1]), .A0_f (new_AGEMA_signal_3406), .A1_t (new_AGEMA_signal_3407), .A1_f (new_AGEMA_signal_3408), .B0_t (keySBIn[1]), .B0_f (new_AGEMA_signal_3409), .B1_t (new_AGEMA_signal_3410), .B1_f (new_AGEMA_signal_3411), .Z0_t (KeyArray_S03reg_gff_1_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_3412), .Z1_t (new_AGEMA_signal_3413), .Z1_f (new_AGEMA_signal_3414) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S03reg_gff_1_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_3412), .B1_t (new_AGEMA_signal_3413), .B1_f (new_AGEMA_signal_3414), .Z0_t (KeyArray_S03reg_gff_1_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_4262), .Z1_t (new_AGEMA_signal_4263), .Z1_f (new_AGEMA_signal_4264) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S03reg_gff_1_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_4262), .A1_t (new_AGEMA_signal_4263), .A1_f (new_AGEMA_signal_4264), .B0_t (KeyArray_outS10ser[1]), .B0_f (new_AGEMA_signal_3406), .B1_t (new_AGEMA_signal_3407), .B1_f (new_AGEMA_signal_3408), .Z0_t (KeyArray_S03reg_gff_1_SFF_1_QD), .Z0_f (new_AGEMA_signal_4752), .Z1_t (new_AGEMA_signal_4753), .Z1_f (new_AGEMA_signal_4754) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S03reg_gff_1_SFF_2_U3 ( .A0_t (KeyArray_S03reg_gff_1_SFF_2_n2), .A0_f (new_AGEMA_signal_6550), .A1_t (new_AGEMA_signal_6551), .A1_f (new_AGEMA_signal_6552), .B0_t (KeyArray_S03reg_gff_1_SFF_2_n1), .B0_f (new_AGEMA_signal_6547), .B1_t (new_AGEMA_signal_6548), .B1_f (new_AGEMA_signal_6549), .Z0_t (KeyArray_outS03ser[2]), .Z0_f (new_AGEMA_signal_3343), .Z1_t (new_AGEMA_signal_3344), .Z1_f (new_AGEMA_signal_3345) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_2_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS03ser[2]), .B0_f (new_AGEMA_signal_3343), .B1_t (new_AGEMA_signal_3344), .B1_f (new_AGEMA_signal_3345), .Z0_t (KeyArray_S03reg_gff_1_SFF_2_n1), .Z0_f (new_AGEMA_signal_6547), .Z1_t (new_AGEMA_signal_6548), .Z1_f (new_AGEMA_signal_6549) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_2_U1 ( .A0_t (KeyArray_S03reg_gff_1_SFF_2_QD), .A0_f (new_AGEMA_signal_4755), .A1_t (new_AGEMA_signal_4756), .A1_f (new_AGEMA_signal_4757), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S03reg_gff_1_SFF_2_n2), .Z0_f (new_AGEMA_signal_6550), .Z1_t (new_AGEMA_signal_6551), .Z1_f (new_AGEMA_signal_6552) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS10ser[2]), .A0_f (new_AGEMA_signal_3415), .A1_t (new_AGEMA_signal_3416), .A1_f (new_AGEMA_signal_3417), .B0_t (keySBIn[2]), .B0_f (new_AGEMA_signal_3418), .B1_t (new_AGEMA_signal_3419), .B1_f (new_AGEMA_signal_3420), .Z0_t (KeyArray_S03reg_gff_1_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_3421), .Z1_t (new_AGEMA_signal_3422), .Z1_f (new_AGEMA_signal_3423) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S03reg_gff_1_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_3421), .B1_t (new_AGEMA_signal_3422), .B1_f (new_AGEMA_signal_3423), .Z0_t (KeyArray_S03reg_gff_1_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_4265), .Z1_t (new_AGEMA_signal_4266), .Z1_f (new_AGEMA_signal_4267) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S03reg_gff_1_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_4265), .A1_t (new_AGEMA_signal_4266), .A1_f (new_AGEMA_signal_4267), .B0_t (KeyArray_outS10ser[2]), .B0_f (new_AGEMA_signal_3415), .B1_t (new_AGEMA_signal_3416), .B1_f (new_AGEMA_signal_3417), .Z0_t (KeyArray_S03reg_gff_1_SFF_2_QD), .Z0_f (new_AGEMA_signal_4755), .Z1_t (new_AGEMA_signal_4756), .Z1_f (new_AGEMA_signal_4757) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S03reg_gff_1_SFF_3_U3 ( .A0_t (KeyArray_S03reg_gff_1_SFF_3_n2), .A0_f (new_AGEMA_signal_6556), .A1_t (new_AGEMA_signal_6557), .A1_f (new_AGEMA_signal_6558), .B0_t (KeyArray_S03reg_gff_1_SFF_3_n1), .B0_f (new_AGEMA_signal_6553), .B1_t (new_AGEMA_signal_6554), .B1_f (new_AGEMA_signal_6555), .Z0_t (KeyArray_outS03ser[3]), .Z0_f (new_AGEMA_signal_3352), .Z1_t (new_AGEMA_signal_3353), .Z1_f (new_AGEMA_signal_3354) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_3_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS03ser[3]), .B0_f (new_AGEMA_signal_3352), .B1_t (new_AGEMA_signal_3353), .B1_f (new_AGEMA_signal_3354), .Z0_t (KeyArray_S03reg_gff_1_SFF_3_n1), .Z0_f (new_AGEMA_signal_6553), .Z1_t (new_AGEMA_signal_6554), .Z1_f (new_AGEMA_signal_6555) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_3_U1 ( .A0_t (KeyArray_S03reg_gff_1_SFF_3_QD), .A0_f (new_AGEMA_signal_4758), .A1_t (new_AGEMA_signal_4759), .A1_f (new_AGEMA_signal_4760), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S03reg_gff_1_SFF_3_n2), .Z0_f (new_AGEMA_signal_6556), .Z1_t (new_AGEMA_signal_6557), .Z1_f (new_AGEMA_signal_6558) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS10ser[3]), .A0_f (new_AGEMA_signal_3424), .A1_t (new_AGEMA_signal_3425), .A1_f (new_AGEMA_signal_3426), .B0_t (keySBIn[3]), .B0_f (new_AGEMA_signal_3427), .B1_t (new_AGEMA_signal_3428), .B1_f (new_AGEMA_signal_3429), .Z0_t (KeyArray_S03reg_gff_1_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_3430), .Z1_t (new_AGEMA_signal_3431), .Z1_f (new_AGEMA_signal_3432) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S03reg_gff_1_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_3430), .B1_t (new_AGEMA_signal_3431), .B1_f (new_AGEMA_signal_3432), .Z0_t (KeyArray_S03reg_gff_1_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_4268), .Z1_t (new_AGEMA_signal_4269), .Z1_f (new_AGEMA_signal_4270) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S03reg_gff_1_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_4268), .A1_t (new_AGEMA_signal_4269), .A1_f (new_AGEMA_signal_4270), .B0_t (KeyArray_outS10ser[3]), .B0_f (new_AGEMA_signal_3424), .B1_t (new_AGEMA_signal_3425), .B1_f (new_AGEMA_signal_3426), .Z0_t (KeyArray_S03reg_gff_1_SFF_3_QD), .Z0_f (new_AGEMA_signal_4758), .Z1_t (new_AGEMA_signal_4759), .Z1_f (new_AGEMA_signal_4760) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S03reg_gff_1_SFF_4_U3 ( .A0_t (KeyArray_S03reg_gff_1_SFF_4_n2), .A0_f (new_AGEMA_signal_6562), .A1_t (new_AGEMA_signal_6563), .A1_f (new_AGEMA_signal_6564), .B0_t (KeyArray_S03reg_gff_1_SFF_4_n1), .B0_f (new_AGEMA_signal_6559), .B1_t (new_AGEMA_signal_6560), .B1_f (new_AGEMA_signal_6561), .Z0_t (KeyArray_outS03ser[4]), .Z0_f (new_AGEMA_signal_3361), .Z1_t (new_AGEMA_signal_3362), .Z1_f (new_AGEMA_signal_3363) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_4_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS03ser[4]), .B0_f (new_AGEMA_signal_3361), .B1_t (new_AGEMA_signal_3362), .B1_f (new_AGEMA_signal_3363), .Z0_t (KeyArray_S03reg_gff_1_SFF_4_n1), .Z0_f (new_AGEMA_signal_6559), .Z1_t (new_AGEMA_signal_6560), .Z1_f (new_AGEMA_signal_6561) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_4_U1 ( .A0_t (KeyArray_S03reg_gff_1_SFF_4_QD), .A0_f (new_AGEMA_signal_4761), .A1_t (new_AGEMA_signal_4762), .A1_f (new_AGEMA_signal_4763), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S03reg_gff_1_SFF_4_n2), .Z0_f (new_AGEMA_signal_6562), .Z1_t (new_AGEMA_signal_6563), .Z1_f (new_AGEMA_signal_6564) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS10ser[4]), .A0_f (new_AGEMA_signal_3433), .A1_t (new_AGEMA_signal_3434), .A1_f (new_AGEMA_signal_3435), .B0_t (keySBIn[4]), .B0_f (new_AGEMA_signal_3436), .B1_t (new_AGEMA_signal_3437), .B1_f (new_AGEMA_signal_3438), .Z0_t (KeyArray_S03reg_gff_1_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_3439), .Z1_t (new_AGEMA_signal_3440), .Z1_f (new_AGEMA_signal_3441) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S03reg_gff_1_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_3439), .B1_t (new_AGEMA_signal_3440), .B1_f (new_AGEMA_signal_3441), .Z0_t (KeyArray_S03reg_gff_1_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_4271), .Z1_t (new_AGEMA_signal_4272), .Z1_f (new_AGEMA_signal_4273) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S03reg_gff_1_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_4271), .A1_t (new_AGEMA_signal_4272), .A1_f (new_AGEMA_signal_4273), .B0_t (KeyArray_outS10ser[4]), .B0_f (new_AGEMA_signal_3433), .B1_t (new_AGEMA_signal_3434), .B1_f (new_AGEMA_signal_3435), .Z0_t (KeyArray_S03reg_gff_1_SFF_4_QD), .Z0_f (new_AGEMA_signal_4761), .Z1_t (new_AGEMA_signal_4762), .Z1_f (new_AGEMA_signal_4763) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S03reg_gff_1_SFF_5_U3 ( .A0_t (KeyArray_S03reg_gff_1_SFF_5_n2), .A0_f (new_AGEMA_signal_6568), .A1_t (new_AGEMA_signal_6569), .A1_f (new_AGEMA_signal_6570), .B0_t (KeyArray_S03reg_gff_1_SFF_5_n1), .B0_f (new_AGEMA_signal_6565), .B1_t (new_AGEMA_signal_6566), .B1_f (new_AGEMA_signal_6567), .Z0_t (KeyArray_outS03ser[5]), .Z0_f (new_AGEMA_signal_3370), .Z1_t (new_AGEMA_signal_3371), .Z1_f (new_AGEMA_signal_3372) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_5_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS03ser[5]), .B0_f (new_AGEMA_signal_3370), .B1_t (new_AGEMA_signal_3371), .B1_f (new_AGEMA_signal_3372), .Z0_t (KeyArray_S03reg_gff_1_SFF_5_n1), .Z0_f (new_AGEMA_signal_6565), .Z1_t (new_AGEMA_signal_6566), .Z1_f (new_AGEMA_signal_6567) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_5_U1 ( .A0_t (KeyArray_S03reg_gff_1_SFF_5_QD), .A0_f (new_AGEMA_signal_4764), .A1_t (new_AGEMA_signal_4765), .A1_f (new_AGEMA_signal_4766), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S03reg_gff_1_SFF_5_n2), .Z0_f (new_AGEMA_signal_6568), .Z1_t (new_AGEMA_signal_6569), .Z1_f (new_AGEMA_signal_6570) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS10ser[5]), .A0_f (new_AGEMA_signal_3442), .A1_t (new_AGEMA_signal_3443), .A1_f (new_AGEMA_signal_3444), .B0_t (keySBIn[5]), .B0_f (new_AGEMA_signal_3445), .B1_t (new_AGEMA_signal_3446), .B1_f (new_AGEMA_signal_3447), .Z0_t (KeyArray_S03reg_gff_1_SFF_5_MUXInst_X), .Z0_f (new_AGEMA_signal_3448), .Z1_t (new_AGEMA_signal_3449), .Z1_f (new_AGEMA_signal_3450) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S03reg_gff_1_SFF_5_MUXInst_X), .B0_f (new_AGEMA_signal_3448), .B1_t (new_AGEMA_signal_3449), .B1_f (new_AGEMA_signal_3450), .Z0_t (KeyArray_S03reg_gff_1_SFF_5_MUXInst_Y), .Z0_f (new_AGEMA_signal_4274), .Z1_t (new_AGEMA_signal_4275), .Z1_f (new_AGEMA_signal_4276) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S03reg_gff_1_SFF_5_MUXInst_Y), .A0_f (new_AGEMA_signal_4274), .A1_t (new_AGEMA_signal_4275), .A1_f (new_AGEMA_signal_4276), .B0_t (KeyArray_outS10ser[5]), .B0_f (new_AGEMA_signal_3442), .B1_t (new_AGEMA_signal_3443), .B1_f (new_AGEMA_signal_3444), .Z0_t (KeyArray_S03reg_gff_1_SFF_5_QD), .Z0_f (new_AGEMA_signal_4764), .Z1_t (new_AGEMA_signal_4765), .Z1_f (new_AGEMA_signal_4766) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S03reg_gff_1_SFF_6_U3 ( .A0_t (KeyArray_S03reg_gff_1_SFF_6_n2), .A0_f (new_AGEMA_signal_6574), .A1_t (new_AGEMA_signal_6575), .A1_f (new_AGEMA_signal_6576), .B0_t (KeyArray_S03reg_gff_1_SFF_6_n1), .B0_f (new_AGEMA_signal_6571), .B1_t (new_AGEMA_signal_6572), .B1_f (new_AGEMA_signal_6573), .Z0_t (KeyArray_outS03ser[6]), .Z0_f (new_AGEMA_signal_3379), .Z1_t (new_AGEMA_signal_3380), .Z1_f (new_AGEMA_signal_3381) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_6_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS03ser[6]), .B0_f (new_AGEMA_signal_3379), .B1_t (new_AGEMA_signal_3380), .B1_f (new_AGEMA_signal_3381), .Z0_t (KeyArray_S03reg_gff_1_SFF_6_n1), .Z0_f (new_AGEMA_signal_6571), .Z1_t (new_AGEMA_signal_6572), .Z1_f (new_AGEMA_signal_6573) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_6_U1 ( .A0_t (KeyArray_S03reg_gff_1_SFF_6_QD), .A0_f (new_AGEMA_signal_4767), .A1_t (new_AGEMA_signal_4768), .A1_f (new_AGEMA_signal_4769), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S03reg_gff_1_SFF_6_n2), .Z0_f (new_AGEMA_signal_6574), .Z1_t (new_AGEMA_signal_6575), .Z1_f (new_AGEMA_signal_6576) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS10ser[6]), .A0_f (new_AGEMA_signal_3451), .A1_t (new_AGEMA_signal_3452), .A1_f (new_AGEMA_signal_3453), .B0_t (keySBIn[6]), .B0_f (new_AGEMA_signal_3454), .B1_t (new_AGEMA_signal_3455), .B1_f (new_AGEMA_signal_3456), .Z0_t (KeyArray_S03reg_gff_1_SFF_6_MUXInst_X), .Z0_f (new_AGEMA_signal_3457), .Z1_t (new_AGEMA_signal_3458), .Z1_f (new_AGEMA_signal_3459) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S03reg_gff_1_SFF_6_MUXInst_X), .B0_f (new_AGEMA_signal_3457), .B1_t (new_AGEMA_signal_3458), .B1_f (new_AGEMA_signal_3459), .Z0_t (KeyArray_S03reg_gff_1_SFF_6_MUXInst_Y), .Z0_f (new_AGEMA_signal_4277), .Z1_t (new_AGEMA_signal_4278), .Z1_f (new_AGEMA_signal_4279) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S03reg_gff_1_SFF_6_MUXInst_Y), .A0_f (new_AGEMA_signal_4277), .A1_t (new_AGEMA_signal_4278), .A1_f (new_AGEMA_signal_4279), .B0_t (KeyArray_outS10ser[6]), .B0_f (new_AGEMA_signal_3451), .B1_t (new_AGEMA_signal_3452), .B1_f (new_AGEMA_signal_3453), .Z0_t (KeyArray_S03reg_gff_1_SFF_6_QD), .Z0_f (new_AGEMA_signal_4767), .Z1_t (new_AGEMA_signal_4768), .Z1_f (new_AGEMA_signal_4769) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S03reg_gff_1_SFF_7_U3 ( .A0_t (KeyArray_S03reg_gff_1_SFF_7_n2), .A0_f (new_AGEMA_signal_6580), .A1_t (new_AGEMA_signal_6581), .A1_f (new_AGEMA_signal_6582), .B0_t (KeyArray_S03reg_gff_1_SFF_7_n1), .B0_f (new_AGEMA_signal_6577), .B1_t (new_AGEMA_signal_6578), .B1_f (new_AGEMA_signal_6579), .Z0_t (KeyArray_outS03ser[7]), .Z0_f (new_AGEMA_signal_3388), .Z1_t (new_AGEMA_signal_3389), .Z1_f (new_AGEMA_signal_3390) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_7_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS03ser[7]), .B0_f (new_AGEMA_signal_3388), .B1_t (new_AGEMA_signal_3389), .B1_f (new_AGEMA_signal_3390), .Z0_t (KeyArray_S03reg_gff_1_SFF_7_n1), .Z0_f (new_AGEMA_signal_6577), .Z1_t (new_AGEMA_signal_6578), .Z1_f (new_AGEMA_signal_6579) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_7_U1 ( .A0_t (KeyArray_S03reg_gff_1_SFF_7_QD), .A0_f (new_AGEMA_signal_4770), .A1_t (new_AGEMA_signal_4771), .A1_f (new_AGEMA_signal_4772), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S03reg_gff_1_SFF_7_n2), .Z0_f (new_AGEMA_signal_6580), .Z1_t (new_AGEMA_signal_6581), .Z1_f (new_AGEMA_signal_6582) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS10ser[7]), .A0_f (new_AGEMA_signal_3460), .A1_t (new_AGEMA_signal_3461), .A1_f (new_AGEMA_signal_3462), .B0_t (keySBIn[7]), .B0_f (new_AGEMA_signal_3463), .B1_t (new_AGEMA_signal_3464), .B1_f (new_AGEMA_signal_3465), .Z0_t (KeyArray_S03reg_gff_1_SFF_7_MUXInst_X), .Z0_f (new_AGEMA_signal_3466), .Z1_t (new_AGEMA_signal_3467), .Z1_f (new_AGEMA_signal_3468) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S03reg_gff_1_SFF_7_MUXInst_X), .B0_f (new_AGEMA_signal_3466), .B1_t (new_AGEMA_signal_3467), .B1_f (new_AGEMA_signal_3468), .Z0_t (KeyArray_S03reg_gff_1_SFF_7_MUXInst_Y), .Z0_f (new_AGEMA_signal_4280), .Z1_t (new_AGEMA_signal_4281), .Z1_f (new_AGEMA_signal_4282) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S03reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S03reg_gff_1_SFF_7_MUXInst_Y), .A0_f (new_AGEMA_signal_4280), .A1_t (new_AGEMA_signal_4281), .A1_f (new_AGEMA_signal_4282), .B0_t (KeyArray_outS10ser[7]), .B0_f (new_AGEMA_signal_3460), .B1_t (new_AGEMA_signal_3461), .B1_f (new_AGEMA_signal_3462), .Z0_t (KeyArray_S03reg_gff_1_SFF_7_QD), .Z0_f (new_AGEMA_signal_4770), .Z1_t (new_AGEMA_signal_4771), .Z1_f (new_AGEMA_signal_4772) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S10reg_gff_1_SFF_0_U3 ( .A0_t (KeyArray_S10reg_gff_1_SFF_0_n2), .A0_f (new_AGEMA_signal_6586), .A1_t (new_AGEMA_signal_6587), .A1_f (new_AGEMA_signal_6588), .B0_t (KeyArray_S10reg_gff_1_SFF_0_n1), .B0_f (new_AGEMA_signal_6583), .B1_t (new_AGEMA_signal_6584), .B1_f (new_AGEMA_signal_6585), .Z0_t (KeyArray_outS10ser[0]), .Z0_f (new_AGEMA_signal_3397), .Z1_t (new_AGEMA_signal_3398), .Z1_f (new_AGEMA_signal_3399) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_0_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS10ser[0]), .B0_f (new_AGEMA_signal_3397), .B1_t (new_AGEMA_signal_3398), .B1_f (new_AGEMA_signal_3399), .Z0_t (KeyArray_S10reg_gff_1_SFF_0_n1), .Z0_f (new_AGEMA_signal_6583), .Z1_t (new_AGEMA_signal_6584), .Z1_f (new_AGEMA_signal_6585) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_0_U1 ( .A0_t (KeyArray_S10reg_gff_1_SFF_0_QD), .A0_f (new_AGEMA_signal_4773), .A1_t (new_AGEMA_signal_4774), .A1_f (new_AGEMA_signal_4775), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S10reg_gff_1_SFF_0_n2), .Z0_f (new_AGEMA_signal_6586), .Z1_t (new_AGEMA_signal_6587), .Z1_f (new_AGEMA_signal_6588) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS11ser[0]), .A0_f (new_AGEMA_signal_3256), .A1_t (new_AGEMA_signal_3257), .A1_f (new_AGEMA_signal_3258), .B0_t (KeyArray_outS20ser[0]), .B0_f (new_AGEMA_signal_3469), .B1_t (new_AGEMA_signal_3470), .B1_f (new_AGEMA_signal_3471), .Z0_t (KeyArray_S10reg_gff_1_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_3472), .Z1_t (new_AGEMA_signal_3473), .Z1_f (new_AGEMA_signal_3474) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S10reg_gff_1_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_3472), .B1_t (new_AGEMA_signal_3473), .B1_f (new_AGEMA_signal_3474), .Z0_t (KeyArray_S10reg_gff_1_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_4283), .Z1_t (new_AGEMA_signal_4284), .Z1_f (new_AGEMA_signal_4285) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S10reg_gff_1_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_4283), .A1_t (new_AGEMA_signal_4284), .A1_f (new_AGEMA_signal_4285), .B0_t (KeyArray_outS11ser[0]), .B0_f (new_AGEMA_signal_3256), .B1_t (new_AGEMA_signal_3257), .B1_f (new_AGEMA_signal_3258), .Z0_t (KeyArray_S10reg_gff_1_SFF_0_QD), .Z0_f (new_AGEMA_signal_4773), .Z1_t (new_AGEMA_signal_4774), .Z1_f (new_AGEMA_signal_4775) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S10reg_gff_1_SFF_1_U3 ( .A0_t (KeyArray_S10reg_gff_1_SFF_1_n2), .A0_f (new_AGEMA_signal_6592), .A1_t (new_AGEMA_signal_6593), .A1_f (new_AGEMA_signal_6594), .B0_t (KeyArray_S10reg_gff_1_SFF_1_n1), .B0_f (new_AGEMA_signal_6589), .B1_t (new_AGEMA_signal_6590), .B1_f (new_AGEMA_signal_6591), .Z0_t (KeyArray_outS10ser[1]), .Z0_f (new_AGEMA_signal_3406), .Z1_t (new_AGEMA_signal_3407), .Z1_f (new_AGEMA_signal_3408) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_1_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS10ser[1]), .B0_f (new_AGEMA_signal_3406), .B1_t (new_AGEMA_signal_3407), .B1_f (new_AGEMA_signal_3408), .Z0_t (KeyArray_S10reg_gff_1_SFF_1_n1), .Z0_f (new_AGEMA_signal_6589), .Z1_t (new_AGEMA_signal_6590), .Z1_f (new_AGEMA_signal_6591) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_1_U1 ( .A0_t (KeyArray_S10reg_gff_1_SFF_1_QD), .A0_f (new_AGEMA_signal_4776), .A1_t (new_AGEMA_signal_4777), .A1_f (new_AGEMA_signal_4778), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S10reg_gff_1_SFF_1_n2), .Z0_f (new_AGEMA_signal_6592), .Z1_t (new_AGEMA_signal_6593), .Z1_f (new_AGEMA_signal_6594) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS11ser[1]), .A0_f (new_AGEMA_signal_3265), .A1_t (new_AGEMA_signal_3266), .A1_f (new_AGEMA_signal_3267), .B0_t (KeyArray_outS20ser[1]), .B0_f (new_AGEMA_signal_3475), .B1_t (new_AGEMA_signal_3476), .B1_f (new_AGEMA_signal_3477), .Z0_t (KeyArray_S10reg_gff_1_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_3478), .Z1_t (new_AGEMA_signal_3479), .Z1_f (new_AGEMA_signal_3480) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S10reg_gff_1_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_3478), .B1_t (new_AGEMA_signal_3479), .B1_f (new_AGEMA_signal_3480), .Z0_t (KeyArray_S10reg_gff_1_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_4286), .Z1_t (new_AGEMA_signal_4287), .Z1_f (new_AGEMA_signal_4288) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S10reg_gff_1_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_4286), .A1_t (new_AGEMA_signal_4287), .A1_f (new_AGEMA_signal_4288), .B0_t (KeyArray_outS11ser[1]), .B0_f (new_AGEMA_signal_3265), .B1_t (new_AGEMA_signal_3266), .B1_f (new_AGEMA_signal_3267), .Z0_t (KeyArray_S10reg_gff_1_SFF_1_QD), .Z0_f (new_AGEMA_signal_4776), .Z1_t (new_AGEMA_signal_4777), .Z1_f (new_AGEMA_signal_4778) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S10reg_gff_1_SFF_2_U3 ( .A0_t (KeyArray_S10reg_gff_1_SFF_2_n2), .A0_f (new_AGEMA_signal_6598), .A1_t (new_AGEMA_signal_6599), .A1_f (new_AGEMA_signal_6600), .B0_t (KeyArray_S10reg_gff_1_SFF_2_n1), .B0_f (new_AGEMA_signal_6595), .B1_t (new_AGEMA_signal_6596), .B1_f (new_AGEMA_signal_6597), .Z0_t (KeyArray_outS10ser[2]), .Z0_f (new_AGEMA_signal_3415), .Z1_t (new_AGEMA_signal_3416), .Z1_f (new_AGEMA_signal_3417) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_2_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS10ser[2]), .B0_f (new_AGEMA_signal_3415), .B1_t (new_AGEMA_signal_3416), .B1_f (new_AGEMA_signal_3417), .Z0_t (KeyArray_S10reg_gff_1_SFF_2_n1), .Z0_f (new_AGEMA_signal_6595), .Z1_t (new_AGEMA_signal_6596), .Z1_f (new_AGEMA_signal_6597) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_2_U1 ( .A0_t (KeyArray_S10reg_gff_1_SFF_2_QD), .A0_f (new_AGEMA_signal_4779), .A1_t (new_AGEMA_signal_4780), .A1_f (new_AGEMA_signal_4781), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S10reg_gff_1_SFF_2_n2), .Z0_f (new_AGEMA_signal_6598), .Z1_t (new_AGEMA_signal_6599), .Z1_f (new_AGEMA_signal_6600) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS11ser[2]), .A0_f (new_AGEMA_signal_3274), .A1_t (new_AGEMA_signal_3275), .A1_f (new_AGEMA_signal_3276), .B0_t (KeyArray_outS20ser[2]), .B0_f (new_AGEMA_signal_3481), .B1_t (new_AGEMA_signal_3482), .B1_f (new_AGEMA_signal_3483), .Z0_t (KeyArray_S10reg_gff_1_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_3484), .Z1_t (new_AGEMA_signal_3485), .Z1_f (new_AGEMA_signal_3486) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S10reg_gff_1_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_3484), .B1_t (new_AGEMA_signal_3485), .B1_f (new_AGEMA_signal_3486), .Z0_t (KeyArray_S10reg_gff_1_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_4289), .Z1_t (new_AGEMA_signal_4290), .Z1_f (new_AGEMA_signal_4291) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S10reg_gff_1_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_4289), .A1_t (new_AGEMA_signal_4290), .A1_f (new_AGEMA_signal_4291), .B0_t (KeyArray_outS11ser[2]), .B0_f (new_AGEMA_signal_3274), .B1_t (new_AGEMA_signal_3275), .B1_f (new_AGEMA_signal_3276), .Z0_t (KeyArray_S10reg_gff_1_SFF_2_QD), .Z0_f (new_AGEMA_signal_4779), .Z1_t (new_AGEMA_signal_4780), .Z1_f (new_AGEMA_signal_4781) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S10reg_gff_1_SFF_3_U3 ( .A0_t (KeyArray_S10reg_gff_1_SFF_3_n2), .A0_f (new_AGEMA_signal_6604), .A1_t (new_AGEMA_signal_6605), .A1_f (new_AGEMA_signal_6606), .B0_t (KeyArray_S10reg_gff_1_SFF_3_n1), .B0_f (new_AGEMA_signal_6601), .B1_t (new_AGEMA_signal_6602), .B1_f (new_AGEMA_signal_6603), .Z0_t (KeyArray_outS10ser[3]), .Z0_f (new_AGEMA_signal_3424), .Z1_t (new_AGEMA_signal_3425), .Z1_f (new_AGEMA_signal_3426) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_3_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS10ser[3]), .B0_f (new_AGEMA_signal_3424), .B1_t (new_AGEMA_signal_3425), .B1_f (new_AGEMA_signal_3426), .Z0_t (KeyArray_S10reg_gff_1_SFF_3_n1), .Z0_f (new_AGEMA_signal_6601), .Z1_t (new_AGEMA_signal_6602), .Z1_f (new_AGEMA_signal_6603) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_3_U1 ( .A0_t (KeyArray_S10reg_gff_1_SFF_3_QD), .A0_f (new_AGEMA_signal_4782), .A1_t (new_AGEMA_signal_4783), .A1_f (new_AGEMA_signal_4784), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S10reg_gff_1_SFF_3_n2), .Z0_f (new_AGEMA_signal_6604), .Z1_t (new_AGEMA_signal_6605), .Z1_f (new_AGEMA_signal_6606) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS11ser[3]), .A0_f (new_AGEMA_signal_3283), .A1_t (new_AGEMA_signal_3284), .A1_f (new_AGEMA_signal_3285), .B0_t (KeyArray_outS20ser[3]), .B0_f (new_AGEMA_signal_3487), .B1_t (new_AGEMA_signal_3488), .B1_f (new_AGEMA_signal_3489), .Z0_t (KeyArray_S10reg_gff_1_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_3490), .Z1_t (new_AGEMA_signal_3491), .Z1_f (new_AGEMA_signal_3492) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S10reg_gff_1_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_3490), .B1_t (new_AGEMA_signal_3491), .B1_f (new_AGEMA_signal_3492), .Z0_t (KeyArray_S10reg_gff_1_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_4292), .Z1_t (new_AGEMA_signal_4293), .Z1_f (new_AGEMA_signal_4294) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S10reg_gff_1_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_4292), .A1_t (new_AGEMA_signal_4293), .A1_f (new_AGEMA_signal_4294), .B0_t (KeyArray_outS11ser[3]), .B0_f (new_AGEMA_signal_3283), .B1_t (new_AGEMA_signal_3284), .B1_f (new_AGEMA_signal_3285), .Z0_t (KeyArray_S10reg_gff_1_SFF_3_QD), .Z0_f (new_AGEMA_signal_4782), .Z1_t (new_AGEMA_signal_4783), .Z1_f (new_AGEMA_signal_4784) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S10reg_gff_1_SFF_4_U3 ( .A0_t (KeyArray_S10reg_gff_1_SFF_4_n2), .A0_f (new_AGEMA_signal_6610), .A1_t (new_AGEMA_signal_6611), .A1_f (new_AGEMA_signal_6612), .B0_t (KeyArray_S10reg_gff_1_SFF_4_n1), .B0_f (new_AGEMA_signal_6607), .B1_t (new_AGEMA_signal_6608), .B1_f (new_AGEMA_signal_6609), .Z0_t (KeyArray_outS10ser[4]), .Z0_f (new_AGEMA_signal_3433), .Z1_t (new_AGEMA_signal_3434), .Z1_f (new_AGEMA_signal_3435) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_4_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS10ser[4]), .B0_f (new_AGEMA_signal_3433), .B1_t (new_AGEMA_signal_3434), .B1_f (new_AGEMA_signal_3435), .Z0_t (KeyArray_S10reg_gff_1_SFF_4_n1), .Z0_f (new_AGEMA_signal_6607), .Z1_t (new_AGEMA_signal_6608), .Z1_f (new_AGEMA_signal_6609) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_4_U1 ( .A0_t (KeyArray_S10reg_gff_1_SFF_4_QD), .A0_f (new_AGEMA_signal_4785), .A1_t (new_AGEMA_signal_4786), .A1_f (new_AGEMA_signal_4787), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S10reg_gff_1_SFF_4_n2), .Z0_f (new_AGEMA_signal_6610), .Z1_t (new_AGEMA_signal_6611), .Z1_f (new_AGEMA_signal_6612) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS11ser[4]), .A0_f (new_AGEMA_signal_3292), .A1_t (new_AGEMA_signal_3293), .A1_f (new_AGEMA_signal_3294), .B0_t (KeyArray_outS20ser[4]), .B0_f (new_AGEMA_signal_3493), .B1_t (new_AGEMA_signal_3494), .B1_f (new_AGEMA_signal_3495), .Z0_t (KeyArray_S10reg_gff_1_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_3496), .Z1_t (new_AGEMA_signal_3497), .Z1_f (new_AGEMA_signal_3498) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S10reg_gff_1_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_3496), .B1_t (new_AGEMA_signal_3497), .B1_f (new_AGEMA_signal_3498), .Z0_t (KeyArray_S10reg_gff_1_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_4295), .Z1_t (new_AGEMA_signal_4296), .Z1_f (new_AGEMA_signal_4297) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S10reg_gff_1_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_4295), .A1_t (new_AGEMA_signal_4296), .A1_f (new_AGEMA_signal_4297), .B0_t (KeyArray_outS11ser[4]), .B0_f (new_AGEMA_signal_3292), .B1_t (new_AGEMA_signal_3293), .B1_f (new_AGEMA_signal_3294), .Z0_t (KeyArray_S10reg_gff_1_SFF_4_QD), .Z0_f (new_AGEMA_signal_4785), .Z1_t (new_AGEMA_signal_4786), .Z1_f (new_AGEMA_signal_4787) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S10reg_gff_1_SFF_5_U3 ( .A0_t (KeyArray_S10reg_gff_1_SFF_5_n2), .A0_f (new_AGEMA_signal_6616), .A1_t (new_AGEMA_signal_6617), .A1_f (new_AGEMA_signal_6618), .B0_t (KeyArray_S10reg_gff_1_SFF_5_n1), .B0_f (new_AGEMA_signal_6613), .B1_t (new_AGEMA_signal_6614), .B1_f (new_AGEMA_signal_6615), .Z0_t (KeyArray_outS10ser[5]), .Z0_f (new_AGEMA_signal_3442), .Z1_t (new_AGEMA_signal_3443), .Z1_f (new_AGEMA_signal_3444) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_5_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS10ser[5]), .B0_f (new_AGEMA_signal_3442), .B1_t (new_AGEMA_signal_3443), .B1_f (new_AGEMA_signal_3444), .Z0_t (KeyArray_S10reg_gff_1_SFF_5_n1), .Z0_f (new_AGEMA_signal_6613), .Z1_t (new_AGEMA_signal_6614), .Z1_f (new_AGEMA_signal_6615) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_5_U1 ( .A0_t (KeyArray_S10reg_gff_1_SFF_5_QD), .A0_f (new_AGEMA_signal_4788), .A1_t (new_AGEMA_signal_4789), .A1_f (new_AGEMA_signal_4790), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S10reg_gff_1_SFF_5_n2), .Z0_f (new_AGEMA_signal_6616), .Z1_t (new_AGEMA_signal_6617), .Z1_f (new_AGEMA_signal_6618) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS11ser[5]), .A0_f (new_AGEMA_signal_3301), .A1_t (new_AGEMA_signal_3302), .A1_f (new_AGEMA_signal_3303), .B0_t (KeyArray_outS20ser[5]), .B0_f (new_AGEMA_signal_3499), .B1_t (new_AGEMA_signal_3500), .B1_f (new_AGEMA_signal_3501), .Z0_t (KeyArray_S10reg_gff_1_SFF_5_MUXInst_X), .Z0_f (new_AGEMA_signal_3502), .Z1_t (new_AGEMA_signal_3503), .Z1_f (new_AGEMA_signal_3504) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S10reg_gff_1_SFF_5_MUXInst_X), .B0_f (new_AGEMA_signal_3502), .B1_t (new_AGEMA_signal_3503), .B1_f (new_AGEMA_signal_3504), .Z0_t (KeyArray_S10reg_gff_1_SFF_5_MUXInst_Y), .Z0_f (new_AGEMA_signal_4298), .Z1_t (new_AGEMA_signal_4299), .Z1_f (new_AGEMA_signal_4300) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S10reg_gff_1_SFF_5_MUXInst_Y), .A0_f (new_AGEMA_signal_4298), .A1_t (new_AGEMA_signal_4299), .A1_f (new_AGEMA_signal_4300), .B0_t (KeyArray_outS11ser[5]), .B0_f (new_AGEMA_signal_3301), .B1_t (new_AGEMA_signal_3302), .B1_f (new_AGEMA_signal_3303), .Z0_t (KeyArray_S10reg_gff_1_SFF_5_QD), .Z0_f (new_AGEMA_signal_4788), .Z1_t (new_AGEMA_signal_4789), .Z1_f (new_AGEMA_signal_4790) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S10reg_gff_1_SFF_6_U3 ( .A0_t (KeyArray_S10reg_gff_1_SFF_6_n2), .A0_f (new_AGEMA_signal_6622), .A1_t (new_AGEMA_signal_6623), .A1_f (new_AGEMA_signal_6624), .B0_t (KeyArray_S10reg_gff_1_SFF_6_n1), .B0_f (new_AGEMA_signal_6619), .B1_t (new_AGEMA_signal_6620), .B1_f (new_AGEMA_signal_6621), .Z0_t (KeyArray_outS10ser[6]), .Z0_f (new_AGEMA_signal_3451), .Z1_t (new_AGEMA_signal_3452), .Z1_f (new_AGEMA_signal_3453) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_6_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS10ser[6]), .B0_f (new_AGEMA_signal_3451), .B1_t (new_AGEMA_signal_3452), .B1_f (new_AGEMA_signal_3453), .Z0_t (KeyArray_S10reg_gff_1_SFF_6_n1), .Z0_f (new_AGEMA_signal_6619), .Z1_t (new_AGEMA_signal_6620), .Z1_f (new_AGEMA_signal_6621) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_6_U1 ( .A0_t (KeyArray_S10reg_gff_1_SFF_6_QD), .A0_f (new_AGEMA_signal_4791), .A1_t (new_AGEMA_signal_4792), .A1_f (new_AGEMA_signal_4793), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S10reg_gff_1_SFF_6_n2), .Z0_f (new_AGEMA_signal_6622), .Z1_t (new_AGEMA_signal_6623), .Z1_f (new_AGEMA_signal_6624) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS11ser[6]), .A0_f (new_AGEMA_signal_3310), .A1_t (new_AGEMA_signal_3311), .A1_f (new_AGEMA_signal_3312), .B0_t (KeyArray_outS20ser[6]), .B0_f (new_AGEMA_signal_3505), .B1_t (new_AGEMA_signal_3506), .B1_f (new_AGEMA_signal_3507), .Z0_t (KeyArray_S10reg_gff_1_SFF_6_MUXInst_X), .Z0_f (new_AGEMA_signal_3508), .Z1_t (new_AGEMA_signal_3509), .Z1_f (new_AGEMA_signal_3510) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S10reg_gff_1_SFF_6_MUXInst_X), .B0_f (new_AGEMA_signal_3508), .B1_t (new_AGEMA_signal_3509), .B1_f (new_AGEMA_signal_3510), .Z0_t (KeyArray_S10reg_gff_1_SFF_6_MUXInst_Y), .Z0_f (new_AGEMA_signal_4301), .Z1_t (new_AGEMA_signal_4302), .Z1_f (new_AGEMA_signal_4303) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S10reg_gff_1_SFF_6_MUXInst_Y), .A0_f (new_AGEMA_signal_4301), .A1_t (new_AGEMA_signal_4302), .A1_f (new_AGEMA_signal_4303), .B0_t (KeyArray_outS11ser[6]), .B0_f (new_AGEMA_signal_3310), .B1_t (new_AGEMA_signal_3311), .B1_f (new_AGEMA_signal_3312), .Z0_t (KeyArray_S10reg_gff_1_SFF_6_QD), .Z0_f (new_AGEMA_signal_4791), .Z1_t (new_AGEMA_signal_4792), .Z1_f (new_AGEMA_signal_4793) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S10reg_gff_1_SFF_7_U3 ( .A0_t (KeyArray_S10reg_gff_1_SFF_7_n2), .A0_f (new_AGEMA_signal_6628), .A1_t (new_AGEMA_signal_6629), .A1_f (new_AGEMA_signal_6630), .B0_t (KeyArray_S10reg_gff_1_SFF_7_n1), .B0_f (new_AGEMA_signal_6625), .B1_t (new_AGEMA_signal_6626), .B1_f (new_AGEMA_signal_6627), .Z0_t (KeyArray_outS10ser[7]), .Z0_f (new_AGEMA_signal_3460), .Z1_t (new_AGEMA_signal_3461), .Z1_f (new_AGEMA_signal_3462) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_7_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS10ser[7]), .B0_f (new_AGEMA_signal_3460), .B1_t (new_AGEMA_signal_3461), .B1_f (new_AGEMA_signal_3462), .Z0_t (KeyArray_S10reg_gff_1_SFF_7_n1), .Z0_f (new_AGEMA_signal_6625), .Z1_t (new_AGEMA_signal_6626), .Z1_f (new_AGEMA_signal_6627) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_7_U1 ( .A0_t (KeyArray_S10reg_gff_1_SFF_7_QD), .A0_f (new_AGEMA_signal_4794), .A1_t (new_AGEMA_signal_4795), .A1_f (new_AGEMA_signal_4796), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S10reg_gff_1_SFF_7_n2), .Z0_f (new_AGEMA_signal_6628), .Z1_t (new_AGEMA_signal_6629), .Z1_f (new_AGEMA_signal_6630) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS11ser[7]), .A0_f (new_AGEMA_signal_3319), .A1_t (new_AGEMA_signal_3320), .A1_f (new_AGEMA_signal_3321), .B0_t (KeyArray_outS20ser[7]), .B0_f (new_AGEMA_signal_3511), .B1_t (new_AGEMA_signal_3512), .B1_f (new_AGEMA_signal_3513), .Z0_t (KeyArray_S10reg_gff_1_SFF_7_MUXInst_X), .Z0_f (new_AGEMA_signal_3514), .Z1_t (new_AGEMA_signal_3515), .Z1_f (new_AGEMA_signal_3516) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S10reg_gff_1_SFF_7_MUXInst_X), .B0_f (new_AGEMA_signal_3514), .B1_t (new_AGEMA_signal_3515), .B1_f (new_AGEMA_signal_3516), .Z0_t (KeyArray_S10reg_gff_1_SFF_7_MUXInst_Y), .Z0_f (new_AGEMA_signal_4304), .Z1_t (new_AGEMA_signal_4305), .Z1_f (new_AGEMA_signal_4306) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S10reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S10reg_gff_1_SFF_7_MUXInst_Y), .A0_f (new_AGEMA_signal_4304), .A1_t (new_AGEMA_signal_4305), .A1_f (new_AGEMA_signal_4306), .B0_t (KeyArray_outS11ser[7]), .B0_f (new_AGEMA_signal_3319), .B1_t (new_AGEMA_signal_3320), .B1_f (new_AGEMA_signal_3321), .Z0_t (KeyArray_S10reg_gff_1_SFF_7_QD), .Z0_f (new_AGEMA_signal_4794), .Z1_t (new_AGEMA_signal_4795), .Z1_f (new_AGEMA_signal_4796) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S11reg_gff_1_SFF_0_U3 ( .A0_t (KeyArray_S11reg_gff_1_SFF_0_n2), .A0_f (new_AGEMA_signal_6634), .A1_t (new_AGEMA_signal_6635), .A1_f (new_AGEMA_signal_6636), .B0_t (KeyArray_S11reg_gff_1_SFF_0_n1), .B0_f (new_AGEMA_signal_6631), .B1_t (new_AGEMA_signal_6632), .B1_f (new_AGEMA_signal_6633), .Z0_t (KeyArray_outS11ser[0]), .Z0_f (new_AGEMA_signal_3256), .Z1_t (new_AGEMA_signal_3257), .Z1_f (new_AGEMA_signal_3258) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_0_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS11ser[0]), .B0_f (new_AGEMA_signal_3256), .B1_t (new_AGEMA_signal_3257), .B1_f (new_AGEMA_signal_3258), .Z0_t (KeyArray_S11reg_gff_1_SFF_0_n1), .Z0_f (new_AGEMA_signal_6631), .Z1_t (new_AGEMA_signal_6632), .Z1_f (new_AGEMA_signal_6633) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_0_U1 ( .A0_t (KeyArray_S11reg_gff_1_SFF_0_QD), .A0_f (new_AGEMA_signal_4797), .A1_t (new_AGEMA_signal_4798), .A1_f (new_AGEMA_signal_4799), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S11reg_gff_1_SFF_0_n2), .Z0_f (new_AGEMA_signal_6634), .Z1_t (new_AGEMA_signal_6635), .Z1_f (new_AGEMA_signal_6636) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS12ser[0]), .A0_f (new_AGEMA_signal_3328), .A1_t (new_AGEMA_signal_3329), .A1_f (new_AGEMA_signal_3330), .B0_t (KeyArray_outS21ser[0]), .B0_f (new_AGEMA_signal_3517), .B1_t (new_AGEMA_signal_3518), .B1_f (new_AGEMA_signal_3519), .Z0_t (KeyArray_S11reg_gff_1_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_3520), .Z1_t (new_AGEMA_signal_3521), .Z1_f (new_AGEMA_signal_3522) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S11reg_gff_1_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_3520), .B1_t (new_AGEMA_signal_3521), .B1_f (new_AGEMA_signal_3522), .Z0_t (KeyArray_S11reg_gff_1_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_4307), .Z1_t (new_AGEMA_signal_4308), .Z1_f (new_AGEMA_signal_4309) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S11reg_gff_1_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_4307), .A1_t (new_AGEMA_signal_4308), .A1_f (new_AGEMA_signal_4309), .B0_t (KeyArray_outS12ser[0]), .B0_f (new_AGEMA_signal_3328), .B1_t (new_AGEMA_signal_3329), .B1_f (new_AGEMA_signal_3330), .Z0_t (KeyArray_S11reg_gff_1_SFF_0_QD), .Z0_f (new_AGEMA_signal_4797), .Z1_t (new_AGEMA_signal_4798), .Z1_f (new_AGEMA_signal_4799) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S11reg_gff_1_SFF_1_U3 ( .A0_t (KeyArray_S11reg_gff_1_SFF_1_n2), .A0_f (new_AGEMA_signal_6640), .A1_t (new_AGEMA_signal_6641), .A1_f (new_AGEMA_signal_6642), .B0_t (KeyArray_S11reg_gff_1_SFF_1_n1), .B0_f (new_AGEMA_signal_6637), .B1_t (new_AGEMA_signal_6638), .B1_f (new_AGEMA_signal_6639), .Z0_t (KeyArray_outS11ser[1]), .Z0_f (new_AGEMA_signal_3265), .Z1_t (new_AGEMA_signal_3266), .Z1_f (new_AGEMA_signal_3267) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_1_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS11ser[1]), .B0_f (new_AGEMA_signal_3265), .B1_t (new_AGEMA_signal_3266), .B1_f (new_AGEMA_signal_3267), .Z0_t (KeyArray_S11reg_gff_1_SFF_1_n1), .Z0_f (new_AGEMA_signal_6637), .Z1_t (new_AGEMA_signal_6638), .Z1_f (new_AGEMA_signal_6639) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_1_U1 ( .A0_t (KeyArray_S11reg_gff_1_SFF_1_QD), .A0_f (new_AGEMA_signal_4800), .A1_t (new_AGEMA_signal_4801), .A1_f (new_AGEMA_signal_4802), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S11reg_gff_1_SFF_1_n2), .Z0_f (new_AGEMA_signal_6640), .Z1_t (new_AGEMA_signal_6641), .Z1_f (new_AGEMA_signal_6642) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS12ser[1]), .A0_f (new_AGEMA_signal_3337), .A1_t (new_AGEMA_signal_3338), .A1_f (new_AGEMA_signal_3339), .B0_t (KeyArray_outS21ser[1]), .B0_f (new_AGEMA_signal_3523), .B1_t (new_AGEMA_signal_3524), .B1_f (new_AGEMA_signal_3525), .Z0_t (KeyArray_S11reg_gff_1_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_3526), .Z1_t (new_AGEMA_signal_3527), .Z1_f (new_AGEMA_signal_3528) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S11reg_gff_1_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_3526), .B1_t (new_AGEMA_signal_3527), .B1_f (new_AGEMA_signal_3528), .Z0_t (KeyArray_S11reg_gff_1_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_4310), .Z1_t (new_AGEMA_signal_4311), .Z1_f (new_AGEMA_signal_4312) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S11reg_gff_1_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_4310), .A1_t (new_AGEMA_signal_4311), .A1_f (new_AGEMA_signal_4312), .B0_t (KeyArray_outS12ser[1]), .B0_f (new_AGEMA_signal_3337), .B1_t (new_AGEMA_signal_3338), .B1_f (new_AGEMA_signal_3339), .Z0_t (KeyArray_S11reg_gff_1_SFF_1_QD), .Z0_f (new_AGEMA_signal_4800), .Z1_t (new_AGEMA_signal_4801), .Z1_f (new_AGEMA_signal_4802) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S11reg_gff_1_SFF_2_U3 ( .A0_t (KeyArray_S11reg_gff_1_SFF_2_n2), .A0_f (new_AGEMA_signal_6646), .A1_t (new_AGEMA_signal_6647), .A1_f (new_AGEMA_signal_6648), .B0_t (KeyArray_S11reg_gff_1_SFF_2_n1), .B0_f (new_AGEMA_signal_6643), .B1_t (new_AGEMA_signal_6644), .B1_f (new_AGEMA_signal_6645), .Z0_t (KeyArray_outS11ser[2]), .Z0_f (new_AGEMA_signal_3274), .Z1_t (new_AGEMA_signal_3275), .Z1_f (new_AGEMA_signal_3276) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_2_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS11ser[2]), .B0_f (new_AGEMA_signal_3274), .B1_t (new_AGEMA_signal_3275), .B1_f (new_AGEMA_signal_3276), .Z0_t (KeyArray_S11reg_gff_1_SFF_2_n1), .Z0_f (new_AGEMA_signal_6643), .Z1_t (new_AGEMA_signal_6644), .Z1_f (new_AGEMA_signal_6645) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_2_U1 ( .A0_t (KeyArray_S11reg_gff_1_SFF_2_QD), .A0_f (new_AGEMA_signal_4803), .A1_t (new_AGEMA_signal_4804), .A1_f (new_AGEMA_signal_4805), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S11reg_gff_1_SFF_2_n2), .Z0_f (new_AGEMA_signal_6646), .Z1_t (new_AGEMA_signal_6647), .Z1_f (new_AGEMA_signal_6648) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS12ser[2]), .A0_f (new_AGEMA_signal_3346), .A1_t (new_AGEMA_signal_3347), .A1_f (new_AGEMA_signal_3348), .B0_t (KeyArray_outS21ser[2]), .B0_f (new_AGEMA_signal_3529), .B1_t (new_AGEMA_signal_3530), .B1_f (new_AGEMA_signal_3531), .Z0_t (KeyArray_S11reg_gff_1_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_3532), .Z1_t (new_AGEMA_signal_3533), .Z1_f (new_AGEMA_signal_3534) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S11reg_gff_1_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_3532), .B1_t (new_AGEMA_signal_3533), .B1_f (new_AGEMA_signal_3534), .Z0_t (KeyArray_S11reg_gff_1_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_4313), .Z1_t (new_AGEMA_signal_4314), .Z1_f (new_AGEMA_signal_4315) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S11reg_gff_1_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_4313), .A1_t (new_AGEMA_signal_4314), .A1_f (new_AGEMA_signal_4315), .B0_t (KeyArray_outS12ser[2]), .B0_f (new_AGEMA_signal_3346), .B1_t (new_AGEMA_signal_3347), .B1_f (new_AGEMA_signal_3348), .Z0_t (KeyArray_S11reg_gff_1_SFF_2_QD), .Z0_f (new_AGEMA_signal_4803), .Z1_t (new_AGEMA_signal_4804), .Z1_f (new_AGEMA_signal_4805) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S11reg_gff_1_SFF_3_U3 ( .A0_t (KeyArray_S11reg_gff_1_SFF_3_n2), .A0_f (new_AGEMA_signal_6652), .A1_t (new_AGEMA_signal_6653), .A1_f (new_AGEMA_signal_6654), .B0_t (KeyArray_S11reg_gff_1_SFF_3_n1), .B0_f (new_AGEMA_signal_6649), .B1_t (new_AGEMA_signal_6650), .B1_f (new_AGEMA_signal_6651), .Z0_t (KeyArray_outS11ser[3]), .Z0_f (new_AGEMA_signal_3283), .Z1_t (new_AGEMA_signal_3284), .Z1_f (new_AGEMA_signal_3285) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_3_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS11ser[3]), .B0_f (new_AGEMA_signal_3283), .B1_t (new_AGEMA_signal_3284), .B1_f (new_AGEMA_signal_3285), .Z0_t (KeyArray_S11reg_gff_1_SFF_3_n1), .Z0_f (new_AGEMA_signal_6649), .Z1_t (new_AGEMA_signal_6650), .Z1_f (new_AGEMA_signal_6651) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_3_U1 ( .A0_t (KeyArray_S11reg_gff_1_SFF_3_QD), .A0_f (new_AGEMA_signal_4806), .A1_t (new_AGEMA_signal_4807), .A1_f (new_AGEMA_signal_4808), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S11reg_gff_1_SFF_3_n2), .Z0_f (new_AGEMA_signal_6652), .Z1_t (new_AGEMA_signal_6653), .Z1_f (new_AGEMA_signal_6654) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS12ser[3]), .A0_f (new_AGEMA_signal_3355), .A1_t (new_AGEMA_signal_3356), .A1_f (new_AGEMA_signal_3357), .B0_t (KeyArray_outS21ser[3]), .B0_f (new_AGEMA_signal_3535), .B1_t (new_AGEMA_signal_3536), .B1_f (new_AGEMA_signal_3537), .Z0_t (KeyArray_S11reg_gff_1_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_3538), .Z1_t (new_AGEMA_signal_3539), .Z1_f (new_AGEMA_signal_3540) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S11reg_gff_1_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_3538), .B1_t (new_AGEMA_signal_3539), .B1_f (new_AGEMA_signal_3540), .Z0_t (KeyArray_S11reg_gff_1_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_4316), .Z1_t (new_AGEMA_signal_4317), .Z1_f (new_AGEMA_signal_4318) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S11reg_gff_1_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_4316), .A1_t (new_AGEMA_signal_4317), .A1_f (new_AGEMA_signal_4318), .B0_t (KeyArray_outS12ser[3]), .B0_f (new_AGEMA_signal_3355), .B1_t (new_AGEMA_signal_3356), .B1_f (new_AGEMA_signal_3357), .Z0_t (KeyArray_S11reg_gff_1_SFF_3_QD), .Z0_f (new_AGEMA_signal_4806), .Z1_t (new_AGEMA_signal_4807), .Z1_f (new_AGEMA_signal_4808) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S11reg_gff_1_SFF_4_U3 ( .A0_t (KeyArray_S11reg_gff_1_SFF_4_n2), .A0_f (new_AGEMA_signal_6658), .A1_t (new_AGEMA_signal_6659), .A1_f (new_AGEMA_signal_6660), .B0_t (KeyArray_S11reg_gff_1_SFF_4_n1), .B0_f (new_AGEMA_signal_6655), .B1_t (new_AGEMA_signal_6656), .B1_f (new_AGEMA_signal_6657), .Z0_t (KeyArray_outS11ser[4]), .Z0_f (new_AGEMA_signal_3292), .Z1_t (new_AGEMA_signal_3293), .Z1_f (new_AGEMA_signal_3294) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_4_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS11ser[4]), .B0_f (new_AGEMA_signal_3292), .B1_t (new_AGEMA_signal_3293), .B1_f (new_AGEMA_signal_3294), .Z0_t (KeyArray_S11reg_gff_1_SFF_4_n1), .Z0_f (new_AGEMA_signal_6655), .Z1_t (new_AGEMA_signal_6656), .Z1_f (new_AGEMA_signal_6657) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_4_U1 ( .A0_t (KeyArray_S11reg_gff_1_SFF_4_QD), .A0_f (new_AGEMA_signal_4809), .A1_t (new_AGEMA_signal_4810), .A1_f (new_AGEMA_signal_4811), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S11reg_gff_1_SFF_4_n2), .Z0_f (new_AGEMA_signal_6658), .Z1_t (new_AGEMA_signal_6659), .Z1_f (new_AGEMA_signal_6660) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS12ser[4]), .A0_f (new_AGEMA_signal_3364), .A1_t (new_AGEMA_signal_3365), .A1_f (new_AGEMA_signal_3366), .B0_t (KeyArray_outS21ser[4]), .B0_f (new_AGEMA_signal_3541), .B1_t (new_AGEMA_signal_3542), .B1_f (new_AGEMA_signal_3543), .Z0_t (KeyArray_S11reg_gff_1_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_3544), .Z1_t (new_AGEMA_signal_3545), .Z1_f (new_AGEMA_signal_3546) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S11reg_gff_1_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_3544), .B1_t (new_AGEMA_signal_3545), .B1_f (new_AGEMA_signal_3546), .Z0_t (KeyArray_S11reg_gff_1_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_4319), .Z1_t (new_AGEMA_signal_4320), .Z1_f (new_AGEMA_signal_4321) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S11reg_gff_1_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_4319), .A1_t (new_AGEMA_signal_4320), .A1_f (new_AGEMA_signal_4321), .B0_t (KeyArray_outS12ser[4]), .B0_f (new_AGEMA_signal_3364), .B1_t (new_AGEMA_signal_3365), .B1_f (new_AGEMA_signal_3366), .Z0_t (KeyArray_S11reg_gff_1_SFF_4_QD), .Z0_f (new_AGEMA_signal_4809), .Z1_t (new_AGEMA_signal_4810), .Z1_f (new_AGEMA_signal_4811) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S11reg_gff_1_SFF_5_U3 ( .A0_t (KeyArray_S11reg_gff_1_SFF_5_n2), .A0_f (new_AGEMA_signal_6664), .A1_t (new_AGEMA_signal_6665), .A1_f (new_AGEMA_signal_6666), .B0_t (KeyArray_S11reg_gff_1_SFF_5_n1), .B0_f (new_AGEMA_signal_6661), .B1_t (new_AGEMA_signal_6662), .B1_f (new_AGEMA_signal_6663), .Z0_t (KeyArray_outS11ser[5]), .Z0_f (new_AGEMA_signal_3301), .Z1_t (new_AGEMA_signal_3302), .Z1_f (new_AGEMA_signal_3303) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_5_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS11ser[5]), .B0_f (new_AGEMA_signal_3301), .B1_t (new_AGEMA_signal_3302), .B1_f (new_AGEMA_signal_3303), .Z0_t (KeyArray_S11reg_gff_1_SFF_5_n1), .Z0_f (new_AGEMA_signal_6661), .Z1_t (new_AGEMA_signal_6662), .Z1_f (new_AGEMA_signal_6663) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_5_U1 ( .A0_t (KeyArray_S11reg_gff_1_SFF_5_QD), .A0_f (new_AGEMA_signal_4812), .A1_t (new_AGEMA_signal_4813), .A1_f (new_AGEMA_signal_4814), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S11reg_gff_1_SFF_5_n2), .Z0_f (new_AGEMA_signal_6664), .Z1_t (new_AGEMA_signal_6665), .Z1_f (new_AGEMA_signal_6666) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS12ser[5]), .A0_f (new_AGEMA_signal_3373), .A1_t (new_AGEMA_signal_3374), .A1_f (new_AGEMA_signal_3375), .B0_t (KeyArray_outS21ser[5]), .B0_f (new_AGEMA_signal_3547), .B1_t (new_AGEMA_signal_3548), .B1_f (new_AGEMA_signal_3549), .Z0_t (KeyArray_S11reg_gff_1_SFF_5_MUXInst_X), .Z0_f (new_AGEMA_signal_3550), .Z1_t (new_AGEMA_signal_3551), .Z1_f (new_AGEMA_signal_3552) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S11reg_gff_1_SFF_5_MUXInst_X), .B0_f (new_AGEMA_signal_3550), .B1_t (new_AGEMA_signal_3551), .B1_f (new_AGEMA_signal_3552), .Z0_t (KeyArray_S11reg_gff_1_SFF_5_MUXInst_Y), .Z0_f (new_AGEMA_signal_4322), .Z1_t (new_AGEMA_signal_4323), .Z1_f (new_AGEMA_signal_4324) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S11reg_gff_1_SFF_5_MUXInst_Y), .A0_f (new_AGEMA_signal_4322), .A1_t (new_AGEMA_signal_4323), .A1_f (new_AGEMA_signal_4324), .B0_t (KeyArray_outS12ser[5]), .B0_f (new_AGEMA_signal_3373), .B1_t (new_AGEMA_signal_3374), .B1_f (new_AGEMA_signal_3375), .Z0_t (KeyArray_S11reg_gff_1_SFF_5_QD), .Z0_f (new_AGEMA_signal_4812), .Z1_t (new_AGEMA_signal_4813), .Z1_f (new_AGEMA_signal_4814) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S11reg_gff_1_SFF_6_U3 ( .A0_t (KeyArray_S11reg_gff_1_SFF_6_n2), .A0_f (new_AGEMA_signal_6670), .A1_t (new_AGEMA_signal_6671), .A1_f (new_AGEMA_signal_6672), .B0_t (KeyArray_S11reg_gff_1_SFF_6_n1), .B0_f (new_AGEMA_signal_6667), .B1_t (new_AGEMA_signal_6668), .B1_f (new_AGEMA_signal_6669), .Z0_t (KeyArray_outS11ser[6]), .Z0_f (new_AGEMA_signal_3310), .Z1_t (new_AGEMA_signal_3311), .Z1_f (new_AGEMA_signal_3312) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_6_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS11ser[6]), .B0_f (new_AGEMA_signal_3310), .B1_t (new_AGEMA_signal_3311), .B1_f (new_AGEMA_signal_3312), .Z0_t (KeyArray_S11reg_gff_1_SFF_6_n1), .Z0_f (new_AGEMA_signal_6667), .Z1_t (new_AGEMA_signal_6668), .Z1_f (new_AGEMA_signal_6669) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_6_U1 ( .A0_t (KeyArray_S11reg_gff_1_SFF_6_QD), .A0_f (new_AGEMA_signal_4815), .A1_t (new_AGEMA_signal_4816), .A1_f (new_AGEMA_signal_4817), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S11reg_gff_1_SFF_6_n2), .Z0_f (new_AGEMA_signal_6670), .Z1_t (new_AGEMA_signal_6671), .Z1_f (new_AGEMA_signal_6672) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS12ser[6]), .A0_f (new_AGEMA_signal_3382), .A1_t (new_AGEMA_signal_3383), .A1_f (new_AGEMA_signal_3384), .B0_t (KeyArray_outS21ser[6]), .B0_f (new_AGEMA_signal_3553), .B1_t (new_AGEMA_signal_3554), .B1_f (new_AGEMA_signal_3555), .Z0_t (KeyArray_S11reg_gff_1_SFF_6_MUXInst_X), .Z0_f (new_AGEMA_signal_3556), .Z1_t (new_AGEMA_signal_3557), .Z1_f (new_AGEMA_signal_3558) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S11reg_gff_1_SFF_6_MUXInst_X), .B0_f (new_AGEMA_signal_3556), .B1_t (new_AGEMA_signal_3557), .B1_f (new_AGEMA_signal_3558), .Z0_t (KeyArray_S11reg_gff_1_SFF_6_MUXInst_Y), .Z0_f (new_AGEMA_signal_4325), .Z1_t (new_AGEMA_signal_4326), .Z1_f (new_AGEMA_signal_4327) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S11reg_gff_1_SFF_6_MUXInst_Y), .A0_f (new_AGEMA_signal_4325), .A1_t (new_AGEMA_signal_4326), .A1_f (new_AGEMA_signal_4327), .B0_t (KeyArray_outS12ser[6]), .B0_f (new_AGEMA_signal_3382), .B1_t (new_AGEMA_signal_3383), .B1_f (new_AGEMA_signal_3384), .Z0_t (KeyArray_S11reg_gff_1_SFF_6_QD), .Z0_f (new_AGEMA_signal_4815), .Z1_t (new_AGEMA_signal_4816), .Z1_f (new_AGEMA_signal_4817) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S11reg_gff_1_SFF_7_U3 ( .A0_t (KeyArray_S11reg_gff_1_SFF_7_n2), .A0_f (new_AGEMA_signal_6676), .A1_t (new_AGEMA_signal_6677), .A1_f (new_AGEMA_signal_6678), .B0_t (KeyArray_S11reg_gff_1_SFF_7_n1), .B0_f (new_AGEMA_signal_6673), .B1_t (new_AGEMA_signal_6674), .B1_f (new_AGEMA_signal_6675), .Z0_t (KeyArray_outS11ser[7]), .Z0_f (new_AGEMA_signal_3319), .Z1_t (new_AGEMA_signal_3320), .Z1_f (new_AGEMA_signal_3321) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_7_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS11ser[7]), .B0_f (new_AGEMA_signal_3319), .B1_t (new_AGEMA_signal_3320), .B1_f (new_AGEMA_signal_3321), .Z0_t (KeyArray_S11reg_gff_1_SFF_7_n1), .Z0_f (new_AGEMA_signal_6673), .Z1_t (new_AGEMA_signal_6674), .Z1_f (new_AGEMA_signal_6675) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_7_U1 ( .A0_t (KeyArray_S11reg_gff_1_SFF_7_QD), .A0_f (new_AGEMA_signal_4818), .A1_t (new_AGEMA_signal_4819), .A1_f (new_AGEMA_signal_4820), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S11reg_gff_1_SFF_7_n2), .Z0_f (new_AGEMA_signal_6676), .Z1_t (new_AGEMA_signal_6677), .Z1_f (new_AGEMA_signal_6678) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS12ser[7]), .A0_f (new_AGEMA_signal_3391), .A1_t (new_AGEMA_signal_3392), .A1_f (new_AGEMA_signal_3393), .B0_t (KeyArray_outS21ser[7]), .B0_f (new_AGEMA_signal_3559), .B1_t (new_AGEMA_signal_3560), .B1_f (new_AGEMA_signal_3561), .Z0_t (KeyArray_S11reg_gff_1_SFF_7_MUXInst_X), .Z0_f (new_AGEMA_signal_3562), .Z1_t (new_AGEMA_signal_3563), .Z1_f (new_AGEMA_signal_3564) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S11reg_gff_1_SFF_7_MUXInst_X), .B0_f (new_AGEMA_signal_3562), .B1_t (new_AGEMA_signal_3563), .B1_f (new_AGEMA_signal_3564), .Z0_t (KeyArray_S11reg_gff_1_SFF_7_MUXInst_Y), .Z0_f (new_AGEMA_signal_4328), .Z1_t (new_AGEMA_signal_4329), .Z1_f (new_AGEMA_signal_4330) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S11reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S11reg_gff_1_SFF_7_MUXInst_Y), .A0_f (new_AGEMA_signal_4328), .A1_t (new_AGEMA_signal_4329), .A1_f (new_AGEMA_signal_4330), .B0_t (KeyArray_outS12ser[7]), .B0_f (new_AGEMA_signal_3391), .B1_t (new_AGEMA_signal_3392), .B1_f (new_AGEMA_signal_3393), .Z0_t (KeyArray_S11reg_gff_1_SFF_7_QD), .Z0_f (new_AGEMA_signal_4818), .Z1_t (new_AGEMA_signal_4819), .Z1_f (new_AGEMA_signal_4820) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S12reg_gff_1_SFF_0_U3 ( .A0_t (KeyArray_S12reg_gff_1_SFF_0_n2), .A0_f (new_AGEMA_signal_6682), .A1_t (new_AGEMA_signal_6683), .A1_f (new_AGEMA_signal_6684), .B0_t (KeyArray_S12reg_gff_1_SFF_0_n1), .B0_f (new_AGEMA_signal_6679), .B1_t (new_AGEMA_signal_6680), .B1_f (new_AGEMA_signal_6681), .Z0_t (KeyArray_outS12ser[0]), .Z0_f (new_AGEMA_signal_3328), .Z1_t (new_AGEMA_signal_3329), .Z1_f (new_AGEMA_signal_3330) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_0_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS12ser[0]), .B0_f (new_AGEMA_signal_3328), .B1_t (new_AGEMA_signal_3329), .B1_f (new_AGEMA_signal_3330), .Z0_t (KeyArray_S12reg_gff_1_SFF_0_n1), .Z0_f (new_AGEMA_signal_6679), .Z1_t (new_AGEMA_signal_6680), .Z1_f (new_AGEMA_signal_6681) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_0_U1 ( .A0_t (KeyArray_S12reg_gff_1_SFF_0_QD), .A0_f (new_AGEMA_signal_4821), .A1_t (new_AGEMA_signal_4822), .A1_f (new_AGEMA_signal_4823), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S12reg_gff_1_SFF_0_n2), .Z0_f (new_AGEMA_signal_6682), .Z1_t (new_AGEMA_signal_6683), .Z1_f (new_AGEMA_signal_6684) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (keySBIn[0]), .A0_f (new_AGEMA_signal_3400), .A1_t (new_AGEMA_signal_3401), .A1_f (new_AGEMA_signal_3402), .B0_t (KeyArray_outS22ser[0]), .B0_f (new_AGEMA_signal_3565), .B1_t (new_AGEMA_signal_3566), .B1_f (new_AGEMA_signal_3567), .Z0_t (KeyArray_S12reg_gff_1_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_3568), .Z1_t (new_AGEMA_signal_3569), .Z1_f (new_AGEMA_signal_3570) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S12reg_gff_1_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_3568), .B1_t (new_AGEMA_signal_3569), .B1_f (new_AGEMA_signal_3570), .Z0_t (KeyArray_S12reg_gff_1_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_4331), .Z1_t (new_AGEMA_signal_4332), .Z1_f (new_AGEMA_signal_4333) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S12reg_gff_1_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_4331), .A1_t (new_AGEMA_signal_4332), .A1_f (new_AGEMA_signal_4333), .B0_t (keySBIn[0]), .B0_f (new_AGEMA_signal_3400), .B1_t (new_AGEMA_signal_3401), .B1_f (new_AGEMA_signal_3402), .Z0_t (KeyArray_S12reg_gff_1_SFF_0_QD), .Z0_f (new_AGEMA_signal_4821), .Z1_t (new_AGEMA_signal_4822), .Z1_f (new_AGEMA_signal_4823) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S12reg_gff_1_SFF_1_U3 ( .A0_t (KeyArray_S12reg_gff_1_SFF_1_n2), .A0_f (new_AGEMA_signal_6688), .A1_t (new_AGEMA_signal_6689), .A1_f (new_AGEMA_signal_6690), .B0_t (KeyArray_S12reg_gff_1_SFF_1_n1), .B0_f (new_AGEMA_signal_6685), .B1_t (new_AGEMA_signal_6686), .B1_f (new_AGEMA_signal_6687), .Z0_t (KeyArray_outS12ser[1]), .Z0_f (new_AGEMA_signal_3337), .Z1_t (new_AGEMA_signal_3338), .Z1_f (new_AGEMA_signal_3339) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_1_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS12ser[1]), .B0_f (new_AGEMA_signal_3337), .B1_t (new_AGEMA_signal_3338), .B1_f (new_AGEMA_signal_3339), .Z0_t (KeyArray_S12reg_gff_1_SFF_1_n1), .Z0_f (new_AGEMA_signal_6685), .Z1_t (new_AGEMA_signal_6686), .Z1_f (new_AGEMA_signal_6687) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_1_U1 ( .A0_t (KeyArray_S12reg_gff_1_SFF_1_QD), .A0_f (new_AGEMA_signal_4824), .A1_t (new_AGEMA_signal_4825), .A1_f (new_AGEMA_signal_4826), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S12reg_gff_1_SFF_1_n2), .Z0_f (new_AGEMA_signal_6688), .Z1_t (new_AGEMA_signal_6689), .Z1_f (new_AGEMA_signal_6690) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (keySBIn[1]), .A0_f (new_AGEMA_signal_3409), .A1_t (new_AGEMA_signal_3410), .A1_f (new_AGEMA_signal_3411), .B0_t (KeyArray_outS22ser[1]), .B0_f (new_AGEMA_signal_3571), .B1_t (new_AGEMA_signal_3572), .B1_f (new_AGEMA_signal_3573), .Z0_t (KeyArray_S12reg_gff_1_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_3574), .Z1_t (new_AGEMA_signal_3575), .Z1_f (new_AGEMA_signal_3576) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S12reg_gff_1_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_3574), .B1_t (new_AGEMA_signal_3575), .B1_f (new_AGEMA_signal_3576), .Z0_t (KeyArray_S12reg_gff_1_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_4334), .Z1_t (new_AGEMA_signal_4335), .Z1_f (new_AGEMA_signal_4336) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S12reg_gff_1_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_4334), .A1_t (new_AGEMA_signal_4335), .A1_f (new_AGEMA_signal_4336), .B0_t (keySBIn[1]), .B0_f (new_AGEMA_signal_3409), .B1_t (new_AGEMA_signal_3410), .B1_f (new_AGEMA_signal_3411), .Z0_t (KeyArray_S12reg_gff_1_SFF_1_QD), .Z0_f (new_AGEMA_signal_4824), .Z1_t (new_AGEMA_signal_4825), .Z1_f (new_AGEMA_signal_4826) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S12reg_gff_1_SFF_2_U3 ( .A0_t (KeyArray_S12reg_gff_1_SFF_2_n2), .A0_f (new_AGEMA_signal_6694), .A1_t (new_AGEMA_signal_6695), .A1_f (new_AGEMA_signal_6696), .B0_t (KeyArray_S12reg_gff_1_SFF_2_n1), .B0_f (new_AGEMA_signal_6691), .B1_t (new_AGEMA_signal_6692), .B1_f (new_AGEMA_signal_6693), .Z0_t (KeyArray_outS12ser[2]), .Z0_f (new_AGEMA_signal_3346), .Z1_t (new_AGEMA_signal_3347), .Z1_f (new_AGEMA_signal_3348) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_2_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS12ser[2]), .B0_f (new_AGEMA_signal_3346), .B1_t (new_AGEMA_signal_3347), .B1_f (new_AGEMA_signal_3348), .Z0_t (KeyArray_S12reg_gff_1_SFF_2_n1), .Z0_f (new_AGEMA_signal_6691), .Z1_t (new_AGEMA_signal_6692), .Z1_f (new_AGEMA_signal_6693) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_2_U1 ( .A0_t (KeyArray_S12reg_gff_1_SFF_2_QD), .A0_f (new_AGEMA_signal_4827), .A1_t (new_AGEMA_signal_4828), .A1_f (new_AGEMA_signal_4829), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S12reg_gff_1_SFF_2_n2), .Z0_f (new_AGEMA_signal_6694), .Z1_t (new_AGEMA_signal_6695), .Z1_f (new_AGEMA_signal_6696) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (keySBIn[2]), .A0_f (new_AGEMA_signal_3418), .A1_t (new_AGEMA_signal_3419), .A1_f (new_AGEMA_signal_3420), .B0_t (KeyArray_outS22ser[2]), .B0_f (new_AGEMA_signal_3577), .B1_t (new_AGEMA_signal_3578), .B1_f (new_AGEMA_signal_3579), .Z0_t (KeyArray_S12reg_gff_1_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_3580), .Z1_t (new_AGEMA_signal_3581), .Z1_f (new_AGEMA_signal_3582) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S12reg_gff_1_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_3580), .B1_t (new_AGEMA_signal_3581), .B1_f (new_AGEMA_signal_3582), .Z0_t (KeyArray_S12reg_gff_1_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_4337), .Z1_t (new_AGEMA_signal_4338), .Z1_f (new_AGEMA_signal_4339) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S12reg_gff_1_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_4337), .A1_t (new_AGEMA_signal_4338), .A1_f (new_AGEMA_signal_4339), .B0_t (keySBIn[2]), .B0_f (new_AGEMA_signal_3418), .B1_t (new_AGEMA_signal_3419), .B1_f (new_AGEMA_signal_3420), .Z0_t (KeyArray_S12reg_gff_1_SFF_2_QD), .Z0_f (new_AGEMA_signal_4827), .Z1_t (new_AGEMA_signal_4828), .Z1_f (new_AGEMA_signal_4829) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S12reg_gff_1_SFF_3_U3 ( .A0_t (KeyArray_S12reg_gff_1_SFF_3_n2), .A0_f (new_AGEMA_signal_6700), .A1_t (new_AGEMA_signal_6701), .A1_f (new_AGEMA_signal_6702), .B0_t (KeyArray_S12reg_gff_1_SFF_3_n1), .B0_f (new_AGEMA_signal_6697), .B1_t (new_AGEMA_signal_6698), .B1_f (new_AGEMA_signal_6699), .Z0_t (KeyArray_outS12ser[3]), .Z0_f (new_AGEMA_signal_3355), .Z1_t (new_AGEMA_signal_3356), .Z1_f (new_AGEMA_signal_3357) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_3_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS12ser[3]), .B0_f (new_AGEMA_signal_3355), .B1_t (new_AGEMA_signal_3356), .B1_f (new_AGEMA_signal_3357), .Z0_t (KeyArray_S12reg_gff_1_SFF_3_n1), .Z0_f (new_AGEMA_signal_6697), .Z1_t (new_AGEMA_signal_6698), .Z1_f (new_AGEMA_signal_6699) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_3_U1 ( .A0_t (KeyArray_S12reg_gff_1_SFF_3_QD), .A0_f (new_AGEMA_signal_4830), .A1_t (new_AGEMA_signal_4831), .A1_f (new_AGEMA_signal_4832), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S12reg_gff_1_SFF_3_n2), .Z0_f (new_AGEMA_signal_6700), .Z1_t (new_AGEMA_signal_6701), .Z1_f (new_AGEMA_signal_6702) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (keySBIn[3]), .A0_f (new_AGEMA_signal_3427), .A1_t (new_AGEMA_signal_3428), .A1_f (new_AGEMA_signal_3429), .B0_t (KeyArray_outS22ser[3]), .B0_f (new_AGEMA_signal_3583), .B1_t (new_AGEMA_signal_3584), .B1_f (new_AGEMA_signal_3585), .Z0_t (KeyArray_S12reg_gff_1_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_3586), .Z1_t (new_AGEMA_signal_3587), .Z1_f (new_AGEMA_signal_3588) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S12reg_gff_1_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_3586), .B1_t (new_AGEMA_signal_3587), .B1_f (new_AGEMA_signal_3588), .Z0_t (KeyArray_S12reg_gff_1_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_4340), .Z1_t (new_AGEMA_signal_4341), .Z1_f (new_AGEMA_signal_4342) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S12reg_gff_1_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_4340), .A1_t (new_AGEMA_signal_4341), .A1_f (new_AGEMA_signal_4342), .B0_t (keySBIn[3]), .B0_f (new_AGEMA_signal_3427), .B1_t (new_AGEMA_signal_3428), .B1_f (new_AGEMA_signal_3429), .Z0_t (KeyArray_S12reg_gff_1_SFF_3_QD), .Z0_f (new_AGEMA_signal_4830), .Z1_t (new_AGEMA_signal_4831), .Z1_f (new_AGEMA_signal_4832) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S12reg_gff_1_SFF_4_U3 ( .A0_t (KeyArray_S12reg_gff_1_SFF_4_n2), .A0_f (new_AGEMA_signal_6706), .A1_t (new_AGEMA_signal_6707), .A1_f (new_AGEMA_signal_6708), .B0_t (KeyArray_S12reg_gff_1_SFF_4_n1), .B0_f (new_AGEMA_signal_6703), .B1_t (new_AGEMA_signal_6704), .B1_f (new_AGEMA_signal_6705), .Z0_t (KeyArray_outS12ser[4]), .Z0_f (new_AGEMA_signal_3364), .Z1_t (new_AGEMA_signal_3365), .Z1_f (new_AGEMA_signal_3366) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_4_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS12ser[4]), .B0_f (new_AGEMA_signal_3364), .B1_t (new_AGEMA_signal_3365), .B1_f (new_AGEMA_signal_3366), .Z0_t (KeyArray_S12reg_gff_1_SFF_4_n1), .Z0_f (new_AGEMA_signal_6703), .Z1_t (new_AGEMA_signal_6704), .Z1_f (new_AGEMA_signal_6705) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_4_U1 ( .A0_t (KeyArray_S12reg_gff_1_SFF_4_QD), .A0_f (new_AGEMA_signal_4833), .A1_t (new_AGEMA_signal_4834), .A1_f (new_AGEMA_signal_4835), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S12reg_gff_1_SFF_4_n2), .Z0_f (new_AGEMA_signal_6706), .Z1_t (new_AGEMA_signal_6707), .Z1_f (new_AGEMA_signal_6708) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (keySBIn[4]), .A0_f (new_AGEMA_signal_3436), .A1_t (new_AGEMA_signal_3437), .A1_f (new_AGEMA_signal_3438), .B0_t (KeyArray_outS22ser[4]), .B0_f (new_AGEMA_signal_3589), .B1_t (new_AGEMA_signal_3590), .B1_f (new_AGEMA_signal_3591), .Z0_t (KeyArray_S12reg_gff_1_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_3592), .Z1_t (new_AGEMA_signal_3593), .Z1_f (new_AGEMA_signal_3594) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S12reg_gff_1_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_3592), .B1_t (new_AGEMA_signal_3593), .B1_f (new_AGEMA_signal_3594), .Z0_t (KeyArray_S12reg_gff_1_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_4343), .Z1_t (new_AGEMA_signal_4344), .Z1_f (new_AGEMA_signal_4345) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S12reg_gff_1_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_4343), .A1_t (new_AGEMA_signal_4344), .A1_f (new_AGEMA_signal_4345), .B0_t (keySBIn[4]), .B0_f (new_AGEMA_signal_3436), .B1_t (new_AGEMA_signal_3437), .B1_f (new_AGEMA_signal_3438), .Z0_t (KeyArray_S12reg_gff_1_SFF_4_QD), .Z0_f (new_AGEMA_signal_4833), .Z1_t (new_AGEMA_signal_4834), .Z1_f (new_AGEMA_signal_4835) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S12reg_gff_1_SFF_5_U3 ( .A0_t (KeyArray_S12reg_gff_1_SFF_5_n2), .A0_f (new_AGEMA_signal_6712), .A1_t (new_AGEMA_signal_6713), .A1_f (new_AGEMA_signal_6714), .B0_t (KeyArray_S12reg_gff_1_SFF_5_n1), .B0_f (new_AGEMA_signal_6709), .B1_t (new_AGEMA_signal_6710), .B1_f (new_AGEMA_signal_6711), .Z0_t (KeyArray_outS12ser[5]), .Z0_f (new_AGEMA_signal_3373), .Z1_t (new_AGEMA_signal_3374), .Z1_f (new_AGEMA_signal_3375) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_5_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS12ser[5]), .B0_f (new_AGEMA_signal_3373), .B1_t (new_AGEMA_signal_3374), .B1_f (new_AGEMA_signal_3375), .Z0_t (KeyArray_S12reg_gff_1_SFF_5_n1), .Z0_f (new_AGEMA_signal_6709), .Z1_t (new_AGEMA_signal_6710), .Z1_f (new_AGEMA_signal_6711) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_5_U1 ( .A0_t (KeyArray_S12reg_gff_1_SFF_5_QD), .A0_f (new_AGEMA_signal_4836), .A1_t (new_AGEMA_signal_4837), .A1_f (new_AGEMA_signal_4838), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S12reg_gff_1_SFF_5_n2), .Z0_f (new_AGEMA_signal_6712), .Z1_t (new_AGEMA_signal_6713), .Z1_f (new_AGEMA_signal_6714) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (keySBIn[5]), .A0_f (new_AGEMA_signal_3445), .A1_t (new_AGEMA_signal_3446), .A1_f (new_AGEMA_signal_3447), .B0_t (KeyArray_outS22ser[5]), .B0_f (new_AGEMA_signal_3595), .B1_t (new_AGEMA_signal_3596), .B1_f (new_AGEMA_signal_3597), .Z0_t (KeyArray_S12reg_gff_1_SFF_5_MUXInst_X), .Z0_f (new_AGEMA_signal_3598), .Z1_t (new_AGEMA_signal_3599), .Z1_f (new_AGEMA_signal_3600) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S12reg_gff_1_SFF_5_MUXInst_X), .B0_f (new_AGEMA_signal_3598), .B1_t (new_AGEMA_signal_3599), .B1_f (new_AGEMA_signal_3600), .Z0_t (KeyArray_S12reg_gff_1_SFF_5_MUXInst_Y), .Z0_f (new_AGEMA_signal_4346), .Z1_t (new_AGEMA_signal_4347), .Z1_f (new_AGEMA_signal_4348) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S12reg_gff_1_SFF_5_MUXInst_Y), .A0_f (new_AGEMA_signal_4346), .A1_t (new_AGEMA_signal_4347), .A1_f (new_AGEMA_signal_4348), .B0_t (keySBIn[5]), .B0_f (new_AGEMA_signal_3445), .B1_t (new_AGEMA_signal_3446), .B1_f (new_AGEMA_signal_3447), .Z0_t (KeyArray_S12reg_gff_1_SFF_5_QD), .Z0_f (new_AGEMA_signal_4836), .Z1_t (new_AGEMA_signal_4837), .Z1_f (new_AGEMA_signal_4838) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S12reg_gff_1_SFF_6_U3 ( .A0_t (KeyArray_S12reg_gff_1_SFF_6_n2), .A0_f (new_AGEMA_signal_6718), .A1_t (new_AGEMA_signal_6719), .A1_f (new_AGEMA_signal_6720), .B0_t (KeyArray_S12reg_gff_1_SFF_6_n1), .B0_f (new_AGEMA_signal_6715), .B1_t (new_AGEMA_signal_6716), .B1_f (new_AGEMA_signal_6717), .Z0_t (KeyArray_outS12ser[6]), .Z0_f (new_AGEMA_signal_3382), .Z1_t (new_AGEMA_signal_3383), .Z1_f (new_AGEMA_signal_3384) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_6_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS12ser[6]), .B0_f (new_AGEMA_signal_3382), .B1_t (new_AGEMA_signal_3383), .B1_f (new_AGEMA_signal_3384), .Z0_t (KeyArray_S12reg_gff_1_SFF_6_n1), .Z0_f (new_AGEMA_signal_6715), .Z1_t (new_AGEMA_signal_6716), .Z1_f (new_AGEMA_signal_6717) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_6_U1 ( .A0_t (KeyArray_S12reg_gff_1_SFF_6_QD), .A0_f (new_AGEMA_signal_4839), .A1_t (new_AGEMA_signal_4840), .A1_f (new_AGEMA_signal_4841), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S12reg_gff_1_SFF_6_n2), .Z0_f (new_AGEMA_signal_6718), .Z1_t (new_AGEMA_signal_6719), .Z1_f (new_AGEMA_signal_6720) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (keySBIn[6]), .A0_f (new_AGEMA_signal_3454), .A1_t (new_AGEMA_signal_3455), .A1_f (new_AGEMA_signal_3456), .B0_t (KeyArray_outS22ser[6]), .B0_f (new_AGEMA_signal_3601), .B1_t (new_AGEMA_signal_3602), .B1_f (new_AGEMA_signal_3603), .Z0_t (KeyArray_S12reg_gff_1_SFF_6_MUXInst_X), .Z0_f (new_AGEMA_signal_3604), .Z1_t (new_AGEMA_signal_3605), .Z1_f (new_AGEMA_signal_3606) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S12reg_gff_1_SFF_6_MUXInst_X), .B0_f (new_AGEMA_signal_3604), .B1_t (new_AGEMA_signal_3605), .B1_f (new_AGEMA_signal_3606), .Z0_t (KeyArray_S12reg_gff_1_SFF_6_MUXInst_Y), .Z0_f (new_AGEMA_signal_4349), .Z1_t (new_AGEMA_signal_4350), .Z1_f (new_AGEMA_signal_4351) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S12reg_gff_1_SFF_6_MUXInst_Y), .A0_f (new_AGEMA_signal_4349), .A1_t (new_AGEMA_signal_4350), .A1_f (new_AGEMA_signal_4351), .B0_t (keySBIn[6]), .B0_f (new_AGEMA_signal_3454), .B1_t (new_AGEMA_signal_3455), .B1_f (new_AGEMA_signal_3456), .Z0_t (KeyArray_S12reg_gff_1_SFF_6_QD), .Z0_f (new_AGEMA_signal_4839), .Z1_t (new_AGEMA_signal_4840), .Z1_f (new_AGEMA_signal_4841) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S12reg_gff_1_SFF_7_U3 ( .A0_t (KeyArray_S12reg_gff_1_SFF_7_n2), .A0_f (new_AGEMA_signal_6724), .A1_t (new_AGEMA_signal_6725), .A1_f (new_AGEMA_signal_6726), .B0_t (KeyArray_S12reg_gff_1_SFF_7_n1), .B0_f (new_AGEMA_signal_6721), .B1_t (new_AGEMA_signal_6722), .B1_f (new_AGEMA_signal_6723), .Z0_t (KeyArray_outS12ser[7]), .Z0_f (new_AGEMA_signal_3391), .Z1_t (new_AGEMA_signal_3392), .Z1_f (new_AGEMA_signal_3393) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_7_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS12ser[7]), .B0_f (new_AGEMA_signal_3391), .B1_t (new_AGEMA_signal_3392), .B1_f (new_AGEMA_signal_3393), .Z0_t (KeyArray_S12reg_gff_1_SFF_7_n1), .Z0_f (new_AGEMA_signal_6721), .Z1_t (new_AGEMA_signal_6722), .Z1_f (new_AGEMA_signal_6723) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_7_U1 ( .A0_t (KeyArray_S12reg_gff_1_SFF_7_QD), .A0_f (new_AGEMA_signal_4842), .A1_t (new_AGEMA_signal_4843), .A1_f (new_AGEMA_signal_4844), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S12reg_gff_1_SFF_7_n2), .Z0_f (new_AGEMA_signal_6724), .Z1_t (new_AGEMA_signal_6725), .Z1_f (new_AGEMA_signal_6726) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (keySBIn[7]), .A0_f (new_AGEMA_signal_3463), .A1_t (new_AGEMA_signal_3464), .A1_f (new_AGEMA_signal_3465), .B0_t (KeyArray_outS22ser[7]), .B0_f (new_AGEMA_signal_3607), .B1_t (new_AGEMA_signal_3608), .B1_f (new_AGEMA_signal_3609), .Z0_t (KeyArray_S12reg_gff_1_SFF_7_MUXInst_X), .Z0_f (new_AGEMA_signal_3610), .Z1_t (new_AGEMA_signal_3611), .Z1_f (new_AGEMA_signal_3612) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S12reg_gff_1_SFF_7_MUXInst_X), .B0_f (new_AGEMA_signal_3610), .B1_t (new_AGEMA_signal_3611), .B1_f (new_AGEMA_signal_3612), .Z0_t (KeyArray_S12reg_gff_1_SFF_7_MUXInst_Y), .Z0_f (new_AGEMA_signal_4352), .Z1_t (new_AGEMA_signal_4353), .Z1_f (new_AGEMA_signal_4354) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S12reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S12reg_gff_1_SFF_7_MUXInst_Y), .A0_f (new_AGEMA_signal_4352), .A1_t (new_AGEMA_signal_4353), .A1_f (new_AGEMA_signal_4354), .B0_t (keySBIn[7]), .B0_f (new_AGEMA_signal_3463), .B1_t (new_AGEMA_signal_3464), .B1_f (new_AGEMA_signal_3465), .Z0_t (KeyArray_S12reg_gff_1_SFF_7_QD), .Z0_f (new_AGEMA_signal_4842), .Z1_t (new_AGEMA_signal_4843), .Z1_f (new_AGEMA_signal_4844) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S13reg_gff_1_SFF_0_U3 ( .A0_t (KeyArray_S13reg_gff_1_SFF_0_n2), .A0_f (new_AGEMA_signal_6730), .A1_t (new_AGEMA_signal_6731), .A1_f (new_AGEMA_signal_6732), .B0_t (KeyArray_S13reg_gff_1_SFF_0_n1), .B0_f (new_AGEMA_signal_6727), .B1_t (new_AGEMA_signal_6728), .B1_f (new_AGEMA_signal_6729), .Z0_t (keySBIn[0]), .Z0_f (new_AGEMA_signal_3400), .Z1_t (new_AGEMA_signal_3401), .Z1_f (new_AGEMA_signal_3402) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_0_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (keySBIn[0]), .B0_f (new_AGEMA_signal_3400), .B1_t (new_AGEMA_signal_3401), .B1_f (new_AGEMA_signal_3402), .Z0_t (KeyArray_S13reg_gff_1_SFF_0_n1), .Z0_f (new_AGEMA_signal_6727), .Z1_t (new_AGEMA_signal_6728), .Z1_f (new_AGEMA_signal_6729) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_0_U1 ( .A0_t (KeyArray_S13reg_gff_1_SFF_0_QD), .A0_f (new_AGEMA_signal_4845), .A1_t (new_AGEMA_signal_4846), .A1_f (new_AGEMA_signal_4847), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S13reg_gff_1_SFF_0_n2), .Z0_f (new_AGEMA_signal_6730), .Z1_t (new_AGEMA_signal_6731), .Z1_f (new_AGEMA_signal_6732) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS20ser[0]), .A0_f (new_AGEMA_signal_3469), .A1_t (new_AGEMA_signal_3470), .A1_f (new_AGEMA_signal_3471), .B0_t (KeyArray_outS23ser[0]), .B0_f (new_AGEMA_signal_3613), .B1_t (new_AGEMA_signal_3614), .B1_f (new_AGEMA_signal_3615), .Z0_t (KeyArray_S13reg_gff_1_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_3616), .Z1_t (new_AGEMA_signal_3617), .Z1_f (new_AGEMA_signal_3618) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S13reg_gff_1_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_3616), .B1_t (new_AGEMA_signal_3617), .B1_f (new_AGEMA_signal_3618), .Z0_t (KeyArray_S13reg_gff_1_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_4355), .Z1_t (new_AGEMA_signal_4356), .Z1_f (new_AGEMA_signal_4357) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S13reg_gff_1_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_4355), .A1_t (new_AGEMA_signal_4356), .A1_f (new_AGEMA_signal_4357), .B0_t (KeyArray_outS20ser[0]), .B0_f (new_AGEMA_signal_3469), .B1_t (new_AGEMA_signal_3470), .B1_f (new_AGEMA_signal_3471), .Z0_t (KeyArray_S13reg_gff_1_SFF_0_QD), .Z0_f (new_AGEMA_signal_4845), .Z1_t (new_AGEMA_signal_4846), .Z1_f (new_AGEMA_signal_4847) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S13reg_gff_1_SFF_1_U3 ( .A0_t (KeyArray_S13reg_gff_1_SFF_1_n2), .A0_f (new_AGEMA_signal_6736), .A1_t (new_AGEMA_signal_6737), .A1_f (new_AGEMA_signal_6738), .B0_t (KeyArray_S13reg_gff_1_SFF_1_n1), .B0_f (new_AGEMA_signal_6733), .B1_t (new_AGEMA_signal_6734), .B1_f (new_AGEMA_signal_6735), .Z0_t (keySBIn[1]), .Z0_f (new_AGEMA_signal_3409), .Z1_t (new_AGEMA_signal_3410), .Z1_f (new_AGEMA_signal_3411) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_1_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (keySBIn[1]), .B0_f (new_AGEMA_signal_3409), .B1_t (new_AGEMA_signal_3410), .B1_f (new_AGEMA_signal_3411), .Z0_t (KeyArray_S13reg_gff_1_SFF_1_n1), .Z0_f (new_AGEMA_signal_6733), .Z1_t (new_AGEMA_signal_6734), .Z1_f (new_AGEMA_signal_6735) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_1_U1 ( .A0_t (KeyArray_S13reg_gff_1_SFF_1_QD), .A0_f (new_AGEMA_signal_4848), .A1_t (new_AGEMA_signal_4849), .A1_f (new_AGEMA_signal_4850), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S13reg_gff_1_SFF_1_n2), .Z0_f (new_AGEMA_signal_6736), .Z1_t (new_AGEMA_signal_6737), .Z1_f (new_AGEMA_signal_6738) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS20ser[1]), .A0_f (new_AGEMA_signal_3475), .A1_t (new_AGEMA_signal_3476), .A1_f (new_AGEMA_signal_3477), .B0_t (KeyArray_outS23ser[1]), .B0_f (new_AGEMA_signal_3619), .B1_t (new_AGEMA_signal_3620), .B1_f (new_AGEMA_signal_3621), .Z0_t (KeyArray_S13reg_gff_1_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_3622), .Z1_t (new_AGEMA_signal_3623), .Z1_f (new_AGEMA_signal_3624) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S13reg_gff_1_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_3622), .B1_t (new_AGEMA_signal_3623), .B1_f (new_AGEMA_signal_3624), .Z0_t (KeyArray_S13reg_gff_1_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_4358), .Z1_t (new_AGEMA_signal_4359), .Z1_f (new_AGEMA_signal_4360) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S13reg_gff_1_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_4358), .A1_t (new_AGEMA_signal_4359), .A1_f (new_AGEMA_signal_4360), .B0_t (KeyArray_outS20ser[1]), .B0_f (new_AGEMA_signal_3475), .B1_t (new_AGEMA_signal_3476), .B1_f (new_AGEMA_signal_3477), .Z0_t (KeyArray_S13reg_gff_1_SFF_1_QD), .Z0_f (new_AGEMA_signal_4848), .Z1_t (new_AGEMA_signal_4849), .Z1_f (new_AGEMA_signal_4850) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S13reg_gff_1_SFF_2_U3 ( .A0_t (KeyArray_S13reg_gff_1_SFF_2_n2), .A0_f (new_AGEMA_signal_6742), .A1_t (new_AGEMA_signal_6743), .A1_f (new_AGEMA_signal_6744), .B0_t (KeyArray_S13reg_gff_1_SFF_2_n1), .B0_f (new_AGEMA_signal_6739), .B1_t (new_AGEMA_signal_6740), .B1_f (new_AGEMA_signal_6741), .Z0_t (keySBIn[2]), .Z0_f (new_AGEMA_signal_3418), .Z1_t (new_AGEMA_signal_3419), .Z1_f (new_AGEMA_signal_3420) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_2_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (keySBIn[2]), .B0_f (new_AGEMA_signal_3418), .B1_t (new_AGEMA_signal_3419), .B1_f (new_AGEMA_signal_3420), .Z0_t (KeyArray_S13reg_gff_1_SFF_2_n1), .Z0_f (new_AGEMA_signal_6739), .Z1_t (new_AGEMA_signal_6740), .Z1_f (new_AGEMA_signal_6741) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_2_U1 ( .A0_t (KeyArray_S13reg_gff_1_SFF_2_QD), .A0_f (new_AGEMA_signal_4851), .A1_t (new_AGEMA_signal_4852), .A1_f (new_AGEMA_signal_4853), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S13reg_gff_1_SFF_2_n2), .Z0_f (new_AGEMA_signal_6742), .Z1_t (new_AGEMA_signal_6743), .Z1_f (new_AGEMA_signal_6744) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS20ser[2]), .A0_f (new_AGEMA_signal_3481), .A1_t (new_AGEMA_signal_3482), .A1_f (new_AGEMA_signal_3483), .B0_t (KeyArray_outS23ser[2]), .B0_f (new_AGEMA_signal_3625), .B1_t (new_AGEMA_signal_3626), .B1_f (new_AGEMA_signal_3627), .Z0_t (KeyArray_S13reg_gff_1_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_3628), .Z1_t (new_AGEMA_signal_3629), .Z1_f (new_AGEMA_signal_3630) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S13reg_gff_1_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_3628), .B1_t (new_AGEMA_signal_3629), .B1_f (new_AGEMA_signal_3630), .Z0_t (KeyArray_S13reg_gff_1_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_4361), .Z1_t (new_AGEMA_signal_4362), .Z1_f (new_AGEMA_signal_4363) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S13reg_gff_1_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_4361), .A1_t (new_AGEMA_signal_4362), .A1_f (new_AGEMA_signal_4363), .B0_t (KeyArray_outS20ser[2]), .B0_f (new_AGEMA_signal_3481), .B1_t (new_AGEMA_signal_3482), .B1_f (new_AGEMA_signal_3483), .Z0_t (KeyArray_S13reg_gff_1_SFF_2_QD), .Z0_f (new_AGEMA_signal_4851), .Z1_t (new_AGEMA_signal_4852), .Z1_f (new_AGEMA_signal_4853) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S13reg_gff_1_SFF_3_U3 ( .A0_t (KeyArray_S13reg_gff_1_SFF_3_n2), .A0_f (new_AGEMA_signal_6748), .A1_t (new_AGEMA_signal_6749), .A1_f (new_AGEMA_signal_6750), .B0_t (KeyArray_S13reg_gff_1_SFF_3_n1), .B0_f (new_AGEMA_signal_6745), .B1_t (new_AGEMA_signal_6746), .B1_f (new_AGEMA_signal_6747), .Z0_t (keySBIn[3]), .Z0_f (new_AGEMA_signal_3427), .Z1_t (new_AGEMA_signal_3428), .Z1_f (new_AGEMA_signal_3429) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_3_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (keySBIn[3]), .B0_f (new_AGEMA_signal_3427), .B1_t (new_AGEMA_signal_3428), .B1_f (new_AGEMA_signal_3429), .Z0_t (KeyArray_S13reg_gff_1_SFF_3_n1), .Z0_f (new_AGEMA_signal_6745), .Z1_t (new_AGEMA_signal_6746), .Z1_f (new_AGEMA_signal_6747) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_3_U1 ( .A0_t (KeyArray_S13reg_gff_1_SFF_3_QD), .A0_f (new_AGEMA_signal_4854), .A1_t (new_AGEMA_signal_4855), .A1_f (new_AGEMA_signal_4856), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S13reg_gff_1_SFF_3_n2), .Z0_f (new_AGEMA_signal_6748), .Z1_t (new_AGEMA_signal_6749), .Z1_f (new_AGEMA_signal_6750) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS20ser[3]), .A0_f (new_AGEMA_signal_3487), .A1_t (new_AGEMA_signal_3488), .A1_f (new_AGEMA_signal_3489), .B0_t (KeyArray_outS23ser[3]), .B0_f (new_AGEMA_signal_3631), .B1_t (new_AGEMA_signal_3632), .B1_f (new_AGEMA_signal_3633), .Z0_t (KeyArray_S13reg_gff_1_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_3634), .Z1_t (new_AGEMA_signal_3635), .Z1_f (new_AGEMA_signal_3636) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S13reg_gff_1_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_3634), .B1_t (new_AGEMA_signal_3635), .B1_f (new_AGEMA_signal_3636), .Z0_t (KeyArray_S13reg_gff_1_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_4364), .Z1_t (new_AGEMA_signal_4365), .Z1_f (new_AGEMA_signal_4366) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S13reg_gff_1_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_4364), .A1_t (new_AGEMA_signal_4365), .A1_f (new_AGEMA_signal_4366), .B0_t (KeyArray_outS20ser[3]), .B0_f (new_AGEMA_signal_3487), .B1_t (new_AGEMA_signal_3488), .B1_f (new_AGEMA_signal_3489), .Z0_t (KeyArray_S13reg_gff_1_SFF_3_QD), .Z0_f (new_AGEMA_signal_4854), .Z1_t (new_AGEMA_signal_4855), .Z1_f (new_AGEMA_signal_4856) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S13reg_gff_1_SFF_4_U3 ( .A0_t (KeyArray_S13reg_gff_1_SFF_4_n2), .A0_f (new_AGEMA_signal_6754), .A1_t (new_AGEMA_signal_6755), .A1_f (new_AGEMA_signal_6756), .B0_t (KeyArray_S13reg_gff_1_SFF_4_n1), .B0_f (new_AGEMA_signal_6751), .B1_t (new_AGEMA_signal_6752), .B1_f (new_AGEMA_signal_6753), .Z0_t (keySBIn[4]), .Z0_f (new_AGEMA_signal_3436), .Z1_t (new_AGEMA_signal_3437), .Z1_f (new_AGEMA_signal_3438) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_4_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (keySBIn[4]), .B0_f (new_AGEMA_signal_3436), .B1_t (new_AGEMA_signal_3437), .B1_f (new_AGEMA_signal_3438), .Z0_t (KeyArray_S13reg_gff_1_SFF_4_n1), .Z0_f (new_AGEMA_signal_6751), .Z1_t (new_AGEMA_signal_6752), .Z1_f (new_AGEMA_signal_6753) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_4_U1 ( .A0_t (KeyArray_S13reg_gff_1_SFF_4_QD), .A0_f (new_AGEMA_signal_4857), .A1_t (new_AGEMA_signal_4858), .A1_f (new_AGEMA_signal_4859), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S13reg_gff_1_SFF_4_n2), .Z0_f (new_AGEMA_signal_6754), .Z1_t (new_AGEMA_signal_6755), .Z1_f (new_AGEMA_signal_6756) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS20ser[4]), .A0_f (new_AGEMA_signal_3493), .A1_t (new_AGEMA_signal_3494), .A1_f (new_AGEMA_signal_3495), .B0_t (KeyArray_outS23ser[4]), .B0_f (new_AGEMA_signal_3637), .B1_t (new_AGEMA_signal_3638), .B1_f (new_AGEMA_signal_3639), .Z0_t (KeyArray_S13reg_gff_1_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_3640), .Z1_t (new_AGEMA_signal_3641), .Z1_f (new_AGEMA_signal_3642) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S13reg_gff_1_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_3640), .B1_t (new_AGEMA_signal_3641), .B1_f (new_AGEMA_signal_3642), .Z0_t (KeyArray_S13reg_gff_1_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_4367), .Z1_t (new_AGEMA_signal_4368), .Z1_f (new_AGEMA_signal_4369) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S13reg_gff_1_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_4367), .A1_t (new_AGEMA_signal_4368), .A1_f (new_AGEMA_signal_4369), .B0_t (KeyArray_outS20ser[4]), .B0_f (new_AGEMA_signal_3493), .B1_t (new_AGEMA_signal_3494), .B1_f (new_AGEMA_signal_3495), .Z0_t (KeyArray_S13reg_gff_1_SFF_4_QD), .Z0_f (new_AGEMA_signal_4857), .Z1_t (new_AGEMA_signal_4858), .Z1_f (new_AGEMA_signal_4859) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S13reg_gff_1_SFF_5_U3 ( .A0_t (KeyArray_S13reg_gff_1_SFF_5_n2), .A0_f (new_AGEMA_signal_6760), .A1_t (new_AGEMA_signal_6761), .A1_f (new_AGEMA_signal_6762), .B0_t (KeyArray_S13reg_gff_1_SFF_5_n1), .B0_f (new_AGEMA_signal_6757), .B1_t (new_AGEMA_signal_6758), .B1_f (new_AGEMA_signal_6759), .Z0_t (keySBIn[5]), .Z0_f (new_AGEMA_signal_3445), .Z1_t (new_AGEMA_signal_3446), .Z1_f (new_AGEMA_signal_3447) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_5_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (keySBIn[5]), .B0_f (new_AGEMA_signal_3445), .B1_t (new_AGEMA_signal_3446), .B1_f (new_AGEMA_signal_3447), .Z0_t (KeyArray_S13reg_gff_1_SFF_5_n1), .Z0_f (new_AGEMA_signal_6757), .Z1_t (new_AGEMA_signal_6758), .Z1_f (new_AGEMA_signal_6759) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_5_U1 ( .A0_t (KeyArray_S13reg_gff_1_SFF_5_QD), .A0_f (new_AGEMA_signal_4860), .A1_t (new_AGEMA_signal_4861), .A1_f (new_AGEMA_signal_4862), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S13reg_gff_1_SFF_5_n2), .Z0_f (new_AGEMA_signal_6760), .Z1_t (new_AGEMA_signal_6761), .Z1_f (new_AGEMA_signal_6762) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS20ser[5]), .A0_f (new_AGEMA_signal_3499), .A1_t (new_AGEMA_signal_3500), .A1_f (new_AGEMA_signal_3501), .B0_t (KeyArray_outS23ser[5]), .B0_f (new_AGEMA_signal_3643), .B1_t (new_AGEMA_signal_3644), .B1_f (new_AGEMA_signal_3645), .Z0_t (KeyArray_S13reg_gff_1_SFF_5_MUXInst_X), .Z0_f (new_AGEMA_signal_3646), .Z1_t (new_AGEMA_signal_3647), .Z1_f (new_AGEMA_signal_3648) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S13reg_gff_1_SFF_5_MUXInst_X), .B0_f (new_AGEMA_signal_3646), .B1_t (new_AGEMA_signal_3647), .B1_f (new_AGEMA_signal_3648), .Z0_t (KeyArray_S13reg_gff_1_SFF_5_MUXInst_Y), .Z0_f (new_AGEMA_signal_4370), .Z1_t (new_AGEMA_signal_4371), .Z1_f (new_AGEMA_signal_4372) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S13reg_gff_1_SFF_5_MUXInst_Y), .A0_f (new_AGEMA_signal_4370), .A1_t (new_AGEMA_signal_4371), .A1_f (new_AGEMA_signal_4372), .B0_t (KeyArray_outS20ser[5]), .B0_f (new_AGEMA_signal_3499), .B1_t (new_AGEMA_signal_3500), .B1_f (new_AGEMA_signal_3501), .Z0_t (KeyArray_S13reg_gff_1_SFF_5_QD), .Z0_f (new_AGEMA_signal_4860), .Z1_t (new_AGEMA_signal_4861), .Z1_f (new_AGEMA_signal_4862) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S13reg_gff_1_SFF_6_U3 ( .A0_t (KeyArray_S13reg_gff_1_SFF_6_n2), .A0_f (new_AGEMA_signal_6766), .A1_t (new_AGEMA_signal_6767), .A1_f (new_AGEMA_signal_6768), .B0_t (KeyArray_S13reg_gff_1_SFF_6_n1), .B0_f (new_AGEMA_signal_6763), .B1_t (new_AGEMA_signal_6764), .B1_f (new_AGEMA_signal_6765), .Z0_t (keySBIn[6]), .Z0_f (new_AGEMA_signal_3454), .Z1_t (new_AGEMA_signal_3455), .Z1_f (new_AGEMA_signal_3456) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_6_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (keySBIn[6]), .B0_f (new_AGEMA_signal_3454), .B1_t (new_AGEMA_signal_3455), .B1_f (new_AGEMA_signal_3456), .Z0_t (KeyArray_S13reg_gff_1_SFF_6_n1), .Z0_f (new_AGEMA_signal_6763), .Z1_t (new_AGEMA_signal_6764), .Z1_f (new_AGEMA_signal_6765) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_6_U1 ( .A0_t (KeyArray_S13reg_gff_1_SFF_6_QD), .A0_f (new_AGEMA_signal_4863), .A1_t (new_AGEMA_signal_4864), .A1_f (new_AGEMA_signal_4865), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S13reg_gff_1_SFF_6_n2), .Z0_f (new_AGEMA_signal_6766), .Z1_t (new_AGEMA_signal_6767), .Z1_f (new_AGEMA_signal_6768) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS20ser[6]), .A0_f (new_AGEMA_signal_3505), .A1_t (new_AGEMA_signal_3506), .A1_f (new_AGEMA_signal_3507), .B0_t (KeyArray_outS23ser[6]), .B0_f (new_AGEMA_signal_3649), .B1_t (new_AGEMA_signal_3650), .B1_f (new_AGEMA_signal_3651), .Z0_t (KeyArray_S13reg_gff_1_SFF_6_MUXInst_X), .Z0_f (new_AGEMA_signal_3652), .Z1_t (new_AGEMA_signal_3653), .Z1_f (new_AGEMA_signal_3654) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S13reg_gff_1_SFF_6_MUXInst_X), .B0_f (new_AGEMA_signal_3652), .B1_t (new_AGEMA_signal_3653), .B1_f (new_AGEMA_signal_3654), .Z0_t (KeyArray_S13reg_gff_1_SFF_6_MUXInst_Y), .Z0_f (new_AGEMA_signal_4373), .Z1_t (new_AGEMA_signal_4374), .Z1_f (new_AGEMA_signal_4375) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S13reg_gff_1_SFF_6_MUXInst_Y), .A0_f (new_AGEMA_signal_4373), .A1_t (new_AGEMA_signal_4374), .A1_f (new_AGEMA_signal_4375), .B0_t (KeyArray_outS20ser[6]), .B0_f (new_AGEMA_signal_3505), .B1_t (new_AGEMA_signal_3506), .B1_f (new_AGEMA_signal_3507), .Z0_t (KeyArray_S13reg_gff_1_SFF_6_QD), .Z0_f (new_AGEMA_signal_4863), .Z1_t (new_AGEMA_signal_4864), .Z1_f (new_AGEMA_signal_4865) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S13reg_gff_1_SFF_7_U3 ( .A0_t (KeyArray_S13reg_gff_1_SFF_7_n2), .A0_f (new_AGEMA_signal_6772), .A1_t (new_AGEMA_signal_6773), .A1_f (new_AGEMA_signal_6774), .B0_t (KeyArray_S13reg_gff_1_SFF_7_n1), .B0_f (new_AGEMA_signal_6769), .B1_t (new_AGEMA_signal_6770), .B1_f (new_AGEMA_signal_6771), .Z0_t (keySBIn[7]), .Z0_f (new_AGEMA_signal_3463), .Z1_t (new_AGEMA_signal_3464), .Z1_f (new_AGEMA_signal_3465) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_7_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (keySBIn[7]), .B0_f (new_AGEMA_signal_3463), .B1_t (new_AGEMA_signal_3464), .B1_f (new_AGEMA_signal_3465), .Z0_t (KeyArray_S13reg_gff_1_SFF_7_n1), .Z0_f (new_AGEMA_signal_6769), .Z1_t (new_AGEMA_signal_6770), .Z1_f (new_AGEMA_signal_6771) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_7_U1 ( .A0_t (KeyArray_S13reg_gff_1_SFF_7_QD), .A0_f (new_AGEMA_signal_4866), .A1_t (new_AGEMA_signal_4867), .A1_f (new_AGEMA_signal_4868), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S13reg_gff_1_SFF_7_n2), .Z0_f (new_AGEMA_signal_6772), .Z1_t (new_AGEMA_signal_6773), .Z1_f (new_AGEMA_signal_6774) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS20ser[7]), .A0_f (new_AGEMA_signal_3511), .A1_t (new_AGEMA_signal_3512), .A1_f (new_AGEMA_signal_3513), .B0_t (KeyArray_outS23ser[7]), .B0_f (new_AGEMA_signal_3655), .B1_t (new_AGEMA_signal_3656), .B1_f (new_AGEMA_signal_3657), .Z0_t (KeyArray_S13reg_gff_1_SFF_7_MUXInst_X), .Z0_f (new_AGEMA_signal_3658), .Z1_t (new_AGEMA_signal_3659), .Z1_f (new_AGEMA_signal_3660) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S13reg_gff_1_SFF_7_MUXInst_X), .B0_f (new_AGEMA_signal_3658), .B1_t (new_AGEMA_signal_3659), .B1_f (new_AGEMA_signal_3660), .Z0_t (KeyArray_S13reg_gff_1_SFF_7_MUXInst_Y), .Z0_f (new_AGEMA_signal_4376), .Z1_t (new_AGEMA_signal_4377), .Z1_f (new_AGEMA_signal_4378) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S13reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S13reg_gff_1_SFF_7_MUXInst_Y), .A0_f (new_AGEMA_signal_4376), .A1_t (new_AGEMA_signal_4377), .A1_f (new_AGEMA_signal_4378), .B0_t (KeyArray_outS20ser[7]), .B0_f (new_AGEMA_signal_3511), .B1_t (new_AGEMA_signal_3512), .B1_f (new_AGEMA_signal_3513), .Z0_t (KeyArray_S13reg_gff_1_SFF_7_QD), .Z0_f (new_AGEMA_signal_4866), .Z1_t (new_AGEMA_signal_4867), .Z1_f (new_AGEMA_signal_4868) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S20reg_gff_1_SFF_0_U3 ( .A0_t (KeyArray_S20reg_gff_1_SFF_0_n2), .A0_f (new_AGEMA_signal_6778), .A1_t (new_AGEMA_signal_6779), .A1_f (new_AGEMA_signal_6780), .B0_t (KeyArray_S20reg_gff_1_SFF_0_n1), .B0_f (new_AGEMA_signal_6775), .B1_t (new_AGEMA_signal_6776), .B1_f (new_AGEMA_signal_6777), .Z0_t (KeyArray_outS20ser[0]), .Z0_f (new_AGEMA_signal_3469), .Z1_t (new_AGEMA_signal_3470), .Z1_f (new_AGEMA_signal_3471) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_0_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS20ser[0]), .B0_f (new_AGEMA_signal_3469), .B1_t (new_AGEMA_signal_3470), .B1_f (new_AGEMA_signal_3471), .Z0_t (KeyArray_S20reg_gff_1_SFF_0_n1), .Z0_f (new_AGEMA_signal_6775), .Z1_t (new_AGEMA_signal_6776), .Z1_f (new_AGEMA_signal_6777) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_0_U1 ( .A0_t (KeyArray_S20reg_gff_1_SFF_0_QD), .A0_f (new_AGEMA_signal_4869), .A1_t (new_AGEMA_signal_4870), .A1_f (new_AGEMA_signal_4871), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S20reg_gff_1_SFF_0_n2), .Z0_f (new_AGEMA_signal_6778), .Z1_t (new_AGEMA_signal_6779), .Z1_f (new_AGEMA_signal_6780) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS21ser[0]), .A0_f (new_AGEMA_signal_3517), .A1_t (new_AGEMA_signal_3518), .A1_f (new_AGEMA_signal_3519), .B0_t (KeyArray_outS30ser[0]), .B0_f (new_AGEMA_signal_3661), .B1_t (new_AGEMA_signal_3662), .B1_f (new_AGEMA_signal_3663), .Z0_t (KeyArray_S20reg_gff_1_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_3664), .Z1_t (new_AGEMA_signal_3665), .Z1_f (new_AGEMA_signal_3666) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S20reg_gff_1_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_3664), .B1_t (new_AGEMA_signal_3665), .B1_f (new_AGEMA_signal_3666), .Z0_t (KeyArray_S20reg_gff_1_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_4379), .Z1_t (new_AGEMA_signal_4380), .Z1_f (new_AGEMA_signal_4381) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S20reg_gff_1_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_4379), .A1_t (new_AGEMA_signal_4380), .A1_f (new_AGEMA_signal_4381), .B0_t (KeyArray_outS21ser[0]), .B0_f (new_AGEMA_signal_3517), .B1_t (new_AGEMA_signal_3518), .B1_f (new_AGEMA_signal_3519), .Z0_t (KeyArray_S20reg_gff_1_SFF_0_QD), .Z0_f (new_AGEMA_signal_4869), .Z1_t (new_AGEMA_signal_4870), .Z1_f (new_AGEMA_signal_4871) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S20reg_gff_1_SFF_1_U3 ( .A0_t (KeyArray_S20reg_gff_1_SFF_1_n2), .A0_f (new_AGEMA_signal_6784), .A1_t (new_AGEMA_signal_6785), .A1_f (new_AGEMA_signal_6786), .B0_t (KeyArray_S20reg_gff_1_SFF_1_n1), .B0_f (new_AGEMA_signal_6781), .B1_t (new_AGEMA_signal_6782), .B1_f (new_AGEMA_signal_6783), .Z0_t (KeyArray_outS20ser[1]), .Z0_f (new_AGEMA_signal_3475), .Z1_t (new_AGEMA_signal_3476), .Z1_f (new_AGEMA_signal_3477) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_1_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS20ser[1]), .B0_f (new_AGEMA_signal_3475), .B1_t (new_AGEMA_signal_3476), .B1_f (new_AGEMA_signal_3477), .Z0_t (KeyArray_S20reg_gff_1_SFF_1_n1), .Z0_f (new_AGEMA_signal_6781), .Z1_t (new_AGEMA_signal_6782), .Z1_f (new_AGEMA_signal_6783) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_1_U1 ( .A0_t (KeyArray_S20reg_gff_1_SFF_1_QD), .A0_f (new_AGEMA_signal_4872), .A1_t (new_AGEMA_signal_4873), .A1_f (new_AGEMA_signal_4874), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S20reg_gff_1_SFF_1_n2), .Z0_f (new_AGEMA_signal_6784), .Z1_t (new_AGEMA_signal_6785), .Z1_f (new_AGEMA_signal_6786) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS21ser[1]), .A0_f (new_AGEMA_signal_3523), .A1_t (new_AGEMA_signal_3524), .A1_f (new_AGEMA_signal_3525), .B0_t (KeyArray_outS30ser[1]), .B0_f (new_AGEMA_signal_3667), .B1_t (new_AGEMA_signal_3668), .B1_f (new_AGEMA_signal_3669), .Z0_t (KeyArray_S20reg_gff_1_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_3670), .Z1_t (new_AGEMA_signal_3671), .Z1_f (new_AGEMA_signal_3672) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S20reg_gff_1_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_3670), .B1_t (new_AGEMA_signal_3671), .B1_f (new_AGEMA_signal_3672), .Z0_t (KeyArray_S20reg_gff_1_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_4382), .Z1_t (new_AGEMA_signal_4383), .Z1_f (new_AGEMA_signal_4384) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S20reg_gff_1_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_4382), .A1_t (new_AGEMA_signal_4383), .A1_f (new_AGEMA_signal_4384), .B0_t (KeyArray_outS21ser[1]), .B0_f (new_AGEMA_signal_3523), .B1_t (new_AGEMA_signal_3524), .B1_f (new_AGEMA_signal_3525), .Z0_t (KeyArray_S20reg_gff_1_SFF_1_QD), .Z0_f (new_AGEMA_signal_4872), .Z1_t (new_AGEMA_signal_4873), .Z1_f (new_AGEMA_signal_4874) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S20reg_gff_1_SFF_2_U3 ( .A0_t (KeyArray_S20reg_gff_1_SFF_2_n2), .A0_f (new_AGEMA_signal_6790), .A1_t (new_AGEMA_signal_6791), .A1_f (new_AGEMA_signal_6792), .B0_t (KeyArray_S20reg_gff_1_SFF_2_n1), .B0_f (new_AGEMA_signal_6787), .B1_t (new_AGEMA_signal_6788), .B1_f (new_AGEMA_signal_6789), .Z0_t (KeyArray_outS20ser[2]), .Z0_f (new_AGEMA_signal_3481), .Z1_t (new_AGEMA_signal_3482), .Z1_f (new_AGEMA_signal_3483) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_2_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS20ser[2]), .B0_f (new_AGEMA_signal_3481), .B1_t (new_AGEMA_signal_3482), .B1_f (new_AGEMA_signal_3483), .Z0_t (KeyArray_S20reg_gff_1_SFF_2_n1), .Z0_f (new_AGEMA_signal_6787), .Z1_t (new_AGEMA_signal_6788), .Z1_f (new_AGEMA_signal_6789) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_2_U1 ( .A0_t (KeyArray_S20reg_gff_1_SFF_2_QD), .A0_f (new_AGEMA_signal_4875), .A1_t (new_AGEMA_signal_4876), .A1_f (new_AGEMA_signal_4877), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S20reg_gff_1_SFF_2_n2), .Z0_f (new_AGEMA_signal_6790), .Z1_t (new_AGEMA_signal_6791), .Z1_f (new_AGEMA_signal_6792) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS21ser[2]), .A0_f (new_AGEMA_signal_3529), .A1_t (new_AGEMA_signal_3530), .A1_f (new_AGEMA_signal_3531), .B0_t (KeyArray_outS30ser[2]), .B0_f (new_AGEMA_signal_3673), .B1_t (new_AGEMA_signal_3674), .B1_f (new_AGEMA_signal_3675), .Z0_t (KeyArray_S20reg_gff_1_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_3676), .Z1_t (new_AGEMA_signal_3677), .Z1_f (new_AGEMA_signal_3678) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S20reg_gff_1_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_3676), .B1_t (new_AGEMA_signal_3677), .B1_f (new_AGEMA_signal_3678), .Z0_t (KeyArray_S20reg_gff_1_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_4385), .Z1_t (new_AGEMA_signal_4386), .Z1_f (new_AGEMA_signal_4387) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S20reg_gff_1_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_4385), .A1_t (new_AGEMA_signal_4386), .A1_f (new_AGEMA_signal_4387), .B0_t (KeyArray_outS21ser[2]), .B0_f (new_AGEMA_signal_3529), .B1_t (new_AGEMA_signal_3530), .B1_f (new_AGEMA_signal_3531), .Z0_t (KeyArray_S20reg_gff_1_SFF_2_QD), .Z0_f (new_AGEMA_signal_4875), .Z1_t (new_AGEMA_signal_4876), .Z1_f (new_AGEMA_signal_4877) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S20reg_gff_1_SFF_3_U3 ( .A0_t (KeyArray_S20reg_gff_1_SFF_3_n2), .A0_f (new_AGEMA_signal_6796), .A1_t (new_AGEMA_signal_6797), .A1_f (new_AGEMA_signal_6798), .B0_t (KeyArray_S20reg_gff_1_SFF_3_n1), .B0_f (new_AGEMA_signal_6793), .B1_t (new_AGEMA_signal_6794), .B1_f (new_AGEMA_signal_6795), .Z0_t (KeyArray_outS20ser[3]), .Z0_f (new_AGEMA_signal_3487), .Z1_t (new_AGEMA_signal_3488), .Z1_f (new_AGEMA_signal_3489) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_3_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS20ser[3]), .B0_f (new_AGEMA_signal_3487), .B1_t (new_AGEMA_signal_3488), .B1_f (new_AGEMA_signal_3489), .Z0_t (KeyArray_S20reg_gff_1_SFF_3_n1), .Z0_f (new_AGEMA_signal_6793), .Z1_t (new_AGEMA_signal_6794), .Z1_f (new_AGEMA_signal_6795) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_3_U1 ( .A0_t (KeyArray_S20reg_gff_1_SFF_3_QD), .A0_f (new_AGEMA_signal_4878), .A1_t (new_AGEMA_signal_4879), .A1_f (new_AGEMA_signal_4880), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S20reg_gff_1_SFF_3_n2), .Z0_f (new_AGEMA_signal_6796), .Z1_t (new_AGEMA_signal_6797), .Z1_f (new_AGEMA_signal_6798) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS21ser[3]), .A0_f (new_AGEMA_signal_3535), .A1_t (new_AGEMA_signal_3536), .A1_f (new_AGEMA_signal_3537), .B0_t (KeyArray_outS30ser[3]), .B0_f (new_AGEMA_signal_3679), .B1_t (new_AGEMA_signal_3680), .B1_f (new_AGEMA_signal_3681), .Z0_t (KeyArray_S20reg_gff_1_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_3682), .Z1_t (new_AGEMA_signal_3683), .Z1_f (new_AGEMA_signal_3684) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S20reg_gff_1_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_3682), .B1_t (new_AGEMA_signal_3683), .B1_f (new_AGEMA_signal_3684), .Z0_t (KeyArray_S20reg_gff_1_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_4388), .Z1_t (new_AGEMA_signal_4389), .Z1_f (new_AGEMA_signal_4390) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S20reg_gff_1_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_4388), .A1_t (new_AGEMA_signal_4389), .A1_f (new_AGEMA_signal_4390), .B0_t (KeyArray_outS21ser[3]), .B0_f (new_AGEMA_signal_3535), .B1_t (new_AGEMA_signal_3536), .B1_f (new_AGEMA_signal_3537), .Z0_t (KeyArray_S20reg_gff_1_SFF_3_QD), .Z0_f (new_AGEMA_signal_4878), .Z1_t (new_AGEMA_signal_4879), .Z1_f (new_AGEMA_signal_4880) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S20reg_gff_1_SFF_4_U3 ( .A0_t (KeyArray_S20reg_gff_1_SFF_4_n2), .A0_f (new_AGEMA_signal_6802), .A1_t (new_AGEMA_signal_6803), .A1_f (new_AGEMA_signal_6804), .B0_t (KeyArray_S20reg_gff_1_SFF_4_n1), .B0_f (new_AGEMA_signal_6799), .B1_t (new_AGEMA_signal_6800), .B1_f (new_AGEMA_signal_6801), .Z0_t (KeyArray_outS20ser[4]), .Z0_f (new_AGEMA_signal_3493), .Z1_t (new_AGEMA_signal_3494), .Z1_f (new_AGEMA_signal_3495) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_4_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS20ser[4]), .B0_f (new_AGEMA_signal_3493), .B1_t (new_AGEMA_signal_3494), .B1_f (new_AGEMA_signal_3495), .Z0_t (KeyArray_S20reg_gff_1_SFF_4_n1), .Z0_f (new_AGEMA_signal_6799), .Z1_t (new_AGEMA_signal_6800), .Z1_f (new_AGEMA_signal_6801) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_4_U1 ( .A0_t (KeyArray_S20reg_gff_1_SFF_4_QD), .A0_f (new_AGEMA_signal_4881), .A1_t (new_AGEMA_signal_4882), .A1_f (new_AGEMA_signal_4883), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S20reg_gff_1_SFF_4_n2), .Z0_f (new_AGEMA_signal_6802), .Z1_t (new_AGEMA_signal_6803), .Z1_f (new_AGEMA_signal_6804) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS21ser[4]), .A0_f (new_AGEMA_signal_3541), .A1_t (new_AGEMA_signal_3542), .A1_f (new_AGEMA_signal_3543), .B0_t (KeyArray_outS30ser[4]), .B0_f (new_AGEMA_signal_3685), .B1_t (new_AGEMA_signal_3686), .B1_f (new_AGEMA_signal_3687), .Z0_t (KeyArray_S20reg_gff_1_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_3688), .Z1_t (new_AGEMA_signal_3689), .Z1_f (new_AGEMA_signal_3690) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S20reg_gff_1_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_3688), .B1_t (new_AGEMA_signal_3689), .B1_f (new_AGEMA_signal_3690), .Z0_t (KeyArray_S20reg_gff_1_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_4391), .Z1_t (new_AGEMA_signal_4392), .Z1_f (new_AGEMA_signal_4393) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S20reg_gff_1_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_4391), .A1_t (new_AGEMA_signal_4392), .A1_f (new_AGEMA_signal_4393), .B0_t (KeyArray_outS21ser[4]), .B0_f (new_AGEMA_signal_3541), .B1_t (new_AGEMA_signal_3542), .B1_f (new_AGEMA_signal_3543), .Z0_t (KeyArray_S20reg_gff_1_SFF_4_QD), .Z0_f (new_AGEMA_signal_4881), .Z1_t (new_AGEMA_signal_4882), .Z1_f (new_AGEMA_signal_4883) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S20reg_gff_1_SFF_5_U3 ( .A0_t (KeyArray_S20reg_gff_1_SFF_5_n2), .A0_f (new_AGEMA_signal_6808), .A1_t (new_AGEMA_signal_6809), .A1_f (new_AGEMA_signal_6810), .B0_t (KeyArray_S20reg_gff_1_SFF_5_n1), .B0_f (new_AGEMA_signal_6805), .B1_t (new_AGEMA_signal_6806), .B1_f (new_AGEMA_signal_6807), .Z0_t (KeyArray_outS20ser[5]), .Z0_f (new_AGEMA_signal_3499), .Z1_t (new_AGEMA_signal_3500), .Z1_f (new_AGEMA_signal_3501) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_5_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS20ser[5]), .B0_f (new_AGEMA_signal_3499), .B1_t (new_AGEMA_signal_3500), .B1_f (new_AGEMA_signal_3501), .Z0_t (KeyArray_S20reg_gff_1_SFF_5_n1), .Z0_f (new_AGEMA_signal_6805), .Z1_t (new_AGEMA_signal_6806), .Z1_f (new_AGEMA_signal_6807) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_5_U1 ( .A0_t (KeyArray_S20reg_gff_1_SFF_5_QD), .A0_f (new_AGEMA_signal_4884), .A1_t (new_AGEMA_signal_4885), .A1_f (new_AGEMA_signal_4886), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S20reg_gff_1_SFF_5_n2), .Z0_f (new_AGEMA_signal_6808), .Z1_t (new_AGEMA_signal_6809), .Z1_f (new_AGEMA_signal_6810) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS21ser[5]), .A0_f (new_AGEMA_signal_3547), .A1_t (new_AGEMA_signal_3548), .A1_f (new_AGEMA_signal_3549), .B0_t (KeyArray_outS30ser[5]), .B0_f (new_AGEMA_signal_3691), .B1_t (new_AGEMA_signal_3692), .B1_f (new_AGEMA_signal_3693), .Z0_t (KeyArray_S20reg_gff_1_SFF_5_MUXInst_X), .Z0_f (new_AGEMA_signal_3694), .Z1_t (new_AGEMA_signal_3695), .Z1_f (new_AGEMA_signal_3696) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S20reg_gff_1_SFF_5_MUXInst_X), .B0_f (new_AGEMA_signal_3694), .B1_t (new_AGEMA_signal_3695), .B1_f (new_AGEMA_signal_3696), .Z0_t (KeyArray_S20reg_gff_1_SFF_5_MUXInst_Y), .Z0_f (new_AGEMA_signal_4394), .Z1_t (new_AGEMA_signal_4395), .Z1_f (new_AGEMA_signal_4396) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S20reg_gff_1_SFF_5_MUXInst_Y), .A0_f (new_AGEMA_signal_4394), .A1_t (new_AGEMA_signal_4395), .A1_f (new_AGEMA_signal_4396), .B0_t (KeyArray_outS21ser[5]), .B0_f (new_AGEMA_signal_3547), .B1_t (new_AGEMA_signal_3548), .B1_f (new_AGEMA_signal_3549), .Z0_t (KeyArray_S20reg_gff_1_SFF_5_QD), .Z0_f (new_AGEMA_signal_4884), .Z1_t (new_AGEMA_signal_4885), .Z1_f (new_AGEMA_signal_4886) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S20reg_gff_1_SFF_6_U3 ( .A0_t (KeyArray_S20reg_gff_1_SFF_6_n2), .A0_f (new_AGEMA_signal_6814), .A1_t (new_AGEMA_signal_6815), .A1_f (new_AGEMA_signal_6816), .B0_t (KeyArray_S20reg_gff_1_SFF_6_n1), .B0_f (new_AGEMA_signal_6811), .B1_t (new_AGEMA_signal_6812), .B1_f (new_AGEMA_signal_6813), .Z0_t (KeyArray_outS20ser[6]), .Z0_f (new_AGEMA_signal_3505), .Z1_t (new_AGEMA_signal_3506), .Z1_f (new_AGEMA_signal_3507) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_6_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS20ser[6]), .B0_f (new_AGEMA_signal_3505), .B1_t (new_AGEMA_signal_3506), .B1_f (new_AGEMA_signal_3507), .Z0_t (KeyArray_S20reg_gff_1_SFF_6_n1), .Z0_f (new_AGEMA_signal_6811), .Z1_t (new_AGEMA_signal_6812), .Z1_f (new_AGEMA_signal_6813) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_6_U1 ( .A0_t (KeyArray_S20reg_gff_1_SFF_6_QD), .A0_f (new_AGEMA_signal_4887), .A1_t (new_AGEMA_signal_4888), .A1_f (new_AGEMA_signal_4889), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S20reg_gff_1_SFF_6_n2), .Z0_f (new_AGEMA_signal_6814), .Z1_t (new_AGEMA_signal_6815), .Z1_f (new_AGEMA_signal_6816) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS21ser[6]), .A0_f (new_AGEMA_signal_3553), .A1_t (new_AGEMA_signal_3554), .A1_f (new_AGEMA_signal_3555), .B0_t (KeyArray_outS30ser[6]), .B0_f (new_AGEMA_signal_3697), .B1_t (new_AGEMA_signal_3698), .B1_f (new_AGEMA_signal_3699), .Z0_t (KeyArray_S20reg_gff_1_SFF_6_MUXInst_X), .Z0_f (new_AGEMA_signal_3700), .Z1_t (new_AGEMA_signal_3701), .Z1_f (new_AGEMA_signal_3702) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S20reg_gff_1_SFF_6_MUXInst_X), .B0_f (new_AGEMA_signal_3700), .B1_t (new_AGEMA_signal_3701), .B1_f (new_AGEMA_signal_3702), .Z0_t (KeyArray_S20reg_gff_1_SFF_6_MUXInst_Y), .Z0_f (new_AGEMA_signal_4397), .Z1_t (new_AGEMA_signal_4398), .Z1_f (new_AGEMA_signal_4399) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S20reg_gff_1_SFF_6_MUXInst_Y), .A0_f (new_AGEMA_signal_4397), .A1_t (new_AGEMA_signal_4398), .A1_f (new_AGEMA_signal_4399), .B0_t (KeyArray_outS21ser[6]), .B0_f (new_AGEMA_signal_3553), .B1_t (new_AGEMA_signal_3554), .B1_f (new_AGEMA_signal_3555), .Z0_t (KeyArray_S20reg_gff_1_SFF_6_QD), .Z0_f (new_AGEMA_signal_4887), .Z1_t (new_AGEMA_signal_4888), .Z1_f (new_AGEMA_signal_4889) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S20reg_gff_1_SFF_7_U3 ( .A0_t (KeyArray_S20reg_gff_1_SFF_7_n2), .A0_f (new_AGEMA_signal_6820), .A1_t (new_AGEMA_signal_6821), .A1_f (new_AGEMA_signal_6822), .B0_t (KeyArray_S20reg_gff_1_SFF_7_n1), .B0_f (new_AGEMA_signal_6817), .B1_t (new_AGEMA_signal_6818), .B1_f (new_AGEMA_signal_6819), .Z0_t (KeyArray_outS20ser[7]), .Z0_f (new_AGEMA_signal_3511), .Z1_t (new_AGEMA_signal_3512), .Z1_f (new_AGEMA_signal_3513) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_7_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS20ser[7]), .B0_f (new_AGEMA_signal_3511), .B1_t (new_AGEMA_signal_3512), .B1_f (new_AGEMA_signal_3513), .Z0_t (KeyArray_S20reg_gff_1_SFF_7_n1), .Z0_f (new_AGEMA_signal_6817), .Z1_t (new_AGEMA_signal_6818), .Z1_f (new_AGEMA_signal_6819) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_7_U1 ( .A0_t (KeyArray_S20reg_gff_1_SFF_7_QD), .A0_f (new_AGEMA_signal_4890), .A1_t (new_AGEMA_signal_4891), .A1_f (new_AGEMA_signal_4892), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S20reg_gff_1_SFF_7_n2), .Z0_f (new_AGEMA_signal_6820), .Z1_t (new_AGEMA_signal_6821), .Z1_f (new_AGEMA_signal_6822) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS21ser[7]), .A0_f (new_AGEMA_signal_3559), .A1_t (new_AGEMA_signal_3560), .A1_f (new_AGEMA_signal_3561), .B0_t (KeyArray_outS30ser[7]), .B0_f (new_AGEMA_signal_3703), .B1_t (new_AGEMA_signal_3704), .B1_f (new_AGEMA_signal_3705), .Z0_t (KeyArray_S20reg_gff_1_SFF_7_MUXInst_X), .Z0_f (new_AGEMA_signal_3706), .Z1_t (new_AGEMA_signal_3707), .Z1_f (new_AGEMA_signal_3708) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S20reg_gff_1_SFF_7_MUXInst_X), .B0_f (new_AGEMA_signal_3706), .B1_t (new_AGEMA_signal_3707), .B1_f (new_AGEMA_signal_3708), .Z0_t (KeyArray_S20reg_gff_1_SFF_7_MUXInst_Y), .Z0_f (new_AGEMA_signal_4400), .Z1_t (new_AGEMA_signal_4401), .Z1_f (new_AGEMA_signal_4402) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S20reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S20reg_gff_1_SFF_7_MUXInst_Y), .A0_f (new_AGEMA_signal_4400), .A1_t (new_AGEMA_signal_4401), .A1_f (new_AGEMA_signal_4402), .B0_t (KeyArray_outS21ser[7]), .B0_f (new_AGEMA_signal_3559), .B1_t (new_AGEMA_signal_3560), .B1_f (new_AGEMA_signal_3561), .Z0_t (KeyArray_S20reg_gff_1_SFF_7_QD), .Z0_f (new_AGEMA_signal_4890), .Z1_t (new_AGEMA_signal_4891), .Z1_f (new_AGEMA_signal_4892) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S21reg_gff_1_SFF_0_U3 ( .A0_t (KeyArray_S21reg_gff_1_SFF_0_n2), .A0_f (new_AGEMA_signal_6826), .A1_t (new_AGEMA_signal_6827), .A1_f (new_AGEMA_signal_6828), .B0_t (KeyArray_S21reg_gff_1_SFF_0_n1), .B0_f (new_AGEMA_signal_6823), .B1_t (new_AGEMA_signal_6824), .B1_f (new_AGEMA_signal_6825), .Z0_t (KeyArray_outS21ser[0]), .Z0_f (new_AGEMA_signal_3517), .Z1_t (new_AGEMA_signal_3518), .Z1_f (new_AGEMA_signal_3519) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_0_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS21ser[0]), .B0_f (new_AGEMA_signal_3517), .B1_t (new_AGEMA_signal_3518), .B1_f (new_AGEMA_signal_3519), .Z0_t (KeyArray_S21reg_gff_1_SFF_0_n1), .Z0_f (new_AGEMA_signal_6823), .Z1_t (new_AGEMA_signal_6824), .Z1_f (new_AGEMA_signal_6825) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_0_U1 ( .A0_t (KeyArray_S21reg_gff_1_SFF_0_QD), .A0_f (new_AGEMA_signal_4893), .A1_t (new_AGEMA_signal_4894), .A1_f (new_AGEMA_signal_4895), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S21reg_gff_1_SFF_0_n2), .Z0_f (new_AGEMA_signal_6826), .Z1_t (new_AGEMA_signal_6827), .Z1_f (new_AGEMA_signal_6828) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS22ser[0]), .A0_f (new_AGEMA_signal_3565), .A1_t (new_AGEMA_signal_3566), .A1_f (new_AGEMA_signal_3567), .B0_t (KeyArray_outS31ser[0]), .B0_f (new_AGEMA_signal_3709), .B1_t (new_AGEMA_signal_3710), .B1_f (new_AGEMA_signal_3711), .Z0_t (KeyArray_S21reg_gff_1_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_3712), .Z1_t (new_AGEMA_signal_3713), .Z1_f (new_AGEMA_signal_3714) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S21reg_gff_1_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_3712), .B1_t (new_AGEMA_signal_3713), .B1_f (new_AGEMA_signal_3714), .Z0_t (KeyArray_S21reg_gff_1_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_4403), .Z1_t (new_AGEMA_signal_4404), .Z1_f (new_AGEMA_signal_4405) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S21reg_gff_1_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_4403), .A1_t (new_AGEMA_signal_4404), .A1_f (new_AGEMA_signal_4405), .B0_t (KeyArray_outS22ser[0]), .B0_f (new_AGEMA_signal_3565), .B1_t (new_AGEMA_signal_3566), .B1_f (new_AGEMA_signal_3567), .Z0_t (KeyArray_S21reg_gff_1_SFF_0_QD), .Z0_f (new_AGEMA_signal_4893), .Z1_t (new_AGEMA_signal_4894), .Z1_f (new_AGEMA_signal_4895) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S21reg_gff_1_SFF_1_U3 ( .A0_t (KeyArray_S21reg_gff_1_SFF_1_n2), .A0_f (new_AGEMA_signal_6832), .A1_t (new_AGEMA_signal_6833), .A1_f (new_AGEMA_signal_6834), .B0_t (KeyArray_S21reg_gff_1_SFF_1_n1), .B0_f (new_AGEMA_signal_6829), .B1_t (new_AGEMA_signal_6830), .B1_f (new_AGEMA_signal_6831), .Z0_t (KeyArray_outS21ser[1]), .Z0_f (new_AGEMA_signal_3523), .Z1_t (new_AGEMA_signal_3524), .Z1_f (new_AGEMA_signal_3525) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_1_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS21ser[1]), .B0_f (new_AGEMA_signal_3523), .B1_t (new_AGEMA_signal_3524), .B1_f (new_AGEMA_signal_3525), .Z0_t (KeyArray_S21reg_gff_1_SFF_1_n1), .Z0_f (new_AGEMA_signal_6829), .Z1_t (new_AGEMA_signal_6830), .Z1_f (new_AGEMA_signal_6831) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_1_U1 ( .A0_t (KeyArray_S21reg_gff_1_SFF_1_QD), .A0_f (new_AGEMA_signal_4896), .A1_t (new_AGEMA_signal_4897), .A1_f (new_AGEMA_signal_4898), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S21reg_gff_1_SFF_1_n2), .Z0_f (new_AGEMA_signal_6832), .Z1_t (new_AGEMA_signal_6833), .Z1_f (new_AGEMA_signal_6834) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS22ser[1]), .A0_f (new_AGEMA_signal_3571), .A1_t (new_AGEMA_signal_3572), .A1_f (new_AGEMA_signal_3573), .B0_t (KeyArray_outS31ser[1]), .B0_f (new_AGEMA_signal_3715), .B1_t (new_AGEMA_signal_3716), .B1_f (new_AGEMA_signal_3717), .Z0_t (KeyArray_S21reg_gff_1_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_3718), .Z1_t (new_AGEMA_signal_3719), .Z1_f (new_AGEMA_signal_3720) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S21reg_gff_1_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_3718), .B1_t (new_AGEMA_signal_3719), .B1_f (new_AGEMA_signal_3720), .Z0_t (KeyArray_S21reg_gff_1_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_4406), .Z1_t (new_AGEMA_signal_4407), .Z1_f (new_AGEMA_signal_4408) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S21reg_gff_1_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_4406), .A1_t (new_AGEMA_signal_4407), .A1_f (new_AGEMA_signal_4408), .B0_t (KeyArray_outS22ser[1]), .B0_f (new_AGEMA_signal_3571), .B1_t (new_AGEMA_signal_3572), .B1_f (new_AGEMA_signal_3573), .Z0_t (KeyArray_S21reg_gff_1_SFF_1_QD), .Z0_f (new_AGEMA_signal_4896), .Z1_t (new_AGEMA_signal_4897), .Z1_f (new_AGEMA_signal_4898) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S21reg_gff_1_SFF_2_U3 ( .A0_t (KeyArray_S21reg_gff_1_SFF_2_n2), .A0_f (new_AGEMA_signal_6838), .A1_t (new_AGEMA_signal_6839), .A1_f (new_AGEMA_signal_6840), .B0_t (KeyArray_S21reg_gff_1_SFF_2_n1), .B0_f (new_AGEMA_signal_6835), .B1_t (new_AGEMA_signal_6836), .B1_f (new_AGEMA_signal_6837), .Z0_t (KeyArray_outS21ser[2]), .Z0_f (new_AGEMA_signal_3529), .Z1_t (new_AGEMA_signal_3530), .Z1_f (new_AGEMA_signal_3531) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_2_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS21ser[2]), .B0_f (new_AGEMA_signal_3529), .B1_t (new_AGEMA_signal_3530), .B1_f (new_AGEMA_signal_3531), .Z0_t (KeyArray_S21reg_gff_1_SFF_2_n1), .Z0_f (new_AGEMA_signal_6835), .Z1_t (new_AGEMA_signal_6836), .Z1_f (new_AGEMA_signal_6837) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_2_U1 ( .A0_t (KeyArray_S21reg_gff_1_SFF_2_QD), .A0_f (new_AGEMA_signal_4899), .A1_t (new_AGEMA_signal_4900), .A1_f (new_AGEMA_signal_4901), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S21reg_gff_1_SFF_2_n2), .Z0_f (new_AGEMA_signal_6838), .Z1_t (new_AGEMA_signal_6839), .Z1_f (new_AGEMA_signal_6840) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS22ser[2]), .A0_f (new_AGEMA_signal_3577), .A1_t (new_AGEMA_signal_3578), .A1_f (new_AGEMA_signal_3579), .B0_t (KeyArray_outS31ser[2]), .B0_f (new_AGEMA_signal_3721), .B1_t (new_AGEMA_signal_3722), .B1_f (new_AGEMA_signal_3723), .Z0_t (KeyArray_S21reg_gff_1_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_3724), .Z1_t (new_AGEMA_signal_3725), .Z1_f (new_AGEMA_signal_3726) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S21reg_gff_1_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_3724), .B1_t (new_AGEMA_signal_3725), .B1_f (new_AGEMA_signal_3726), .Z0_t (KeyArray_S21reg_gff_1_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_4409), .Z1_t (new_AGEMA_signal_4410), .Z1_f (new_AGEMA_signal_4411) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S21reg_gff_1_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_4409), .A1_t (new_AGEMA_signal_4410), .A1_f (new_AGEMA_signal_4411), .B0_t (KeyArray_outS22ser[2]), .B0_f (new_AGEMA_signal_3577), .B1_t (new_AGEMA_signal_3578), .B1_f (new_AGEMA_signal_3579), .Z0_t (KeyArray_S21reg_gff_1_SFF_2_QD), .Z0_f (new_AGEMA_signal_4899), .Z1_t (new_AGEMA_signal_4900), .Z1_f (new_AGEMA_signal_4901) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S21reg_gff_1_SFF_3_U3 ( .A0_t (KeyArray_S21reg_gff_1_SFF_3_n2), .A0_f (new_AGEMA_signal_6844), .A1_t (new_AGEMA_signal_6845), .A1_f (new_AGEMA_signal_6846), .B0_t (KeyArray_S21reg_gff_1_SFF_3_n1), .B0_f (new_AGEMA_signal_6841), .B1_t (new_AGEMA_signal_6842), .B1_f (new_AGEMA_signal_6843), .Z0_t (KeyArray_outS21ser[3]), .Z0_f (new_AGEMA_signal_3535), .Z1_t (new_AGEMA_signal_3536), .Z1_f (new_AGEMA_signal_3537) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_3_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS21ser[3]), .B0_f (new_AGEMA_signal_3535), .B1_t (new_AGEMA_signal_3536), .B1_f (new_AGEMA_signal_3537), .Z0_t (KeyArray_S21reg_gff_1_SFF_3_n1), .Z0_f (new_AGEMA_signal_6841), .Z1_t (new_AGEMA_signal_6842), .Z1_f (new_AGEMA_signal_6843) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_3_U1 ( .A0_t (KeyArray_S21reg_gff_1_SFF_3_QD), .A0_f (new_AGEMA_signal_4902), .A1_t (new_AGEMA_signal_4903), .A1_f (new_AGEMA_signal_4904), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S21reg_gff_1_SFF_3_n2), .Z0_f (new_AGEMA_signal_6844), .Z1_t (new_AGEMA_signal_6845), .Z1_f (new_AGEMA_signal_6846) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS22ser[3]), .A0_f (new_AGEMA_signal_3583), .A1_t (new_AGEMA_signal_3584), .A1_f (new_AGEMA_signal_3585), .B0_t (KeyArray_outS31ser[3]), .B0_f (new_AGEMA_signal_3727), .B1_t (new_AGEMA_signal_3728), .B1_f (new_AGEMA_signal_3729), .Z0_t (KeyArray_S21reg_gff_1_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_3730), .Z1_t (new_AGEMA_signal_3731), .Z1_f (new_AGEMA_signal_3732) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S21reg_gff_1_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_3730), .B1_t (new_AGEMA_signal_3731), .B1_f (new_AGEMA_signal_3732), .Z0_t (KeyArray_S21reg_gff_1_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_4412), .Z1_t (new_AGEMA_signal_4413), .Z1_f (new_AGEMA_signal_4414) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S21reg_gff_1_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_4412), .A1_t (new_AGEMA_signal_4413), .A1_f (new_AGEMA_signal_4414), .B0_t (KeyArray_outS22ser[3]), .B0_f (new_AGEMA_signal_3583), .B1_t (new_AGEMA_signal_3584), .B1_f (new_AGEMA_signal_3585), .Z0_t (KeyArray_S21reg_gff_1_SFF_3_QD), .Z0_f (new_AGEMA_signal_4902), .Z1_t (new_AGEMA_signal_4903), .Z1_f (new_AGEMA_signal_4904) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S21reg_gff_1_SFF_4_U3 ( .A0_t (KeyArray_S21reg_gff_1_SFF_4_n2), .A0_f (new_AGEMA_signal_6850), .A1_t (new_AGEMA_signal_6851), .A1_f (new_AGEMA_signal_6852), .B0_t (KeyArray_S21reg_gff_1_SFF_4_n1), .B0_f (new_AGEMA_signal_6847), .B1_t (new_AGEMA_signal_6848), .B1_f (new_AGEMA_signal_6849), .Z0_t (KeyArray_outS21ser[4]), .Z0_f (new_AGEMA_signal_3541), .Z1_t (new_AGEMA_signal_3542), .Z1_f (new_AGEMA_signal_3543) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_4_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS21ser[4]), .B0_f (new_AGEMA_signal_3541), .B1_t (new_AGEMA_signal_3542), .B1_f (new_AGEMA_signal_3543), .Z0_t (KeyArray_S21reg_gff_1_SFF_4_n1), .Z0_f (new_AGEMA_signal_6847), .Z1_t (new_AGEMA_signal_6848), .Z1_f (new_AGEMA_signal_6849) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_4_U1 ( .A0_t (KeyArray_S21reg_gff_1_SFF_4_QD), .A0_f (new_AGEMA_signal_4905), .A1_t (new_AGEMA_signal_4906), .A1_f (new_AGEMA_signal_4907), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S21reg_gff_1_SFF_4_n2), .Z0_f (new_AGEMA_signal_6850), .Z1_t (new_AGEMA_signal_6851), .Z1_f (new_AGEMA_signal_6852) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS22ser[4]), .A0_f (new_AGEMA_signal_3589), .A1_t (new_AGEMA_signal_3590), .A1_f (new_AGEMA_signal_3591), .B0_t (KeyArray_outS31ser[4]), .B0_f (new_AGEMA_signal_3733), .B1_t (new_AGEMA_signal_3734), .B1_f (new_AGEMA_signal_3735), .Z0_t (KeyArray_S21reg_gff_1_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_3736), .Z1_t (new_AGEMA_signal_3737), .Z1_f (new_AGEMA_signal_3738) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S21reg_gff_1_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_3736), .B1_t (new_AGEMA_signal_3737), .B1_f (new_AGEMA_signal_3738), .Z0_t (KeyArray_S21reg_gff_1_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_4415), .Z1_t (new_AGEMA_signal_4416), .Z1_f (new_AGEMA_signal_4417) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S21reg_gff_1_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_4415), .A1_t (new_AGEMA_signal_4416), .A1_f (new_AGEMA_signal_4417), .B0_t (KeyArray_outS22ser[4]), .B0_f (new_AGEMA_signal_3589), .B1_t (new_AGEMA_signal_3590), .B1_f (new_AGEMA_signal_3591), .Z0_t (KeyArray_S21reg_gff_1_SFF_4_QD), .Z0_f (new_AGEMA_signal_4905), .Z1_t (new_AGEMA_signal_4906), .Z1_f (new_AGEMA_signal_4907) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S21reg_gff_1_SFF_5_U3 ( .A0_t (KeyArray_S21reg_gff_1_SFF_5_n2), .A0_f (new_AGEMA_signal_6856), .A1_t (new_AGEMA_signal_6857), .A1_f (new_AGEMA_signal_6858), .B0_t (KeyArray_S21reg_gff_1_SFF_5_n1), .B0_f (new_AGEMA_signal_6853), .B1_t (new_AGEMA_signal_6854), .B1_f (new_AGEMA_signal_6855), .Z0_t (KeyArray_outS21ser[5]), .Z0_f (new_AGEMA_signal_3547), .Z1_t (new_AGEMA_signal_3548), .Z1_f (new_AGEMA_signal_3549) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_5_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS21ser[5]), .B0_f (new_AGEMA_signal_3547), .B1_t (new_AGEMA_signal_3548), .B1_f (new_AGEMA_signal_3549), .Z0_t (KeyArray_S21reg_gff_1_SFF_5_n1), .Z0_f (new_AGEMA_signal_6853), .Z1_t (new_AGEMA_signal_6854), .Z1_f (new_AGEMA_signal_6855) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_5_U1 ( .A0_t (KeyArray_S21reg_gff_1_SFF_5_QD), .A0_f (new_AGEMA_signal_4908), .A1_t (new_AGEMA_signal_4909), .A1_f (new_AGEMA_signal_4910), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S21reg_gff_1_SFF_5_n2), .Z0_f (new_AGEMA_signal_6856), .Z1_t (new_AGEMA_signal_6857), .Z1_f (new_AGEMA_signal_6858) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS22ser[5]), .A0_f (new_AGEMA_signal_3595), .A1_t (new_AGEMA_signal_3596), .A1_f (new_AGEMA_signal_3597), .B0_t (KeyArray_outS31ser[5]), .B0_f (new_AGEMA_signal_3739), .B1_t (new_AGEMA_signal_3740), .B1_f (new_AGEMA_signal_3741), .Z0_t (KeyArray_S21reg_gff_1_SFF_5_MUXInst_X), .Z0_f (new_AGEMA_signal_3742), .Z1_t (new_AGEMA_signal_3743), .Z1_f (new_AGEMA_signal_3744) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S21reg_gff_1_SFF_5_MUXInst_X), .B0_f (new_AGEMA_signal_3742), .B1_t (new_AGEMA_signal_3743), .B1_f (new_AGEMA_signal_3744), .Z0_t (KeyArray_S21reg_gff_1_SFF_5_MUXInst_Y), .Z0_f (new_AGEMA_signal_4418), .Z1_t (new_AGEMA_signal_4419), .Z1_f (new_AGEMA_signal_4420) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S21reg_gff_1_SFF_5_MUXInst_Y), .A0_f (new_AGEMA_signal_4418), .A1_t (new_AGEMA_signal_4419), .A1_f (new_AGEMA_signal_4420), .B0_t (KeyArray_outS22ser[5]), .B0_f (new_AGEMA_signal_3595), .B1_t (new_AGEMA_signal_3596), .B1_f (new_AGEMA_signal_3597), .Z0_t (KeyArray_S21reg_gff_1_SFF_5_QD), .Z0_f (new_AGEMA_signal_4908), .Z1_t (new_AGEMA_signal_4909), .Z1_f (new_AGEMA_signal_4910) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S21reg_gff_1_SFF_6_U3 ( .A0_t (KeyArray_S21reg_gff_1_SFF_6_n2), .A0_f (new_AGEMA_signal_6862), .A1_t (new_AGEMA_signal_6863), .A1_f (new_AGEMA_signal_6864), .B0_t (KeyArray_S21reg_gff_1_SFF_6_n1), .B0_f (new_AGEMA_signal_6859), .B1_t (new_AGEMA_signal_6860), .B1_f (new_AGEMA_signal_6861), .Z0_t (KeyArray_outS21ser[6]), .Z0_f (new_AGEMA_signal_3553), .Z1_t (new_AGEMA_signal_3554), .Z1_f (new_AGEMA_signal_3555) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_6_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS21ser[6]), .B0_f (new_AGEMA_signal_3553), .B1_t (new_AGEMA_signal_3554), .B1_f (new_AGEMA_signal_3555), .Z0_t (KeyArray_S21reg_gff_1_SFF_6_n1), .Z0_f (new_AGEMA_signal_6859), .Z1_t (new_AGEMA_signal_6860), .Z1_f (new_AGEMA_signal_6861) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_6_U1 ( .A0_t (KeyArray_S21reg_gff_1_SFF_6_QD), .A0_f (new_AGEMA_signal_4911), .A1_t (new_AGEMA_signal_4912), .A1_f (new_AGEMA_signal_4913), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S21reg_gff_1_SFF_6_n2), .Z0_f (new_AGEMA_signal_6862), .Z1_t (new_AGEMA_signal_6863), .Z1_f (new_AGEMA_signal_6864) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS22ser[6]), .A0_f (new_AGEMA_signal_3601), .A1_t (new_AGEMA_signal_3602), .A1_f (new_AGEMA_signal_3603), .B0_t (KeyArray_outS31ser[6]), .B0_f (new_AGEMA_signal_3745), .B1_t (new_AGEMA_signal_3746), .B1_f (new_AGEMA_signal_3747), .Z0_t (KeyArray_S21reg_gff_1_SFF_6_MUXInst_X), .Z0_f (new_AGEMA_signal_3748), .Z1_t (new_AGEMA_signal_3749), .Z1_f (new_AGEMA_signal_3750) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S21reg_gff_1_SFF_6_MUXInst_X), .B0_f (new_AGEMA_signal_3748), .B1_t (new_AGEMA_signal_3749), .B1_f (new_AGEMA_signal_3750), .Z0_t (KeyArray_S21reg_gff_1_SFF_6_MUXInst_Y), .Z0_f (new_AGEMA_signal_4421), .Z1_t (new_AGEMA_signal_4422), .Z1_f (new_AGEMA_signal_4423) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S21reg_gff_1_SFF_6_MUXInst_Y), .A0_f (new_AGEMA_signal_4421), .A1_t (new_AGEMA_signal_4422), .A1_f (new_AGEMA_signal_4423), .B0_t (KeyArray_outS22ser[6]), .B0_f (new_AGEMA_signal_3601), .B1_t (new_AGEMA_signal_3602), .B1_f (new_AGEMA_signal_3603), .Z0_t (KeyArray_S21reg_gff_1_SFF_6_QD), .Z0_f (new_AGEMA_signal_4911), .Z1_t (new_AGEMA_signal_4912), .Z1_f (new_AGEMA_signal_4913) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S21reg_gff_1_SFF_7_U3 ( .A0_t (KeyArray_S21reg_gff_1_SFF_7_n2), .A0_f (new_AGEMA_signal_6868), .A1_t (new_AGEMA_signal_6869), .A1_f (new_AGEMA_signal_6870), .B0_t (KeyArray_S21reg_gff_1_SFF_7_n1), .B0_f (new_AGEMA_signal_6865), .B1_t (new_AGEMA_signal_6866), .B1_f (new_AGEMA_signal_6867), .Z0_t (KeyArray_outS21ser[7]), .Z0_f (new_AGEMA_signal_3559), .Z1_t (new_AGEMA_signal_3560), .Z1_f (new_AGEMA_signal_3561) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_7_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS21ser[7]), .B0_f (new_AGEMA_signal_3559), .B1_t (new_AGEMA_signal_3560), .B1_f (new_AGEMA_signal_3561), .Z0_t (KeyArray_S21reg_gff_1_SFF_7_n1), .Z0_f (new_AGEMA_signal_6865), .Z1_t (new_AGEMA_signal_6866), .Z1_f (new_AGEMA_signal_6867) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_7_U1 ( .A0_t (KeyArray_S21reg_gff_1_SFF_7_QD), .A0_f (new_AGEMA_signal_4914), .A1_t (new_AGEMA_signal_4915), .A1_f (new_AGEMA_signal_4916), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S21reg_gff_1_SFF_7_n2), .Z0_f (new_AGEMA_signal_6868), .Z1_t (new_AGEMA_signal_6869), .Z1_f (new_AGEMA_signal_6870) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS22ser[7]), .A0_f (new_AGEMA_signal_3607), .A1_t (new_AGEMA_signal_3608), .A1_f (new_AGEMA_signal_3609), .B0_t (KeyArray_outS31ser[7]), .B0_f (new_AGEMA_signal_3751), .B1_t (new_AGEMA_signal_3752), .B1_f (new_AGEMA_signal_3753), .Z0_t (KeyArray_S21reg_gff_1_SFF_7_MUXInst_X), .Z0_f (new_AGEMA_signal_3754), .Z1_t (new_AGEMA_signal_3755), .Z1_f (new_AGEMA_signal_3756) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S21reg_gff_1_SFF_7_MUXInst_X), .B0_f (new_AGEMA_signal_3754), .B1_t (new_AGEMA_signal_3755), .B1_f (new_AGEMA_signal_3756), .Z0_t (KeyArray_S21reg_gff_1_SFF_7_MUXInst_Y), .Z0_f (new_AGEMA_signal_4424), .Z1_t (new_AGEMA_signal_4425), .Z1_f (new_AGEMA_signal_4426) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S21reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S21reg_gff_1_SFF_7_MUXInst_Y), .A0_f (new_AGEMA_signal_4424), .A1_t (new_AGEMA_signal_4425), .A1_f (new_AGEMA_signal_4426), .B0_t (KeyArray_outS22ser[7]), .B0_f (new_AGEMA_signal_3607), .B1_t (new_AGEMA_signal_3608), .B1_f (new_AGEMA_signal_3609), .Z0_t (KeyArray_S21reg_gff_1_SFF_7_QD), .Z0_f (new_AGEMA_signal_4914), .Z1_t (new_AGEMA_signal_4915), .Z1_f (new_AGEMA_signal_4916) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S22reg_gff_1_SFF_0_U3 ( .A0_t (KeyArray_S22reg_gff_1_SFF_0_n2), .A0_f (new_AGEMA_signal_6874), .A1_t (new_AGEMA_signal_6875), .A1_f (new_AGEMA_signal_6876), .B0_t (KeyArray_S22reg_gff_1_SFF_0_n1), .B0_f (new_AGEMA_signal_6871), .B1_t (new_AGEMA_signal_6872), .B1_f (new_AGEMA_signal_6873), .Z0_t (KeyArray_outS22ser[0]), .Z0_f (new_AGEMA_signal_3565), .Z1_t (new_AGEMA_signal_3566), .Z1_f (new_AGEMA_signal_3567) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_0_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS22ser[0]), .B0_f (new_AGEMA_signal_3565), .B1_t (new_AGEMA_signal_3566), .B1_f (new_AGEMA_signal_3567), .Z0_t (KeyArray_S22reg_gff_1_SFF_0_n1), .Z0_f (new_AGEMA_signal_6871), .Z1_t (new_AGEMA_signal_6872), .Z1_f (new_AGEMA_signal_6873) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_0_U1 ( .A0_t (KeyArray_S22reg_gff_1_SFF_0_QD), .A0_f (new_AGEMA_signal_4917), .A1_t (new_AGEMA_signal_4918), .A1_f (new_AGEMA_signal_4919), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S22reg_gff_1_SFF_0_n2), .Z0_f (new_AGEMA_signal_6874), .Z1_t (new_AGEMA_signal_6875), .Z1_f (new_AGEMA_signal_6876) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS23ser[0]), .A0_f (new_AGEMA_signal_3613), .A1_t (new_AGEMA_signal_3614), .A1_f (new_AGEMA_signal_3615), .B0_t (KeyArray_outS32ser[0]), .B0_f (new_AGEMA_signal_3757), .B1_t (new_AGEMA_signal_3758), .B1_f (new_AGEMA_signal_3759), .Z0_t (KeyArray_S22reg_gff_1_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_3760), .Z1_t (new_AGEMA_signal_3761), .Z1_f (new_AGEMA_signal_3762) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S22reg_gff_1_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_3760), .B1_t (new_AGEMA_signal_3761), .B1_f (new_AGEMA_signal_3762), .Z0_t (KeyArray_S22reg_gff_1_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_4427), .Z1_t (new_AGEMA_signal_4428), .Z1_f (new_AGEMA_signal_4429) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S22reg_gff_1_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_4427), .A1_t (new_AGEMA_signal_4428), .A1_f (new_AGEMA_signal_4429), .B0_t (KeyArray_outS23ser[0]), .B0_f (new_AGEMA_signal_3613), .B1_t (new_AGEMA_signal_3614), .B1_f (new_AGEMA_signal_3615), .Z0_t (KeyArray_S22reg_gff_1_SFF_0_QD), .Z0_f (new_AGEMA_signal_4917), .Z1_t (new_AGEMA_signal_4918), .Z1_f (new_AGEMA_signal_4919) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S22reg_gff_1_SFF_1_U3 ( .A0_t (KeyArray_S22reg_gff_1_SFF_1_n2), .A0_f (new_AGEMA_signal_6880), .A1_t (new_AGEMA_signal_6881), .A1_f (new_AGEMA_signal_6882), .B0_t (KeyArray_S22reg_gff_1_SFF_1_n1), .B0_f (new_AGEMA_signal_6877), .B1_t (new_AGEMA_signal_6878), .B1_f (new_AGEMA_signal_6879), .Z0_t (KeyArray_outS22ser[1]), .Z0_f (new_AGEMA_signal_3571), .Z1_t (new_AGEMA_signal_3572), .Z1_f (new_AGEMA_signal_3573) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_1_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS22ser[1]), .B0_f (new_AGEMA_signal_3571), .B1_t (new_AGEMA_signal_3572), .B1_f (new_AGEMA_signal_3573), .Z0_t (KeyArray_S22reg_gff_1_SFF_1_n1), .Z0_f (new_AGEMA_signal_6877), .Z1_t (new_AGEMA_signal_6878), .Z1_f (new_AGEMA_signal_6879) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_1_U1 ( .A0_t (KeyArray_S22reg_gff_1_SFF_1_QD), .A0_f (new_AGEMA_signal_4920), .A1_t (new_AGEMA_signal_4921), .A1_f (new_AGEMA_signal_4922), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S22reg_gff_1_SFF_1_n2), .Z0_f (new_AGEMA_signal_6880), .Z1_t (new_AGEMA_signal_6881), .Z1_f (new_AGEMA_signal_6882) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS23ser[1]), .A0_f (new_AGEMA_signal_3619), .A1_t (new_AGEMA_signal_3620), .A1_f (new_AGEMA_signal_3621), .B0_t (KeyArray_outS32ser[1]), .B0_f (new_AGEMA_signal_3763), .B1_t (new_AGEMA_signal_3764), .B1_f (new_AGEMA_signal_3765), .Z0_t (KeyArray_S22reg_gff_1_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_3766), .Z1_t (new_AGEMA_signal_3767), .Z1_f (new_AGEMA_signal_3768) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S22reg_gff_1_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_3766), .B1_t (new_AGEMA_signal_3767), .B1_f (new_AGEMA_signal_3768), .Z0_t (KeyArray_S22reg_gff_1_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_4430), .Z1_t (new_AGEMA_signal_4431), .Z1_f (new_AGEMA_signal_4432) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S22reg_gff_1_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_4430), .A1_t (new_AGEMA_signal_4431), .A1_f (new_AGEMA_signal_4432), .B0_t (KeyArray_outS23ser[1]), .B0_f (new_AGEMA_signal_3619), .B1_t (new_AGEMA_signal_3620), .B1_f (new_AGEMA_signal_3621), .Z0_t (KeyArray_S22reg_gff_1_SFF_1_QD), .Z0_f (new_AGEMA_signal_4920), .Z1_t (new_AGEMA_signal_4921), .Z1_f (new_AGEMA_signal_4922) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S22reg_gff_1_SFF_2_U3 ( .A0_t (KeyArray_S22reg_gff_1_SFF_2_n2), .A0_f (new_AGEMA_signal_6886), .A1_t (new_AGEMA_signal_6887), .A1_f (new_AGEMA_signal_6888), .B0_t (KeyArray_S22reg_gff_1_SFF_2_n1), .B0_f (new_AGEMA_signal_6883), .B1_t (new_AGEMA_signal_6884), .B1_f (new_AGEMA_signal_6885), .Z0_t (KeyArray_outS22ser[2]), .Z0_f (new_AGEMA_signal_3577), .Z1_t (new_AGEMA_signal_3578), .Z1_f (new_AGEMA_signal_3579) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_2_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS22ser[2]), .B0_f (new_AGEMA_signal_3577), .B1_t (new_AGEMA_signal_3578), .B1_f (new_AGEMA_signal_3579), .Z0_t (KeyArray_S22reg_gff_1_SFF_2_n1), .Z0_f (new_AGEMA_signal_6883), .Z1_t (new_AGEMA_signal_6884), .Z1_f (new_AGEMA_signal_6885) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_2_U1 ( .A0_t (KeyArray_S22reg_gff_1_SFF_2_QD), .A0_f (new_AGEMA_signal_4923), .A1_t (new_AGEMA_signal_4924), .A1_f (new_AGEMA_signal_4925), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S22reg_gff_1_SFF_2_n2), .Z0_f (new_AGEMA_signal_6886), .Z1_t (new_AGEMA_signal_6887), .Z1_f (new_AGEMA_signal_6888) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS23ser[2]), .A0_f (new_AGEMA_signal_3625), .A1_t (new_AGEMA_signal_3626), .A1_f (new_AGEMA_signal_3627), .B0_t (KeyArray_outS32ser[2]), .B0_f (new_AGEMA_signal_3769), .B1_t (new_AGEMA_signal_3770), .B1_f (new_AGEMA_signal_3771), .Z0_t (KeyArray_S22reg_gff_1_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_3772), .Z1_t (new_AGEMA_signal_3773), .Z1_f (new_AGEMA_signal_3774) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S22reg_gff_1_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_3772), .B1_t (new_AGEMA_signal_3773), .B1_f (new_AGEMA_signal_3774), .Z0_t (KeyArray_S22reg_gff_1_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_4433), .Z1_t (new_AGEMA_signal_4434), .Z1_f (new_AGEMA_signal_4435) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S22reg_gff_1_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_4433), .A1_t (new_AGEMA_signal_4434), .A1_f (new_AGEMA_signal_4435), .B0_t (KeyArray_outS23ser[2]), .B0_f (new_AGEMA_signal_3625), .B1_t (new_AGEMA_signal_3626), .B1_f (new_AGEMA_signal_3627), .Z0_t (KeyArray_S22reg_gff_1_SFF_2_QD), .Z0_f (new_AGEMA_signal_4923), .Z1_t (new_AGEMA_signal_4924), .Z1_f (new_AGEMA_signal_4925) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S22reg_gff_1_SFF_3_U3 ( .A0_t (KeyArray_S22reg_gff_1_SFF_3_n2), .A0_f (new_AGEMA_signal_6892), .A1_t (new_AGEMA_signal_6893), .A1_f (new_AGEMA_signal_6894), .B0_t (KeyArray_S22reg_gff_1_SFF_3_n1), .B0_f (new_AGEMA_signal_6889), .B1_t (new_AGEMA_signal_6890), .B1_f (new_AGEMA_signal_6891), .Z0_t (KeyArray_outS22ser[3]), .Z0_f (new_AGEMA_signal_3583), .Z1_t (new_AGEMA_signal_3584), .Z1_f (new_AGEMA_signal_3585) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_3_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS22ser[3]), .B0_f (new_AGEMA_signal_3583), .B1_t (new_AGEMA_signal_3584), .B1_f (new_AGEMA_signal_3585), .Z0_t (KeyArray_S22reg_gff_1_SFF_3_n1), .Z0_f (new_AGEMA_signal_6889), .Z1_t (new_AGEMA_signal_6890), .Z1_f (new_AGEMA_signal_6891) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_3_U1 ( .A0_t (KeyArray_S22reg_gff_1_SFF_3_QD), .A0_f (new_AGEMA_signal_4926), .A1_t (new_AGEMA_signal_4927), .A1_f (new_AGEMA_signal_4928), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S22reg_gff_1_SFF_3_n2), .Z0_f (new_AGEMA_signal_6892), .Z1_t (new_AGEMA_signal_6893), .Z1_f (new_AGEMA_signal_6894) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS23ser[3]), .A0_f (new_AGEMA_signal_3631), .A1_t (new_AGEMA_signal_3632), .A1_f (new_AGEMA_signal_3633), .B0_t (KeyArray_outS32ser[3]), .B0_f (new_AGEMA_signal_3775), .B1_t (new_AGEMA_signal_3776), .B1_f (new_AGEMA_signal_3777), .Z0_t (KeyArray_S22reg_gff_1_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_3778), .Z1_t (new_AGEMA_signal_3779), .Z1_f (new_AGEMA_signal_3780) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S22reg_gff_1_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_3778), .B1_t (new_AGEMA_signal_3779), .B1_f (new_AGEMA_signal_3780), .Z0_t (KeyArray_S22reg_gff_1_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_4436), .Z1_t (new_AGEMA_signal_4437), .Z1_f (new_AGEMA_signal_4438) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S22reg_gff_1_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_4436), .A1_t (new_AGEMA_signal_4437), .A1_f (new_AGEMA_signal_4438), .B0_t (KeyArray_outS23ser[3]), .B0_f (new_AGEMA_signal_3631), .B1_t (new_AGEMA_signal_3632), .B1_f (new_AGEMA_signal_3633), .Z0_t (KeyArray_S22reg_gff_1_SFF_3_QD), .Z0_f (new_AGEMA_signal_4926), .Z1_t (new_AGEMA_signal_4927), .Z1_f (new_AGEMA_signal_4928) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S22reg_gff_1_SFF_4_U3 ( .A0_t (KeyArray_S22reg_gff_1_SFF_4_n2), .A0_f (new_AGEMA_signal_6898), .A1_t (new_AGEMA_signal_6899), .A1_f (new_AGEMA_signal_6900), .B0_t (KeyArray_S22reg_gff_1_SFF_4_n1), .B0_f (new_AGEMA_signal_6895), .B1_t (new_AGEMA_signal_6896), .B1_f (new_AGEMA_signal_6897), .Z0_t (KeyArray_outS22ser[4]), .Z0_f (new_AGEMA_signal_3589), .Z1_t (new_AGEMA_signal_3590), .Z1_f (new_AGEMA_signal_3591) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_4_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS22ser[4]), .B0_f (new_AGEMA_signal_3589), .B1_t (new_AGEMA_signal_3590), .B1_f (new_AGEMA_signal_3591), .Z0_t (KeyArray_S22reg_gff_1_SFF_4_n1), .Z0_f (new_AGEMA_signal_6895), .Z1_t (new_AGEMA_signal_6896), .Z1_f (new_AGEMA_signal_6897) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_4_U1 ( .A0_t (KeyArray_S22reg_gff_1_SFF_4_QD), .A0_f (new_AGEMA_signal_4929), .A1_t (new_AGEMA_signal_4930), .A1_f (new_AGEMA_signal_4931), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S22reg_gff_1_SFF_4_n2), .Z0_f (new_AGEMA_signal_6898), .Z1_t (new_AGEMA_signal_6899), .Z1_f (new_AGEMA_signal_6900) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS23ser[4]), .A0_f (new_AGEMA_signal_3637), .A1_t (new_AGEMA_signal_3638), .A1_f (new_AGEMA_signal_3639), .B0_t (KeyArray_outS32ser[4]), .B0_f (new_AGEMA_signal_3781), .B1_t (new_AGEMA_signal_3782), .B1_f (new_AGEMA_signal_3783), .Z0_t (KeyArray_S22reg_gff_1_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_3784), .Z1_t (new_AGEMA_signal_3785), .Z1_f (new_AGEMA_signal_3786) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S22reg_gff_1_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_3784), .B1_t (new_AGEMA_signal_3785), .B1_f (new_AGEMA_signal_3786), .Z0_t (KeyArray_S22reg_gff_1_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_4439), .Z1_t (new_AGEMA_signal_4440), .Z1_f (new_AGEMA_signal_4441) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S22reg_gff_1_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_4439), .A1_t (new_AGEMA_signal_4440), .A1_f (new_AGEMA_signal_4441), .B0_t (KeyArray_outS23ser[4]), .B0_f (new_AGEMA_signal_3637), .B1_t (new_AGEMA_signal_3638), .B1_f (new_AGEMA_signal_3639), .Z0_t (KeyArray_S22reg_gff_1_SFF_4_QD), .Z0_f (new_AGEMA_signal_4929), .Z1_t (new_AGEMA_signal_4930), .Z1_f (new_AGEMA_signal_4931) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S22reg_gff_1_SFF_5_U3 ( .A0_t (KeyArray_S22reg_gff_1_SFF_5_n2), .A0_f (new_AGEMA_signal_6904), .A1_t (new_AGEMA_signal_6905), .A1_f (new_AGEMA_signal_6906), .B0_t (KeyArray_S22reg_gff_1_SFF_5_n1), .B0_f (new_AGEMA_signal_6901), .B1_t (new_AGEMA_signal_6902), .B1_f (new_AGEMA_signal_6903), .Z0_t (KeyArray_outS22ser[5]), .Z0_f (new_AGEMA_signal_3595), .Z1_t (new_AGEMA_signal_3596), .Z1_f (new_AGEMA_signal_3597) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_5_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS22ser[5]), .B0_f (new_AGEMA_signal_3595), .B1_t (new_AGEMA_signal_3596), .B1_f (new_AGEMA_signal_3597), .Z0_t (KeyArray_S22reg_gff_1_SFF_5_n1), .Z0_f (new_AGEMA_signal_6901), .Z1_t (new_AGEMA_signal_6902), .Z1_f (new_AGEMA_signal_6903) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_5_U1 ( .A0_t (KeyArray_S22reg_gff_1_SFF_5_QD), .A0_f (new_AGEMA_signal_4932), .A1_t (new_AGEMA_signal_4933), .A1_f (new_AGEMA_signal_4934), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S22reg_gff_1_SFF_5_n2), .Z0_f (new_AGEMA_signal_6904), .Z1_t (new_AGEMA_signal_6905), .Z1_f (new_AGEMA_signal_6906) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS23ser[5]), .A0_f (new_AGEMA_signal_3643), .A1_t (new_AGEMA_signal_3644), .A1_f (new_AGEMA_signal_3645), .B0_t (KeyArray_outS32ser[5]), .B0_f (new_AGEMA_signal_3787), .B1_t (new_AGEMA_signal_3788), .B1_f (new_AGEMA_signal_3789), .Z0_t (KeyArray_S22reg_gff_1_SFF_5_MUXInst_X), .Z0_f (new_AGEMA_signal_3790), .Z1_t (new_AGEMA_signal_3791), .Z1_f (new_AGEMA_signal_3792) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S22reg_gff_1_SFF_5_MUXInst_X), .B0_f (new_AGEMA_signal_3790), .B1_t (new_AGEMA_signal_3791), .B1_f (new_AGEMA_signal_3792), .Z0_t (KeyArray_S22reg_gff_1_SFF_5_MUXInst_Y), .Z0_f (new_AGEMA_signal_4442), .Z1_t (new_AGEMA_signal_4443), .Z1_f (new_AGEMA_signal_4444) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S22reg_gff_1_SFF_5_MUXInst_Y), .A0_f (new_AGEMA_signal_4442), .A1_t (new_AGEMA_signal_4443), .A1_f (new_AGEMA_signal_4444), .B0_t (KeyArray_outS23ser[5]), .B0_f (new_AGEMA_signal_3643), .B1_t (new_AGEMA_signal_3644), .B1_f (new_AGEMA_signal_3645), .Z0_t (KeyArray_S22reg_gff_1_SFF_5_QD), .Z0_f (new_AGEMA_signal_4932), .Z1_t (new_AGEMA_signal_4933), .Z1_f (new_AGEMA_signal_4934) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S22reg_gff_1_SFF_6_U3 ( .A0_t (KeyArray_S22reg_gff_1_SFF_6_n2), .A0_f (new_AGEMA_signal_6910), .A1_t (new_AGEMA_signal_6911), .A1_f (new_AGEMA_signal_6912), .B0_t (KeyArray_S22reg_gff_1_SFF_6_n1), .B0_f (new_AGEMA_signal_6907), .B1_t (new_AGEMA_signal_6908), .B1_f (new_AGEMA_signal_6909), .Z0_t (KeyArray_outS22ser[6]), .Z0_f (new_AGEMA_signal_3601), .Z1_t (new_AGEMA_signal_3602), .Z1_f (new_AGEMA_signal_3603) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_6_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS22ser[6]), .B0_f (new_AGEMA_signal_3601), .B1_t (new_AGEMA_signal_3602), .B1_f (new_AGEMA_signal_3603), .Z0_t (KeyArray_S22reg_gff_1_SFF_6_n1), .Z0_f (new_AGEMA_signal_6907), .Z1_t (new_AGEMA_signal_6908), .Z1_f (new_AGEMA_signal_6909) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_6_U1 ( .A0_t (KeyArray_S22reg_gff_1_SFF_6_QD), .A0_f (new_AGEMA_signal_4935), .A1_t (new_AGEMA_signal_4936), .A1_f (new_AGEMA_signal_4937), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S22reg_gff_1_SFF_6_n2), .Z0_f (new_AGEMA_signal_6910), .Z1_t (new_AGEMA_signal_6911), .Z1_f (new_AGEMA_signal_6912) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS23ser[6]), .A0_f (new_AGEMA_signal_3649), .A1_t (new_AGEMA_signal_3650), .A1_f (new_AGEMA_signal_3651), .B0_t (KeyArray_outS32ser[6]), .B0_f (new_AGEMA_signal_3793), .B1_t (new_AGEMA_signal_3794), .B1_f (new_AGEMA_signal_3795), .Z0_t (KeyArray_S22reg_gff_1_SFF_6_MUXInst_X), .Z0_f (new_AGEMA_signal_3796), .Z1_t (new_AGEMA_signal_3797), .Z1_f (new_AGEMA_signal_3798) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S22reg_gff_1_SFF_6_MUXInst_X), .B0_f (new_AGEMA_signal_3796), .B1_t (new_AGEMA_signal_3797), .B1_f (new_AGEMA_signal_3798), .Z0_t (KeyArray_S22reg_gff_1_SFF_6_MUXInst_Y), .Z0_f (new_AGEMA_signal_4445), .Z1_t (new_AGEMA_signal_4446), .Z1_f (new_AGEMA_signal_4447) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S22reg_gff_1_SFF_6_MUXInst_Y), .A0_f (new_AGEMA_signal_4445), .A1_t (new_AGEMA_signal_4446), .A1_f (new_AGEMA_signal_4447), .B0_t (KeyArray_outS23ser[6]), .B0_f (new_AGEMA_signal_3649), .B1_t (new_AGEMA_signal_3650), .B1_f (new_AGEMA_signal_3651), .Z0_t (KeyArray_S22reg_gff_1_SFF_6_QD), .Z0_f (new_AGEMA_signal_4935), .Z1_t (new_AGEMA_signal_4936), .Z1_f (new_AGEMA_signal_4937) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S22reg_gff_1_SFF_7_U3 ( .A0_t (KeyArray_S22reg_gff_1_SFF_7_n2), .A0_f (new_AGEMA_signal_6916), .A1_t (new_AGEMA_signal_6917), .A1_f (new_AGEMA_signal_6918), .B0_t (KeyArray_S22reg_gff_1_SFF_7_n1), .B0_f (new_AGEMA_signal_6913), .B1_t (new_AGEMA_signal_6914), .B1_f (new_AGEMA_signal_6915), .Z0_t (KeyArray_outS22ser[7]), .Z0_f (new_AGEMA_signal_3607), .Z1_t (new_AGEMA_signal_3608), .Z1_f (new_AGEMA_signal_3609) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_7_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS22ser[7]), .B0_f (new_AGEMA_signal_3607), .B1_t (new_AGEMA_signal_3608), .B1_f (new_AGEMA_signal_3609), .Z0_t (KeyArray_S22reg_gff_1_SFF_7_n1), .Z0_f (new_AGEMA_signal_6913), .Z1_t (new_AGEMA_signal_6914), .Z1_f (new_AGEMA_signal_6915) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_7_U1 ( .A0_t (KeyArray_S22reg_gff_1_SFF_7_QD), .A0_f (new_AGEMA_signal_4938), .A1_t (new_AGEMA_signal_4939), .A1_f (new_AGEMA_signal_4940), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S22reg_gff_1_SFF_7_n2), .Z0_f (new_AGEMA_signal_6916), .Z1_t (new_AGEMA_signal_6917), .Z1_f (new_AGEMA_signal_6918) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS23ser[7]), .A0_f (new_AGEMA_signal_3655), .A1_t (new_AGEMA_signal_3656), .A1_f (new_AGEMA_signal_3657), .B0_t (KeyArray_outS32ser[7]), .B0_f (new_AGEMA_signal_3799), .B1_t (new_AGEMA_signal_3800), .B1_f (new_AGEMA_signal_3801), .Z0_t (KeyArray_S22reg_gff_1_SFF_7_MUXInst_X), .Z0_f (new_AGEMA_signal_3802), .Z1_t (new_AGEMA_signal_3803), .Z1_f (new_AGEMA_signal_3804) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S22reg_gff_1_SFF_7_MUXInst_X), .B0_f (new_AGEMA_signal_3802), .B1_t (new_AGEMA_signal_3803), .B1_f (new_AGEMA_signal_3804), .Z0_t (KeyArray_S22reg_gff_1_SFF_7_MUXInst_Y), .Z0_f (new_AGEMA_signal_4448), .Z1_t (new_AGEMA_signal_4449), .Z1_f (new_AGEMA_signal_4450) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S22reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S22reg_gff_1_SFF_7_MUXInst_Y), .A0_f (new_AGEMA_signal_4448), .A1_t (new_AGEMA_signal_4449), .A1_f (new_AGEMA_signal_4450), .B0_t (KeyArray_outS23ser[7]), .B0_f (new_AGEMA_signal_3655), .B1_t (new_AGEMA_signal_3656), .B1_f (new_AGEMA_signal_3657), .Z0_t (KeyArray_S22reg_gff_1_SFF_7_QD), .Z0_f (new_AGEMA_signal_4938), .Z1_t (new_AGEMA_signal_4939), .Z1_f (new_AGEMA_signal_4940) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S23reg_gff_1_SFF_0_U3 ( .A0_t (KeyArray_S23reg_gff_1_SFF_0_n2), .A0_f (new_AGEMA_signal_6922), .A1_t (new_AGEMA_signal_6923), .A1_f (new_AGEMA_signal_6924), .B0_t (KeyArray_S23reg_gff_1_SFF_0_n1), .B0_f (new_AGEMA_signal_6919), .B1_t (new_AGEMA_signal_6920), .B1_f (new_AGEMA_signal_6921), .Z0_t (KeyArray_outS23ser[0]), .Z0_f (new_AGEMA_signal_3613), .Z1_t (new_AGEMA_signal_3614), .Z1_f (new_AGEMA_signal_3615) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_0_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS23ser[0]), .B0_f (new_AGEMA_signal_3613), .B1_t (new_AGEMA_signal_3614), .B1_f (new_AGEMA_signal_3615), .Z0_t (KeyArray_S23reg_gff_1_SFF_0_n1), .Z0_f (new_AGEMA_signal_6919), .Z1_t (new_AGEMA_signal_6920), .Z1_f (new_AGEMA_signal_6921) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_0_U1 ( .A0_t (KeyArray_S23reg_gff_1_SFF_0_QD), .A0_f (new_AGEMA_signal_4941), .A1_t (new_AGEMA_signal_4942), .A1_f (new_AGEMA_signal_4943), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S23reg_gff_1_SFF_0_n2), .Z0_f (new_AGEMA_signal_6922), .Z1_t (new_AGEMA_signal_6923), .Z1_f (new_AGEMA_signal_6924) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS30ser[0]), .A0_f (new_AGEMA_signal_3661), .A1_t (new_AGEMA_signal_3662), .A1_f (new_AGEMA_signal_3663), .B0_t (KeyArray_outS33ser[0]), .B0_f (new_AGEMA_signal_3805), .B1_t (new_AGEMA_signal_3806), .B1_f (new_AGEMA_signal_3807), .Z0_t (KeyArray_S23reg_gff_1_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_3808), .Z1_t (new_AGEMA_signal_3809), .Z1_f (new_AGEMA_signal_3810) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S23reg_gff_1_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_3808), .B1_t (new_AGEMA_signal_3809), .B1_f (new_AGEMA_signal_3810), .Z0_t (KeyArray_S23reg_gff_1_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_4451), .Z1_t (new_AGEMA_signal_4452), .Z1_f (new_AGEMA_signal_4453) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S23reg_gff_1_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_4451), .A1_t (new_AGEMA_signal_4452), .A1_f (new_AGEMA_signal_4453), .B0_t (KeyArray_outS30ser[0]), .B0_f (new_AGEMA_signal_3661), .B1_t (new_AGEMA_signal_3662), .B1_f (new_AGEMA_signal_3663), .Z0_t (KeyArray_S23reg_gff_1_SFF_0_QD), .Z0_f (new_AGEMA_signal_4941), .Z1_t (new_AGEMA_signal_4942), .Z1_f (new_AGEMA_signal_4943) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S23reg_gff_1_SFF_1_U3 ( .A0_t (KeyArray_S23reg_gff_1_SFF_1_n2), .A0_f (new_AGEMA_signal_6928), .A1_t (new_AGEMA_signal_6929), .A1_f (new_AGEMA_signal_6930), .B0_t (KeyArray_S23reg_gff_1_SFF_1_n1), .B0_f (new_AGEMA_signal_6925), .B1_t (new_AGEMA_signal_6926), .B1_f (new_AGEMA_signal_6927), .Z0_t (KeyArray_outS23ser[1]), .Z0_f (new_AGEMA_signal_3619), .Z1_t (new_AGEMA_signal_3620), .Z1_f (new_AGEMA_signal_3621) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_1_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS23ser[1]), .B0_f (new_AGEMA_signal_3619), .B1_t (new_AGEMA_signal_3620), .B1_f (new_AGEMA_signal_3621), .Z0_t (KeyArray_S23reg_gff_1_SFF_1_n1), .Z0_f (new_AGEMA_signal_6925), .Z1_t (new_AGEMA_signal_6926), .Z1_f (new_AGEMA_signal_6927) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_1_U1 ( .A0_t (KeyArray_S23reg_gff_1_SFF_1_QD), .A0_f (new_AGEMA_signal_4944), .A1_t (new_AGEMA_signal_4945), .A1_f (new_AGEMA_signal_4946), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S23reg_gff_1_SFF_1_n2), .Z0_f (new_AGEMA_signal_6928), .Z1_t (new_AGEMA_signal_6929), .Z1_f (new_AGEMA_signal_6930) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS30ser[1]), .A0_f (new_AGEMA_signal_3667), .A1_t (new_AGEMA_signal_3668), .A1_f (new_AGEMA_signal_3669), .B0_t (KeyArray_outS33ser[1]), .B0_f (new_AGEMA_signal_3811), .B1_t (new_AGEMA_signal_3812), .B1_f (new_AGEMA_signal_3813), .Z0_t (KeyArray_S23reg_gff_1_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_3814), .Z1_t (new_AGEMA_signal_3815), .Z1_f (new_AGEMA_signal_3816) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S23reg_gff_1_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_3814), .B1_t (new_AGEMA_signal_3815), .B1_f (new_AGEMA_signal_3816), .Z0_t (KeyArray_S23reg_gff_1_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_4454), .Z1_t (new_AGEMA_signal_4455), .Z1_f (new_AGEMA_signal_4456) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S23reg_gff_1_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_4454), .A1_t (new_AGEMA_signal_4455), .A1_f (new_AGEMA_signal_4456), .B0_t (KeyArray_outS30ser[1]), .B0_f (new_AGEMA_signal_3667), .B1_t (new_AGEMA_signal_3668), .B1_f (new_AGEMA_signal_3669), .Z0_t (KeyArray_S23reg_gff_1_SFF_1_QD), .Z0_f (new_AGEMA_signal_4944), .Z1_t (new_AGEMA_signal_4945), .Z1_f (new_AGEMA_signal_4946) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S23reg_gff_1_SFF_2_U3 ( .A0_t (KeyArray_S23reg_gff_1_SFF_2_n2), .A0_f (new_AGEMA_signal_6934), .A1_t (new_AGEMA_signal_6935), .A1_f (new_AGEMA_signal_6936), .B0_t (KeyArray_S23reg_gff_1_SFF_2_n1), .B0_f (new_AGEMA_signal_6931), .B1_t (new_AGEMA_signal_6932), .B1_f (new_AGEMA_signal_6933), .Z0_t (KeyArray_outS23ser[2]), .Z0_f (new_AGEMA_signal_3625), .Z1_t (new_AGEMA_signal_3626), .Z1_f (new_AGEMA_signal_3627) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_2_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS23ser[2]), .B0_f (new_AGEMA_signal_3625), .B1_t (new_AGEMA_signal_3626), .B1_f (new_AGEMA_signal_3627), .Z0_t (KeyArray_S23reg_gff_1_SFF_2_n1), .Z0_f (new_AGEMA_signal_6931), .Z1_t (new_AGEMA_signal_6932), .Z1_f (new_AGEMA_signal_6933) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_2_U1 ( .A0_t (KeyArray_S23reg_gff_1_SFF_2_QD), .A0_f (new_AGEMA_signal_4947), .A1_t (new_AGEMA_signal_4948), .A1_f (new_AGEMA_signal_4949), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S23reg_gff_1_SFF_2_n2), .Z0_f (new_AGEMA_signal_6934), .Z1_t (new_AGEMA_signal_6935), .Z1_f (new_AGEMA_signal_6936) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS30ser[2]), .A0_f (new_AGEMA_signal_3673), .A1_t (new_AGEMA_signal_3674), .A1_f (new_AGEMA_signal_3675), .B0_t (KeyArray_outS33ser[2]), .B0_f (new_AGEMA_signal_3817), .B1_t (new_AGEMA_signal_3818), .B1_f (new_AGEMA_signal_3819), .Z0_t (KeyArray_S23reg_gff_1_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_3820), .Z1_t (new_AGEMA_signal_3821), .Z1_f (new_AGEMA_signal_3822) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S23reg_gff_1_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_3820), .B1_t (new_AGEMA_signal_3821), .B1_f (new_AGEMA_signal_3822), .Z0_t (KeyArray_S23reg_gff_1_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_4457), .Z1_t (new_AGEMA_signal_4458), .Z1_f (new_AGEMA_signal_4459) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S23reg_gff_1_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_4457), .A1_t (new_AGEMA_signal_4458), .A1_f (new_AGEMA_signal_4459), .B0_t (KeyArray_outS30ser[2]), .B0_f (new_AGEMA_signal_3673), .B1_t (new_AGEMA_signal_3674), .B1_f (new_AGEMA_signal_3675), .Z0_t (KeyArray_S23reg_gff_1_SFF_2_QD), .Z0_f (new_AGEMA_signal_4947), .Z1_t (new_AGEMA_signal_4948), .Z1_f (new_AGEMA_signal_4949) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S23reg_gff_1_SFF_3_U3 ( .A0_t (KeyArray_S23reg_gff_1_SFF_3_n2), .A0_f (new_AGEMA_signal_6940), .A1_t (new_AGEMA_signal_6941), .A1_f (new_AGEMA_signal_6942), .B0_t (KeyArray_S23reg_gff_1_SFF_3_n1), .B0_f (new_AGEMA_signal_6937), .B1_t (new_AGEMA_signal_6938), .B1_f (new_AGEMA_signal_6939), .Z0_t (KeyArray_outS23ser[3]), .Z0_f (new_AGEMA_signal_3631), .Z1_t (new_AGEMA_signal_3632), .Z1_f (new_AGEMA_signal_3633) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_3_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS23ser[3]), .B0_f (new_AGEMA_signal_3631), .B1_t (new_AGEMA_signal_3632), .B1_f (new_AGEMA_signal_3633), .Z0_t (KeyArray_S23reg_gff_1_SFF_3_n1), .Z0_f (new_AGEMA_signal_6937), .Z1_t (new_AGEMA_signal_6938), .Z1_f (new_AGEMA_signal_6939) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_3_U1 ( .A0_t (KeyArray_S23reg_gff_1_SFF_3_QD), .A0_f (new_AGEMA_signal_4950), .A1_t (new_AGEMA_signal_4951), .A1_f (new_AGEMA_signal_4952), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S23reg_gff_1_SFF_3_n2), .Z0_f (new_AGEMA_signal_6940), .Z1_t (new_AGEMA_signal_6941), .Z1_f (new_AGEMA_signal_6942) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS30ser[3]), .A0_f (new_AGEMA_signal_3679), .A1_t (new_AGEMA_signal_3680), .A1_f (new_AGEMA_signal_3681), .B0_t (KeyArray_outS33ser[3]), .B0_f (new_AGEMA_signal_3823), .B1_t (new_AGEMA_signal_3824), .B1_f (new_AGEMA_signal_3825), .Z0_t (KeyArray_S23reg_gff_1_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_3826), .Z1_t (new_AGEMA_signal_3827), .Z1_f (new_AGEMA_signal_3828) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S23reg_gff_1_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_3826), .B1_t (new_AGEMA_signal_3827), .B1_f (new_AGEMA_signal_3828), .Z0_t (KeyArray_S23reg_gff_1_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_4460), .Z1_t (new_AGEMA_signal_4461), .Z1_f (new_AGEMA_signal_4462) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S23reg_gff_1_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_4460), .A1_t (new_AGEMA_signal_4461), .A1_f (new_AGEMA_signal_4462), .B0_t (KeyArray_outS30ser[3]), .B0_f (new_AGEMA_signal_3679), .B1_t (new_AGEMA_signal_3680), .B1_f (new_AGEMA_signal_3681), .Z0_t (KeyArray_S23reg_gff_1_SFF_3_QD), .Z0_f (new_AGEMA_signal_4950), .Z1_t (new_AGEMA_signal_4951), .Z1_f (new_AGEMA_signal_4952) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S23reg_gff_1_SFF_4_U3 ( .A0_t (KeyArray_S23reg_gff_1_SFF_4_n2), .A0_f (new_AGEMA_signal_6946), .A1_t (new_AGEMA_signal_6947), .A1_f (new_AGEMA_signal_6948), .B0_t (KeyArray_S23reg_gff_1_SFF_4_n1), .B0_f (new_AGEMA_signal_6943), .B1_t (new_AGEMA_signal_6944), .B1_f (new_AGEMA_signal_6945), .Z0_t (KeyArray_outS23ser[4]), .Z0_f (new_AGEMA_signal_3637), .Z1_t (new_AGEMA_signal_3638), .Z1_f (new_AGEMA_signal_3639) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_4_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS23ser[4]), .B0_f (new_AGEMA_signal_3637), .B1_t (new_AGEMA_signal_3638), .B1_f (new_AGEMA_signal_3639), .Z0_t (KeyArray_S23reg_gff_1_SFF_4_n1), .Z0_f (new_AGEMA_signal_6943), .Z1_t (new_AGEMA_signal_6944), .Z1_f (new_AGEMA_signal_6945) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_4_U1 ( .A0_t (KeyArray_S23reg_gff_1_SFF_4_QD), .A0_f (new_AGEMA_signal_4953), .A1_t (new_AGEMA_signal_4954), .A1_f (new_AGEMA_signal_4955), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S23reg_gff_1_SFF_4_n2), .Z0_f (new_AGEMA_signal_6946), .Z1_t (new_AGEMA_signal_6947), .Z1_f (new_AGEMA_signal_6948) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS30ser[4]), .A0_f (new_AGEMA_signal_3685), .A1_t (new_AGEMA_signal_3686), .A1_f (new_AGEMA_signal_3687), .B0_t (KeyArray_outS33ser[4]), .B0_f (new_AGEMA_signal_3829), .B1_t (new_AGEMA_signal_3830), .B1_f (new_AGEMA_signal_3831), .Z0_t (KeyArray_S23reg_gff_1_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_3832), .Z1_t (new_AGEMA_signal_3833), .Z1_f (new_AGEMA_signal_3834) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S23reg_gff_1_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_3832), .B1_t (new_AGEMA_signal_3833), .B1_f (new_AGEMA_signal_3834), .Z0_t (KeyArray_S23reg_gff_1_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_4463), .Z1_t (new_AGEMA_signal_4464), .Z1_f (new_AGEMA_signal_4465) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S23reg_gff_1_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_4463), .A1_t (new_AGEMA_signal_4464), .A1_f (new_AGEMA_signal_4465), .B0_t (KeyArray_outS30ser[4]), .B0_f (new_AGEMA_signal_3685), .B1_t (new_AGEMA_signal_3686), .B1_f (new_AGEMA_signal_3687), .Z0_t (KeyArray_S23reg_gff_1_SFF_4_QD), .Z0_f (new_AGEMA_signal_4953), .Z1_t (new_AGEMA_signal_4954), .Z1_f (new_AGEMA_signal_4955) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S23reg_gff_1_SFF_5_U3 ( .A0_t (KeyArray_S23reg_gff_1_SFF_5_n2), .A0_f (new_AGEMA_signal_6952), .A1_t (new_AGEMA_signal_6953), .A1_f (new_AGEMA_signal_6954), .B0_t (KeyArray_S23reg_gff_1_SFF_5_n1), .B0_f (new_AGEMA_signal_6949), .B1_t (new_AGEMA_signal_6950), .B1_f (new_AGEMA_signal_6951), .Z0_t (KeyArray_outS23ser[5]), .Z0_f (new_AGEMA_signal_3643), .Z1_t (new_AGEMA_signal_3644), .Z1_f (new_AGEMA_signal_3645) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_5_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS23ser[5]), .B0_f (new_AGEMA_signal_3643), .B1_t (new_AGEMA_signal_3644), .B1_f (new_AGEMA_signal_3645), .Z0_t (KeyArray_S23reg_gff_1_SFF_5_n1), .Z0_f (new_AGEMA_signal_6949), .Z1_t (new_AGEMA_signal_6950), .Z1_f (new_AGEMA_signal_6951) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_5_U1 ( .A0_t (KeyArray_S23reg_gff_1_SFF_5_QD), .A0_f (new_AGEMA_signal_4956), .A1_t (new_AGEMA_signal_4957), .A1_f (new_AGEMA_signal_4958), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S23reg_gff_1_SFF_5_n2), .Z0_f (new_AGEMA_signal_6952), .Z1_t (new_AGEMA_signal_6953), .Z1_f (new_AGEMA_signal_6954) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS30ser[5]), .A0_f (new_AGEMA_signal_3691), .A1_t (new_AGEMA_signal_3692), .A1_f (new_AGEMA_signal_3693), .B0_t (KeyArray_outS33ser[5]), .B0_f (new_AGEMA_signal_3835), .B1_t (new_AGEMA_signal_3836), .B1_f (new_AGEMA_signal_3837), .Z0_t (KeyArray_S23reg_gff_1_SFF_5_MUXInst_X), .Z0_f (new_AGEMA_signal_3838), .Z1_t (new_AGEMA_signal_3839), .Z1_f (new_AGEMA_signal_3840) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S23reg_gff_1_SFF_5_MUXInst_X), .B0_f (new_AGEMA_signal_3838), .B1_t (new_AGEMA_signal_3839), .B1_f (new_AGEMA_signal_3840), .Z0_t (KeyArray_S23reg_gff_1_SFF_5_MUXInst_Y), .Z0_f (new_AGEMA_signal_4466), .Z1_t (new_AGEMA_signal_4467), .Z1_f (new_AGEMA_signal_4468) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S23reg_gff_1_SFF_5_MUXInst_Y), .A0_f (new_AGEMA_signal_4466), .A1_t (new_AGEMA_signal_4467), .A1_f (new_AGEMA_signal_4468), .B0_t (KeyArray_outS30ser[5]), .B0_f (new_AGEMA_signal_3691), .B1_t (new_AGEMA_signal_3692), .B1_f (new_AGEMA_signal_3693), .Z0_t (KeyArray_S23reg_gff_1_SFF_5_QD), .Z0_f (new_AGEMA_signal_4956), .Z1_t (new_AGEMA_signal_4957), .Z1_f (new_AGEMA_signal_4958) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S23reg_gff_1_SFF_6_U3 ( .A0_t (KeyArray_S23reg_gff_1_SFF_6_n2), .A0_f (new_AGEMA_signal_6958), .A1_t (new_AGEMA_signal_6959), .A1_f (new_AGEMA_signal_6960), .B0_t (KeyArray_S23reg_gff_1_SFF_6_n1), .B0_f (new_AGEMA_signal_6955), .B1_t (new_AGEMA_signal_6956), .B1_f (new_AGEMA_signal_6957), .Z0_t (KeyArray_outS23ser[6]), .Z0_f (new_AGEMA_signal_3649), .Z1_t (new_AGEMA_signal_3650), .Z1_f (new_AGEMA_signal_3651) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_6_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS23ser[6]), .B0_f (new_AGEMA_signal_3649), .B1_t (new_AGEMA_signal_3650), .B1_f (new_AGEMA_signal_3651), .Z0_t (KeyArray_S23reg_gff_1_SFF_6_n1), .Z0_f (new_AGEMA_signal_6955), .Z1_t (new_AGEMA_signal_6956), .Z1_f (new_AGEMA_signal_6957) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_6_U1 ( .A0_t (KeyArray_S23reg_gff_1_SFF_6_QD), .A0_f (new_AGEMA_signal_4959), .A1_t (new_AGEMA_signal_4960), .A1_f (new_AGEMA_signal_4961), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S23reg_gff_1_SFF_6_n2), .Z0_f (new_AGEMA_signal_6958), .Z1_t (new_AGEMA_signal_6959), .Z1_f (new_AGEMA_signal_6960) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS30ser[6]), .A0_f (new_AGEMA_signal_3697), .A1_t (new_AGEMA_signal_3698), .A1_f (new_AGEMA_signal_3699), .B0_t (KeyArray_outS33ser[6]), .B0_f (new_AGEMA_signal_3841), .B1_t (new_AGEMA_signal_3842), .B1_f (new_AGEMA_signal_3843), .Z0_t (KeyArray_S23reg_gff_1_SFF_6_MUXInst_X), .Z0_f (new_AGEMA_signal_3844), .Z1_t (new_AGEMA_signal_3845), .Z1_f (new_AGEMA_signal_3846) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S23reg_gff_1_SFF_6_MUXInst_X), .B0_f (new_AGEMA_signal_3844), .B1_t (new_AGEMA_signal_3845), .B1_f (new_AGEMA_signal_3846), .Z0_t (KeyArray_S23reg_gff_1_SFF_6_MUXInst_Y), .Z0_f (new_AGEMA_signal_4469), .Z1_t (new_AGEMA_signal_4470), .Z1_f (new_AGEMA_signal_4471) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S23reg_gff_1_SFF_6_MUXInst_Y), .A0_f (new_AGEMA_signal_4469), .A1_t (new_AGEMA_signal_4470), .A1_f (new_AGEMA_signal_4471), .B0_t (KeyArray_outS30ser[6]), .B0_f (new_AGEMA_signal_3697), .B1_t (new_AGEMA_signal_3698), .B1_f (new_AGEMA_signal_3699), .Z0_t (KeyArray_S23reg_gff_1_SFF_6_QD), .Z0_f (new_AGEMA_signal_4959), .Z1_t (new_AGEMA_signal_4960), .Z1_f (new_AGEMA_signal_4961) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S23reg_gff_1_SFF_7_U3 ( .A0_t (KeyArray_S23reg_gff_1_SFF_7_n2), .A0_f (new_AGEMA_signal_6964), .A1_t (new_AGEMA_signal_6965), .A1_f (new_AGEMA_signal_6966), .B0_t (KeyArray_S23reg_gff_1_SFF_7_n1), .B0_f (new_AGEMA_signal_6961), .B1_t (new_AGEMA_signal_6962), .B1_f (new_AGEMA_signal_6963), .Z0_t (KeyArray_outS23ser[7]), .Z0_f (new_AGEMA_signal_3655), .Z1_t (new_AGEMA_signal_3656), .Z1_f (new_AGEMA_signal_3657) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_7_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS23ser[7]), .B0_f (new_AGEMA_signal_3655), .B1_t (new_AGEMA_signal_3656), .B1_f (new_AGEMA_signal_3657), .Z0_t (KeyArray_S23reg_gff_1_SFF_7_n1), .Z0_f (new_AGEMA_signal_6961), .Z1_t (new_AGEMA_signal_6962), .Z1_f (new_AGEMA_signal_6963) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_7_U1 ( .A0_t (KeyArray_S23reg_gff_1_SFF_7_QD), .A0_f (new_AGEMA_signal_4962), .A1_t (new_AGEMA_signal_4963), .A1_f (new_AGEMA_signal_4964), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S23reg_gff_1_SFF_7_n2), .Z0_f (new_AGEMA_signal_6964), .Z1_t (new_AGEMA_signal_6965), .Z1_f (new_AGEMA_signal_6966) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS30ser[7]), .A0_f (new_AGEMA_signal_3703), .A1_t (new_AGEMA_signal_3704), .A1_f (new_AGEMA_signal_3705), .B0_t (KeyArray_outS33ser[7]), .B0_f (new_AGEMA_signal_3847), .B1_t (new_AGEMA_signal_3848), .B1_f (new_AGEMA_signal_3849), .Z0_t (KeyArray_S23reg_gff_1_SFF_7_MUXInst_X), .Z0_f (new_AGEMA_signal_3850), .Z1_t (new_AGEMA_signal_3851), .Z1_f (new_AGEMA_signal_3852) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S23reg_gff_1_SFF_7_MUXInst_X), .B0_f (new_AGEMA_signal_3850), .B1_t (new_AGEMA_signal_3851), .B1_f (new_AGEMA_signal_3852), .Z0_t (KeyArray_S23reg_gff_1_SFF_7_MUXInst_Y), .Z0_f (new_AGEMA_signal_4472), .Z1_t (new_AGEMA_signal_4473), .Z1_f (new_AGEMA_signal_4474) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S23reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S23reg_gff_1_SFF_7_MUXInst_Y), .A0_f (new_AGEMA_signal_4472), .A1_t (new_AGEMA_signal_4473), .A1_f (new_AGEMA_signal_4474), .B0_t (KeyArray_outS30ser[7]), .B0_f (new_AGEMA_signal_3703), .B1_t (new_AGEMA_signal_3704), .B1_f (new_AGEMA_signal_3705), .Z0_t (KeyArray_S23reg_gff_1_SFF_7_QD), .Z0_f (new_AGEMA_signal_4962), .Z1_t (new_AGEMA_signal_4963), .Z1_f (new_AGEMA_signal_4964) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S30reg_gff_1_SFF_0_U3 ( .A0_t (KeyArray_S30reg_gff_1_SFF_0_n2), .A0_f (new_AGEMA_signal_7748), .A1_t (new_AGEMA_signal_7749), .A1_f (new_AGEMA_signal_7750), .B0_t (KeyArray_S30reg_gff_1_SFF_0_n1), .B0_f (new_AGEMA_signal_6967), .B1_t (new_AGEMA_signal_6968), .B1_f (new_AGEMA_signal_6969), .Z0_t (KeyArray_outS30ser[0]), .Z0_f (new_AGEMA_signal_3661), .Z1_t (new_AGEMA_signal_3662), .Z1_f (new_AGEMA_signal_3663) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_0_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS30ser[0]), .B0_f (new_AGEMA_signal_3661), .B1_t (new_AGEMA_signal_3662), .B1_f (new_AGEMA_signal_3663), .Z0_t (KeyArray_S30reg_gff_1_SFF_0_n1), .Z0_f (new_AGEMA_signal_6967), .Z1_t (new_AGEMA_signal_6968), .Z1_f (new_AGEMA_signal_6969) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_0_U1 ( .A0_t (KeyArray_S30reg_gff_1_SFF_0_QD), .A0_f (new_AGEMA_signal_7700), .A1_t (new_AGEMA_signal_7701), .A1_f (new_AGEMA_signal_7702), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S30reg_gff_1_SFF_0_n2), .Z0_f (new_AGEMA_signal_7748), .Z1_t (new_AGEMA_signal_7749), .Z1_f (new_AGEMA_signal_7750) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS31ser[0]), .A0_f (new_AGEMA_signal_3709), .A1_t (new_AGEMA_signal_3710), .A1_f (new_AGEMA_signal_3711), .B0_t (KeyArray_inS30par[0]), .B0_f (new_AGEMA_signal_7577), .B1_t (new_AGEMA_signal_7578), .B1_f (new_AGEMA_signal_7579), .Z0_t (KeyArray_S30reg_gff_1_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_7625), .Z1_t (new_AGEMA_signal_7626), .Z1_f (new_AGEMA_signal_7627) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S30reg_gff_1_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_7625), .B1_t (new_AGEMA_signal_7626), .B1_f (new_AGEMA_signal_7627), .Z0_t (KeyArray_S30reg_gff_1_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_7652), .Z1_t (new_AGEMA_signal_7653), .Z1_f (new_AGEMA_signal_7654) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S30reg_gff_1_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_7652), .A1_t (new_AGEMA_signal_7653), .A1_f (new_AGEMA_signal_7654), .B0_t (KeyArray_outS31ser[0]), .B0_f (new_AGEMA_signal_3709), .B1_t (new_AGEMA_signal_3710), .B1_f (new_AGEMA_signal_3711), .Z0_t (KeyArray_S30reg_gff_1_SFF_0_QD), .Z0_f (new_AGEMA_signal_7700), .Z1_t (new_AGEMA_signal_7701), .Z1_f (new_AGEMA_signal_7702) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S30reg_gff_1_SFF_1_U3 ( .A0_t (KeyArray_S30reg_gff_1_SFF_1_n2), .A0_f (new_AGEMA_signal_7799), .A1_t (new_AGEMA_signal_7800), .A1_f (new_AGEMA_signal_7801), .B0_t (KeyArray_S30reg_gff_1_SFF_1_n1), .B0_f (new_AGEMA_signal_6970), .B1_t (new_AGEMA_signal_6971), .B1_f (new_AGEMA_signal_6972), .Z0_t (KeyArray_outS30ser[1]), .Z0_f (new_AGEMA_signal_3667), .Z1_t (new_AGEMA_signal_3668), .Z1_f (new_AGEMA_signal_3669) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_1_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS30ser[1]), .B0_f (new_AGEMA_signal_3667), .B1_t (new_AGEMA_signal_3668), .B1_f (new_AGEMA_signal_3669), .Z0_t (KeyArray_S30reg_gff_1_SFF_1_n1), .Z0_f (new_AGEMA_signal_6970), .Z1_t (new_AGEMA_signal_6971), .Z1_f (new_AGEMA_signal_6972) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_1_U1 ( .A0_t (KeyArray_S30reg_gff_1_SFF_1_QD), .A0_f (new_AGEMA_signal_7751), .A1_t (new_AGEMA_signal_7752), .A1_f (new_AGEMA_signal_7753), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S30reg_gff_1_SFF_1_n2), .Z0_f (new_AGEMA_signal_7799), .Z1_t (new_AGEMA_signal_7800), .Z1_f (new_AGEMA_signal_7801) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS31ser[1]), .A0_f (new_AGEMA_signal_3715), .A1_t (new_AGEMA_signal_3716), .A1_f (new_AGEMA_signal_3717), .B0_t (KeyArray_inS30par[1]), .B0_f (new_AGEMA_signal_7622), .B1_t (new_AGEMA_signal_7623), .B1_f (new_AGEMA_signal_7624), .Z0_t (KeyArray_S30reg_gff_1_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_7655), .Z1_t (new_AGEMA_signal_7656), .Z1_f (new_AGEMA_signal_7657) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S30reg_gff_1_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_7655), .B1_t (new_AGEMA_signal_7656), .B1_f (new_AGEMA_signal_7657), .Z0_t (KeyArray_S30reg_gff_1_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_7703), .Z1_t (new_AGEMA_signal_7704), .Z1_f (new_AGEMA_signal_7705) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S30reg_gff_1_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_7703), .A1_t (new_AGEMA_signal_7704), .A1_f (new_AGEMA_signal_7705), .B0_t (KeyArray_outS31ser[1]), .B0_f (new_AGEMA_signal_3715), .B1_t (new_AGEMA_signal_3716), .B1_f (new_AGEMA_signal_3717), .Z0_t (KeyArray_S30reg_gff_1_SFF_1_QD), .Z0_f (new_AGEMA_signal_7751), .Z1_t (new_AGEMA_signal_7752), .Z1_f (new_AGEMA_signal_7753) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S30reg_gff_1_SFF_2_U3 ( .A0_t (KeyArray_S30reg_gff_1_SFF_2_n2), .A0_f (new_AGEMA_signal_7802), .A1_t (new_AGEMA_signal_7803), .A1_f (new_AGEMA_signal_7804), .B0_t (KeyArray_S30reg_gff_1_SFF_2_n1), .B0_f (new_AGEMA_signal_6973), .B1_t (new_AGEMA_signal_6974), .B1_f (new_AGEMA_signal_6975), .Z0_t (KeyArray_outS30ser[2]), .Z0_f (new_AGEMA_signal_3673), .Z1_t (new_AGEMA_signal_3674), .Z1_f (new_AGEMA_signal_3675) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_2_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS30ser[2]), .B0_f (new_AGEMA_signal_3673), .B1_t (new_AGEMA_signal_3674), .B1_f (new_AGEMA_signal_3675), .Z0_t (KeyArray_S30reg_gff_1_SFF_2_n1), .Z0_f (new_AGEMA_signal_6973), .Z1_t (new_AGEMA_signal_6974), .Z1_f (new_AGEMA_signal_6975) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_2_U1 ( .A0_t (KeyArray_S30reg_gff_1_SFF_2_QD), .A0_f (new_AGEMA_signal_7754), .A1_t (new_AGEMA_signal_7755), .A1_f (new_AGEMA_signal_7756), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S30reg_gff_1_SFF_2_n2), .Z0_f (new_AGEMA_signal_7802), .Z1_t (new_AGEMA_signal_7803), .Z1_f (new_AGEMA_signal_7804) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS31ser[2]), .A0_f (new_AGEMA_signal_3721), .A1_t (new_AGEMA_signal_3722), .A1_f (new_AGEMA_signal_3723), .B0_t (KeyArray_inS30par[2]), .B0_f (new_AGEMA_signal_7619), .B1_t (new_AGEMA_signal_7620), .B1_f (new_AGEMA_signal_7621), .Z0_t (KeyArray_S30reg_gff_1_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_7658), .Z1_t (new_AGEMA_signal_7659), .Z1_f (new_AGEMA_signal_7660) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S30reg_gff_1_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_7658), .B1_t (new_AGEMA_signal_7659), .B1_f (new_AGEMA_signal_7660), .Z0_t (KeyArray_S30reg_gff_1_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_7706), .Z1_t (new_AGEMA_signal_7707), .Z1_f (new_AGEMA_signal_7708) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S30reg_gff_1_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_7706), .A1_t (new_AGEMA_signal_7707), .A1_f (new_AGEMA_signal_7708), .B0_t (KeyArray_outS31ser[2]), .B0_f (new_AGEMA_signal_3721), .B1_t (new_AGEMA_signal_3722), .B1_f (new_AGEMA_signal_3723), .Z0_t (KeyArray_S30reg_gff_1_SFF_2_QD), .Z0_f (new_AGEMA_signal_7754), .Z1_t (new_AGEMA_signal_7755), .Z1_f (new_AGEMA_signal_7756) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S30reg_gff_1_SFF_3_U3 ( .A0_t (KeyArray_S30reg_gff_1_SFF_3_n2), .A0_f (new_AGEMA_signal_7805), .A1_t (new_AGEMA_signal_7806), .A1_f (new_AGEMA_signal_7807), .B0_t (KeyArray_S30reg_gff_1_SFF_3_n1), .B0_f (new_AGEMA_signal_6976), .B1_t (new_AGEMA_signal_6977), .B1_f (new_AGEMA_signal_6978), .Z0_t (KeyArray_outS30ser[3]), .Z0_f (new_AGEMA_signal_3679), .Z1_t (new_AGEMA_signal_3680), .Z1_f (new_AGEMA_signal_3681) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_3_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS30ser[3]), .B0_f (new_AGEMA_signal_3679), .B1_t (new_AGEMA_signal_3680), .B1_f (new_AGEMA_signal_3681), .Z0_t (KeyArray_S30reg_gff_1_SFF_3_n1), .Z0_f (new_AGEMA_signal_6976), .Z1_t (new_AGEMA_signal_6977), .Z1_f (new_AGEMA_signal_6978) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_3_U1 ( .A0_t (KeyArray_S30reg_gff_1_SFF_3_QD), .A0_f (new_AGEMA_signal_7757), .A1_t (new_AGEMA_signal_7758), .A1_f (new_AGEMA_signal_7759), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S30reg_gff_1_SFF_3_n2), .Z0_f (new_AGEMA_signal_7805), .Z1_t (new_AGEMA_signal_7806), .Z1_f (new_AGEMA_signal_7807) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS31ser[3]), .A0_f (new_AGEMA_signal_3727), .A1_t (new_AGEMA_signal_3728), .A1_f (new_AGEMA_signal_3729), .B0_t (KeyArray_inS30par[3]), .B0_f (new_AGEMA_signal_7616), .B1_t (new_AGEMA_signal_7617), .B1_f (new_AGEMA_signal_7618), .Z0_t (KeyArray_S30reg_gff_1_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_7661), .Z1_t (new_AGEMA_signal_7662), .Z1_f (new_AGEMA_signal_7663) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S30reg_gff_1_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_7661), .B1_t (new_AGEMA_signal_7662), .B1_f (new_AGEMA_signal_7663), .Z0_t (KeyArray_S30reg_gff_1_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_7709), .Z1_t (new_AGEMA_signal_7710), .Z1_f (new_AGEMA_signal_7711) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S30reg_gff_1_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_7709), .A1_t (new_AGEMA_signal_7710), .A1_f (new_AGEMA_signal_7711), .B0_t (KeyArray_outS31ser[3]), .B0_f (new_AGEMA_signal_3727), .B1_t (new_AGEMA_signal_3728), .B1_f (new_AGEMA_signal_3729), .Z0_t (KeyArray_S30reg_gff_1_SFF_3_QD), .Z0_f (new_AGEMA_signal_7757), .Z1_t (new_AGEMA_signal_7758), .Z1_f (new_AGEMA_signal_7759) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S30reg_gff_1_SFF_4_U3 ( .A0_t (KeyArray_S30reg_gff_1_SFF_4_n2), .A0_f (new_AGEMA_signal_7808), .A1_t (new_AGEMA_signal_7809), .A1_f (new_AGEMA_signal_7810), .B0_t (KeyArray_S30reg_gff_1_SFF_4_n1), .B0_f (new_AGEMA_signal_6979), .B1_t (new_AGEMA_signal_6980), .B1_f (new_AGEMA_signal_6981), .Z0_t (KeyArray_outS30ser[4]), .Z0_f (new_AGEMA_signal_3685), .Z1_t (new_AGEMA_signal_3686), .Z1_f (new_AGEMA_signal_3687) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_4_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS30ser[4]), .B0_f (new_AGEMA_signal_3685), .B1_t (new_AGEMA_signal_3686), .B1_f (new_AGEMA_signal_3687), .Z0_t (KeyArray_S30reg_gff_1_SFF_4_n1), .Z0_f (new_AGEMA_signal_6979), .Z1_t (new_AGEMA_signal_6980), .Z1_f (new_AGEMA_signal_6981) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_4_U1 ( .A0_t (KeyArray_S30reg_gff_1_SFF_4_QD), .A0_f (new_AGEMA_signal_7760), .A1_t (new_AGEMA_signal_7761), .A1_f (new_AGEMA_signal_7762), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S30reg_gff_1_SFF_4_n2), .Z0_f (new_AGEMA_signal_7808), .Z1_t (new_AGEMA_signal_7809), .Z1_f (new_AGEMA_signal_7810) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS31ser[4]), .A0_f (new_AGEMA_signal_3733), .A1_t (new_AGEMA_signal_3734), .A1_f (new_AGEMA_signal_3735), .B0_t (KeyArray_inS30par[4]), .B0_f (new_AGEMA_signal_7613), .B1_t (new_AGEMA_signal_7614), .B1_f (new_AGEMA_signal_7615), .Z0_t (KeyArray_S30reg_gff_1_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_7664), .Z1_t (new_AGEMA_signal_7665), .Z1_f (new_AGEMA_signal_7666) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S30reg_gff_1_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_7664), .B1_t (new_AGEMA_signal_7665), .B1_f (new_AGEMA_signal_7666), .Z0_t (KeyArray_S30reg_gff_1_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_7712), .Z1_t (new_AGEMA_signal_7713), .Z1_f (new_AGEMA_signal_7714) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S30reg_gff_1_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_7712), .A1_t (new_AGEMA_signal_7713), .A1_f (new_AGEMA_signal_7714), .B0_t (KeyArray_outS31ser[4]), .B0_f (new_AGEMA_signal_3733), .B1_t (new_AGEMA_signal_3734), .B1_f (new_AGEMA_signal_3735), .Z0_t (KeyArray_S30reg_gff_1_SFF_4_QD), .Z0_f (new_AGEMA_signal_7760), .Z1_t (new_AGEMA_signal_7761), .Z1_f (new_AGEMA_signal_7762) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S30reg_gff_1_SFF_5_U3 ( .A0_t (KeyArray_S30reg_gff_1_SFF_5_n2), .A0_f (new_AGEMA_signal_7811), .A1_t (new_AGEMA_signal_7812), .A1_f (new_AGEMA_signal_7813), .B0_t (KeyArray_S30reg_gff_1_SFF_5_n1), .B0_f (new_AGEMA_signal_6982), .B1_t (new_AGEMA_signal_6983), .B1_f (new_AGEMA_signal_6984), .Z0_t (KeyArray_outS30ser[5]), .Z0_f (new_AGEMA_signal_3691), .Z1_t (new_AGEMA_signal_3692), .Z1_f (new_AGEMA_signal_3693) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_5_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS30ser[5]), .B0_f (new_AGEMA_signal_3691), .B1_t (new_AGEMA_signal_3692), .B1_f (new_AGEMA_signal_3693), .Z0_t (KeyArray_S30reg_gff_1_SFF_5_n1), .Z0_f (new_AGEMA_signal_6982), .Z1_t (new_AGEMA_signal_6983), .Z1_f (new_AGEMA_signal_6984) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_5_U1 ( .A0_t (KeyArray_S30reg_gff_1_SFF_5_QD), .A0_f (new_AGEMA_signal_7763), .A1_t (new_AGEMA_signal_7764), .A1_f (new_AGEMA_signal_7765), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S30reg_gff_1_SFF_5_n2), .Z0_f (new_AGEMA_signal_7811), .Z1_t (new_AGEMA_signal_7812), .Z1_f (new_AGEMA_signal_7813) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS31ser[5]), .A0_f (new_AGEMA_signal_3739), .A1_t (new_AGEMA_signal_3740), .A1_f (new_AGEMA_signal_3741), .B0_t (KeyArray_inS30par[5]), .B0_f (new_AGEMA_signal_7610), .B1_t (new_AGEMA_signal_7611), .B1_f (new_AGEMA_signal_7612), .Z0_t (KeyArray_S30reg_gff_1_SFF_5_MUXInst_X), .Z0_f (new_AGEMA_signal_7667), .Z1_t (new_AGEMA_signal_7668), .Z1_f (new_AGEMA_signal_7669) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S30reg_gff_1_SFF_5_MUXInst_X), .B0_f (new_AGEMA_signal_7667), .B1_t (new_AGEMA_signal_7668), .B1_f (new_AGEMA_signal_7669), .Z0_t (KeyArray_S30reg_gff_1_SFF_5_MUXInst_Y), .Z0_f (new_AGEMA_signal_7715), .Z1_t (new_AGEMA_signal_7716), .Z1_f (new_AGEMA_signal_7717) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S30reg_gff_1_SFF_5_MUXInst_Y), .A0_f (new_AGEMA_signal_7715), .A1_t (new_AGEMA_signal_7716), .A1_f (new_AGEMA_signal_7717), .B0_t (KeyArray_outS31ser[5]), .B0_f (new_AGEMA_signal_3739), .B1_t (new_AGEMA_signal_3740), .B1_f (new_AGEMA_signal_3741), .Z0_t (KeyArray_S30reg_gff_1_SFF_5_QD), .Z0_f (new_AGEMA_signal_7763), .Z1_t (new_AGEMA_signal_7764), .Z1_f (new_AGEMA_signal_7765) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S30reg_gff_1_SFF_6_U3 ( .A0_t (KeyArray_S30reg_gff_1_SFF_6_n2), .A0_f (new_AGEMA_signal_7814), .A1_t (new_AGEMA_signal_7815), .A1_f (new_AGEMA_signal_7816), .B0_t (KeyArray_S30reg_gff_1_SFF_6_n1), .B0_f (new_AGEMA_signal_6985), .B1_t (new_AGEMA_signal_6986), .B1_f (new_AGEMA_signal_6987), .Z0_t (KeyArray_outS30ser[6]), .Z0_f (new_AGEMA_signal_3697), .Z1_t (new_AGEMA_signal_3698), .Z1_f (new_AGEMA_signal_3699) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_6_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS30ser[6]), .B0_f (new_AGEMA_signal_3697), .B1_t (new_AGEMA_signal_3698), .B1_f (new_AGEMA_signal_3699), .Z0_t (KeyArray_S30reg_gff_1_SFF_6_n1), .Z0_f (new_AGEMA_signal_6985), .Z1_t (new_AGEMA_signal_6986), .Z1_f (new_AGEMA_signal_6987) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_6_U1 ( .A0_t (KeyArray_S30reg_gff_1_SFF_6_QD), .A0_f (new_AGEMA_signal_7766), .A1_t (new_AGEMA_signal_7767), .A1_f (new_AGEMA_signal_7768), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S30reg_gff_1_SFF_6_n2), .Z0_f (new_AGEMA_signal_7814), .Z1_t (new_AGEMA_signal_7815), .Z1_f (new_AGEMA_signal_7816) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS31ser[6]), .A0_f (new_AGEMA_signal_3745), .A1_t (new_AGEMA_signal_3746), .A1_f (new_AGEMA_signal_3747), .B0_t (KeyArray_inS30par[6]), .B0_f (new_AGEMA_signal_7607), .B1_t (new_AGEMA_signal_7608), .B1_f (new_AGEMA_signal_7609), .Z0_t (KeyArray_S30reg_gff_1_SFF_6_MUXInst_X), .Z0_f (new_AGEMA_signal_7670), .Z1_t (new_AGEMA_signal_7671), .Z1_f (new_AGEMA_signal_7672) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S30reg_gff_1_SFF_6_MUXInst_X), .B0_f (new_AGEMA_signal_7670), .B1_t (new_AGEMA_signal_7671), .B1_f (new_AGEMA_signal_7672), .Z0_t (KeyArray_S30reg_gff_1_SFF_6_MUXInst_Y), .Z0_f (new_AGEMA_signal_7718), .Z1_t (new_AGEMA_signal_7719), .Z1_f (new_AGEMA_signal_7720) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S30reg_gff_1_SFF_6_MUXInst_Y), .A0_f (new_AGEMA_signal_7718), .A1_t (new_AGEMA_signal_7719), .A1_f (new_AGEMA_signal_7720), .B0_t (KeyArray_outS31ser[6]), .B0_f (new_AGEMA_signal_3745), .B1_t (new_AGEMA_signal_3746), .B1_f (new_AGEMA_signal_3747), .Z0_t (KeyArray_S30reg_gff_1_SFF_6_QD), .Z0_f (new_AGEMA_signal_7766), .Z1_t (new_AGEMA_signal_7767), .Z1_f (new_AGEMA_signal_7768) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S30reg_gff_1_SFF_7_U3 ( .A0_t (KeyArray_S30reg_gff_1_SFF_7_n2), .A0_f (new_AGEMA_signal_7817), .A1_t (new_AGEMA_signal_7818), .A1_f (new_AGEMA_signal_7819), .B0_t (KeyArray_S30reg_gff_1_SFF_7_n1), .B0_f (new_AGEMA_signal_6988), .B1_t (new_AGEMA_signal_6989), .B1_f (new_AGEMA_signal_6990), .Z0_t (KeyArray_outS30ser[7]), .Z0_f (new_AGEMA_signal_3703), .Z1_t (new_AGEMA_signal_3704), .Z1_f (new_AGEMA_signal_3705) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_7_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS30ser[7]), .B0_f (new_AGEMA_signal_3703), .B1_t (new_AGEMA_signal_3704), .B1_f (new_AGEMA_signal_3705), .Z0_t (KeyArray_S30reg_gff_1_SFF_7_n1), .Z0_f (new_AGEMA_signal_6988), .Z1_t (new_AGEMA_signal_6989), .Z1_f (new_AGEMA_signal_6990) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_7_U1 ( .A0_t (KeyArray_S30reg_gff_1_SFF_7_QD), .A0_f (new_AGEMA_signal_7769), .A1_t (new_AGEMA_signal_7770), .A1_f (new_AGEMA_signal_7771), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S30reg_gff_1_SFF_7_n2), .Z0_f (new_AGEMA_signal_7817), .Z1_t (new_AGEMA_signal_7818), .Z1_f (new_AGEMA_signal_7819) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS31ser[7]), .A0_f (new_AGEMA_signal_3751), .A1_t (new_AGEMA_signal_3752), .A1_f (new_AGEMA_signal_3753), .B0_t (KeyArray_inS30par[7]), .B0_f (new_AGEMA_signal_7604), .B1_t (new_AGEMA_signal_7605), .B1_f (new_AGEMA_signal_7606), .Z0_t (KeyArray_S30reg_gff_1_SFF_7_MUXInst_X), .Z0_f (new_AGEMA_signal_7673), .Z1_t (new_AGEMA_signal_7674), .Z1_f (new_AGEMA_signal_7675) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S30reg_gff_1_SFF_7_MUXInst_X), .B0_f (new_AGEMA_signal_7673), .B1_t (new_AGEMA_signal_7674), .B1_f (new_AGEMA_signal_7675), .Z0_t (KeyArray_S30reg_gff_1_SFF_7_MUXInst_Y), .Z0_f (new_AGEMA_signal_7721), .Z1_t (new_AGEMA_signal_7722), .Z1_f (new_AGEMA_signal_7723) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S30reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S30reg_gff_1_SFF_7_MUXInst_Y), .A0_f (new_AGEMA_signal_7721), .A1_t (new_AGEMA_signal_7722), .A1_f (new_AGEMA_signal_7723), .B0_t (KeyArray_outS31ser[7]), .B0_f (new_AGEMA_signal_3751), .B1_t (new_AGEMA_signal_3752), .B1_f (new_AGEMA_signal_3753), .Z0_t (KeyArray_S30reg_gff_1_SFF_7_QD), .Z0_f (new_AGEMA_signal_7769), .Z1_t (new_AGEMA_signal_7770), .Z1_f (new_AGEMA_signal_7771) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S31reg_gff_1_SFF_0_U3 ( .A0_t (KeyArray_S31reg_gff_1_SFF_0_n2), .A0_f (new_AGEMA_signal_6994), .A1_t (new_AGEMA_signal_6995), .A1_f (new_AGEMA_signal_6996), .B0_t (KeyArray_S31reg_gff_1_SFF_0_n1), .B0_f (new_AGEMA_signal_6991), .B1_t (new_AGEMA_signal_6992), .B1_f (new_AGEMA_signal_6993), .Z0_t (KeyArray_outS31ser[0]), .Z0_f (new_AGEMA_signal_3709), .Z1_t (new_AGEMA_signal_3710), .Z1_f (new_AGEMA_signal_3711) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_0_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS31ser[0]), .B0_f (new_AGEMA_signal_3709), .B1_t (new_AGEMA_signal_3710), .B1_f (new_AGEMA_signal_3711), .Z0_t (KeyArray_S31reg_gff_1_SFF_0_n1), .Z0_f (new_AGEMA_signal_6991), .Z1_t (new_AGEMA_signal_6992), .Z1_f (new_AGEMA_signal_6993) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_0_U1 ( .A0_t (KeyArray_S31reg_gff_1_SFF_0_QD), .A0_f (new_AGEMA_signal_4965), .A1_t (new_AGEMA_signal_4966), .A1_f (new_AGEMA_signal_4967), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S31reg_gff_1_SFF_0_n2), .Z0_f (new_AGEMA_signal_6994), .Z1_t (new_AGEMA_signal_6995), .Z1_f (new_AGEMA_signal_6996) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS32ser[0]), .A0_f (new_AGEMA_signal_3757), .A1_t (new_AGEMA_signal_3758), .A1_f (new_AGEMA_signal_3759), .B0_t (KeyArray_outS01ser_0_), .B0_f (new_AGEMA_signal_3247), .B1_t (new_AGEMA_signal_3248), .B1_f (new_AGEMA_signal_3249), .Z0_t (KeyArray_S31reg_gff_1_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_3853), .Z1_t (new_AGEMA_signal_3854), .Z1_f (new_AGEMA_signal_3855) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S31reg_gff_1_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_3853), .B1_t (new_AGEMA_signal_3854), .B1_f (new_AGEMA_signal_3855), .Z0_t (KeyArray_S31reg_gff_1_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_4475), .Z1_t (new_AGEMA_signal_4476), .Z1_f (new_AGEMA_signal_4477) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S31reg_gff_1_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_4475), .A1_t (new_AGEMA_signal_4476), .A1_f (new_AGEMA_signal_4477), .B0_t (KeyArray_outS32ser[0]), .B0_f (new_AGEMA_signal_3757), .B1_t (new_AGEMA_signal_3758), .B1_f (new_AGEMA_signal_3759), .Z0_t (KeyArray_S31reg_gff_1_SFF_0_QD), .Z0_f (new_AGEMA_signal_4965), .Z1_t (new_AGEMA_signal_4966), .Z1_f (new_AGEMA_signal_4967) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S31reg_gff_1_SFF_1_U3 ( .A0_t (KeyArray_S31reg_gff_1_SFF_1_n2), .A0_f (new_AGEMA_signal_7000), .A1_t (new_AGEMA_signal_7001), .A1_f (new_AGEMA_signal_7002), .B0_t (KeyArray_S31reg_gff_1_SFF_1_n1), .B0_f (new_AGEMA_signal_6997), .B1_t (new_AGEMA_signal_6998), .B1_f (new_AGEMA_signal_6999), .Z0_t (KeyArray_outS31ser[1]), .Z0_f (new_AGEMA_signal_3715), .Z1_t (new_AGEMA_signal_3716), .Z1_f (new_AGEMA_signal_3717) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_1_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS31ser[1]), .B0_f (new_AGEMA_signal_3715), .B1_t (new_AGEMA_signal_3716), .B1_f (new_AGEMA_signal_3717), .Z0_t (KeyArray_S31reg_gff_1_SFF_1_n1), .Z0_f (new_AGEMA_signal_6997), .Z1_t (new_AGEMA_signal_6998), .Z1_f (new_AGEMA_signal_6999) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_1_U1 ( .A0_t (KeyArray_S31reg_gff_1_SFF_1_QD), .A0_f (new_AGEMA_signal_4968), .A1_t (new_AGEMA_signal_4969), .A1_f (new_AGEMA_signal_4970), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S31reg_gff_1_SFF_1_n2), .Z0_f (new_AGEMA_signal_7000), .Z1_t (new_AGEMA_signal_7001), .Z1_f (new_AGEMA_signal_7002) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS32ser[1]), .A0_f (new_AGEMA_signal_3763), .A1_t (new_AGEMA_signal_3764), .A1_f (new_AGEMA_signal_3765), .B0_t (KeyArray_outS01ser_1_), .B0_f (new_AGEMA_signal_3241), .B1_t (new_AGEMA_signal_3242), .B1_f (new_AGEMA_signal_3243), .Z0_t (KeyArray_S31reg_gff_1_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_3856), .Z1_t (new_AGEMA_signal_3857), .Z1_f (new_AGEMA_signal_3858) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S31reg_gff_1_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_3856), .B1_t (new_AGEMA_signal_3857), .B1_f (new_AGEMA_signal_3858), .Z0_t (KeyArray_S31reg_gff_1_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_4478), .Z1_t (new_AGEMA_signal_4479), .Z1_f (new_AGEMA_signal_4480) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S31reg_gff_1_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_4478), .A1_t (new_AGEMA_signal_4479), .A1_f (new_AGEMA_signal_4480), .B0_t (KeyArray_outS32ser[1]), .B0_f (new_AGEMA_signal_3763), .B1_t (new_AGEMA_signal_3764), .B1_f (new_AGEMA_signal_3765), .Z0_t (KeyArray_S31reg_gff_1_SFF_1_QD), .Z0_f (new_AGEMA_signal_4968), .Z1_t (new_AGEMA_signal_4969), .Z1_f (new_AGEMA_signal_4970) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S31reg_gff_1_SFF_2_U3 ( .A0_t (KeyArray_S31reg_gff_1_SFF_2_n2), .A0_f (new_AGEMA_signal_7006), .A1_t (new_AGEMA_signal_7007), .A1_f (new_AGEMA_signal_7008), .B0_t (KeyArray_S31reg_gff_1_SFF_2_n1), .B0_f (new_AGEMA_signal_7003), .B1_t (new_AGEMA_signal_7004), .B1_f (new_AGEMA_signal_7005), .Z0_t (KeyArray_outS31ser[2]), .Z0_f (new_AGEMA_signal_3721), .Z1_t (new_AGEMA_signal_3722), .Z1_f (new_AGEMA_signal_3723) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_2_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS31ser[2]), .B0_f (new_AGEMA_signal_3721), .B1_t (new_AGEMA_signal_3722), .B1_f (new_AGEMA_signal_3723), .Z0_t (KeyArray_S31reg_gff_1_SFF_2_n1), .Z0_f (new_AGEMA_signal_7003), .Z1_t (new_AGEMA_signal_7004), .Z1_f (new_AGEMA_signal_7005) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_2_U1 ( .A0_t (KeyArray_S31reg_gff_1_SFF_2_QD), .A0_f (new_AGEMA_signal_4971), .A1_t (new_AGEMA_signal_4972), .A1_f (new_AGEMA_signal_4973), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S31reg_gff_1_SFF_2_n2), .Z0_f (new_AGEMA_signal_7006), .Z1_t (new_AGEMA_signal_7007), .Z1_f (new_AGEMA_signal_7008) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS32ser[2]), .A0_f (new_AGEMA_signal_3769), .A1_t (new_AGEMA_signal_3770), .A1_f (new_AGEMA_signal_3771), .B0_t (KeyArray_outS01ser_2_), .B0_f (new_AGEMA_signal_3235), .B1_t (new_AGEMA_signal_3236), .B1_f (new_AGEMA_signal_3237), .Z0_t (KeyArray_S31reg_gff_1_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_3859), .Z1_t (new_AGEMA_signal_3860), .Z1_f (new_AGEMA_signal_3861) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S31reg_gff_1_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_3859), .B1_t (new_AGEMA_signal_3860), .B1_f (new_AGEMA_signal_3861), .Z0_t (KeyArray_S31reg_gff_1_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_4481), .Z1_t (new_AGEMA_signal_4482), .Z1_f (new_AGEMA_signal_4483) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S31reg_gff_1_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_4481), .A1_t (new_AGEMA_signal_4482), .A1_f (new_AGEMA_signal_4483), .B0_t (KeyArray_outS32ser[2]), .B0_f (new_AGEMA_signal_3769), .B1_t (new_AGEMA_signal_3770), .B1_f (new_AGEMA_signal_3771), .Z0_t (KeyArray_S31reg_gff_1_SFF_2_QD), .Z0_f (new_AGEMA_signal_4971), .Z1_t (new_AGEMA_signal_4972), .Z1_f (new_AGEMA_signal_4973) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S31reg_gff_1_SFF_3_U3 ( .A0_t (KeyArray_S31reg_gff_1_SFF_3_n2), .A0_f (new_AGEMA_signal_7012), .A1_t (new_AGEMA_signal_7013), .A1_f (new_AGEMA_signal_7014), .B0_t (KeyArray_S31reg_gff_1_SFF_3_n1), .B0_f (new_AGEMA_signal_7009), .B1_t (new_AGEMA_signal_7010), .B1_f (new_AGEMA_signal_7011), .Z0_t (KeyArray_outS31ser[3]), .Z0_f (new_AGEMA_signal_3727), .Z1_t (new_AGEMA_signal_3728), .Z1_f (new_AGEMA_signal_3729) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_3_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS31ser[3]), .B0_f (new_AGEMA_signal_3727), .B1_t (new_AGEMA_signal_3728), .B1_f (new_AGEMA_signal_3729), .Z0_t (KeyArray_S31reg_gff_1_SFF_3_n1), .Z0_f (new_AGEMA_signal_7009), .Z1_t (new_AGEMA_signal_7010), .Z1_f (new_AGEMA_signal_7011) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_3_U1 ( .A0_t (KeyArray_S31reg_gff_1_SFF_3_QD), .A0_f (new_AGEMA_signal_4974), .A1_t (new_AGEMA_signal_4975), .A1_f (new_AGEMA_signal_4976), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S31reg_gff_1_SFF_3_n2), .Z0_f (new_AGEMA_signal_7012), .Z1_t (new_AGEMA_signal_7013), .Z1_f (new_AGEMA_signal_7014) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS32ser[3]), .A0_f (new_AGEMA_signal_3775), .A1_t (new_AGEMA_signal_3776), .A1_f (new_AGEMA_signal_3777), .B0_t (KeyArray_outS01ser_3_), .B0_f (new_AGEMA_signal_3229), .B1_t (new_AGEMA_signal_3230), .B1_f (new_AGEMA_signal_3231), .Z0_t (KeyArray_S31reg_gff_1_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_3862), .Z1_t (new_AGEMA_signal_3863), .Z1_f (new_AGEMA_signal_3864) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S31reg_gff_1_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_3862), .B1_t (new_AGEMA_signal_3863), .B1_f (new_AGEMA_signal_3864), .Z0_t (KeyArray_S31reg_gff_1_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_4484), .Z1_t (new_AGEMA_signal_4485), .Z1_f (new_AGEMA_signal_4486) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S31reg_gff_1_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_4484), .A1_t (new_AGEMA_signal_4485), .A1_f (new_AGEMA_signal_4486), .B0_t (KeyArray_outS32ser[3]), .B0_f (new_AGEMA_signal_3775), .B1_t (new_AGEMA_signal_3776), .B1_f (new_AGEMA_signal_3777), .Z0_t (KeyArray_S31reg_gff_1_SFF_3_QD), .Z0_f (new_AGEMA_signal_4974), .Z1_t (new_AGEMA_signal_4975), .Z1_f (new_AGEMA_signal_4976) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S31reg_gff_1_SFF_4_U3 ( .A0_t (KeyArray_S31reg_gff_1_SFF_4_n2), .A0_f (new_AGEMA_signal_7018), .A1_t (new_AGEMA_signal_7019), .A1_f (new_AGEMA_signal_7020), .B0_t (KeyArray_S31reg_gff_1_SFF_4_n1), .B0_f (new_AGEMA_signal_7015), .B1_t (new_AGEMA_signal_7016), .B1_f (new_AGEMA_signal_7017), .Z0_t (KeyArray_outS31ser[4]), .Z0_f (new_AGEMA_signal_3733), .Z1_t (new_AGEMA_signal_3734), .Z1_f (new_AGEMA_signal_3735) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_4_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS31ser[4]), .B0_f (new_AGEMA_signal_3733), .B1_t (new_AGEMA_signal_3734), .B1_f (new_AGEMA_signal_3735), .Z0_t (KeyArray_S31reg_gff_1_SFF_4_n1), .Z0_f (new_AGEMA_signal_7015), .Z1_t (new_AGEMA_signal_7016), .Z1_f (new_AGEMA_signal_7017) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_4_U1 ( .A0_t (KeyArray_S31reg_gff_1_SFF_4_QD), .A0_f (new_AGEMA_signal_4977), .A1_t (new_AGEMA_signal_4978), .A1_f (new_AGEMA_signal_4979), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S31reg_gff_1_SFF_4_n2), .Z0_f (new_AGEMA_signal_7018), .Z1_t (new_AGEMA_signal_7019), .Z1_f (new_AGEMA_signal_7020) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS32ser[4]), .A0_f (new_AGEMA_signal_3781), .A1_t (new_AGEMA_signal_3782), .A1_f (new_AGEMA_signal_3783), .B0_t (KeyArray_outS01ser_4_), .B0_f (new_AGEMA_signal_3223), .B1_t (new_AGEMA_signal_3224), .B1_f (new_AGEMA_signal_3225), .Z0_t (KeyArray_S31reg_gff_1_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_3865), .Z1_t (new_AGEMA_signal_3866), .Z1_f (new_AGEMA_signal_3867) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S31reg_gff_1_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_3865), .B1_t (new_AGEMA_signal_3866), .B1_f (new_AGEMA_signal_3867), .Z0_t (KeyArray_S31reg_gff_1_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_4487), .Z1_t (new_AGEMA_signal_4488), .Z1_f (new_AGEMA_signal_4489) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S31reg_gff_1_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_4487), .A1_t (new_AGEMA_signal_4488), .A1_f (new_AGEMA_signal_4489), .B0_t (KeyArray_outS32ser[4]), .B0_f (new_AGEMA_signal_3781), .B1_t (new_AGEMA_signal_3782), .B1_f (new_AGEMA_signal_3783), .Z0_t (KeyArray_S31reg_gff_1_SFF_4_QD), .Z0_f (new_AGEMA_signal_4977), .Z1_t (new_AGEMA_signal_4978), .Z1_f (new_AGEMA_signal_4979) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S31reg_gff_1_SFF_5_U3 ( .A0_t (KeyArray_S31reg_gff_1_SFF_5_n2), .A0_f (new_AGEMA_signal_7024), .A1_t (new_AGEMA_signal_7025), .A1_f (new_AGEMA_signal_7026), .B0_t (KeyArray_S31reg_gff_1_SFF_5_n1), .B0_f (new_AGEMA_signal_7021), .B1_t (new_AGEMA_signal_7022), .B1_f (new_AGEMA_signal_7023), .Z0_t (KeyArray_outS31ser[5]), .Z0_f (new_AGEMA_signal_3739), .Z1_t (new_AGEMA_signal_3740), .Z1_f (new_AGEMA_signal_3741) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_5_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS31ser[5]), .B0_f (new_AGEMA_signal_3739), .B1_t (new_AGEMA_signal_3740), .B1_f (new_AGEMA_signal_3741), .Z0_t (KeyArray_S31reg_gff_1_SFF_5_n1), .Z0_f (new_AGEMA_signal_7021), .Z1_t (new_AGEMA_signal_7022), .Z1_f (new_AGEMA_signal_7023) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_5_U1 ( .A0_t (KeyArray_S31reg_gff_1_SFF_5_QD), .A0_f (new_AGEMA_signal_4980), .A1_t (new_AGEMA_signal_4981), .A1_f (new_AGEMA_signal_4982), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S31reg_gff_1_SFF_5_n2), .Z0_f (new_AGEMA_signal_7024), .Z1_t (new_AGEMA_signal_7025), .Z1_f (new_AGEMA_signal_7026) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS32ser[5]), .A0_f (new_AGEMA_signal_3787), .A1_t (new_AGEMA_signal_3788), .A1_f (new_AGEMA_signal_3789), .B0_t (KeyArray_outS01ser_5_), .B0_f (new_AGEMA_signal_3217), .B1_t (new_AGEMA_signal_3218), .B1_f (new_AGEMA_signal_3219), .Z0_t (KeyArray_S31reg_gff_1_SFF_5_MUXInst_X), .Z0_f (new_AGEMA_signal_3868), .Z1_t (new_AGEMA_signal_3869), .Z1_f (new_AGEMA_signal_3870) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S31reg_gff_1_SFF_5_MUXInst_X), .B0_f (new_AGEMA_signal_3868), .B1_t (new_AGEMA_signal_3869), .B1_f (new_AGEMA_signal_3870), .Z0_t (KeyArray_S31reg_gff_1_SFF_5_MUXInst_Y), .Z0_f (new_AGEMA_signal_4490), .Z1_t (new_AGEMA_signal_4491), .Z1_f (new_AGEMA_signal_4492) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S31reg_gff_1_SFF_5_MUXInst_Y), .A0_f (new_AGEMA_signal_4490), .A1_t (new_AGEMA_signal_4491), .A1_f (new_AGEMA_signal_4492), .B0_t (KeyArray_outS32ser[5]), .B0_f (new_AGEMA_signal_3787), .B1_t (new_AGEMA_signal_3788), .B1_f (new_AGEMA_signal_3789), .Z0_t (KeyArray_S31reg_gff_1_SFF_5_QD), .Z0_f (new_AGEMA_signal_4980), .Z1_t (new_AGEMA_signal_4981), .Z1_f (new_AGEMA_signal_4982) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S31reg_gff_1_SFF_6_U3 ( .A0_t (KeyArray_S31reg_gff_1_SFF_6_n2), .A0_f (new_AGEMA_signal_7030), .A1_t (new_AGEMA_signal_7031), .A1_f (new_AGEMA_signal_7032), .B0_t (KeyArray_S31reg_gff_1_SFF_6_n1), .B0_f (new_AGEMA_signal_7027), .B1_t (new_AGEMA_signal_7028), .B1_f (new_AGEMA_signal_7029), .Z0_t (KeyArray_outS31ser[6]), .Z0_f (new_AGEMA_signal_3745), .Z1_t (new_AGEMA_signal_3746), .Z1_f (new_AGEMA_signal_3747) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_6_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS31ser[6]), .B0_f (new_AGEMA_signal_3745), .B1_t (new_AGEMA_signal_3746), .B1_f (new_AGEMA_signal_3747), .Z0_t (KeyArray_S31reg_gff_1_SFF_6_n1), .Z0_f (new_AGEMA_signal_7027), .Z1_t (new_AGEMA_signal_7028), .Z1_f (new_AGEMA_signal_7029) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_6_U1 ( .A0_t (KeyArray_S31reg_gff_1_SFF_6_QD), .A0_f (new_AGEMA_signal_4983), .A1_t (new_AGEMA_signal_4984), .A1_f (new_AGEMA_signal_4985), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S31reg_gff_1_SFF_6_n2), .Z0_f (new_AGEMA_signal_7030), .Z1_t (new_AGEMA_signal_7031), .Z1_f (new_AGEMA_signal_7032) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS32ser[6]), .A0_f (new_AGEMA_signal_3793), .A1_t (new_AGEMA_signal_3794), .A1_f (new_AGEMA_signal_3795), .B0_t (KeyArray_outS01ser_6_), .B0_f (new_AGEMA_signal_3211), .B1_t (new_AGEMA_signal_3212), .B1_f (new_AGEMA_signal_3213), .Z0_t (KeyArray_S31reg_gff_1_SFF_6_MUXInst_X), .Z0_f (new_AGEMA_signal_3871), .Z1_t (new_AGEMA_signal_3872), .Z1_f (new_AGEMA_signal_3873) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S31reg_gff_1_SFF_6_MUXInst_X), .B0_f (new_AGEMA_signal_3871), .B1_t (new_AGEMA_signal_3872), .B1_f (new_AGEMA_signal_3873), .Z0_t (KeyArray_S31reg_gff_1_SFF_6_MUXInst_Y), .Z0_f (new_AGEMA_signal_4493), .Z1_t (new_AGEMA_signal_4494), .Z1_f (new_AGEMA_signal_4495) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S31reg_gff_1_SFF_6_MUXInst_Y), .A0_f (new_AGEMA_signal_4493), .A1_t (new_AGEMA_signal_4494), .A1_f (new_AGEMA_signal_4495), .B0_t (KeyArray_outS32ser[6]), .B0_f (new_AGEMA_signal_3793), .B1_t (new_AGEMA_signal_3794), .B1_f (new_AGEMA_signal_3795), .Z0_t (KeyArray_S31reg_gff_1_SFF_6_QD), .Z0_f (new_AGEMA_signal_4983), .Z1_t (new_AGEMA_signal_4984), .Z1_f (new_AGEMA_signal_4985) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S31reg_gff_1_SFF_7_U3 ( .A0_t (KeyArray_S31reg_gff_1_SFF_7_n2), .A0_f (new_AGEMA_signal_7036), .A1_t (new_AGEMA_signal_7037), .A1_f (new_AGEMA_signal_7038), .B0_t (KeyArray_S31reg_gff_1_SFF_7_n1), .B0_f (new_AGEMA_signal_7033), .B1_t (new_AGEMA_signal_7034), .B1_f (new_AGEMA_signal_7035), .Z0_t (KeyArray_outS31ser[7]), .Z0_f (new_AGEMA_signal_3751), .Z1_t (new_AGEMA_signal_3752), .Z1_f (new_AGEMA_signal_3753) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_7_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS31ser[7]), .B0_f (new_AGEMA_signal_3751), .B1_t (new_AGEMA_signal_3752), .B1_f (new_AGEMA_signal_3753), .Z0_t (KeyArray_S31reg_gff_1_SFF_7_n1), .Z0_f (new_AGEMA_signal_7033), .Z1_t (new_AGEMA_signal_7034), .Z1_f (new_AGEMA_signal_7035) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_7_U1 ( .A0_t (KeyArray_S31reg_gff_1_SFF_7_QD), .A0_f (new_AGEMA_signal_4986), .A1_t (new_AGEMA_signal_4987), .A1_f (new_AGEMA_signal_4988), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S31reg_gff_1_SFF_7_n2), .Z0_f (new_AGEMA_signal_7036), .Z1_t (new_AGEMA_signal_7037), .Z1_f (new_AGEMA_signal_7038) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS32ser[7]), .A0_f (new_AGEMA_signal_3799), .A1_t (new_AGEMA_signal_3800), .A1_f (new_AGEMA_signal_3801), .B0_t (KeyArray_outS01ser_7_), .B0_f (new_AGEMA_signal_3205), .B1_t (new_AGEMA_signal_3206), .B1_f (new_AGEMA_signal_3207), .Z0_t (KeyArray_S31reg_gff_1_SFF_7_MUXInst_X), .Z0_f (new_AGEMA_signal_3874), .Z1_t (new_AGEMA_signal_3875), .Z1_f (new_AGEMA_signal_3876) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S31reg_gff_1_SFF_7_MUXInst_X), .B0_f (new_AGEMA_signal_3874), .B1_t (new_AGEMA_signal_3875), .B1_f (new_AGEMA_signal_3876), .Z0_t (KeyArray_S31reg_gff_1_SFF_7_MUXInst_Y), .Z0_f (new_AGEMA_signal_4496), .Z1_t (new_AGEMA_signal_4497), .Z1_f (new_AGEMA_signal_4498) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S31reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S31reg_gff_1_SFF_7_MUXInst_Y), .A0_f (new_AGEMA_signal_4496), .A1_t (new_AGEMA_signal_4497), .A1_f (new_AGEMA_signal_4498), .B0_t (KeyArray_outS32ser[7]), .B0_f (new_AGEMA_signal_3799), .B1_t (new_AGEMA_signal_3800), .B1_f (new_AGEMA_signal_3801), .Z0_t (KeyArray_S31reg_gff_1_SFF_7_QD), .Z0_f (new_AGEMA_signal_4986), .Z1_t (new_AGEMA_signal_4987), .Z1_f (new_AGEMA_signal_4988) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S32reg_gff_1_SFF_0_U3 ( .A0_t (KeyArray_S32reg_gff_1_SFF_0_n2), .A0_f (new_AGEMA_signal_7042), .A1_t (new_AGEMA_signal_7043), .A1_f (new_AGEMA_signal_7044), .B0_t (KeyArray_S32reg_gff_1_SFF_0_n1), .B0_f (new_AGEMA_signal_7039), .B1_t (new_AGEMA_signal_7040), .B1_f (new_AGEMA_signal_7041), .Z0_t (KeyArray_outS32ser[0]), .Z0_f (new_AGEMA_signal_3757), .Z1_t (new_AGEMA_signal_3758), .Z1_f (new_AGEMA_signal_3759) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_0_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS32ser[0]), .B0_f (new_AGEMA_signal_3757), .B1_t (new_AGEMA_signal_3758), .B1_f (new_AGEMA_signal_3759), .Z0_t (KeyArray_S32reg_gff_1_SFF_0_n1), .Z0_f (new_AGEMA_signal_7039), .Z1_t (new_AGEMA_signal_7040), .Z1_f (new_AGEMA_signal_7041) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_0_U1 ( .A0_t (KeyArray_S32reg_gff_1_SFF_0_QD), .A0_f (new_AGEMA_signal_4989), .A1_t (new_AGEMA_signal_4990), .A1_f (new_AGEMA_signal_4991), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S32reg_gff_1_SFF_0_n2), .Z0_f (new_AGEMA_signal_7042), .Z1_t (new_AGEMA_signal_7043), .Z1_f (new_AGEMA_signal_7044) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS33ser[0]), .A0_f (new_AGEMA_signal_3805), .A1_t (new_AGEMA_signal_3806), .A1_f (new_AGEMA_signal_3807), .B0_t (KeyArray_outS02ser[0]), .B0_f (new_AGEMA_signal_3253), .B1_t (new_AGEMA_signal_3254), .B1_f (new_AGEMA_signal_3255), .Z0_t (KeyArray_S32reg_gff_1_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_3877), .Z1_t (new_AGEMA_signal_3878), .Z1_f (new_AGEMA_signal_3879) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S32reg_gff_1_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_3877), .B1_t (new_AGEMA_signal_3878), .B1_f (new_AGEMA_signal_3879), .Z0_t (KeyArray_S32reg_gff_1_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_4499), .Z1_t (new_AGEMA_signal_4500), .Z1_f (new_AGEMA_signal_4501) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S32reg_gff_1_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_4499), .A1_t (new_AGEMA_signal_4500), .A1_f (new_AGEMA_signal_4501), .B0_t (KeyArray_outS33ser[0]), .B0_f (new_AGEMA_signal_3805), .B1_t (new_AGEMA_signal_3806), .B1_f (new_AGEMA_signal_3807), .Z0_t (KeyArray_S32reg_gff_1_SFF_0_QD), .Z0_f (new_AGEMA_signal_4989), .Z1_t (new_AGEMA_signal_4990), .Z1_f (new_AGEMA_signal_4991) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S32reg_gff_1_SFF_1_U3 ( .A0_t (KeyArray_S32reg_gff_1_SFF_1_n2), .A0_f (new_AGEMA_signal_7048), .A1_t (new_AGEMA_signal_7049), .A1_f (new_AGEMA_signal_7050), .B0_t (KeyArray_S32reg_gff_1_SFF_1_n1), .B0_f (new_AGEMA_signal_7045), .B1_t (new_AGEMA_signal_7046), .B1_f (new_AGEMA_signal_7047), .Z0_t (KeyArray_outS32ser[1]), .Z0_f (new_AGEMA_signal_3763), .Z1_t (new_AGEMA_signal_3764), .Z1_f (new_AGEMA_signal_3765) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_1_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS32ser[1]), .B0_f (new_AGEMA_signal_3763), .B1_t (new_AGEMA_signal_3764), .B1_f (new_AGEMA_signal_3765), .Z0_t (KeyArray_S32reg_gff_1_SFF_1_n1), .Z0_f (new_AGEMA_signal_7045), .Z1_t (new_AGEMA_signal_7046), .Z1_f (new_AGEMA_signal_7047) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_1_U1 ( .A0_t (KeyArray_S32reg_gff_1_SFF_1_QD), .A0_f (new_AGEMA_signal_4992), .A1_t (new_AGEMA_signal_4993), .A1_f (new_AGEMA_signal_4994), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S32reg_gff_1_SFF_1_n2), .Z0_f (new_AGEMA_signal_7048), .Z1_t (new_AGEMA_signal_7049), .Z1_f (new_AGEMA_signal_7050) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS33ser[1]), .A0_f (new_AGEMA_signal_3811), .A1_t (new_AGEMA_signal_3812), .A1_f (new_AGEMA_signal_3813), .B0_t (KeyArray_outS02ser[1]), .B0_f (new_AGEMA_signal_3262), .B1_t (new_AGEMA_signal_3263), .B1_f (new_AGEMA_signal_3264), .Z0_t (KeyArray_S32reg_gff_1_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_3880), .Z1_t (new_AGEMA_signal_3881), .Z1_f (new_AGEMA_signal_3882) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S32reg_gff_1_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_3880), .B1_t (new_AGEMA_signal_3881), .B1_f (new_AGEMA_signal_3882), .Z0_t (KeyArray_S32reg_gff_1_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_4502), .Z1_t (new_AGEMA_signal_4503), .Z1_f (new_AGEMA_signal_4504) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S32reg_gff_1_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_4502), .A1_t (new_AGEMA_signal_4503), .A1_f (new_AGEMA_signal_4504), .B0_t (KeyArray_outS33ser[1]), .B0_f (new_AGEMA_signal_3811), .B1_t (new_AGEMA_signal_3812), .B1_f (new_AGEMA_signal_3813), .Z0_t (KeyArray_S32reg_gff_1_SFF_1_QD), .Z0_f (new_AGEMA_signal_4992), .Z1_t (new_AGEMA_signal_4993), .Z1_f (new_AGEMA_signal_4994) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S32reg_gff_1_SFF_2_U3 ( .A0_t (KeyArray_S32reg_gff_1_SFF_2_n2), .A0_f (new_AGEMA_signal_7054), .A1_t (new_AGEMA_signal_7055), .A1_f (new_AGEMA_signal_7056), .B0_t (KeyArray_S32reg_gff_1_SFF_2_n1), .B0_f (new_AGEMA_signal_7051), .B1_t (new_AGEMA_signal_7052), .B1_f (new_AGEMA_signal_7053), .Z0_t (KeyArray_outS32ser[2]), .Z0_f (new_AGEMA_signal_3769), .Z1_t (new_AGEMA_signal_3770), .Z1_f (new_AGEMA_signal_3771) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_2_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS32ser[2]), .B0_f (new_AGEMA_signal_3769), .B1_t (new_AGEMA_signal_3770), .B1_f (new_AGEMA_signal_3771), .Z0_t (KeyArray_S32reg_gff_1_SFF_2_n1), .Z0_f (new_AGEMA_signal_7051), .Z1_t (new_AGEMA_signal_7052), .Z1_f (new_AGEMA_signal_7053) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_2_U1 ( .A0_t (KeyArray_S32reg_gff_1_SFF_2_QD), .A0_f (new_AGEMA_signal_4995), .A1_t (new_AGEMA_signal_4996), .A1_f (new_AGEMA_signal_4997), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S32reg_gff_1_SFF_2_n2), .Z0_f (new_AGEMA_signal_7054), .Z1_t (new_AGEMA_signal_7055), .Z1_f (new_AGEMA_signal_7056) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS33ser[2]), .A0_f (new_AGEMA_signal_3817), .A1_t (new_AGEMA_signal_3818), .A1_f (new_AGEMA_signal_3819), .B0_t (KeyArray_outS02ser[2]), .B0_f (new_AGEMA_signal_3271), .B1_t (new_AGEMA_signal_3272), .B1_f (new_AGEMA_signal_3273), .Z0_t (KeyArray_S32reg_gff_1_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_3883), .Z1_t (new_AGEMA_signal_3884), .Z1_f (new_AGEMA_signal_3885) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S32reg_gff_1_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_3883), .B1_t (new_AGEMA_signal_3884), .B1_f (new_AGEMA_signal_3885), .Z0_t (KeyArray_S32reg_gff_1_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_4505), .Z1_t (new_AGEMA_signal_4506), .Z1_f (new_AGEMA_signal_4507) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S32reg_gff_1_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_4505), .A1_t (new_AGEMA_signal_4506), .A1_f (new_AGEMA_signal_4507), .B0_t (KeyArray_outS33ser[2]), .B0_f (new_AGEMA_signal_3817), .B1_t (new_AGEMA_signal_3818), .B1_f (new_AGEMA_signal_3819), .Z0_t (KeyArray_S32reg_gff_1_SFF_2_QD), .Z0_f (new_AGEMA_signal_4995), .Z1_t (new_AGEMA_signal_4996), .Z1_f (new_AGEMA_signal_4997) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S32reg_gff_1_SFF_3_U3 ( .A0_t (KeyArray_S32reg_gff_1_SFF_3_n2), .A0_f (new_AGEMA_signal_7060), .A1_t (new_AGEMA_signal_7061), .A1_f (new_AGEMA_signal_7062), .B0_t (KeyArray_S32reg_gff_1_SFF_3_n1), .B0_f (new_AGEMA_signal_7057), .B1_t (new_AGEMA_signal_7058), .B1_f (new_AGEMA_signal_7059), .Z0_t (KeyArray_outS32ser[3]), .Z0_f (new_AGEMA_signal_3775), .Z1_t (new_AGEMA_signal_3776), .Z1_f (new_AGEMA_signal_3777) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_3_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS32ser[3]), .B0_f (new_AGEMA_signal_3775), .B1_t (new_AGEMA_signal_3776), .B1_f (new_AGEMA_signal_3777), .Z0_t (KeyArray_S32reg_gff_1_SFF_3_n1), .Z0_f (new_AGEMA_signal_7057), .Z1_t (new_AGEMA_signal_7058), .Z1_f (new_AGEMA_signal_7059) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_3_U1 ( .A0_t (KeyArray_S32reg_gff_1_SFF_3_QD), .A0_f (new_AGEMA_signal_4998), .A1_t (new_AGEMA_signal_4999), .A1_f (new_AGEMA_signal_5000), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S32reg_gff_1_SFF_3_n2), .Z0_f (new_AGEMA_signal_7060), .Z1_t (new_AGEMA_signal_7061), .Z1_f (new_AGEMA_signal_7062) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS33ser[3]), .A0_f (new_AGEMA_signal_3823), .A1_t (new_AGEMA_signal_3824), .A1_f (new_AGEMA_signal_3825), .B0_t (KeyArray_outS02ser[3]), .B0_f (new_AGEMA_signal_3280), .B1_t (new_AGEMA_signal_3281), .B1_f (new_AGEMA_signal_3282), .Z0_t (KeyArray_S32reg_gff_1_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_3886), .Z1_t (new_AGEMA_signal_3887), .Z1_f (new_AGEMA_signal_3888) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S32reg_gff_1_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_3886), .B1_t (new_AGEMA_signal_3887), .B1_f (new_AGEMA_signal_3888), .Z0_t (KeyArray_S32reg_gff_1_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_4508), .Z1_t (new_AGEMA_signal_4509), .Z1_f (new_AGEMA_signal_4510) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S32reg_gff_1_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_4508), .A1_t (new_AGEMA_signal_4509), .A1_f (new_AGEMA_signal_4510), .B0_t (KeyArray_outS33ser[3]), .B0_f (new_AGEMA_signal_3823), .B1_t (new_AGEMA_signal_3824), .B1_f (new_AGEMA_signal_3825), .Z0_t (KeyArray_S32reg_gff_1_SFF_3_QD), .Z0_f (new_AGEMA_signal_4998), .Z1_t (new_AGEMA_signal_4999), .Z1_f (new_AGEMA_signal_5000) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S32reg_gff_1_SFF_4_U3 ( .A0_t (KeyArray_S32reg_gff_1_SFF_4_n2), .A0_f (new_AGEMA_signal_7066), .A1_t (new_AGEMA_signal_7067), .A1_f (new_AGEMA_signal_7068), .B0_t (KeyArray_S32reg_gff_1_SFF_4_n1), .B0_f (new_AGEMA_signal_7063), .B1_t (new_AGEMA_signal_7064), .B1_f (new_AGEMA_signal_7065), .Z0_t (KeyArray_outS32ser[4]), .Z0_f (new_AGEMA_signal_3781), .Z1_t (new_AGEMA_signal_3782), .Z1_f (new_AGEMA_signal_3783) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_4_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS32ser[4]), .B0_f (new_AGEMA_signal_3781), .B1_t (new_AGEMA_signal_3782), .B1_f (new_AGEMA_signal_3783), .Z0_t (KeyArray_S32reg_gff_1_SFF_4_n1), .Z0_f (new_AGEMA_signal_7063), .Z1_t (new_AGEMA_signal_7064), .Z1_f (new_AGEMA_signal_7065) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_4_U1 ( .A0_t (KeyArray_S32reg_gff_1_SFF_4_QD), .A0_f (new_AGEMA_signal_5001), .A1_t (new_AGEMA_signal_5002), .A1_f (new_AGEMA_signal_5003), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S32reg_gff_1_SFF_4_n2), .Z0_f (new_AGEMA_signal_7066), .Z1_t (new_AGEMA_signal_7067), .Z1_f (new_AGEMA_signal_7068) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS33ser[4]), .A0_f (new_AGEMA_signal_3829), .A1_t (new_AGEMA_signal_3830), .A1_f (new_AGEMA_signal_3831), .B0_t (KeyArray_outS02ser[4]), .B0_f (new_AGEMA_signal_3289), .B1_t (new_AGEMA_signal_3290), .B1_f (new_AGEMA_signal_3291), .Z0_t (KeyArray_S32reg_gff_1_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_3889), .Z1_t (new_AGEMA_signal_3890), .Z1_f (new_AGEMA_signal_3891) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S32reg_gff_1_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_3889), .B1_t (new_AGEMA_signal_3890), .B1_f (new_AGEMA_signal_3891), .Z0_t (KeyArray_S32reg_gff_1_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_4511), .Z1_t (new_AGEMA_signal_4512), .Z1_f (new_AGEMA_signal_4513) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S32reg_gff_1_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_4511), .A1_t (new_AGEMA_signal_4512), .A1_f (new_AGEMA_signal_4513), .B0_t (KeyArray_outS33ser[4]), .B0_f (new_AGEMA_signal_3829), .B1_t (new_AGEMA_signal_3830), .B1_f (new_AGEMA_signal_3831), .Z0_t (KeyArray_S32reg_gff_1_SFF_4_QD), .Z0_f (new_AGEMA_signal_5001), .Z1_t (new_AGEMA_signal_5002), .Z1_f (new_AGEMA_signal_5003) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S32reg_gff_1_SFF_5_U3 ( .A0_t (KeyArray_S32reg_gff_1_SFF_5_n2), .A0_f (new_AGEMA_signal_7072), .A1_t (new_AGEMA_signal_7073), .A1_f (new_AGEMA_signal_7074), .B0_t (KeyArray_S32reg_gff_1_SFF_5_n1), .B0_f (new_AGEMA_signal_7069), .B1_t (new_AGEMA_signal_7070), .B1_f (new_AGEMA_signal_7071), .Z0_t (KeyArray_outS32ser[5]), .Z0_f (new_AGEMA_signal_3787), .Z1_t (new_AGEMA_signal_3788), .Z1_f (new_AGEMA_signal_3789) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_5_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS32ser[5]), .B0_f (new_AGEMA_signal_3787), .B1_t (new_AGEMA_signal_3788), .B1_f (new_AGEMA_signal_3789), .Z0_t (KeyArray_S32reg_gff_1_SFF_5_n1), .Z0_f (new_AGEMA_signal_7069), .Z1_t (new_AGEMA_signal_7070), .Z1_f (new_AGEMA_signal_7071) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_5_U1 ( .A0_t (KeyArray_S32reg_gff_1_SFF_5_QD), .A0_f (new_AGEMA_signal_5004), .A1_t (new_AGEMA_signal_5005), .A1_f (new_AGEMA_signal_5006), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S32reg_gff_1_SFF_5_n2), .Z0_f (new_AGEMA_signal_7072), .Z1_t (new_AGEMA_signal_7073), .Z1_f (new_AGEMA_signal_7074) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS33ser[5]), .A0_f (new_AGEMA_signal_3835), .A1_t (new_AGEMA_signal_3836), .A1_f (new_AGEMA_signal_3837), .B0_t (KeyArray_outS02ser[5]), .B0_f (new_AGEMA_signal_3298), .B1_t (new_AGEMA_signal_3299), .B1_f (new_AGEMA_signal_3300), .Z0_t (KeyArray_S32reg_gff_1_SFF_5_MUXInst_X), .Z0_f (new_AGEMA_signal_3892), .Z1_t (new_AGEMA_signal_3893), .Z1_f (new_AGEMA_signal_3894) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S32reg_gff_1_SFF_5_MUXInst_X), .B0_f (new_AGEMA_signal_3892), .B1_t (new_AGEMA_signal_3893), .B1_f (new_AGEMA_signal_3894), .Z0_t (KeyArray_S32reg_gff_1_SFF_5_MUXInst_Y), .Z0_f (new_AGEMA_signal_4514), .Z1_t (new_AGEMA_signal_4515), .Z1_f (new_AGEMA_signal_4516) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S32reg_gff_1_SFF_5_MUXInst_Y), .A0_f (new_AGEMA_signal_4514), .A1_t (new_AGEMA_signal_4515), .A1_f (new_AGEMA_signal_4516), .B0_t (KeyArray_outS33ser[5]), .B0_f (new_AGEMA_signal_3835), .B1_t (new_AGEMA_signal_3836), .B1_f (new_AGEMA_signal_3837), .Z0_t (KeyArray_S32reg_gff_1_SFF_5_QD), .Z0_f (new_AGEMA_signal_5004), .Z1_t (new_AGEMA_signal_5005), .Z1_f (new_AGEMA_signal_5006) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S32reg_gff_1_SFF_6_U3 ( .A0_t (KeyArray_S32reg_gff_1_SFF_6_n2), .A0_f (new_AGEMA_signal_7078), .A1_t (new_AGEMA_signal_7079), .A1_f (new_AGEMA_signal_7080), .B0_t (KeyArray_S32reg_gff_1_SFF_6_n1), .B0_f (new_AGEMA_signal_7075), .B1_t (new_AGEMA_signal_7076), .B1_f (new_AGEMA_signal_7077), .Z0_t (KeyArray_outS32ser[6]), .Z0_f (new_AGEMA_signal_3793), .Z1_t (new_AGEMA_signal_3794), .Z1_f (new_AGEMA_signal_3795) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_6_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS32ser[6]), .B0_f (new_AGEMA_signal_3793), .B1_t (new_AGEMA_signal_3794), .B1_f (new_AGEMA_signal_3795), .Z0_t (KeyArray_S32reg_gff_1_SFF_6_n1), .Z0_f (new_AGEMA_signal_7075), .Z1_t (new_AGEMA_signal_7076), .Z1_f (new_AGEMA_signal_7077) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_6_U1 ( .A0_t (KeyArray_S32reg_gff_1_SFF_6_QD), .A0_f (new_AGEMA_signal_5007), .A1_t (new_AGEMA_signal_5008), .A1_f (new_AGEMA_signal_5009), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S32reg_gff_1_SFF_6_n2), .Z0_f (new_AGEMA_signal_7078), .Z1_t (new_AGEMA_signal_7079), .Z1_f (new_AGEMA_signal_7080) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS33ser[6]), .A0_f (new_AGEMA_signal_3841), .A1_t (new_AGEMA_signal_3842), .A1_f (new_AGEMA_signal_3843), .B0_t (KeyArray_outS02ser[6]), .B0_f (new_AGEMA_signal_3307), .B1_t (new_AGEMA_signal_3308), .B1_f (new_AGEMA_signal_3309), .Z0_t (KeyArray_S32reg_gff_1_SFF_6_MUXInst_X), .Z0_f (new_AGEMA_signal_3895), .Z1_t (new_AGEMA_signal_3896), .Z1_f (new_AGEMA_signal_3897) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S32reg_gff_1_SFF_6_MUXInst_X), .B0_f (new_AGEMA_signal_3895), .B1_t (new_AGEMA_signal_3896), .B1_f (new_AGEMA_signal_3897), .Z0_t (KeyArray_S32reg_gff_1_SFF_6_MUXInst_Y), .Z0_f (new_AGEMA_signal_4517), .Z1_t (new_AGEMA_signal_4518), .Z1_f (new_AGEMA_signal_4519) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S32reg_gff_1_SFF_6_MUXInst_Y), .A0_f (new_AGEMA_signal_4517), .A1_t (new_AGEMA_signal_4518), .A1_f (new_AGEMA_signal_4519), .B0_t (KeyArray_outS33ser[6]), .B0_f (new_AGEMA_signal_3841), .B1_t (new_AGEMA_signal_3842), .B1_f (new_AGEMA_signal_3843), .Z0_t (KeyArray_S32reg_gff_1_SFF_6_QD), .Z0_f (new_AGEMA_signal_5007), .Z1_t (new_AGEMA_signal_5008), .Z1_f (new_AGEMA_signal_5009) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S32reg_gff_1_SFF_7_U3 ( .A0_t (KeyArray_S32reg_gff_1_SFF_7_n2), .A0_f (new_AGEMA_signal_7084), .A1_t (new_AGEMA_signal_7085), .A1_f (new_AGEMA_signal_7086), .B0_t (KeyArray_S32reg_gff_1_SFF_7_n1), .B0_f (new_AGEMA_signal_7081), .B1_t (new_AGEMA_signal_7082), .B1_f (new_AGEMA_signal_7083), .Z0_t (KeyArray_outS32ser[7]), .Z0_f (new_AGEMA_signal_3799), .Z1_t (new_AGEMA_signal_3800), .Z1_f (new_AGEMA_signal_3801) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_7_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS32ser[7]), .B0_f (new_AGEMA_signal_3799), .B1_t (new_AGEMA_signal_3800), .B1_f (new_AGEMA_signal_3801), .Z0_t (KeyArray_S32reg_gff_1_SFF_7_n1), .Z0_f (new_AGEMA_signal_7081), .Z1_t (new_AGEMA_signal_7082), .Z1_f (new_AGEMA_signal_7083) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_7_U1 ( .A0_t (KeyArray_S32reg_gff_1_SFF_7_QD), .A0_f (new_AGEMA_signal_5010), .A1_t (new_AGEMA_signal_5011), .A1_f (new_AGEMA_signal_5012), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S32reg_gff_1_SFF_7_n2), .Z0_f (new_AGEMA_signal_7084), .Z1_t (new_AGEMA_signal_7085), .Z1_f (new_AGEMA_signal_7086) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (KeyArray_outS33ser[7]), .A0_f (new_AGEMA_signal_3847), .A1_t (new_AGEMA_signal_3848), .A1_f (new_AGEMA_signal_3849), .B0_t (KeyArray_outS02ser[7]), .B0_f (new_AGEMA_signal_3316), .B1_t (new_AGEMA_signal_3317), .B1_f (new_AGEMA_signal_3318), .Z0_t (KeyArray_S32reg_gff_1_SFF_7_MUXInst_X), .Z0_f (new_AGEMA_signal_3898), .Z1_t (new_AGEMA_signal_3899), .Z1_f (new_AGEMA_signal_3900) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S32reg_gff_1_SFF_7_MUXInst_X), .B0_f (new_AGEMA_signal_3898), .B1_t (new_AGEMA_signal_3899), .B1_f (new_AGEMA_signal_3900), .Z0_t (KeyArray_S32reg_gff_1_SFF_7_MUXInst_Y), .Z0_f (new_AGEMA_signal_4520), .Z1_t (new_AGEMA_signal_4521), .Z1_f (new_AGEMA_signal_4522) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S32reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S32reg_gff_1_SFF_7_MUXInst_Y), .A0_f (new_AGEMA_signal_4520), .A1_t (new_AGEMA_signal_4521), .A1_f (new_AGEMA_signal_4522), .B0_t (KeyArray_outS33ser[7]), .B0_f (new_AGEMA_signal_3847), .B1_t (new_AGEMA_signal_3848), .B1_f (new_AGEMA_signal_3849), .Z0_t (KeyArray_S32reg_gff_1_SFF_7_QD), .Z0_f (new_AGEMA_signal_5010), .Z1_t (new_AGEMA_signal_5011), .Z1_f (new_AGEMA_signal_5012) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S33reg_gff_1_SFF_0_U3 ( .A0_t (KeyArray_S33reg_gff_1_SFF_0_n2), .A0_f (new_AGEMA_signal_7090), .A1_t (new_AGEMA_signal_7091), .A1_f (new_AGEMA_signal_7092), .B0_t (KeyArray_S33reg_gff_1_SFF_0_n1), .B0_f (new_AGEMA_signal_7087), .B1_t (new_AGEMA_signal_7088), .B1_f (new_AGEMA_signal_7089), .Z0_t (KeyArray_outS33ser[0]), .Z0_f (new_AGEMA_signal_3805), .Z1_t (new_AGEMA_signal_3806), .Z1_f (new_AGEMA_signal_3807) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_0_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS33ser[0]), .B0_f (new_AGEMA_signal_3805), .B1_t (new_AGEMA_signal_3806), .B1_f (new_AGEMA_signal_3807), .Z0_t (KeyArray_S33reg_gff_1_SFF_0_n1), .Z0_f (new_AGEMA_signal_7087), .Z1_t (new_AGEMA_signal_7088), .Z1_f (new_AGEMA_signal_7089) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_0_U1 ( .A0_t (KeyArray_S33reg_gff_1_SFF_0_QD), .A0_f (new_AGEMA_signal_5560), .A1_t (new_AGEMA_signal_5561), .A1_f (new_AGEMA_signal_5562), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S33reg_gff_1_SFF_0_n2), .Z0_f (new_AGEMA_signal_7090), .Z1_t (new_AGEMA_signal_7091), .Z1_f (new_AGEMA_signal_7092) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_0_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS33ser[0]), .A0_f (new_AGEMA_signal_5013), .A1_t (new_AGEMA_signal_5014), .A1_f (new_AGEMA_signal_5015), .B0_t (KeyArray_outS03ser[0]), .B0_f (new_AGEMA_signal_3325), .B1_t (new_AGEMA_signal_3326), .B1_f (new_AGEMA_signal_3327), .Z0_t (KeyArray_S33reg_gff_1_SFF_0_MUXInst_X), .Z0_f (new_AGEMA_signal_5223), .Z1_t (new_AGEMA_signal_5224), .Z1_f (new_AGEMA_signal_5225) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_0_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S33reg_gff_1_SFF_0_MUXInst_X), .B0_f (new_AGEMA_signal_5223), .B1_t (new_AGEMA_signal_5224), .B1_f (new_AGEMA_signal_5225), .Z0_t (KeyArray_S33reg_gff_1_SFF_0_MUXInst_Y), .Z0_f (new_AGEMA_signal_5407), .Z1_t (new_AGEMA_signal_5408), .Z1_f (new_AGEMA_signal_5409) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_0_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S33reg_gff_1_SFF_0_MUXInst_Y), .A0_f (new_AGEMA_signal_5407), .A1_t (new_AGEMA_signal_5408), .A1_f (new_AGEMA_signal_5409), .B0_t (KeyArray_inS33ser[0]), .B0_f (new_AGEMA_signal_5013), .B1_t (new_AGEMA_signal_5014), .B1_f (new_AGEMA_signal_5015), .Z0_t (KeyArray_S33reg_gff_1_SFF_0_QD), .Z0_f (new_AGEMA_signal_5560), .Z1_t (new_AGEMA_signal_5561), .Z1_f (new_AGEMA_signal_5562) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S33reg_gff_1_SFF_1_U3 ( .A0_t (KeyArray_S33reg_gff_1_SFF_1_n2), .A0_f (new_AGEMA_signal_7096), .A1_t (new_AGEMA_signal_7097), .A1_f (new_AGEMA_signal_7098), .B0_t (KeyArray_S33reg_gff_1_SFF_1_n1), .B0_f (new_AGEMA_signal_7093), .B1_t (new_AGEMA_signal_7094), .B1_f (new_AGEMA_signal_7095), .Z0_t (KeyArray_outS33ser[1]), .Z0_f (new_AGEMA_signal_3811), .Z1_t (new_AGEMA_signal_3812), .Z1_f (new_AGEMA_signal_3813) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_1_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS33ser[1]), .B0_f (new_AGEMA_signal_3811), .B1_t (new_AGEMA_signal_3812), .B1_f (new_AGEMA_signal_3813), .Z0_t (KeyArray_S33reg_gff_1_SFF_1_n1), .Z0_f (new_AGEMA_signal_7093), .Z1_t (new_AGEMA_signal_7094), .Z1_f (new_AGEMA_signal_7095) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_1_U1 ( .A0_t (KeyArray_S33reg_gff_1_SFF_1_QD), .A0_f (new_AGEMA_signal_5563), .A1_t (new_AGEMA_signal_5564), .A1_f (new_AGEMA_signal_5565), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S33reg_gff_1_SFF_1_n2), .Z0_f (new_AGEMA_signal_7096), .Z1_t (new_AGEMA_signal_7097), .Z1_f (new_AGEMA_signal_7098) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_1_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS33ser[1]), .A0_f (new_AGEMA_signal_5016), .A1_t (new_AGEMA_signal_5017), .A1_f (new_AGEMA_signal_5018), .B0_t (KeyArray_outS03ser[1]), .B0_f (new_AGEMA_signal_3334), .B1_t (new_AGEMA_signal_3335), .B1_f (new_AGEMA_signal_3336), .Z0_t (KeyArray_S33reg_gff_1_SFF_1_MUXInst_X), .Z0_f (new_AGEMA_signal_5226), .Z1_t (new_AGEMA_signal_5227), .Z1_f (new_AGEMA_signal_5228) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_1_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S33reg_gff_1_SFF_1_MUXInst_X), .B0_f (new_AGEMA_signal_5226), .B1_t (new_AGEMA_signal_5227), .B1_f (new_AGEMA_signal_5228), .Z0_t (KeyArray_S33reg_gff_1_SFF_1_MUXInst_Y), .Z0_f (new_AGEMA_signal_5410), .Z1_t (new_AGEMA_signal_5411), .Z1_f (new_AGEMA_signal_5412) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_1_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S33reg_gff_1_SFF_1_MUXInst_Y), .A0_f (new_AGEMA_signal_5410), .A1_t (new_AGEMA_signal_5411), .A1_f (new_AGEMA_signal_5412), .B0_t (KeyArray_inS33ser[1]), .B0_f (new_AGEMA_signal_5016), .B1_t (new_AGEMA_signal_5017), .B1_f (new_AGEMA_signal_5018), .Z0_t (KeyArray_S33reg_gff_1_SFF_1_QD), .Z0_f (new_AGEMA_signal_5563), .Z1_t (new_AGEMA_signal_5564), .Z1_f (new_AGEMA_signal_5565) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S33reg_gff_1_SFF_2_U3 ( .A0_t (KeyArray_S33reg_gff_1_SFF_2_n2), .A0_f (new_AGEMA_signal_7102), .A1_t (new_AGEMA_signal_7103), .A1_f (new_AGEMA_signal_7104), .B0_t (KeyArray_S33reg_gff_1_SFF_2_n1), .B0_f (new_AGEMA_signal_7099), .B1_t (new_AGEMA_signal_7100), .B1_f (new_AGEMA_signal_7101), .Z0_t (KeyArray_outS33ser[2]), .Z0_f (new_AGEMA_signal_3817), .Z1_t (new_AGEMA_signal_3818), .Z1_f (new_AGEMA_signal_3819) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_2_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS33ser[2]), .B0_f (new_AGEMA_signal_3817), .B1_t (new_AGEMA_signal_3818), .B1_f (new_AGEMA_signal_3819), .Z0_t (KeyArray_S33reg_gff_1_SFF_2_n1), .Z0_f (new_AGEMA_signal_7099), .Z1_t (new_AGEMA_signal_7100), .Z1_f (new_AGEMA_signal_7101) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_2_U1 ( .A0_t (KeyArray_S33reg_gff_1_SFF_2_QD), .A0_f (new_AGEMA_signal_5566), .A1_t (new_AGEMA_signal_5567), .A1_f (new_AGEMA_signal_5568), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S33reg_gff_1_SFF_2_n2), .Z0_f (new_AGEMA_signal_7102), .Z1_t (new_AGEMA_signal_7103), .Z1_f (new_AGEMA_signal_7104) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_2_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS33ser[2]), .A0_f (new_AGEMA_signal_5019), .A1_t (new_AGEMA_signal_5020), .A1_f (new_AGEMA_signal_5021), .B0_t (KeyArray_outS03ser[2]), .B0_f (new_AGEMA_signal_3343), .B1_t (new_AGEMA_signal_3344), .B1_f (new_AGEMA_signal_3345), .Z0_t (KeyArray_S33reg_gff_1_SFF_2_MUXInst_X), .Z0_f (new_AGEMA_signal_5229), .Z1_t (new_AGEMA_signal_5230), .Z1_f (new_AGEMA_signal_5231) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_2_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S33reg_gff_1_SFF_2_MUXInst_X), .B0_f (new_AGEMA_signal_5229), .B1_t (new_AGEMA_signal_5230), .B1_f (new_AGEMA_signal_5231), .Z0_t (KeyArray_S33reg_gff_1_SFF_2_MUXInst_Y), .Z0_f (new_AGEMA_signal_5413), .Z1_t (new_AGEMA_signal_5414), .Z1_f (new_AGEMA_signal_5415) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_2_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S33reg_gff_1_SFF_2_MUXInst_Y), .A0_f (new_AGEMA_signal_5413), .A1_t (new_AGEMA_signal_5414), .A1_f (new_AGEMA_signal_5415), .B0_t (KeyArray_inS33ser[2]), .B0_f (new_AGEMA_signal_5019), .B1_t (new_AGEMA_signal_5020), .B1_f (new_AGEMA_signal_5021), .Z0_t (KeyArray_S33reg_gff_1_SFF_2_QD), .Z0_f (new_AGEMA_signal_5566), .Z1_t (new_AGEMA_signal_5567), .Z1_f (new_AGEMA_signal_5568) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S33reg_gff_1_SFF_3_U3 ( .A0_t (KeyArray_S33reg_gff_1_SFF_3_n2), .A0_f (new_AGEMA_signal_7108), .A1_t (new_AGEMA_signal_7109), .A1_f (new_AGEMA_signal_7110), .B0_t (KeyArray_S33reg_gff_1_SFF_3_n1), .B0_f (new_AGEMA_signal_7105), .B1_t (new_AGEMA_signal_7106), .B1_f (new_AGEMA_signal_7107), .Z0_t (KeyArray_outS33ser[3]), .Z0_f (new_AGEMA_signal_3823), .Z1_t (new_AGEMA_signal_3824), .Z1_f (new_AGEMA_signal_3825) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_3_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS33ser[3]), .B0_f (new_AGEMA_signal_3823), .B1_t (new_AGEMA_signal_3824), .B1_f (new_AGEMA_signal_3825), .Z0_t (KeyArray_S33reg_gff_1_SFF_3_n1), .Z0_f (new_AGEMA_signal_7105), .Z1_t (new_AGEMA_signal_7106), .Z1_f (new_AGEMA_signal_7107) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_3_U1 ( .A0_t (KeyArray_S33reg_gff_1_SFF_3_QD), .A0_f (new_AGEMA_signal_5569), .A1_t (new_AGEMA_signal_5570), .A1_f (new_AGEMA_signal_5571), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S33reg_gff_1_SFF_3_n2), .Z0_f (new_AGEMA_signal_7108), .Z1_t (new_AGEMA_signal_7109), .Z1_f (new_AGEMA_signal_7110) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_3_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS33ser[3]), .A0_f (new_AGEMA_signal_5022), .A1_t (new_AGEMA_signal_5023), .A1_f (new_AGEMA_signal_5024), .B0_t (KeyArray_outS03ser[3]), .B0_f (new_AGEMA_signal_3352), .B1_t (new_AGEMA_signal_3353), .B1_f (new_AGEMA_signal_3354), .Z0_t (KeyArray_S33reg_gff_1_SFF_3_MUXInst_X), .Z0_f (new_AGEMA_signal_5232), .Z1_t (new_AGEMA_signal_5233), .Z1_f (new_AGEMA_signal_5234) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_3_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S33reg_gff_1_SFF_3_MUXInst_X), .B0_f (new_AGEMA_signal_5232), .B1_t (new_AGEMA_signal_5233), .B1_f (new_AGEMA_signal_5234), .Z0_t (KeyArray_S33reg_gff_1_SFF_3_MUXInst_Y), .Z0_f (new_AGEMA_signal_5416), .Z1_t (new_AGEMA_signal_5417), .Z1_f (new_AGEMA_signal_5418) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_3_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S33reg_gff_1_SFF_3_MUXInst_Y), .A0_f (new_AGEMA_signal_5416), .A1_t (new_AGEMA_signal_5417), .A1_f (new_AGEMA_signal_5418), .B0_t (KeyArray_inS33ser[3]), .B0_f (new_AGEMA_signal_5022), .B1_t (new_AGEMA_signal_5023), .B1_f (new_AGEMA_signal_5024), .Z0_t (KeyArray_S33reg_gff_1_SFF_3_QD), .Z0_f (new_AGEMA_signal_5569), .Z1_t (new_AGEMA_signal_5570), .Z1_f (new_AGEMA_signal_5571) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S33reg_gff_1_SFF_4_U3 ( .A0_t (KeyArray_S33reg_gff_1_SFF_4_n2), .A0_f (new_AGEMA_signal_7114), .A1_t (new_AGEMA_signal_7115), .A1_f (new_AGEMA_signal_7116), .B0_t (KeyArray_S33reg_gff_1_SFF_4_n1), .B0_f (new_AGEMA_signal_7111), .B1_t (new_AGEMA_signal_7112), .B1_f (new_AGEMA_signal_7113), .Z0_t (KeyArray_outS33ser[4]), .Z0_f (new_AGEMA_signal_3829), .Z1_t (new_AGEMA_signal_3830), .Z1_f (new_AGEMA_signal_3831) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_4_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS33ser[4]), .B0_f (new_AGEMA_signal_3829), .B1_t (new_AGEMA_signal_3830), .B1_f (new_AGEMA_signal_3831), .Z0_t (KeyArray_S33reg_gff_1_SFF_4_n1), .Z0_f (new_AGEMA_signal_7111), .Z1_t (new_AGEMA_signal_7112), .Z1_f (new_AGEMA_signal_7113) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_4_U1 ( .A0_t (KeyArray_S33reg_gff_1_SFF_4_QD), .A0_f (new_AGEMA_signal_5572), .A1_t (new_AGEMA_signal_5573), .A1_f (new_AGEMA_signal_5574), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S33reg_gff_1_SFF_4_n2), .Z0_f (new_AGEMA_signal_7114), .Z1_t (new_AGEMA_signal_7115), .Z1_f (new_AGEMA_signal_7116) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_4_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS33ser[4]), .A0_f (new_AGEMA_signal_5025), .A1_t (new_AGEMA_signal_5026), .A1_f (new_AGEMA_signal_5027), .B0_t (KeyArray_outS03ser[4]), .B0_f (new_AGEMA_signal_3361), .B1_t (new_AGEMA_signal_3362), .B1_f (new_AGEMA_signal_3363), .Z0_t (KeyArray_S33reg_gff_1_SFF_4_MUXInst_X), .Z0_f (new_AGEMA_signal_5235), .Z1_t (new_AGEMA_signal_5236), .Z1_f (new_AGEMA_signal_5237) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_4_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S33reg_gff_1_SFF_4_MUXInst_X), .B0_f (new_AGEMA_signal_5235), .B1_t (new_AGEMA_signal_5236), .B1_f (new_AGEMA_signal_5237), .Z0_t (KeyArray_S33reg_gff_1_SFF_4_MUXInst_Y), .Z0_f (new_AGEMA_signal_5419), .Z1_t (new_AGEMA_signal_5420), .Z1_f (new_AGEMA_signal_5421) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_4_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S33reg_gff_1_SFF_4_MUXInst_Y), .A0_f (new_AGEMA_signal_5419), .A1_t (new_AGEMA_signal_5420), .A1_f (new_AGEMA_signal_5421), .B0_t (KeyArray_inS33ser[4]), .B0_f (new_AGEMA_signal_5025), .B1_t (new_AGEMA_signal_5026), .B1_f (new_AGEMA_signal_5027), .Z0_t (KeyArray_S33reg_gff_1_SFF_4_QD), .Z0_f (new_AGEMA_signal_5572), .Z1_t (new_AGEMA_signal_5573), .Z1_f (new_AGEMA_signal_5574) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S33reg_gff_1_SFF_5_U3 ( .A0_t (KeyArray_S33reg_gff_1_SFF_5_n2), .A0_f (new_AGEMA_signal_7120), .A1_t (new_AGEMA_signal_7121), .A1_f (new_AGEMA_signal_7122), .B0_t (KeyArray_S33reg_gff_1_SFF_5_n1), .B0_f (new_AGEMA_signal_7117), .B1_t (new_AGEMA_signal_7118), .B1_f (new_AGEMA_signal_7119), .Z0_t (KeyArray_outS33ser[5]), .Z0_f (new_AGEMA_signal_3835), .Z1_t (new_AGEMA_signal_3836), .Z1_f (new_AGEMA_signal_3837) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_5_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS33ser[5]), .B0_f (new_AGEMA_signal_3835), .B1_t (new_AGEMA_signal_3836), .B1_f (new_AGEMA_signal_3837), .Z0_t (KeyArray_S33reg_gff_1_SFF_5_n1), .Z0_f (new_AGEMA_signal_7117), .Z1_t (new_AGEMA_signal_7118), .Z1_f (new_AGEMA_signal_7119) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_5_U1 ( .A0_t (KeyArray_S33reg_gff_1_SFF_5_QD), .A0_f (new_AGEMA_signal_5575), .A1_t (new_AGEMA_signal_5576), .A1_f (new_AGEMA_signal_5577), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S33reg_gff_1_SFF_5_n2), .Z0_f (new_AGEMA_signal_7120), .Z1_t (new_AGEMA_signal_7121), .Z1_f (new_AGEMA_signal_7122) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_5_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS33ser[5]), .A0_f (new_AGEMA_signal_5028), .A1_t (new_AGEMA_signal_5029), .A1_f (new_AGEMA_signal_5030), .B0_t (KeyArray_outS03ser[5]), .B0_f (new_AGEMA_signal_3370), .B1_t (new_AGEMA_signal_3371), .B1_f (new_AGEMA_signal_3372), .Z0_t (KeyArray_S33reg_gff_1_SFF_5_MUXInst_X), .Z0_f (new_AGEMA_signal_5238), .Z1_t (new_AGEMA_signal_5239), .Z1_f (new_AGEMA_signal_5240) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_5_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S33reg_gff_1_SFF_5_MUXInst_X), .B0_f (new_AGEMA_signal_5238), .B1_t (new_AGEMA_signal_5239), .B1_f (new_AGEMA_signal_5240), .Z0_t (KeyArray_S33reg_gff_1_SFF_5_MUXInst_Y), .Z0_f (new_AGEMA_signal_5422), .Z1_t (new_AGEMA_signal_5423), .Z1_f (new_AGEMA_signal_5424) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_5_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S33reg_gff_1_SFF_5_MUXInst_Y), .A0_f (new_AGEMA_signal_5422), .A1_t (new_AGEMA_signal_5423), .A1_f (new_AGEMA_signal_5424), .B0_t (KeyArray_inS33ser[5]), .B0_f (new_AGEMA_signal_5028), .B1_t (new_AGEMA_signal_5029), .B1_f (new_AGEMA_signal_5030), .Z0_t (KeyArray_S33reg_gff_1_SFF_5_QD), .Z0_f (new_AGEMA_signal_5575), .Z1_t (new_AGEMA_signal_5576), .Z1_f (new_AGEMA_signal_5577) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S33reg_gff_1_SFF_6_U3 ( .A0_t (KeyArray_S33reg_gff_1_SFF_6_n2), .A0_f (new_AGEMA_signal_7126), .A1_t (new_AGEMA_signal_7127), .A1_f (new_AGEMA_signal_7128), .B0_t (KeyArray_S33reg_gff_1_SFF_6_n1), .B0_f (new_AGEMA_signal_7123), .B1_t (new_AGEMA_signal_7124), .B1_f (new_AGEMA_signal_7125), .Z0_t (KeyArray_outS33ser[6]), .Z0_f (new_AGEMA_signal_3841), .Z1_t (new_AGEMA_signal_3842), .Z1_f (new_AGEMA_signal_3843) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_6_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS33ser[6]), .B0_f (new_AGEMA_signal_3841), .B1_t (new_AGEMA_signal_3842), .B1_f (new_AGEMA_signal_3843), .Z0_t (KeyArray_S33reg_gff_1_SFF_6_n1), .Z0_f (new_AGEMA_signal_7123), .Z1_t (new_AGEMA_signal_7124), .Z1_f (new_AGEMA_signal_7125) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_6_U1 ( .A0_t (KeyArray_S33reg_gff_1_SFF_6_QD), .A0_f (new_AGEMA_signal_5578), .A1_t (new_AGEMA_signal_5579), .A1_f (new_AGEMA_signal_5580), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S33reg_gff_1_SFF_6_n2), .Z0_f (new_AGEMA_signal_7126), .Z1_t (new_AGEMA_signal_7127), .Z1_f (new_AGEMA_signal_7128) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_6_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS33ser[6]), .A0_f (new_AGEMA_signal_5031), .A1_t (new_AGEMA_signal_5032), .A1_f (new_AGEMA_signal_5033), .B0_t (KeyArray_outS03ser[6]), .B0_f (new_AGEMA_signal_3379), .B1_t (new_AGEMA_signal_3380), .B1_f (new_AGEMA_signal_3381), .Z0_t (KeyArray_S33reg_gff_1_SFF_6_MUXInst_X), .Z0_f (new_AGEMA_signal_5241), .Z1_t (new_AGEMA_signal_5242), .Z1_f (new_AGEMA_signal_5243) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_6_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S33reg_gff_1_SFF_6_MUXInst_X), .B0_f (new_AGEMA_signal_5241), .B1_t (new_AGEMA_signal_5242), .B1_f (new_AGEMA_signal_5243), .Z0_t (KeyArray_S33reg_gff_1_SFF_6_MUXInst_Y), .Z0_f (new_AGEMA_signal_5425), .Z1_t (new_AGEMA_signal_5426), .Z1_f (new_AGEMA_signal_5427) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_6_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S33reg_gff_1_SFF_6_MUXInst_Y), .A0_f (new_AGEMA_signal_5425), .A1_t (new_AGEMA_signal_5426), .A1_f (new_AGEMA_signal_5427), .B0_t (KeyArray_inS33ser[6]), .B0_f (new_AGEMA_signal_5031), .B1_t (new_AGEMA_signal_5032), .B1_f (new_AGEMA_signal_5033), .Z0_t (KeyArray_S33reg_gff_1_SFF_6_QD), .Z0_f (new_AGEMA_signal_5578), .Z1_t (new_AGEMA_signal_5579), .Z1_f (new_AGEMA_signal_5580) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1)) KeyArray_S33reg_gff_1_SFF_7_U3 ( .A0_t (KeyArray_S33reg_gff_1_SFF_7_n2), .A0_f (new_AGEMA_signal_7132), .A1_t (new_AGEMA_signal_7133), .A1_f (new_AGEMA_signal_7134), .B0_t (KeyArray_S33reg_gff_1_SFF_7_n1), .B0_f (new_AGEMA_signal_7129), .B1_t (new_AGEMA_signal_7130), .B1_f (new_AGEMA_signal_7131), .Z0_t (KeyArray_outS33ser[7]), .Z0_f (new_AGEMA_signal_3847), .Z1_t (new_AGEMA_signal_3848), .Z1_f (new_AGEMA_signal_3849) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_7_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (enKS), .A1_f (new_AGEMA_signal_5916), .B0_t (KeyArray_outS33ser[7]), .B0_f (new_AGEMA_signal_3847), .B1_t (new_AGEMA_signal_3848), .B1_f (new_AGEMA_signal_3849), .Z0_t (KeyArray_S33reg_gff_1_SFF_7_n1), .Z0_f (new_AGEMA_signal_7129), .Z1_t (new_AGEMA_signal_7130), .Z1_f (new_AGEMA_signal_7131) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_7_U1 ( .A0_t (KeyArray_S33reg_gff_1_SFF_7_QD), .A0_f (new_AGEMA_signal_5581), .A1_t (new_AGEMA_signal_5582), .A1_f (new_AGEMA_signal_5583), .B0_t (1'b0), .B0_f (1'b1), .B1_t (enKS), .B1_f (new_AGEMA_signal_5916), .Z0_t (KeyArray_S33reg_gff_1_SFF_7_n2), .Z0_f (new_AGEMA_signal_7132), .Z1_t (new_AGEMA_signal_7133), .Z1_f (new_AGEMA_signal_7134) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_7_MUXInst_XOR1_U1 ( .A0_t (KeyArray_inS33ser[7]), .A0_f (new_AGEMA_signal_5034), .A1_t (new_AGEMA_signal_5035), .A1_f (new_AGEMA_signal_5036), .B0_t (KeyArray_outS03ser[7]), .B0_f (new_AGEMA_signal_3388), .B1_t (new_AGEMA_signal_3389), .B1_f (new_AGEMA_signal_3390), .Z0_t (KeyArray_S33reg_gff_1_SFF_7_MUXInst_X), .Z0_f (new_AGEMA_signal_5244), .Z1_t (new_AGEMA_signal_5245), .Z1_f (new_AGEMA_signal_5246) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_7_MUXInst_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (KeyArray_S33reg_gff_1_SFF_7_MUXInst_X), .B0_f (new_AGEMA_signal_5244), .B1_t (new_AGEMA_signal_5245), .B1_f (new_AGEMA_signal_5246), .Z0_t (KeyArray_S33reg_gff_1_SFF_7_MUXInst_Y), .Z0_f (new_AGEMA_signal_5428), .Z1_t (new_AGEMA_signal_5429), .Z1_f (new_AGEMA_signal_5430) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_S33reg_gff_1_SFF_7_MUXInst_XOR2_U1 ( .A0_t (KeyArray_S33reg_gff_1_SFF_7_MUXInst_Y), .A0_f (new_AGEMA_signal_5428), .A1_t (new_AGEMA_signal_5429), .A1_f (new_AGEMA_signal_5430), .B0_t (KeyArray_inS33ser[7]), .B0_f (new_AGEMA_signal_5034), .B1_t (new_AGEMA_signal_5035), .B1_f (new_AGEMA_signal_5036), .Z0_t (KeyArray_S33reg_gff_1_SFF_7_QD), .Z0_f (new_AGEMA_signal_5581), .Z1_t (new_AGEMA_signal_5582), .Z1_f (new_AGEMA_signal_5583) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_0_XOR1_U1 ( .A0_t (KeyArray_outS01ser_0_), .A0_f (new_AGEMA_signal_3247), .A1_t (new_AGEMA_signal_3248), .A1_f (new_AGEMA_signal_3249), .B0_t (KeyArray_outS01ser_XOR_00[0]), .B0_f (new_AGEMA_signal_3250), .B1_t (new_AGEMA_signal_3251), .B1_f (new_AGEMA_signal_3252), .Z0_t (KeyArray_MUX_inS00ser_mux_inst_0_X), .Z0_f (new_AGEMA_signal_4523), .Z1_t (new_AGEMA_signal_4524), .Z1_f (new_AGEMA_signal_4525) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_0_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (KeyArray_nReset_selXOR), .A1_f (new_AGEMA_signal_5406), .B0_t (KeyArray_MUX_inS00ser_mux_inst_0_X), .B0_f (new_AGEMA_signal_4523), .B1_t (new_AGEMA_signal_4524), .B1_f (new_AGEMA_signal_4525), .Z0_t (KeyArray_MUX_inS00ser_mux_inst_0_Y), .Z0_f (new_AGEMA_signal_5584), .Z1_t (new_AGEMA_signal_5585), .Z1_f (new_AGEMA_signal_5586) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_0_XOR2_U1 ( .A0_t (KeyArray_MUX_inS00ser_mux_inst_0_Y), .A0_f (new_AGEMA_signal_5584), .A1_t (new_AGEMA_signal_5585), .A1_f (new_AGEMA_signal_5586), .B0_t (KeyArray_outS01ser_0_), .B0_f (new_AGEMA_signal_3247), .B1_t (new_AGEMA_signal_3248), .B1_f (new_AGEMA_signal_3249), .Z0_t (KeyArray_inS00ser[0]), .Z0_f (new_AGEMA_signal_5714), .Z1_t (new_AGEMA_signal_5715), .Z1_f (new_AGEMA_signal_5716) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_1_XOR1_U1 ( .A0_t (KeyArray_outS01ser_1_), .A0_f (new_AGEMA_signal_3241), .A1_t (new_AGEMA_signal_3242), .A1_f (new_AGEMA_signal_3243), .B0_t (KeyArray_outS01ser_XOR_00[1]), .B0_f (new_AGEMA_signal_3244), .B1_t (new_AGEMA_signal_3245), .B1_f (new_AGEMA_signal_3246), .Z0_t (KeyArray_MUX_inS00ser_mux_inst_1_X), .Z0_f (new_AGEMA_signal_4526), .Z1_t (new_AGEMA_signal_4527), .Z1_f (new_AGEMA_signal_4528) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (KeyArray_nReset_selXOR), .A1_f (new_AGEMA_signal_5406), .B0_t (KeyArray_MUX_inS00ser_mux_inst_1_X), .B0_f (new_AGEMA_signal_4526), .B1_t (new_AGEMA_signal_4527), .B1_f (new_AGEMA_signal_4528), .Z0_t (KeyArray_MUX_inS00ser_mux_inst_1_Y), .Z0_f (new_AGEMA_signal_5587), .Z1_t (new_AGEMA_signal_5588), .Z1_f (new_AGEMA_signal_5589) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_1_XOR2_U1 ( .A0_t (KeyArray_MUX_inS00ser_mux_inst_1_Y), .A0_f (new_AGEMA_signal_5587), .A1_t (new_AGEMA_signal_5588), .A1_f (new_AGEMA_signal_5589), .B0_t (KeyArray_outS01ser_1_), .B0_f (new_AGEMA_signal_3241), .B1_t (new_AGEMA_signal_3242), .B1_f (new_AGEMA_signal_3243), .Z0_t (KeyArray_inS00ser[1]), .Z0_f (new_AGEMA_signal_5717), .Z1_t (new_AGEMA_signal_5718), .Z1_f (new_AGEMA_signal_5719) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_2_XOR1_U1 ( .A0_t (KeyArray_outS01ser_2_), .A0_f (new_AGEMA_signal_3235), .A1_t (new_AGEMA_signal_3236), .A1_f (new_AGEMA_signal_3237), .B0_t (KeyArray_outS01ser_XOR_00[2]), .B0_f (new_AGEMA_signal_3238), .B1_t (new_AGEMA_signal_3239), .B1_f (new_AGEMA_signal_3240), .Z0_t (KeyArray_MUX_inS00ser_mux_inst_2_X), .Z0_f (new_AGEMA_signal_4529), .Z1_t (new_AGEMA_signal_4530), .Z1_f (new_AGEMA_signal_4531) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_2_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (KeyArray_nReset_selXOR), .A1_f (new_AGEMA_signal_5406), .B0_t (KeyArray_MUX_inS00ser_mux_inst_2_X), .B0_f (new_AGEMA_signal_4529), .B1_t (new_AGEMA_signal_4530), .B1_f (new_AGEMA_signal_4531), .Z0_t (KeyArray_MUX_inS00ser_mux_inst_2_Y), .Z0_f (new_AGEMA_signal_5590), .Z1_t (new_AGEMA_signal_5591), .Z1_f (new_AGEMA_signal_5592) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_2_XOR2_U1 ( .A0_t (KeyArray_MUX_inS00ser_mux_inst_2_Y), .A0_f (new_AGEMA_signal_5590), .A1_t (new_AGEMA_signal_5591), .A1_f (new_AGEMA_signal_5592), .B0_t (KeyArray_outS01ser_2_), .B0_f (new_AGEMA_signal_3235), .B1_t (new_AGEMA_signal_3236), .B1_f (new_AGEMA_signal_3237), .Z0_t (KeyArray_inS00ser[2]), .Z0_f (new_AGEMA_signal_5720), .Z1_t (new_AGEMA_signal_5721), .Z1_f (new_AGEMA_signal_5722) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_3_XOR1_U1 ( .A0_t (KeyArray_outS01ser_3_), .A0_f (new_AGEMA_signal_3229), .A1_t (new_AGEMA_signal_3230), .A1_f (new_AGEMA_signal_3231), .B0_t (KeyArray_outS01ser_XOR_00[3]), .B0_f (new_AGEMA_signal_3232), .B1_t (new_AGEMA_signal_3233), .B1_f (new_AGEMA_signal_3234), .Z0_t (KeyArray_MUX_inS00ser_mux_inst_3_X), .Z0_f (new_AGEMA_signal_4532), .Z1_t (new_AGEMA_signal_4533), .Z1_f (new_AGEMA_signal_4534) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_3_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (KeyArray_nReset_selXOR), .A1_f (new_AGEMA_signal_5406), .B0_t (KeyArray_MUX_inS00ser_mux_inst_3_X), .B0_f (new_AGEMA_signal_4532), .B1_t (new_AGEMA_signal_4533), .B1_f (new_AGEMA_signal_4534), .Z0_t (KeyArray_MUX_inS00ser_mux_inst_3_Y), .Z0_f (new_AGEMA_signal_5593), .Z1_t (new_AGEMA_signal_5594), .Z1_f (new_AGEMA_signal_5595) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_3_XOR2_U1 ( .A0_t (KeyArray_MUX_inS00ser_mux_inst_3_Y), .A0_f (new_AGEMA_signal_5593), .A1_t (new_AGEMA_signal_5594), .A1_f (new_AGEMA_signal_5595), .B0_t (KeyArray_outS01ser_3_), .B0_f (new_AGEMA_signal_3229), .B1_t (new_AGEMA_signal_3230), .B1_f (new_AGEMA_signal_3231), .Z0_t (KeyArray_inS00ser[3]), .Z0_f (new_AGEMA_signal_5723), .Z1_t (new_AGEMA_signal_5724), .Z1_f (new_AGEMA_signal_5725) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_4_XOR1_U1 ( .A0_t (KeyArray_outS01ser_4_), .A0_f (new_AGEMA_signal_3223), .A1_t (new_AGEMA_signal_3224), .A1_f (new_AGEMA_signal_3225), .B0_t (KeyArray_outS01ser_XOR_00[4]), .B0_f (new_AGEMA_signal_3226), .B1_t (new_AGEMA_signal_3227), .B1_f (new_AGEMA_signal_3228), .Z0_t (KeyArray_MUX_inS00ser_mux_inst_4_X), .Z0_f (new_AGEMA_signal_4535), .Z1_t (new_AGEMA_signal_4536), .Z1_f (new_AGEMA_signal_4537) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_4_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (KeyArray_nReset_selXOR), .A1_f (new_AGEMA_signal_5406), .B0_t (KeyArray_MUX_inS00ser_mux_inst_4_X), .B0_f (new_AGEMA_signal_4535), .B1_t (new_AGEMA_signal_4536), .B1_f (new_AGEMA_signal_4537), .Z0_t (KeyArray_MUX_inS00ser_mux_inst_4_Y), .Z0_f (new_AGEMA_signal_5596), .Z1_t (new_AGEMA_signal_5597), .Z1_f (new_AGEMA_signal_5598) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_4_XOR2_U1 ( .A0_t (KeyArray_MUX_inS00ser_mux_inst_4_Y), .A0_f (new_AGEMA_signal_5596), .A1_t (new_AGEMA_signal_5597), .A1_f (new_AGEMA_signal_5598), .B0_t (KeyArray_outS01ser_4_), .B0_f (new_AGEMA_signal_3223), .B1_t (new_AGEMA_signal_3224), .B1_f (new_AGEMA_signal_3225), .Z0_t (KeyArray_inS00ser[4]), .Z0_f (new_AGEMA_signal_5726), .Z1_t (new_AGEMA_signal_5727), .Z1_f (new_AGEMA_signal_5728) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_5_XOR1_U1 ( .A0_t (KeyArray_outS01ser_5_), .A0_f (new_AGEMA_signal_3217), .A1_t (new_AGEMA_signal_3218), .A1_f (new_AGEMA_signal_3219), .B0_t (KeyArray_outS01ser_XOR_00[5]), .B0_f (new_AGEMA_signal_3220), .B1_t (new_AGEMA_signal_3221), .B1_f (new_AGEMA_signal_3222), .Z0_t (KeyArray_MUX_inS00ser_mux_inst_5_X), .Z0_f (new_AGEMA_signal_4538), .Z1_t (new_AGEMA_signal_4539), .Z1_f (new_AGEMA_signal_4540) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_5_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (KeyArray_nReset_selXOR), .A1_f (new_AGEMA_signal_5406), .B0_t (KeyArray_MUX_inS00ser_mux_inst_5_X), .B0_f (new_AGEMA_signal_4538), .B1_t (new_AGEMA_signal_4539), .B1_f (new_AGEMA_signal_4540), .Z0_t (KeyArray_MUX_inS00ser_mux_inst_5_Y), .Z0_f (new_AGEMA_signal_5599), .Z1_t (new_AGEMA_signal_5600), .Z1_f (new_AGEMA_signal_5601) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_5_XOR2_U1 ( .A0_t (KeyArray_MUX_inS00ser_mux_inst_5_Y), .A0_f (new_AGEMA_signal_5599), .A1_t (new_AGEMA_signal_5600), .A1_f (new_AGEMA_signal_5601), .B0_t (KeyArray_outS01ser_5_), .B0_f (new_AGEMA_signal_3217), .B1_t (new_AGEMA_signal_3218), .B1_f (new_AGEMA_signal_3219), .Z0_t (KeyArray_inS00ser[5]), .Z0_f (new_AGEMA_signal_5729), .Z1_t (new_AGEMA_signal_5730), .Z1_f (new_AGEMA_signal_5731) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_6_XOR1_U1 ( .A0_t (KeyArray_outS01ser_6_), .A0_f (new_AGEMA_signal_3211), .A1_t (new_AGEMA_signal_3212), .A1_f (new_AGEMA_signal_3213), .B0_t (KeyArray_outS01ser_XOR_00[6]), .B0_f (new_AGEMA_signal_3214), .B1_t (new_AGEMA_signal_3215), .B1_f (new_AGEMA_signal_3216), .Z0_t (KeyArray_MUX_inS00ser_mux_inst_6_X), .Z0_f (new_AGEMA_signal_4541), .Z1_t (new_AGEMA_signal_4542), .Z1_f (new_AGEMA_signal_4543) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_6_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (KeyArray_nReset_selXOR), .A1_f (new_AGEMA_signal_5406), .B0_t (KeyArray_MUX_inS00ser_mux_inst_6_X), .B0_f (new_AGEMA_signal_4541), .B1_t (new_AGEMA_signal_4542), .B1_f (new_AGEMA_signal_4543), .Z0_t (KeyArray_MUX_inS00ser_mux_inst_6_Y), .Z0_f (new_AGEMA_signal_5602), .Z1_t (new_AGEMA_signal_5603), .Z1_f (new_AGEMA_signal_5604) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_6_XOR2_U1 ( .A0_t (KeyArray_MUX_inS00ser_mux_inst_6_Y), .A0_f (new_AGEMA_signal_5602), .A1_t (new_AGEMA_signal_5603), .A1_f (new_AGEMA_signal_5604), .B0_t (KeyArray_outS01ser_6_), .B0_f (new_AGEMA_signal_3211), .B1_t (new_AGEMA_signal_3212), .B1_f (new_AGEMA_signal_3213), .Z0_t (KeyArray_inS00ser[6]), .Z0_f (new_AGEMA_signal_5732), .Z1_t (new_AGEMA_signal_5733), .Z1_f (new_AGEMA_signal_5734) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_7_XOR1_U1 ( .A0_t (KeyArray_outS01ser_7_), .A0_f (new_AGEMA_signal_3205), .A1_t (new_AGEMA_signal_3206), .A1_f (new_AGEMA_signal_3207), .B0_t (KeyArray_outS01ser_XOR_00[7]), .B0_f (new_AGEMA_signal_3208), .B1_t (new_AGEMA_signal_3209), .B1_f (new_AGEMA_signal_3210), .Z0_t (KeyArray_MUX_inS00ser_mux_inst_7_X), .Z0_f (new_AGEMA_signal_4544), .Z1_t (new_AGEMA_signal_4545), .Z1_f (new_AGEMA_signal_4546) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_7_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (KeyArray_nReset_selXOR), .A1_f (new_AGEMA_signal_5406), .B0_t (KeyArray_MUX_inS00ser_mux_inst_7_X), .B0_f (new_AGEMA_signal_4544), .B1_t (new_AGEMA_signal_4545), .B1_f (new_AGEMA_signal_4546), .Z0_t (KeyArray_MUX_inS00ser_mux_inst_7_Y), .Z0_f (new_AGEMA_signal_5605), .Z1_t (new_AGEMA_signal_5606), .Z1_f (new_AGEMA_signal_5607) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS00ser_mux_inst_7_XOR2_U1 ( .A0_t (KeyArray_MUX_inS00ser_mux_inst_7_Y), .A0_f (new_AGEMA_signal_5605), .A1_t (new_AGEMA_signal_5606), .A1_f (new_AGEMA_signal_5607), .B0_t (KeyArray_outS01ser_7_), .B0_f (new_AGEMA_signal_3205), .B1_t (new_AGEMA_signal_3206), .B1_f (new_AGEMA_signal_3207), .Z0_t (KeyArray_inS00ser[7]), .Z0_f (new_AGEMA_signal_5735), .Z1_t (new_AGEMA_signal_5736), .Z1_f (new_AGEMA_signal_5737) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_0_XOR1_U1 ( .A0_t (port_out_s0_t[0]), .A0_f (port_out_s0_f[0]), .A1_t (port_out_s1_t[0]), .A1_f (port_out_s1_f[0]), .B0_t (keyStateIn[0]), .B0_f (new_AGEMA_signal_2489), .B1_t (new_AGEMA_signal_2490), .B1_f (new_AGEMA_signal_2491), .Z0_t (KeyArray_MUX_inS33ser_mux_inst_0_X), .Z0_f (new_AGEMA_signal_3901), .Z1_t (new_AGEMA_signal_3902), .Z1_f (new_AGEMA_signal_3903) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_0_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyArray_MUX_inS33ser_mux_inst_0_X), .B0_f (new_AGEMA_signal_3901), .B1_t (new_AGEMA_signal_3902), .B1_f (new_AGEMA_signal_3903), .Z0_t (KeyArray_MUX_inS33ser_mux_inst_0_Y), .Z0_f (new_AGEMA_signal_4547), .Z1_t (new_AGEMA_signal_4548), .Z1_f (new_AGEMA_signal_4549) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_0_XOR2_U1 ( .A0_t (KeyArray_MUX_inS33ser_mux_inst_0_Y), .A0_f (new_AGEMA_signal_4547), .A1_t (new_AGEMA_signal_4548), .A1_f (new_AGEMA_signal_4549), .B0_t (port_out_s0_t[0]), .B0_f (port_out_s0_f[0]), .B1_t (port_out_s1_t[0]), .B1_f (port_out_s1_f[0]), .Z0_t (KeyArray_inS33ser[0]), .Z0_f (new_AGEMA_signal_5013), .Z1_t (new_AGEMA_signal_5014), .Z1_f (new_AGEMA_signal_5015) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_1_XOR1_U1 ( .A0_t (port_out_s0_t[1]), .A0_f (port_out_s0_f[1]), .A1_t (port_out_s1_t[1]), .A1_f (port_out_s1_f[1]), .B0_t (keyStateIn[1]), .B0_f (new_AGEMA_signal_2498), .B1_t (new_AGEMA_signal_2499), .B1_f (new_AGEMA_signal_2500), .Z0_t (KeyArray_MUX_inS33ser_mux_inst_1_X), .Z0_f (new_AGEMA_signal_3904), .Z1_t (new_AGEMA_signal_3905), .Z1_f (new_AGEMA_signal_3906) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyArray_MUX_inS33ser_mux_inst_1_X), .B0_f (new_AGEMA_signal_3904), .B1_t (new_AGEMA_signal_3905), .B1_f (new_AGEMA_signal_3906), .Z0_t (KeyArray_MUX_inS33ser_mux_inst_1_Y), .Z0_f (new_AGEMA_signal_4550), .Z1_t (new_AGEMA_signal_4551), .Z1_f (new_AGEMA_signal_4552) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_1_XOR2_U1 ( .A0_t (KeyArray_MUX_inS33ser_mux_inst_1_Y), .A0_f (new_AGEMA_signal_4550), .A1_t (new_AGEMA_signal_4551), .A1_f (new_AGEMA_signal_4552), .B0_t (port_out_s0_t[1]), .B0_f (port_out_s0_f[1]), .B1_t (port_out_s1_t[1]), .B1_f (port_out_s1_f[1]), .Z0_t (KeyArray_inS33ser[1]), .Z0_f (new_AGEMA_signal_5016), .Z1_t (new_AGEMA_signal_5017), .Z1_f (new_AGEMA_signal_5018) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_2_XOR1_U1 ( .A0_t (port_out_s0_t[2]), .A0_f (port_out_s0_f[2]), .A1_t (port_out_s1_t[2]), .A1_f (port_out_s1_f[2]), .B0_t (keyStateIn[2]), .B0_f (new_AGEMA_signal_2507), .B1_t (new_AGEMA_signal_2508), .B1_f (new_AGEMA_signal_2509), .Z0_t (KeyArray_MUX_inS33ser_mux_inst_2_X), .Z0_f (new_AGEMA_signal_3907), .Z1_t (new_AGEMA_signal_3908), .Z1_f (new_AGEMA_signal_3909) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_2_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyArray_MUX_inS33ser_mux_inst_2_X), .B0_f (new_AGEMA_signal_3907), .B1_t (new_AGEMA_signal_3908), .B1_f (new_AGEMA_signal_3909), .Z0_t (KeyArray_MUX_inS33ser_mux_inst_2_Y), .Z0_f (new_AGEMA_signal_4553), .Z1_t (new_AGEMA_signal_4554), .Z1_f (new_AGEMA_signal_4555) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_2_XOR2_U1 ( .A0_t (KeyArray_MUX_inS33ser_mux_inst_2_Y), .A0_f (new_AGEMA_signal_4553), .A1_t (new_AGEMA_signal_4554), .A1_f (new_AGEMA_signal_4555), .B0_t (port_out_s0_t[2]), .B0_f (port_out_s0_f[2]), .B1_t (port_out_s1_t[2]), .B1_f (port_out_s1_f[2]), .Z0_t (KeyArray_inS33ser[2]), .Z0_f (new_AGEMA_signal_5019), .Z1_t (new_AGEMA_signal_5020), .Z1_f (new_AGEMA_signal_5021) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_3_XOR1_U1 ( .A0_t (port_out_s0_t[3]), .A0_f (port_out_s0_f[3]), .A1_t (port_out_s1_t[3]), .A1_f (port_out_s1_f[3]), .B0_t (keyStateIn[3]), .B0_f (new_AGEMA_signal_2516), .B1_t (new_AGEMA_signal_2517), .B1_f (new_AGEMA_signal_2518), .Z0_t (KeyArray_MUX_inS33ser_mux_inst_3_X), .Z0_f (new_AGEMA_signal_3910), .Z1_t (new_AGEMA_signal_3911), .Z1_f (new_AGEMA_signal_3912) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_3_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyArray_MUX_inS33ser_mux_inst_3_X), .B0_f (new_AGEMA_signal_3910), .B1_t (new_AGEMA_signal_3911), .B1_f (new_AGEMA_signal_3912), .Z0_t (KeyArray_MUX_inS33ser_mux_inst_3_Y), .Z0_f (new_AGEMA_signal_4556), .Z1_t (new_AGEMA_signal_4557), .Z1_f (new_AGEMA_signal_4558) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_3_XOR2_U1 ( .A0_t (KeyArray_MUX_inS33ser_mux_inst_3_Y), .A0_f (new_AGEMA_signal_4556), .A1_t (new_AGEMA_signal_4557), .A1_f (new_AGEMA_signal_4558), .B0_t (port_out_s0_t[3]), .B0_f (port_out_s0_f[3]), .B1_t (port_out_s1_t[3]), .B1_f (port_out_s1_f[3]), .Z0_t (KeyArray_inS33ser[3]), .Z0_f (new_AGEMA_signal_5022), .Z1_t (new_AGEMA_signal_5023), .Z1_f (new_AGEMA_signal_5024) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_4_XOR1_U1 ( .A0_t (port_out_s0_t[4]), .A0_f (port_out_s0_f[4]), .A1_t (port_out_s1_t[4]), .A1_f (port_out_s1_f[4]), .B0_t (keyStateIn[4]), .B0_f (new_AGEMA_signal_2525), .B1_t (new_AGEMA_signal_2526), .B1_f (new_AGEMA_signal_2527), .Z0_t (KeyArray_MUX_inS33ser_mux_inst_4_X), .Z0_f (new_AGEMA_signal_3913), .Z1_t (new_AGEMA_signal_3914), .Z1_f (new_AGEMA_signal_3915) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_4_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyArray_MUX_inS33ser_mux_inst_4_X), .B0_f (new_AGEMA_signal_3913), .B1_t (new_AGEMA_signal_3914), .B1_f (new_AGEMA_signal_3915), .Z0_t (KeyArray_MUX_inS33ser_mux_inst_4_Y), .Z0_f (new_AGEMA_signal_4559), .Z1_t (new_AGEMA_signal_4560), .Z1_f (new_AGEMA_signal_4561) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_4_XOR2_U1 ( .A0_t (KeyArray_MUX_inS33ser_mux_inst_4_Y), .A0_f (new_AGEMA_signal_4559), .A1_t (new_AGEMA_signal_4560), .A1_f (new_AGEMA_signal_4561), .B0_t (port_out_s0_t[4]), .B0_f (port_out_s0_f[4]), .B1_t (port_out_s1_t[4]), .B1_f (port_out_s1_f[4]), .Z0_t (KeyArray_inS33ser[4]), .Z0_f (new_AGEMA_signal_5025), .Z1_t (new_AGEMA_signal_5026), .Z1_f (new_AGEMA_signal_5027) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_5_XOR1_U1 ( .A0_t (port_out_s0_t[5]), .A0_f (port_out_s0_f[5]), .A1_t (port_out_s1_t[5]), .A1_f (port_out_s1_f[5]), .B0_t (keyStateIn[5]), .B0_f (new_AGEMA_signal_2534), .B1_t (new_AGEMA_signal_2535), .B1_f (new_AGEMA_signal_2536), .Z0_t (KeyArray_MUX_inS33ser_mux_inst_5_X), .Z0_f (new_AGEMA_signal_3916), .Z1_t (new_AGEMA_signal_3917), .Z1_f (new_AGEMA_signal_3918) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_5_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyArray_MUX_inS33ser_mux_inst_5_X), .B0_f (new_AGEMA_signal_3916), .B1_t (new_AGEMA_signal_3917), .B1_f (new_AGEMA_signal_3918), .Z0_t (KeyArray_MUX_inS33ser_mux_inst_5_Y), .Z0_f (new_AGEMA_signal_4562), .Z1_t (new_AGEMA_signal_4563), .Z1_f (new_AGEMA_signal_4564) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_5_XOR2_U1 ( .A0_t (KeyArray_MUX_inS33ser_mux_inst_5_Y), .A0_f (new_AGEMA_signal_4562), .A1_t (new_AGEMA_signal_4563), .A1_f (new_AGEMA_signal_4564), .B0_t (port_out_s0_t[5]), .B0_f (port_out_s0_f[5]), .B1_t (port_out_s1_t[5]), .B1_f (port_out_s1_f[5]), .Z0_t (KeyArray_inS33ser[5]), .Z0_f (new_AGEMA_signal_5028), .Z1_t (new_AGEMA_signal_5029), .Z1_f (new_AGEMA_signal_5030) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_6_XOR1_U1 ( .A0_t (port_out_s0_t[6]), .A0_f (port_out_s0_f[6]), .A1_t (port_out_s1_t[6]), .A1_f (port_out_s1_f[6]), .B0_t (keyStateIn[6]), .B0_f (new_AGEMA_signal_2543), .B1_t (new_AGEMA_signal_2544), .B1_f (new_AGEMA_signal_2545), .Z0_t (KeyArray_MUX_inS33ser_mux_inst_6_X), .Z0_f (new_AGEMA_signal_3919), .Z1_t (new_AGEMA_signal_3920), .Z1_f (new_AGEMA_signal_3921) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_6_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyArray_MUX_inS33ser_mux_inst_6_X), .B0_f (new_AGEMA_signal_3919), .B1_t (new_AGEMA_signal_3920), .B1_f (new_AGEMA_signal_3921), .Z0_t (KeyArray_MUX_inS33ser_mux_inst_6_Y), .Z0_f (new_AGEMA_signal_4565), .Z1_t (new_AGEMA_signal_4566), .Z1_f (new_AGEMA_signal_4567) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_6_XOR2_U1 ( .A0_t (KeyArray_MUX_inS33ser_mux_inst_6_Y), .A0_f (new_AGEMA_signal_4565), .A1_t (new_AGEMA_signal_4566), .A1_f (new_AGEMA_signal_4567), .B0_t (port_out_s0_t[6]), .B0_f (port_out_s0_f[6]), .B1_t (port_out_s1_t[6]), .B1_f (port_out_s1_f[6]), .Z0_t (KeyArray_inS33ser[6]), .Z0_f (new_AGEMA_signal_5031), .Z1_t (new_AGEMA_signal_5032), .Z1_f (new_AGEMA_signal_5033) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_7_XOR1_U1 ( .A0_t (port_out_s0_t[7]), .A0_f (port_out_s0_f[7]), .A1_t (port_out_s1_t[7]), .A1_f (port_out_s1_f[7]), .B0_t (keyStateIn[7]), .B0_f (new_AGEMA_signal_2552), .B1_t (new_AGEMA_signal_2553), .B1_f (new_AGEMA_signal_2554), .Z0_t (KeyArray_MUX_inS33ser_mux_inst_7_X), .Z0_f (new_AGEMA_signal_3922), .Z1_t (new_AGEMA_signal_3923), .Z1_f (new_AGEMA_signal_3924) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_7_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (start_t), .A1_f (start_f), .B0_t (KeyArray_MUX_inS33ser_mux_inst_7_X), .B0_f (new_AGEMA_signal_3922), .B1_t (new_AGEMA_signal_3923), .B1_f (new_AGEMA_signal_3924), .Z0_t (KeyArray_MUX_inS33ser_mux_inst_7_Y), .Z0_f (new_AGEMA_signal_4568), .Z1_t (new_AGEMA_signal_4569), .Z1_f (new_AGEMA_signal_4570) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) KeyArray_MUX_inS33ser_mux_inst_7_XOR2_U1 ( .A0_t (KeyArray_MUX_inS33ser_mux_inst_7_Y), .A0_f (new_AGEMA_signal_4568), .A1_t (new_AGEMA_signal_4569), .A1_f (new_AGEMA_signal_4570), .B0_t (port_out_s0_t[7]), .B0_f (port_out_s0_f[7]), .B1_t (port_out_s1_t[7]), .B1_f (port_out_s1_f[7]), .Z0_t (KeyArray_inS33ser[7]), .Z0_f (new_AGEMA_signal_5034), .Z1_t (new_AGEMA_signal_5035), .Z1_f (new_AGEMA_signal_5036) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line0_U24 ( .A0_t (MixColumns_line0_n16), .A0_f (new_AGEMA_signal_4571), .A1_t (new_AGEMA_signal_4572), .A1_f (new_AGEMA_signal_4573), .B0_t (MixColumns_line0_n15), .B0_f (new_AGEMA_signal_3925), .B1_t (new_AGEMA_signal_3926), .B1_f (new_AGEMA_signal_3927), .Z0_t (MCout[31]), .Z0_f (new_AGEMA_signal_5037), .Z1_t (new_AGEMA_signal_5038), .Z1_f (new_AGEMA_signal_5039) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line0_U23 ( .A0_t (MixColumns_line2_S02[0]), .A0_f (new_AGEMA_signal_3031), .A1_t (new_AGEMA_signal_3032), .A1_f (new_AGEMA_signal_3033), .B0_t (MixColumns_line3_S02[0]), .B0_f (new_AGEMA_signal_3175), .B1_t (new_AGEMA_signal_3176), .B1_f (new_AGEMA_signal_3177), .Z0_t (MixColumns_line0_n15), .Z0_f (new_AGEMA_signal_3925), .Z1_t (new_AGEMA_signal_3926), .Z1_f (new_AGEMA_signal_3927) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_U22 ( .A0_t (port_out_s0_t[6]), .A0_f (port_out_s0_f[6]), .A1_t (port_out_s1_t[6]), .A1_f (port_out_s1_f[6]), .B0_t (MixColumns_line0_S13[7]), .B0_f (new_AGEMA_signal_3964), .B1_t (new_AGEMA_signal_3965), .B1_f (new_AGEMA_signal_3966), .Z0_t (MixColumns_line0_n16), .Z0_f (new_AGEMA_signal_4571), .Z1_t (new_AGEMA_signal_4572), .Z1_f (new_AGEMA_signal_4573) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line0_U21 ( .A0_t (MixColumns_line0_n14), .A0_f (new_AGEMA_signal_4574), .A1_t (new_AGEMA_signal_4575), .A1_f (new_AGEMA_signal_4576), .B0_t (MixColumns_line0_n13), .B0_f (new_AGEMA_signal_3928), .B1_t (new_AGEMA_signal_3929), .B1_f (new_AGEMA_signal_3930), .Z0_t (MCout[30]), .Z0_f (new_AGEMA_signal_5040), .Z1_t (new_AGEMA_signal_5041), .Z1_f (new_AGEMA_signal_5042) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line0_U20 ( .A0_t (MixColumns_line2_S02[7]), .A0_f (new_AGEMA_signal_3025), .A1_t (new_AGEMA_signal_3026), .A1_f (new_AGEMA_signal_3027), .B0_t (MixColumns_line3_S02[7]), .B0_f (new_AGEMA_signal_3166), .B1_t (new_AGEMA_signal_3167), .B1_f (new_AGEMA_signal_3168), .Z0_t (MixColumns_line0_n13), .Z0_f (new_AGEMA_signal_3928), .Z1_t (new_AGEMA_signal_3929), .Z1_f (new_AGEMA_signal_3930) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_U19 ( .A0_t (port_out_s0_t[5]), .A0_f (port_out_s0_f[5]), .A1_t (port_out_s1_t[5]), .A1_f (port_out_s1_f[5]), .B0_t (MixColumns_line0_S13[6]), .B0_f (new_AGEMA_signal_3970), .B1_t (new_AGEMA_signal_3971), .B1_f (new_AGEMA_signal_3972), .Z0_t (MixColumns_line0_n14), .Z0_f (new_AGEMA_signal_4574), .Z1_t (new_AGEMA_signal_4575), .Z1_f (new_AGEMA_signal_4576) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line0_U18 ( .A0_t (MixColumns_line0_n12), .A0_f (new_AGEMA_signal_4577), .A1_t (new_AGEMA_signal_4578), .A1_f (new_AGEMA_signal_4579), .B0_t (MixColumns_line0_n11), .B0_f (new_AGEMA_signal_3931), .B1_t (new_AGEMA_signal_3932), .B1_f (new_AGEMA_signal_3933), .Z0_t (MCout[29]), .Z0_f (new_AGEMA_signal_5043), .Z1_t (new_AGEMA_signal_5044), .Z1_f (new_AGEMA_signal_5045) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line0_U17 ( .A0_t (MixColumns_line2_S02[6]), .A0_f (new_AGEMA_signal_3019), .A1_t (new_AGEMA_signal_3020), .A1_f (new_AGEMA_signal_3021), .B0_t (MixColumns_line3_S02[6]), .B0_f (new_AGEMA_signal_3157), .B1_t (new_AGEMA_signal_3158), .B1_f (new_AGEMA_signal_3159), .Z0_t (MixColumns_line0_n11), .Z0_f (new_AGEMA_signal_3931), .Z1_t (new_AGEMA_signal_3932), .Z1_f (new_AGEMA_signal_3933) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_U16 ( .A0_t (port_out_s0_t[4]), .A0_f (port_out_s0_f[4]), .A1_t (port_out_s1_t[4]), .A1_f (port_out_s1_f[4]), .B0_t (MixColumns_line0_S13[5]), .B0_f (new_AGEMA_signal_3976), .B1_t (new_AGEMA_signal_3977), .B1_f (new_AGEMA_signal_3978), .Z0_t (MixColumns_line0_n12), .Z0_f (new_AGEMA_signal_4577), .Z1_t (new_AGEMA_signal_4578), .Z1_f (new_AGEMA_signal_4579) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line0_U15 ( .A0_t (MixColumns_line0_n10), .A0_f (new_AGEMA_signal_5046), .A1_t (new_AGEMA_signal_5047), .A1_f (new_AGEMA_signal_5048), .B0_t (MixColumns_line0_n9), .B0_f (new_AGEMA_signal_3934), .B1_t (new_AGEMA_signal_3935), .B1_f (new_AGEMA_signal_3936), .Z0_t (MCout[28]), .Z0_f (new_AGEMA_signal_5247), .Z1_t (new_AGEMA_signal_5248), .Z1_f (new_AGEMA_signal_5249) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line0_U14 ( .A0_t (MixColumns_line2_S02[5]), .A0_f (new_AGEMA_signal_3013), .A1_t (new_AGEMA_signal_3014), .A1_f (new_AGEMA_signal_3015), .B0_t (MixColumns_line3_S02[5]), .B0_f (new_AGEMA_signal_3148), .B1_t (new_AGEMA_signal_3149), .B1_f (new_AGEMA_signal_3150), .Z0_t (MixColumns_line0_n9), .Z0_f (new_AGEMA_signal_3934), .Z1_t (new_AGEMA_signal_3935), .Z1_f (new_AGEMA_signal_3936) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_U13 ( .A0_t (MixColumns_line0_S02[4]), .A0_f (new_AGEMA_signal_3949), .A1_t (new_AGEMA_signal_3950), .A1_f (new_AGEMA_signal_3951), .B0_t (MixColumns_line0_S13[4]), .B0_f (new_AGEMA_signal_4586), .B1_t (new_AGEMA_signal_4587), .B1_f (new_AGEMA_signal_4588), .Z0_t (MixColumns_line0_n10), .Z0_f (new_AGEMA_signal_5046), .Z1_t (new_AGEMA_signal_5047), .Z1_f (new_AGEMA_signal_5048) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line0_U12 ( .A0_t (MixColumns_line0_n8), .A0_f (new_AGEMA_signal_5049), .A1_t (new_AGEMA_signal_5050), .A1_f (new_AGEMA_signal_5051), .B0_t (MixColumns_line0_n7), .B0_f (new_AGEMA_signal_3937), .B1_t (new_AGEMA_signal_3938), .B1_f (new_AGEMA_signal_3939), .Z0_t (MCout[27]), .Z0_f (new_AGEMA_signal_5250), .Z1_t (new_AGEMA_signal_5251), .Z1_f (new_AGEMA_signal_5252) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line0_U11 ( .A0_t (MCin[11]), .A0_f (new_AGEMA_signal_3007), .A1_t (new_AGEMA_signal_3008), .A1_f (new_AGEMA_signal_3009), .B0_t (MCin[3]), .B0_f (new_AGEMA_signal_3139), .B1_t (new_AGEMA_signal_3140), .B1_f (new_AGEMA_signal_3141), .Z0_t (MixColumns_line0_n7), .Z0_f (new_AGEMA_signal_3937), .Z1_t (new_AGEMA_signal_3938), .Z1_f (new_AGEMA_signal_3939) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_U10 ( .A0_t (MixColumns_line0_S02[3]), .A0_f (new_AGEMA_signal_3952), .A1_t (new_AGEMA_signal_3953), .A1_f (new_AGEMA_signal_3954), .B0_t (MixColumns_line0_S13[3]), .B0_f (new_AGEMA_signal_4589), .B1_t (new_AGEMA_signal_4590), .B1_f (new_AGEMA_signal_4591), .Z0_t (MixColumns_line0_n8), .Z0_f (new_AGEMA_signal_5049), .Z1_t (new_AGEMA_signal_5050), .Z1_f (new_AGEMA_signal_5051) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line0_U9 ( .A0_t (MixColumns_line0_n6), .A0_f (new_AGEMA_signal_4580), .A1_t (new_AGEMA_signal_4581), .A1_f (new_AGEMA_signal_4582), .B0_t (MixColumns_line0_n5), .B0_f (new_AGEMA_signal_3940), .B1_t (new_AGEMA_signal_3941), .B1_f (new_AGEMA_signal_3942), .Z0_t (MCout[26]), .Z0_f (new_AGEMA_signal_5052), .Z1_t (new_AGEMA_signal_5053), .Z1_f (new_AGEMA_signal_5054) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line0_U8 ( .A0_t (MCin[10]), .A0_f (new_AGEMA_signal_3001), .A1_t (new_AGEMA_signal_3002), .A1_f (new_AGEMA_signal_3003), .B0_t (MCin[2]), .B0_f (new_AGEMA_signal_3130), .B1_t (new_AGEMA_signal_3131), .B1_f (new_AGEMA_signal_3132), .Z0_t (MixColumns_line0_n5), .Z0_f (new_AGEMA_signal_3940), .Z1_t (new_AGEMA_signal_3941), .Z1_f (new_AGEMA_signal_3942) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_U7 ( .A0_t (port_out_s0_t[1]), .A0_f (port_out_s0_f[1]), .A1_t (port_out_s1_t[1]), .A1_f (port_out_s1_f[1]), .B0_t (MixColumns_line0_S13[2]), .B0_f (new_AGEMA_signal_3985), .B1_t (new_AGEMA_signal_3986), .B1_f (new_AGEMA_signal_3987), .Z0_t (MixColumns_line0_n6), .Z0_f (new_AGEMA_signal_4580), .Z1_t (new_AGEMA_signal_4581), .Z1_f (new_AGEMA_signal_4582) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line0_U6 ( .A0_t (MixColumns_line0_n4), .A0_f (new_AGEMA_signal_5055), .A1_t (new_AGEMA_signal_5056), .A1_f (new_AGEMA_signal_5057), .B0_t (MixColumns_line0_n3), .B0_f (new_AGEMA_signal_3943), .B1_t (new_AGEMA_signal_3944), .B1_f (new_AGEMA_signal_3945), .Z0_t (MCout[25]), .Z0_f (new_AGEMA_signal_5253), .Z1_t (new_AGEMA_signal_5254), .Z1_f (new_AGEMA_signal_5255) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line0_U5 ( .A0_t (MixColumns_line3_S02[2]), .A0_f (new_AGEMA_signal_3121), .A1_t (new_AGEMA_signal_3122), .A1_f (new_AGEMA_signal_3123), .B0_t (MixColumns_line2_S02[2]), .B0_f (new_AGEMA_signal_2995), .B1_t (new_AGEMA_signal_2996), .B1_f (new_AGEMA_signal_2997), .Z0_t (MixColumns_line0_n3), .Z0_f (new_AGEMA_signal_3943), .Z1_t (new_AGEMA_signal_3944), .Z1_f (new_AGEMA_signal_3945) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_U4 ( .A0_t (MixColumns_line0_S02[1]), .A0_f (new_AGEMA_signal_3955), .A1_t (new_AGEMA_signal_3956), .A1_f (new_AGEMA_signal_3957), .B0_t (MixColumns_line0_S13[1]), .B0_f (new_AGEMA_signal_4592), .B1_t (new_AGEMA_signal_4593), .B1_f (new_AGEMA_signal_4594), .Z0_t (MixColumns_line0_n4), .Z0_f (new_AGEMA_signal_5055), .Z1_t (new_AGEMA_signal_5056), .Z1_f (new_AGEMA_signal_5057) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line0_U3 ( .A0_t (MixColumns_line0_n2), .A0_f (new_AGEMA_signal_4583), .A1_t (new_AGEMA_signal_4584), .A1_f (new_AGEMA_signal_4585), .B0_t (MixColumns_line0_n1), .B0_f (new_AGEMA_signal_3946), .B1_t (new_AGEMA_signal_3947), .B1_f (new_AGEMA_signal_3948), .Z0_t (MCout[24]), .Z0_f (new_AGEMA_signal_5058), .Z1_t (new_AGEMA_signal_5059), .Z1_f (new_AGEMA_signal_5060) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line0_U2 ( .A0_t (MCin[0]), .A0_f (new_AGEMA_signal_3112), .A1_t (new_AGEMA_signal_3113), .A1_f (new_AGEMA_signal_3114), .B0_t (MCin[8]), .B0_f (new_AGEMA_signal_2989), .B1_t (new_AGEMA_signal_2990), .B1_f (new_AGEMA_signal_2991), .Z0_t (MixColumns_line0_n1), .Z0_f (new_AGEMA_signal_3946), .Z1_t (new_AGEMA_signal_3947), .Z1_f (new_AGEMA_signal_3948) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_U1 ( .A0_t (port_out_s0_t[7]), .A0_f (port_out_s0_f[7]), .A1_t (port_out_s1_t[7]), .A1_f (port_out_s1_f[7]), .B0_t (MixColumns_line0_S13[0]), .B0_f (new_AGEMA_signal_3991), .B1_t (new_AGEMA_signal_3992), .B1_f (new_AGEMA_signal_3993), .Z0_t (MixColumns_line0_n2), .Z0_f (new_AGEMA_signal_4583), .Z1_t (new_AGEMA_signal_4584), .Z1_f (new_AGEMA_signal_4585) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_timesTWO_U3 ( .A0_t (port_out_s0_t[7]), .A0_f (port_out_s0_f[7]), .A1_t (port_out_s1_t[7]), .A1_f (port_out_s1_f[7]), .B0_t (port_out_s0_t[3]), .B0_f (port_out_s0_f[3]), .B1_t (port_out_s1_t[3]), .B1_f (port_out_s1_f[3]), .Z0_t (MixColumns_line0_S02[4]), .Z0_f (new_AGEMA_signal_3949), .Z1_t (new_AGEMA_signal_3950), .Z1_f (new_AGEMA_signal_3951) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_timesTWO_U2 ( .A0_t (port_out_s0_t[7]), .A0_f (port_out_s0_f[7]), .A1_t (port_out_s1_t[7]), .A1_f (port_out_s1_f[7]), .B0_t (port_out_s0_t[2]), .B0_f (port_out_s0_f[2]), .B1_t (port_out_s1_t[2]), .B1_f (port_out_s1_f[2]), .Z0_t (MixColumns_line0_S02[3]), .Z0_f (new_AGEMA_signal_3952), .Z1_t (new_AGEMA_signal_3953), .Z1_f (new_AGEMA_signal_3954) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_timesTWO_U1 ( .A0_t (port_out_s0_t[7]), .A0_f (port_out_s0_f[7]), .A1_t (port_out_s1_t[7]), .A1_f (port_out_s1_f[7]), .B0_t (port_out_s0_t[0]), .B0_f (port_out_s0_f[0]), .B1_t (port_out_s1_t[0]), .B1_f (port_out_s1_f[0]), .Z0_t (MixColumns_line0_S02[1]), .Z0_f (new_AGEMA_signal_3955), .Z1_t (new_AGEMA_signal_3956), .Z1_f (new_AGEMA_signal_3957) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_timesTHREE_U8 ( .A0_t (MixColumns_line1_S02[0]), .A0_f (new_AGEMA_signal_3958), .A1_t (new_AGEMA_signal_3959), .A1_f (new_AGEMA_signal_3960), .B0_t (MixColumns_line1_S02[7]), .B0_f (new_AGEMA_signal_3961), .B1_t (new_AGEMA_signal_3962), .B1_f (new_AGEMA_signal_3963), .Z0_t (MixColumns_line0_S13[7]), .Z0_f (new_AGEMA_signal_3964), .Z1_t (new_AGEMA_signal_3965), .Z1_f (new_AGEMA_signal_3966) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_timesTHREE_U7 ( .A0_t (MixColumns_line1_S02[7]), .A0_f (new_AGEMA_signal_3961), .A1_t (new_AGEMA_signal_3962), .A1_f (new_AGEMA_signal_3963), .B0_t (MixColumns_line1_S02[6]), .B0_f (new_AGEMA_signal_3967), .B1_t (new_AGEMA_signal_3968), .B1_f (new_AGEMA_signal_3969), .Z0_t (MixColumns_line0_S13[6]), .Z0_f (new_AGEMA_signal_3970), .Z1_t (new_AGEMA_signal_3971), .Z1_f (new_AGEMA_signal_3972) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_timesTHREE_U6 ( .A0_t (MixColumns_line1_S02[6]), .A0_f (new_AGEMA_signal_3967), .A1_t (new_AGEMA_signal_3968), .A1_f (new_AGEMA_signal_3969), .B0_t (MixColumns_line1_S02[5]), .B0_f (new_AGEMA_signal_3973), .B1_t (new_AGEMA_signal_3974), .B1_f (new_AGEMA_signal_3975), .Z0_t (MixColumns_line0_S13[5]), .Z0_f (new_AGEMA_signal_3976), .Z1_t (new_AGEMA_signal_3977), .Z1_f (new_AGEMA_signal_3978) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_timesTHREE_U5 ( .A0_t (MixColumns_line1_S02[5]), .A0_f (new_AGEMA_signal_3973), .A1_t (new_AGEMA_signal_3974), .A1_f (new_AGEMA_signal_3975), .B0_t (MixColumns_line0_timesTHREE_input2[4]), .B0_f (new_AGEMA_signal_3997), .B1_t (new_AGEMA_signal_3998), .B1_f (new_AGEMA_signal_3999), .Z0_t (MixColumns_line0_S13[4]), .Z0_f (new_AGEMA_signal_4586), .Z1_t (new_AGEMA_signal_4587), .Z1_f (new_AGEMA_signal_4588) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_timesTHREE_U4 ( .A0_t (MCin[19]), .A0_f (new_AGEMA_signal_3994), .A1_t (new_AGEMA_signal_3995), .A1_f (new_AGEMA_signal_3996), .B0_t (MixColumns_line0_timesTHREE_input2[3]), .B0_f (new_AGEMA_signal_4000), .B1_t (new_AGEMA_signal_4001), .B1_f (new_AGEMA_signal_4002), .Z0_t (MixColumns_line0_S13[3]), .Z0_f (new_AGEMA_signal_4589), .Z1_t (new_AGEMA_signal_4590), .Z1_f (new_AGEMA_signal_4591) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_timesTHREE_U3 ( .A0_t (MCin[18]), .A0_f (new_AGEMA_signal_3979), .A1_t (new_AGEMA_signal_3980), .A1_f (new_AGEMA_signal_3981), .B0_t (MixColumns_line1_S02[2]), .B0_f (new_AGEMA_signal_3982), .B1_t (new_AGEMA_signal_3983), .B1_f (new_AGEMA_signal_3984), .Z0_t (MixColumns_line0_S13[2]), .Z0_f (new_AGEMA_signal_3985), .Z1_t (new_AGEMA_signal_3986), .Z1_f (new_AGEMA_signal_3987) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_timesTHREE_U2 ( .A0_t (MixColumns_line1_S02[2]), .A0_f (new_AGEMA_signal_3982), .A1_t (new_AGEMA_signal_3983), .A1_f (new_AGEMA_signal_3984), .B0_t (MixColumns_line0_timesTHREE_input2[1]), .B0_f (new_AGEMA_signal_4003), .B1_t (new_AGEMA_signal_4004), .B1_f (new_AGEMA_signal_4005), .Z0_t (MixColumns_line0_S13[1]), .Z0_f (new_AGEMA_signal_4592), .Z1_t (new_AGEMA_signal_4593), .Z1_f (new_AGEMA_signal_4594) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_timesTHREE_U1 ( .A0_t (MCin[16]), .A0_f (new_AGEMA_signal_3988), .A1_t (new_AGEMA_signal_3989), .A1_f (new_AGEMA_signal_3990), .B0_t (MixColumns_line1_S02[0]), .B0_f (new_AGEMA_signal_3958), .B1_t (new_AGEMA_signal_3959), .B1_f (new_AGEMA_signal_3960), .Z0_t (MixColumns_line0_S13[0]), .Z0_f (new_AGEMA_signal_3991), .Z1_t (new_AGEMA_signal_3992), .Z1_f (new_AGEMA_signal_3993) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_timesTHREE_timesTWO_U3 ( .A0_t (MixColumns_line1_S02[0]), .A0_f (new_AGEMA_signal_3958), .A1_t (new_AGEMA_signal_3959), .A1_f (new_AGEMA_signal_3960), .B0_t (MCin[19]), .B0_f (new_AGEMA_signal_3994), .B1_t (new_AGEMA_signal_3995), .B1_f (new_AGEMA_signal_3996), .Z0_t (MixColumns_line0_timesTHREE_input2[4]), .Z0_f (new_AGEMA_signal_3997), .Z1_t (new_AGEMA_signal_3998), .Z1_f (new_AGEMA_signal_3999) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_timesTHREE_timesTWO_U2 ( .A0_t (MixColumns_line1_S02[0]), .A0_f (new_AGEMA_signal_3958), .A1_t (new_AGEMA_signal_3959), .A1_f (new_AGEMA_signal_3960), .B0_t (MCin[18]), .B0_f (new_AGEMA_signal_3979), .B1_t (new_AGEMA_signal_3980), .B1_f (new_AGEMA_signal_3981), .Z0_t (MixColumns_line0_timesTHREE_input2[3]), .Z0_f (new_AGEMA_signal_4000), .Z1_t (new_AGEMA_signal_4001), .Z1_f (new_AGEMA_signal_4002) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line0_timesTHREE_timesTWO_U1 ( .A0_t (MixColumns_line1_S02[0]), .A0_f (new_AGEMA_signal_3958), .A1_t (new_AGEMA_signal_3959), .A1_f (new_AGEMA_signal_3960), .B0_t (MCin[16]), .B0_f (new_AGEMA_signal_3988), .B1_t (new_AGEMA_signal_3989), .B1_f (new_AGEMA_signal_3990), .Z0_t (MixColumns_line0_timesTHREE_input2[1]), .Z0_f (new_AGEMA_signal_4003), .Z1_t (new_AGEMA_signal_4004), .Z1_f (new_AGEMA_signal_4005) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line1_U24 ( .A0_t (MixColumns_line1_n16), .A0_f (new_AGEMA_signal_4595), .A1_t (new_AGEMA_signal_4596), .A1_f (new_AGEMA_signal_4597), .B0_t (MixColumns_line1_n15), .B0_f (new_AGEMA_signal_4006), .B1_t (new_AGEMA_signal_4007), .B1_f (new_AGEMA_signal_4008), .Z0_t (MCout[23]), .Z0_f (new_AGEMA_signal_5061), .Z1_t (new_AGEMA_signal_5062), .Z1_f (new_AGEMA_signal_5063) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line1_U23 ( .A0_t (MixColumns_line3_S02[0]), .A0_f (new_AGEMA_signal_3175), .A1_t (new_AGEMA_signal_3176), .A1_f (new_AGEMA_signal_3177), .B0_t (port_out_s0_t[7]), .B0_f (port_out_s0_f[7]), .B1_t (port_out_s1_t[7]), .B1_f (port_out_s1_f[7]), .Z0_t (MixColumns_line1_n15), .Z0_f (new_AGEMA_signal_4006), .Z1_t (new_AGEMA_signal_4007), .Z1_f (new_AGEMA_signal_4008) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_U22 ( .A0_t (MixColumns_line1_S02[7]), .A0_f (new_AGEMA_signal_3961), .A1_t (new_AGEMA_signal_3962), .A1_f (new_AGEMA_signal_3963), .B0_t (MixColumns_line1_S13[7]), .B0_f (new_AGEMA_signal_4039), .B1_t (new_AGEMA_signal_4040), .B1_f (new_AGEMA_signal_4041), .Z0_t (MixColumns_line1_n16), .Z0_f (new_AGEMA_signal_4595), .Z1_t (new_AGEMA_signal_4596), .Z1_f (new_AGEMA_signal_4597) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line1_U21 ( .A0_t (MixColumns_line1_n14), .A0_f (new_AGEMA_signal_4598), .A1_t (new_AGEMA_signal_4599), .A1_f (new_AGEMA_signal_4600), .B0_t (MixColumns_line1_n13), .B0_f (new_AGEMA_signal_4009), .B1_t (new_AGEMA_signal_4010), .B1_f (new_AGEMA_signal_4011), .Z0_t (MCout[22]), .Z0_f (new_AGEMA_signal_5064), .Z1_t (new_AGEMA_signal_5065), .Z1_f (new_AGEMA_signal_5066) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line1_U20 ( .A0_t (MixColumns_line3_S02[7]), .A0_f (new_AGEMA_signal_3166), .A1_t (new_AGEMA_signal_3167), .A1_f (new_AGEMA_signal_3168), .B0_t (port_out_s0_t[6]), .B0_f (port_out_s0_f[6]), .B1_t (port_out_s1_t[6]), .B1_f (port_out_s1_f[6]), .Z0_t (MixColumns_line1_n13), .Z0_f (new_AGEMA_signal_4009), .Z1_t (new_AGEMA_signal_4010), .Z1_f (new_AGEMA_signal_4011) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_U19 ( .A0_t (MixColumns_line1_S02[6]), .A0_f (new_AGEMA_signal_3967), .A1_t (new_AGEMA_signal_3968), .A1_f (new_AGEMA_signal_3969), .B0_t (MixColumns_line1_S13[6]), .B0_f (new_AGEMA_signal_4042), .B1_t (new_AGEMA_signal_4043), .B1_f (new_AGEMA_signal_4044), .Z0_t (MixColumns_line1_n14), .Z0_f (new_AGEMA_signal_4598), .Z1_t (new_AGEMA_signal_4599), .Z1_f (new_AGEMA_signal_4600) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line1_U18 ( .A0_t (MixColumns_line1_n12), .A0_f (new_AGEMA_signal_4601), .A1_t (new_AGEMA_signal_4602), .A1_f (new_AGEMA_signal_4603), .B0_t (MixColumns_line1_n11), .B0_f (new_AGEMA_signal_4012), .B1_t (new_AGEMA_signal_4013), .B1_f (new_AGEMA_signal_4014), .Z0_t (MCout[21]), .Z0_f (new_AGEMA_signal_5067), .Z1_t (new_AGEMA_signal_5068), .Z1_f (new_AGEMA_signal_5069) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line1_U17 ( .A0_t (MixColumns_line3_S02[6]), .A0_f (new_AGEMA_signal_3157), .A1_t (new_AGEMA_signal_3158), .A1_f (new_AGEMA_signal_3159), .B0_t (port_out_s0_t[5]), .B0_f (port_out_s0_f[5]), .B1_t (port_out_s1_t[5]), .B1_f (port_out_s1_f[5]), .Z0_t (MixColumns_line1_n11), .Z0_f (new_AGEMA_signal_4012), .Z1_t (new_AGEMA_signal_4013), .Z1_f (new_AGEMA_signal_4014) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_U16 ( .A0_t (MixColumns_line1_S02[5]), .A0_f (new_AGEMA_signal_3973), .A1_t (new_AGEMA_signal_3974), .A1_f (new_AGEMA_signal_3975), .B0_t (MixColumns_line1_S13[5]), .B0_f (new_AGEMA_signal_4045), .B1_t (new_AGEMA_signal_4046), .B1_f (new_AGEMA_signal_4047), .Z0_t (MixColumns_line1_n12), .Z0_f (new_AGEMA_signal_4601), .Z1_t (new_AGEMA_signal_4602), .Z1_f (new_AGEMA_signal_4603) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line1_U15 ( .A0_t (MixColumns_line1_n10), .A0_f (new_AGEMA_signal_5070), .A1_t (new_AGEMA_signal_5071), .A1_f (new_AGEMA_signal_5072), .B0_t (MixColumns_line1_n9), .B0_f (new_AGEMA_signal_4015), .B1_t (new_AGEMA_signal_4016), .B1_f (new_AGEMA_signal_4017), .Z0_t (MCout[20]), .Z0_f (new_AGEMA_signal_5256), .Z1_t (new_AGEMA_signal_5257), .Z1_f (new_AGEMA_signal_5258) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line1_U14 ( .A0_t (MixColumns_line3_S02[5]), .A0_f (new_AGEMA_signal_3148), .A1_t (new_AGEMA_signal_3149), .A1_f (new_AGEMA_signal_3150), .B0_t (port_out_s0_t[4]), .B0_f (port_out_s0_f[4]), .B1_t (port_out_s1_t[4]), .B1_f (port_out_s1_f[4]), .Z0_t (MixColumns_line1_n9), .Z0_f (new_AGEMA_signal_4015), .Z1_t (new_AGEMA_signal_4016), .Z1_f (new_AGEMA_signal_4017) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_U13 ( .A0_t (MixColumns_line1_S02[4]), .A0_f (new_AGEMA_signal_4030), .A1_t (new_AGEMA_signal_4031), .A1_f (new_AGEMA_signal_4032), .B0_t (MixColumns_line1_S13[4]), .B0_f (new_AGEMA_signal_4610), .B1_t (new_AGEMA_signal_4611), .B1_f (new_AGEMA_signal_4612), .Z0_t (MixColumns_line1_n10), .Z0_f (new_AGEMA_signal_5070), .Z1_t (new_AGEMA_signal_5071), .Z1_f (new_AGEMA_signal_5072) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line1_U12 ( .A0_t (MixColumns_line1_n8), .A0_f (new_AGEMA_signal_5073), .A1_t (new_AGEMA_signal_5074), .A1_f (new_AGEMA_signal_5075), .B0_t (MixColumns_line1_n7), .B0_f (new_AGEMA_signal_4018), .B1_t (new_AGEMA_signal_4019), .B1_f (new_AGEMA_signal_4020), .Z0_t (MCout[19]), .Z0_f (new_AGEMA_signal_5259), .Z1_t (new_AGEMA_signal_5260), .Z1_f (new_AGEMA_signal_5261) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line1_U11 ( .A0_t (MCin[3]), .A0_f (new_AGEMA_signal_3139), .A1_t (new_AGEMA_signal_3140), .A1_f (new_AGEMA_signal_3141), .B0_t (port_out_s0_t[3]), .B0_f (port_out_s0_f[3]), .B1_t (port_out_s1_t[3]), .B1_f (port_out_s1_f[3]), .Z0_t (MixColumns_line1_n7), .Z0_f (new_AGEMA_signal_4018), .Z1_t (new_AGEMA_signal_4019), .Z1_f (new_AGEMA_signal_4020) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_U10 ( .A0_t (MixColumns_line1_S02[3]), .A0_f (new_AGEMA_signal_4033), .A1_t (new_AGEMA_signal_4034), .A1_f (new_AGEMA_signal_4035), .B0_t (MixColumns_line1_S13[3]), .B0_f (new_AGEMA_signal_4613), .B1_t (new_AGEMA_signal_4614), .B1_f (new_AGEMA_signal_4615), .Z0_t (MixColumns_line1_n8), .Z0_f (new_AGEMA_signal_5073), .Z1_t (new_AGEMA_signal_5074), .Z1_f (new_AGEMA_signal_5075) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line1_U9 ( .A0_t (MixColumns_line1_n6), .A0_f (new_AGEMA_signal_4604), .A1_t (new_AGEMA_signal_4605), .A1_f (new_AGEMA_signal_4606), .B0_t (MixColumns_line1_n5), .B0_f (new_AGEMA_signal_4021), .B1_t (new_AGEMA_signal_4022), .B1_f (new_AGEMA_signal_4023), .Z0_t (MCout[18]), .Z0_f (new_AGEMA_signal_5076), .Z1_t (new_AGEMA_signal_5077), .Z1_f (new_AGEMA_signal_5078) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line1_U8 ( .A0_t (MCin[2]), .A0_f (new_AGEMA_signal_3130), .A1_t (new_AGEMA_signal_3131), .A1_f (new_AGEMA_signal_3132), .B0_t (port_out_s0_t[2]), .B0_f (port_out_s0_f[2]), .B1_t (port_out_s1_t[2]), .B1_f (port_out_s1_f[2]), .Z0_t (MixColumns_line1_n5), .Z0_f (new_AGEMA_signal_4021), .Z1_t (new_AGEMA_signal_4022), .Z1_f (new_AGEMA_signal_4023) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_U7 ( .A0_t (MixColumns_line1_S02[2]), .A0_f (new_AGEMA_signal_3982), .A1_t (new_AGEMA_signal_3983), .A1_f (new_AGEMA_signal_3984), .B0_t (MixColumns_line1_S13[2]), .B0_f (new_AGEMA_signal_4048), .B1_t (new_AGEMA_signal_4049), .B1_f (new_AGEMA_signal_4050), .Z0_t (MixColumns_line1_n6), .Z0_f (new_AGEMA_signal_4604), .Z1_t (new_AGEMA_signal_4605), .Z1_f (new_AGEMA_signal_4606) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line1_U6 ( .A0_t (MixColumns_line1_n4), .A0_f (new_AGEMA_signal_5079), .A1_t (new_AGEMA_signal_5080), .A1_f (new_AGEMA_signal_5081), .B0_t (MixColumns_line1_n3), .B0_f (new_AGEMA_signal_4024), .B1_t (new_AGEMA_signal_4025), .B1_f (new_AGEMA_signal_4026), .Z0_t (MCout[17]), .Z0_f (new_AGEMA_signal_5262), .Z1_t (new_AGEMA_signal_5263), .Z1_f (new_AGEMA_signal_5264) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line1_U5 ( .A0_t (port_out_s0_t[1]), .A0_f (port_out_s0_f[1]), .A1_t (port_out_s1_t[1]), .A1_f (port_out_s1_f[1]), .B0_t (MixColumns_line3_S02[2]), .B0_f (new_AGEMA_signal_3121), .B1_t (new_AGEMA_signal_3122), .B1_f (new_AGEMA_signal_3123), .Z0_t (MixColumns_line1_n3), .Z0_f (new_AGEMA_signal_4024), .Z1_t (new_AGEMA_signal_4025), .Z1_f (new_AGEMA_signal_4026) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_U4 ( .A0_t (MixColumns_line1_S02[1]), .A0_f (new_AGEMA_signal_4036), .A1_t (new_AGEMA_signal_4037), .A1_f (new_AGEMA_signal_4038), .B0_t (MixColumns_line1_S13[1]), .B0_f (new_AGEMA_signal_4616), .B1_t (new_AGEMA_signal_4617), .B1_f (new_AGEMA_signal_4618), .Z0_t (MixColumns_line1_n4), .Z0_f (new_AGEMA_signal_5079), .Z1_t (new_AGEMA_signal_5080), .Z1_f (new_AGEMA_signal_5081) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line1_U3 ( .A0_t (MixColumns_line1_n2), .A0_f (new_AGEMA_signal_4607), .A1_t (new_AGEMA_signal_4608), .A1_f (new_AGEMA_signal_4609), .B0_t (MixColumns_line1_n1), .B0_f (new_AGEMA_signal_4027), .B1_t (new_AGEMA_signal_4028), .B1_f (new_AGEMA_signal_4029), .Z0_t (MCout[16]), .Z0_f (new_AGEMA_signal_5082), .Z1_t (new_AGEMA_signal_5083), .Z1_f (new_AGEMA_signal_5084) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line1_U2 ( .A0_t (port_out_s0_t[0]), .A0_f (port_out_s0_f[0]), .A1_t (port_out_s1_t[0]), .A1_f (port_out_s1_f[0]), .B0_t (MCin[0]), .B0_f (new_AGEMA_signal_3112), .B1_t (new_AGEMA_signal_3113), .B1_f (new_AGEMA_signal_3114), .Z0_t (MixColumns_line1_n1), .Z0_f (new_AGEMA_signal_4027), .Z1_t (new_AGEMA_signal_4028), .Z1_f (new_AGEMA_signal_4029) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_U1 ( .A0_t (MixColumns_line1_S02[0]), .A0_f (new_AGEMA_signal_3958), .A1_t (new_AGEMA_signal_3959), .A1_f (new_AGEMA_signal_3960), .B0_t (MixColumns_line1_S13[0]), .B0_f (new_AGEMA_signal_4051), .B1_t (new_AGEMA_signal_4052), .B1_f (new_AGEMA_signal_4053), .Z0_t (MixColumns_line1_n2), .Z0_f (new_AGEMA_signal_4607), .Z1_t (new_AGEMA_signal_4608), .Z1_f (new_AGEMA_signal_4609) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_timesTWO_U3 ( .A0_t (MixColumns_line1_S02[0]), .A0_f (new_AGEMA_signal_3958), .A1_t (new_AGEMA_signal_3959), .A1_f (new_AGEMA_signal_3960), .B0_t (MCin[19]), .B0_f (new_AGEMA_signal_3994), .B1_t (new_AGEMA_signal_3995), .B1_f (new_AGEMA_signal_3996), .Z0_t (MixColumns_line1_S02[4]), .Z0_f (new_AGEMA_signal_4030), .Z1_t (new_AGEMA_signal_4031), .Z1_f (new_AGEMA_signal_4032) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_timesTWO_U2 ( .A0_t (MixColumns_line1_S02[0]), .A0_f (new_AGEMA_signal_3958), .A1_t (new_AGEMA_signal_3959), .A1_f (new_AGEMA_signal_3960), .B0_t (MCin[18]), .B0_f (new_AGEMA_signal_3979), .B1_t (new_AGEMA_signal_3980), .B1_f (new_AGEMA_signal_3981), .Z0_t (MixColumns_line1_S02[3]), .Z0_f (new_AGEMA_signal_4033), .Z1_t (new_AGEMA_signal_4034), .Z1_f (new_AGEMA_signal_4035) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_timesTWO_U1 ( .A0_t (MixColumns_line1_S02[0]), .A0_f (new_AGEMA_signal_3958), .A1_t (new_AGEMA_signal_3959), .A1_f (new_AGEMA_signal_3960), .B0_t (MCin[16]), .B0_f (new_AGEMA_signal_3988), .B1_t (new_AGEMA_signal_3989), .B1_f (new_AGEMA_signal_3990), .Z0_t (MixColumns_line1_S02[1]), .Z0_f (new_AGEMA_signal_4036), .Z1_t (new_AGEMA_signal_4037), .Z1_f (new_AGEMA_signal_4038) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_timesTHREE_U8 ( .A0_t (MixColumns_line2_S02[0]), .A0_f (new_AGEMA_signal_3031), .A1_t (new_AGEMA_signal_3032), .A1_f (new_AGEMA_signal_3033), .B0_t (MixColumns_line2_S02[7]), .B0_f (new_AGEMA_signal_3025), .B1_t (new_AGEMA_signal_3026), .B1_f (new_AGEMA_signal_3027), .Z0_t (MixColumns_line1_S13[7]), .Z0_f (new_AGEMA_signal_4039), .Z1_t (new_AGEMA_signal_4040), .Z1_f (new_AGEMA_signal_4041) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_timesTHREE_U7 ( .A0_t (MixColumns_line2_S02[7]), .A0_f (new_AGEMA_signal_3025), .A1_t (new_AGEMA_signal_3026), .A1_f (new_AGEMA_signal_3027), .B0_t (MixColumns_line2_S02[6]), .B0_f (new_AGEMA_signal_3019), .B1_t (new_AGEMA_signal_3020), .B1_f (new_AGEMA_signal_3021), .Z0_t (MixColumns_line1_S13[6]), .Z0_f (new_AGEMA_signal_4042), .Z1_t (new_AGEMA_signal_4043), .Z1_f (new_AGEMA_signal_4044) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_timesTHREE_U6 ( .A0_t (MixColumns_line2_S02[6]), .A0_f (new_AGEMA_signal_3019), .A1_t (new_AGEMA_signal_3020), .A1_f (new_AGEMA_signal_3021), .B0_t (MixColumns_line2_S02[5]), .B0_f (new_AGEMA_signal_3013), .B1_t (new_AGEMA_signal_3014), .B1_f (new_AGEMA_signal_3015), .Z0_t (MixColumns_line1_S13[5]), .Z0_f (new_AGEMA_signal_4045), .Z1_t (new_AGEMA_signal_4046), .Z1_f (new_AGEMA_signal_4047) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_timesTHREE_U5 ( .A0_t (MixColumns_line2_S02[5]), .A0_f (new_AGEMA_signal_3013), .A1_t (new_AGEMA_signal_3014), .A1_f (new_AGEMA_signal_3015), .B0_t (MixColumns_line1_timesTHREE_input2[4]), .B0_f (new_AGEMA_signal_4054), .B1_t (new_AGEMA_signal_4055), .B1_f (new_AGEMA_signal_4056), .Z0_t (MixColumns_line1_S13[4]), .Z0_f (new_AGEMA_signal_4610), .Z1_t (new_AGEMA_signal_4611), .Z1_f (new_AGEMA_signal_4612) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_timesTHREE_U4 ( .A0_t (MCin[11]), .A0_f (new_AGEMA_signal_3007), .A1_t (new_AGEMA_signal_3008), .A1_f (new_AGEMA_signal_3009), .B0_t (MixColumns_line1_timesTHREE_input2[3]), .B0_f (new_AGEMA_signal_4057), .B1_t (new_AGEMA_signal_4058), .B1_f (new_AGEMA_signal_4059), .Z0_t (MixColumns_line1_S13[3]), .Z0_f (new_AGEMA_signal_4613), .Z1_t (new_AGEMA_signal_4614), .Z1_f (new_AGEMA_signal_4615) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_timesTHREE_U3 ( .A0_t (MCin[10]), .A0_f (new_AGEMA_signal_3001), .A1_t (new_AGEMA_signal_3002), .A1_f (new_AGEMA_signal_3003), .B0_t (MixColumns_line2_S02[2]), .B0_f (new_AGEMA_signal_2995), .B1_t (new_AGEMA_signal_2996), .B1_f (new_AGEMA_signal_2997), .Z0_t (MixColumns_line1_S13[2]), .Z0_f (new_AGEMA_signal_4048), .Z1_t (new_AGEMA_signal_4049), .Z1_f (new_AGEMA_signal_4050) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_timesTHREE_U2 ( .A0_t (MixColumns_line2_S02[2]), .A0_f (new_AGEMA_signal_2995), .A1_t (new_AGEMA_signal_2996), .A1_f (new_AGEMA_signal_2997), .B0_t (MixColumns_line1_timesTHREE_input2[1]), .B0_f (new_AGEMA_signal_4060), .B1_t (new_AGEMA_signal_4061), .B1_f (new_AGEMA_signal_4062), .Z0_t (MixColumns_line1_S13[1]), .Z0_f (new_AGEMA_signal_4616), .Z1_t (new_AGEMA_signal_4617), .Z1_f (new_AGEMA_signal_4618) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_timesTHREE_U1 ( .A0_t (MCin[8]), .A0_f (new_AGEMA_signal_2989), .A1_t (new_AGEMA_signal_2990), .A1_f (new_AGEMA_signal_2991), .B0_t (MixColumns_line2_S02[0]), .B0_f (new_AGEMA_signal_3031), .B1_t (new_AGEMA_signal_3032), .B1_f (new_AGEMA_signal_3033), .Z0_t (MixColumns_line1_S13[0]), .Z0_f (new_AGEMA_signal_4051), .Z1_t (new_AGEMA_signal_4052), .Z1_f (new_AGEMA_signal_4053) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_timesTHREE_timesTWO_U3 ( .A0_t (MixColumns_line2_S02[0]), .A0_f (new_AGEMA_signal_3031), .A1_t (new_AGEMA_signal_3032), .A1_f (new_AGEMA_signal_3033), .B0_t (MCin[11]), .B0_f (new_AGEMA_signal_3007), .B1_t (new_AGEMA_signal_3008), .B1_f (new_AGEMA_signal_3009), .Z0_t (MixColumns_line1_timesTHREE_input2[4]), .Z0_f (new_AGEMA_signal_4054), .Z1_t (new_AGEMA_signal_4055), .Z1_f (new_AGEMA_signal_4056) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_timesTHREE_timesTWO_U2 ( .A0_t (MixColumns_line2_S02[0]), .A0_f (new_AGEMA_signal_3031), .A1_t (new_AGEMA_signal_3032), .A1_f (new_AGEMA_signal_3033), .B0_t (MCin[10]), .B0_f (new_AGEMA_signal_3001), .B1_t (new_AGEMA_signal_3002), .B1_f (new_AGEMA_signal_3003), .Z0_t (MixColumns_line1_timesTHREE_input2[3]), .Z0_f (new_AGEMA_signal_4057), .Z1_t (new_AGEMA_signal_4058), .Z1_f (new_AGEMA_signal_4059) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line1_timesTHREE_timesTWO_U1 ( .A0_t (MixColumns_line2_S02[0]), .A0_f (new_AGEMA_signal_3031), .A1_t (new_AGEMA_signal_3032), .A1_f (new_AGEMA_signal_3033), .B0_t (MCin[8]), .B0_f (new_AGEMA_signal_2989), .B1_t (new_AGEMA_signal_2990), .B1_f (new_AGEMA_signal_2991), .Z0_t (MixColumns_line1_timesTHREE_input2[1]), .Z0_f (new_AGEMA_signal_4060), .Z1_t (new_AGEMA_signal_4061), .Z1_f (new_AGEMA_signal_4062) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line2_U24 ( .A0_t (MixColumns_line2_n16), .A0_f (new_AGEMA_signal_4619), .A1_t (new_AGEMA_signal_4620), .A1_f (new_AGEMA_signal_4621), .B0_t (MixColumns_line2_n15), .B0_f (new_AGEMA_signal_4063), .B1_t (new_AGEMA_signal_4064), .B1_f (new_AGEMA_signal_4065), .Z0_t (MCout[15]), .Z0_f (new_AGEMA_signal_5085), .Z1_t (new_AGEMA_signal_5086), .Z1_f (new_AGEMA_signal_5087) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line2_U23 ( .A0_t (port_out_s0_t[7]), .A0_f (port_out_s0_f[7]), .A1_t (port_out_s1_t[7]), .A1_f (port_out_s1_f[7]), .B0_t (MixColumns_line1_S02[0]), .B0_f (new_AGEMA_signal_3958), .B1_t (new_AGEMA_signal_3959), .B1_f (new_AGEMA_signal_3960), .Z0_t (MixColumns_line2_n15), .Z0_f (new_AGEMA_signal_4063), .Z1_t (new_AGEMA_signal_4064), .Z1_f (new_AGEMA_signal_4065) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_U22 ( .A0_t (MixColumns_line2_S02[7]), .A0_f (new_AGEMA_signal_3025), .A1_t (new_AGEMA_signal_3026), .A1_f (new_AGEMA_signal_3027), .B0_t (MixColumns_line2_S13[7]), .B0_f (new_AGEMA_signal_4096), .B1_t (new_AGEMA_signal_4097), .B1_f (new_AGEMA_signal_4098), .Z0_t (MixColumns_line2_n16), .Z0_f (new_AGEMA_signal_4619), .Z1_t (new_AGEMA_signal_4620), .Z1_f (new_AGEMA_signal_4621) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line2_U21 ( .A0_t (MixColumns_line2_n14), .A0_f (new_AGEMA_signal_4622), .A1_t (new_AGEMA_signal_4623), .A1_f (new_AGEMA_signal_4624), .B0_t (MixColumns_line2_n13), .B0_f (new_AGEMA_signal_4066), .B1_t (new_AGEMA_signal_4067), .B1_f (new_AGEMA_signal_4068), .Z0_t (MCout[14]), .Z0_f (new_AGEMA_signal_5088), .Z1_t (new_AGEMA_signal_5089), .Z1_f (new_AGEMA_signal_5090) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line2_U20 ( .A0_t (port_out_s0_t[6]), .A0_f (port_out_s0_f[6]), .A1_t (port_out_s1_t[6]), .A1_f (port_out_s1_f[6]), .B0_t (MixColumns_line1_S02[7]), .B0_f (new_AGEMA_signal_3961), .B1_t (new_AGEMA_signal_3962), .B1_f (new_AGEMA_signal_3963), .Z0_t (MixColumns_line2_n13), .Z0_f (new_AGEMA_signal_4066), .Z1_t (new_AGEMA_signal_4067), .Z1_f (new_AGEMA_signal_4068) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_U19 ( .A0_t (MixColumns_line2_S02[6]), .A0_f (new_AGEMA_signal_3019), .A1_t (new_AGEMA_signal_3020), .A1_f (new_AGEMA_signal_3021), .B0_t (MixColumns_line2_S13[6]), .B0_f (new_AGEMA_signal_4099), .B1_t (new_AGEMA_signal_4100), .B1_f (new_AGEMA_signal_4101), .Z0_t (MixColumns_line2_n14), .Z0_f (new_AGEMA_signal_4622), .Z1_t (new_AGEMA_signal_4623), .Z1_f (new_AGEMA_signal_4624) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line2_U18 ( .A0_t (MixColumns_line2_n12), .A0_f (new_AGEMA_signal_4625), .A1_t (new_AGEMA_signal_4626), .A1_f (new_AGEMA_signal_4627), .B0_t (MixColumns_line2_n11), .B0_f (new_AGEMA_signal_4069), .B1_t (new_AGEMA_signal_4070), .B1_f (new_AGEMA_signal_4071), .Z0_t (MCout[13]), .Z0_f (new_AGEMA_signal_5091), .Z1_t (new_AGEMA_signal_5092), .Z1_f (new_AGEMA_signal_5093) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line2_U17 ( .A0_t (port_out_s0_t[5]), .A0_f (port_out_s0_f[5]), .A1_t (port_out_s1_t[5]), .A1_f (port_out_s1_f[5]), .B0_t (MixColumns_line1_S02[6]), .B0_f (new_AGEMA_signal_3967), .B1_t (new_AGEMA_signal_3968), .B1_f (new_AGEMA_signal_3969), .Z0_t (MixColumns_line2_n11), .Z0_f (new_AGEMA_signal_4069), .Z1_t (new_AGEMA_signal_4070), .Z1_f (new_AGEMA_signal_4071) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_U16 ( .A0_t (MixColumns_line2_S02[5]), .A0_f (new_AGEMA_signal_3013), .A1_t (new_AGEMA_signal_3014), .A1_f (new_AGEMA_signal_3015), .B0_t (MixColumns_line2_S13[5]), .B0_f (new_AGEMA_signal_4102), .B1_t (new_AGEMA_signal_4103), .B1_f (new_AGEMA_signal_4104), .Z0_t (MixColumns_line2_n12), .Z0_f (new_AGEMA_signal_4625), .Z1_t (new_AGEMA_signal_4626), .Z1_f (new_AGEMA_signal_4627) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line2_U15 ( .A0_t (MixColumns_line2_n10), .A0_f (new_AGEMA_signal_5094), .A1_t (new_AGEMA_signal_5095), .A1_f (new_AGEMA_signal_5096), .B0_t (MixColumns_line2_n9), .B0_f (new_AGEMA_signal_4072), .B1_t (new_AGEMA_signal_4073), .B1_f (new_AGEMA_signal_4074), .Z0_t (MCout[12]), .Z0_f (new_AGEMA_signal_5265), .Z1_t (new_AGEMA_signal_5266), .Z1_f (new_AGEMA_signal_5267) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line2_U14 ( .A0_t (port_out_s0_t[4]), .A0_f (port_out_s0_f[4]), .A1_t (port_out_s1_t[4]), .A1_f (port_out_s1_f[4]), .B0_t (MixColumns_line1_S02[5]), .B0_f (new_AGEMA_signal_3973), .B1_t (new_AGEMA_signal_3974), .B1_f (new_AGEMA_signal_3975), .Z0_t (MixColumns_line2_n9), .Z0_f (new_AGEMA_signal_4072), .Z1_t (new_AGEMA_signal_4073), .Z1_f (new_AGEMA_signal_4074) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_U13 ( .A0_t (MixColumns_line2_S02[4]), .A0_f (new_AGEMA_signal_4087), .A1_t (new_AGEMA_signal_4088), .A1_f (new_AGEMA_signal_4089), .B0_t (MixColumns_line2_S13[4]), .B0_f (new_AGEMA_signal_4634), .B1_t (new_AGEMA_signal_4635), .B1_f (new_AGEMA_signal_4636), .Z0_t (MixColumns_line2_n10), .Z0_f (new_AGEMA_signal_5094), .Z1_t (new_AGEMA_signal_5095), .Z1_f (new_AGEMA_signal_5096) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line2_U12 ( .A0_t (MixColumns_line2_n8), .A0_f (new_AGEMA_signal_5097), .A1_t (new_AGEMA_signal_5098), .A1_f (new_AGEMA_signal_5099), .B0_t (MixColumns_line2_n7), .B0_f (new_AGEMA_signal_4075), .B1_t (new_AGEMA_signal_4076), .B1_f (new_AGEMA_signal_4077), .Z0_t (MCout[11]), .Z0_f (new_AGEMA_signal_5268), .Z1_t (new_AGEMA_signal_5269), .Z1_f (new_AGEMA_signal_5270) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line2_U11 ( .A0_t (port_out_s0_t[3]), .A0_f (port_out_s0_f[3]), .A1_t (port_out_s1_t[3]), .A1_f (port_out_s1_f[3]), .B0_t (MCin[19]), .B0_f (new_AGEMA_signal_3994), .B1_t (new_AGEMA_signal_3995), .B1_f (new_AGEMA_signal_3996), .Z0_t (MixColumns_line2_n7), .Z0_f (new_AGEMA_signal_4075), .Z1_t (new_AGEMA_signal_4076), .Z1_f (new_AGEMA_signal_4077) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_U10 ( .A0_t (MixColumns_line2_S02[3]), .A0_f (new_AGEMA_signal_4090), .A1_t (new_AGEMA_signal_4091), .A1_f (new_AGEMA_signal_4092), .B0_t (MixColumns_line2_S13[3]), .B0_f (new_AGEMA_signal_4637), .B1_t (new_AGEMA_signal_4638), .B1_f (new_AGEMA_signal_4639), .Z0_t (MixColumns_line2_n8), .Z0_f (new_AGEMA_signal_5097), .Z1_t (new_AGEMA_signal_5098), .Z1_f (new_AGEMA_signal_5099) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line2_U9 ( .A0_t (MixColumns_line2_n6), .A0_f (new_AGEMA_signal_4628), .A1_t (new_AGEMA_signal_4629), .A1_f (new_AGEMA_signal_4630), .B0_t (MixColumns_line2_n5), .B0_f (new_AGEMA_signal_4078), .B1_t (new_AGEMA_signal_4079), .B1_f (new_AGEMA_signal_4080), .Z0_t (MCout[10]), .Z0_f (new_AGEMA_signal_5100), .Z1_t (new_AGEMA_signal_5101), .Z1_f (new_AGEMA_signal_5102) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line2_U8 ( .A0_t (port_out_s0_t[2]), .A0_f (port_out_s0_f[2]), .A1_t (port_out_s1_t[2]), .A1_f (port_out_s1_f[2]), .B0_t (MCin[18]), .B0_f (new_AGEMA_signal_3979), .B1_t (new_AGEMA_signal_3980), .B1_f (new_AGEMA_signal_3981), .Z0_t (MixColumns_line2_n5), .Z0_f (new_AGEMA_signal_4078), .Z1_t (new_AGEMA_signal_4079), .Z1_f (new_AGEMA_signal_4080) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_U7 ( .A0_t (MixColumns_line2_S02[2]), .A0_f (new_AGEMA_signal_2995), .A1_t (new_AGEMA_signal_2996), .A1_f (new_AGEMA_signal_2997), .B0_t (MixColumns_line2_S13[2]), .B0_f (new_AGEMA_signal_4105), .B1_t (new_AGEMA_signal_4106), .B1_f (new_AGEMA_signal_4107), .Z0_t (MixColumns_line2_n6), .Z0_f (new_AGEMA_signal_4628), .Z1_t (new_AGEMA_signal_4629), .Z1_f (new_AGEMA_signal_4630) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line2_U6 ( .A0_t (MixColumns_line2_n4), .A0_f (new_AGEMA_signal_5103), .A1_t (new_AGEMA_signal_5104), .A1_f (new_AGEMA_signal_5105), .B0_t (MixColumns_line2_n3), .B0_f (new_AGEMA_signal_4081), .B1_t (new_AGEMA_signal_4082), .B1_f (new_AGEMA_signal_4083), .Z0_t (MCout[9]), .Z0_f (new_AGEMA_signal_5271), .Z1_t (new_AGEMA_signal_5272), .Z1_f (new_AGEMA_signal_5273) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line2_U5 ( .A0_t (MixColumns_line1_S02[2]), .A0_f (new_AGEMA_signal_3982), .A1_t (new_AGEMA_signal_3983), .A1_f (new_AGEMA_signal_3984), .B0_t (port_out_s0_t[1]), .B0_f (port_out_s0_f[1]), .B1_t (port_out_s1_t[1]), .B1_f (port_out_s1_f[1]), .Z0_t (MixColumns_line2_n3), .Z0_f (new_AGEMA_signal_4081), .Z1_t (new_AGEMA_signal_4082), .Z1_f (new_AGEMA_signal_4083) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_U4 ( .A0_t (MixColumns_line2_S02[1]), .A0_f (new_AGEMA_signal_4093), .A1_t (new_AGEMA_signal_4094), .A1_f (new_AGEMA_signal_4095), .B0_t (MixColumns_line2_S13[1]), .B0_f (new_AGEMA_signal_4640), .B1_t (new_AGEMA_signal_4641), .B1_f (new_AGEMA_signal_4642), .Z0_t (MixColumns_line2_n4), .Z0_f (new_AGEMA_signal_5103), .Z1_t (new_AGEMA_signal_5104), .Z1_f (new_AGEMA_signal_5105) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line2_U3 ( .A0_t (MixColumns_line2_n2), .A0_f (new_AGEMA_signal_4631), .A1_t (new_AGEMA_signal_4632), .A1_f (new_AGEMA_signal_4633), .B0_t (MixColumns_line2_n1), .B0_f (new_AGEMA_signal_4084), .B1_t (new_AGEMA_signal_4085), .B1_f (new_AGEMA_signal_4086), .Z0_t (MCout[8]), .Z0_f (new_AGEMA_signal_5106), .Z1_t (new_AGEMA_signal_5107), .Z1_f (new_AGEMA_signal_5108) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line2_U2 ( .A0_t (MCin[16]), .A0_f (new_AGEMA_signal_3988), .A1_t (new_AGEMA_signal_3989), .A1_f (new_AGEMA_signal_3990), .B0_t (port_out_s0_t[0]), .B0_f (port_out_s0_f[0]), .B1_t (port_out_s1_t[0]), .B1_f (port_out_s1_f[0]), .Z0_t (MixColumns_line2_n1), .Z0_f (new_AGEMA_signal_4084), .Z1_t (new_AGEMA_signal_4085), .Z1_f (new_AGEMA_signal_4086) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_U1 ( .A0_t (MixColumns_line2_S02[0]), .A0_f (new_AGEMA_signal_3031), .A1_t (new_AGEMA_signal_3032), .A1_f (new_AGEMA_signal_3033), .B0_t (MixColumns_line2_S13[0]), .B0_f (new_AGEMA_signal_4108), .B1_t (new_AGEMA_signal_4109), .B1_f (new_AGEMA_signal_4110), .Z0_t (MixColumns_line2_n2), .Z0_f (new_AGEMA_signal_4631), .Z1_t (new_AGEMA_signal_4632), .Z1_f (new_AGEMA_signal_4633) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_timesTWO_U3 ( .A0_t (MixColumns_line2_S02[0]), .A0_f (new_AGEMA_signal_3031), .A1_t (new_AGEMA_signal_3032), .A1_f (new_AGEMA_signal_3033), .B0_t (MCin[11]), .B0_f (new_AGEMA_signal_3007), .B1_t (new_AGEMA_signal_3008), .B1_f (new_AGEMA_signal_3009), .Z0_t (MixColumns_line2_S02[4]), .Z0_f (new_AGEMA_signal_4087), .Z1_t (new_AGEMA_signal_4088), .Z1_f (new_AGEMA_signal_4089) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_timesTWO_U2 ( .A0_t (MixColumns_line2_S02[0]), .A0_f (new_AGEMA_signal_3031), .A1_t (new_AGEMA_signal_3032), .A1_f (new_AGEMA_signal_3033), .B0_t (MCin[10]), .B0_f (new_AGEMA_signal_3001), .B1_t (new_AGEMA_signal_3002), .B1_f (new_AGEMA_signal_3003), .Z0_t (MixColumns_line2_S02[3]), .Z0_f (new_AGEMA_signal_4090), .Z1_t (new_AGEMA_signal_4091), .Z1_f (new_AGEMA_signal_4092) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_timesTWO_U1 ( .A0_t (MixColumns_line2_S02[0]), .A0_f (new_AGEMA_signal_3031), .A1_t (new_AGEMA_signal_3032), .A1_f (new_AGEMA_signal_3033), .B0_t (MCin[8]), .B0_f (new_AGEMA_signal_2989), .B1_t (new_AGEMA_signal_2990), .B1_f (new_AGEMA_signal_2991), .Z0_t (MixColumns_line2_S02[1]), .Z0_f (new_AGEMA_signal_4093), .Z1_t (new_AGEMA_signal_4094), .Z1_f (new_AGEMA_signal_4095) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_timesTHREE_U8 ( .A0_t (MixColumns_line3_S02[0]), .A0_f (new_AGEMA_signal_3175), .A1_t (new_AGEMA_signal_3176), .A1_f (new_AGEMA_signal_3177), .B0_t (MixColumns_line3_S02[7]), .B0_f (new_AGEMA_signal_3166), .B1_t (new_AGEMA_signal_3167), .B1_f (new_AGEMA_signal_3168), .Z0_t (MixColumns_line2_S13[7]), .Z0_f (new_AGEMA_signal_4096), .Z1_t (new_AGEMA_signal_4097), .Z1_f (new_AGEMA_signal_4098) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_timesTHREE_U7 ( .A0_t (MixColumns_line3_S02[7]), .A0_f (new_AGEMA_signal_3166), .A1_t (new_AGEMA_signal_3167), .A1_f (new_AGEMA_signal_3168), .B0_t (MixColumns_line3_S02[6]), .B0_f (new_AGEMA_signal_3157), .B1_t (new_AGEMA_signal_3158), .B1_f (new_AGEMA_signal_3159), .Z0_t (MixColumns_line2_S13[6]), .Z0_f (new_AGEMA_signal_4099), .Z1_t (new_AGEMA_signal_4100), .Z1_f (new_AGEMA_signal_4101) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_timesTHREE_U6 ( .A0_t (MixColumns_line3_S02[6]), .A0_f (new_AGEMA_signal_3157), .A1_t (new_AGEMA_signal_3158), .A1_f (new_AGEMA_signal_3159), .B0_t (MixColumns_line3_S02[5]), .B0_f (new_AGEMA_signal_3148), .B1_t (new_AGEMA_signal_3149), .B1_f (new_AGEMA_signal_3150), .Z0_t (MixColumns_line2_S13[5]), .Z0_f (new_AGEMA_signal_4102), .Z1_t (new_AGEMA_signal_4103), .Z1_f (new_AGEMA_signal_4104) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_timesTHREE_U5 ( .A0_t (MixColumns_line3_S02[5]), .A0_f (new_AGEMA_signal_3148), .A1_t (new_AGEMA_signal_3149), .A1_f (new_AGEMA_signal_3150), .B0_t (MixColumns_line2_timesTHREE_input2[4]), .B0_f (new_AGEMA_signal_4111), .B1_t (new_AGEMA_signal_4112), .B1_f (new_AGEMA_signal_4113), .Z0_t (MixColumns_line2_S13[4]), .Z0_f (new_AGEMA_signal_4634), .Z1_t (new_AGEMA_signal_4635), .Z1_f (new_AGEMA_signal_4636) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_timesTHREE_U4 ( .A0_t (MCin[3]), .A0_f (new_AGEMA_signal_3139), .A1_t (new_AGEMA_signal_3140), .A1_f (new_AGEMA_signal_3141), .B0_t (MixColumns_line2_timesTHREE_input2[3]), .B0_f (new_AGEMA_signal_4114), .B1_t (new_AGEMA_signal_4115), .B1_f (new_AGEMA_signal_4116), .Z0_t (MixColumns_line2_S13[3]), .Z0_f (new_AGEMA_signal_4637), .Z1_t (new_AGEMA_signal_4638), .Z1_f (new_AGEMA_signal_4639) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_timesTHREE_U3 ( .A0_t (MCin[2]), .A0_f (new_AGEMA_signal_3130), .A1_t (new_AGEMA_signal_3131), .A1_f (new_AGEMA_signal_3132), .B0_t (MixColumns_line3_S02[2]), .B0_f (new_AGEMA_signal_3121), .B1_t (new_AGEMA_signal_3122), .B1_f (new_AGEMA_signal_3123), .Z0_t (MixColumns_line2_S13[2]), .Z0_f (new_AGEMA_signal_4105), .Z1_t (new_AGEMA_signal_4106), .Z1_f (new_AGEMA_signal_4107) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_timesTHREE_U2 ( .A0_t (MixColumns_line3_S02[2]), .A0_f (new_AGEMA_signal_3121), .A1_t (new_AGEMA_signal_3122), .A1_f (new_AGEMA_signal_3123), .B0_t (MixColumns_line2_timesTHREE_input2[1]), .B0_f (new_AGEMA_signal_4117), .B1_t (new_AGEMA_signal_4118), .B1_f (new_AGEMA_signal_4119), .Z0_t (MixColumns_line2_S13[1]), .Z0_f (new_AGEMA_signal_4640), .Z1_t (new_AGEMA_signal_4641), .Z1_f (new_AGEMA_signal_4642) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_timesTHREE_U1 ( .A0_t (MCin[0]), .A0_f (new_AGEMA_signal_3112), .A1_t (new_AGEMA_signal_3113), .A1_f (new_AGEMA_signal_3114), .B0_t (MixColumns_line3_S02[0]), .B0_f (new_AGEMA_signal_3175), .B1_t (new_AGEMA_signal_3176), .B1_f (new_AGEMA_signal_3177), .Z0_t (MixColumns_line2_S13[0]), .Z0_f (new_AGEMA_signal_4108), .Z1_t (new_AGEMA_signal_4109), .Z1_f (new_AGEMA_signal_4110) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_timesTHREE_timesTWO_U3 ( .A0_t (MixColumns_line3_S02[0]), .A0_f (new_AGEMA_signal_3175), .A1_t (new_AGEMA_signal_3176), .A1_f (new_AGEMA_signal_3177), .B0_t (MCin[3]), .B0_f (new_AGEMA_signal_3139), .B1_t (new_AGEMA_signal_3140), .B1_f (new_AGEMA_signal_3141), .Z0_t (MixColumns_line2_timesTHREE_input2[4]), .Z0_f (new_AGEMA_signal_4111), .Z1_t (new_AGEMA_signal_4112), .Z1_f (new_AGEMA_signal_4113) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_timesTHREE_timesTWO_U2 ( .A0_t (MixColumns_line3_S02[0]), .A0_f (new_AGEMA_signal_3175), .A1_t (new_AGEMA_signal_3176), .A1_f (new_AGEMA_signal_3177), .B0_t (MCin[2]), .B0_f (new_AGEMA_signal_3130), .B1_t (new_AGEMA_signal_3131), .B1_f (new_AGEMA_signal_3132), .Z0_t (MixColumns_line2_timesTHREE_input2[3]), .Z0_f (new_AGEMA_signal_4114), .Z1_t (new_AGEMA_signal_4115), .Z1_f (new_AGEMA_signal_4116) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line2_timesTHREE_timesTWO_U1 ( .A0_t (MixColumns_line3_S02[0]), .A0_f (new_AGEMA_signal_3175), .A1_t (new_AGEMA_signal_3176), .A1_f (new_AGEMA_signal_3177), .B0_t (MCin[0]), .B0_f (new_AGEMA_signal_3112), .B1_t (new_AGEMA_signal_3113), .B1_f (new_AGEMA_signal_3114), .Z0_t (MixColumns_line2_timesTHREE_input2[1]), .Z0_f (new_AGEMA_signal_4117), .Z1_t (new_AGEMA_signal_4118), .Z1_f (new_AGEMA_signal_4119) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line3_U24 ( .A0_t (MixColumns_line3_n16), .A0_f (new_AGEMA_signal_4643), .A1_t (new_AGEMA_signal_4644), .A1_f (new_AGEMA_signal_4645), .B0_t (MixColumns_line3_n15), .B0_f (new_AGEMA_signal_4120), .B1_t (new_AGEMA_signal_4121), .B1_f (new_AGEMA_signal_4122), .Z0_t (MCout[7]), .Z0_f (new_AGEMA_signal_5109), .Z1_t (new_AGEMA_signal_5110), .Z1_f (new_AGEMA_signal_5111) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line3_U23 ( .A0_t (MixColumns_line1_S02[0]), .A0_f (new_AGEMA_signal_3958), .A1_t (new_AGEMA_signal_3959), .A1_f (new_AGEMA_signal_3960), .B0_t (MixColumns_line2_S02[0]), .B0_f (new_AGEMA_signal_3031), .B1_t (new_AGEMA_signal_3032), .B1_f (new_AGEMA_signal_3033), .Z0_t (MixColumns_line3_n15), .Z0_f (new_AGEMA_signal_4120), .Z1_t (new_AGEMA_signal_4121), .Z1_f (new_AGEMA_signal_4122) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_U22 ( .A0_t (MixColumns_line3_S02[7]), .A0_f (new_AGEMA_signal_3166), .A1_t (new_AGEMA_signal_3167), .A1_f (new_AGEMA_signal_3168), .B0_t (MixColumns_line3_S13[7]), .B0_f (new_AGEMA_signal_4153), .B1_t (new_AGEMA_signal_4154), .B1_f (new_AGEMA_signal_4155), .Z0_t (MixColumns_line3_n16), .Z0_f (new_AGEMA_signal_4643), .Z1_t (new_AGEMA_signal_4644), .Z1_f (new_AGEMA_signal_4645) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line3_U21 ( .A0_t (MixColumns_line3_n14), .A0_f (new_AGEMA_signal_4646), .A1_t (new_AGEMA_signal_4647), .A1_f (new_AGEMA_signal_4648), .B0_t (MixColumns_line3_n13), .B0_f (new_AGEMA_signal_4123), .B1_t (new_AGEMA_signal_4124), .B1_f (new_AGEMA_signal_4125), .Z0_t (MCout[6]), .Z0_f (new_AGEMA_signal_5112), .Z1_t (new_AGEMA_signal_5113), .Z1_f (new_AGEMA_signal_5114) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line3_U20 ( .A0_t (MixColumns_line1_S02[7]), .A0_f (new_AGEMA_signal_3961), .A1_t (new_AGEMA_signal_3962), .A1_f (new_AGEMA_signal_3963), .B0_t (MixColumns_line2_S02[7]), .B0_f (new_AGEMA_signal_3025), .B1_t (new_AGEMA_signal_3026), .B1_f (new_AGEMA_signal_3027), .Z0_t (MixColumns_line3_n13), .Z0_f (new_AGEMA_signal_4123), .Z1_t (new_AGEMA_signal_4124), .Z1_f (new_AGEMA_signal_4125) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_U19 ( .A0_t (MixColumns_line3_S02[6]), .A0_f (new_AGEMA_signal_3157), .A1_t (new_AGEMA_signal_3158), .A1_f (new_AGEMA_signal_3159), .B0_t (MixColumns_line3_S13[6]), .B0_f (new_AGEMA_signal_4156), .B1_t (new_AGEMA_signal_4157), .B1_f (new_AGEMA_signal_4158), .Z0_t (MixColumns_line3_n14), .Z0_f (new_AGEMA_signal_4646), .Z1_t (new_AGEMA_signal_4647), .Z1_f (new_AGEMA_signal_4648) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line3_U18 ( .A0_t (MixColumns_line3_n12), .A0_f (new_AGEMA_signal_4649), .A1_t (new_AGEMA_signal_4650), .A1_f (new_AGEMA_signal_4651), .B0_t (MixColumns_line3_n11), .B0_f (new_AGEMA_signal_4126), .B1_t (new_AGEMA_signal_4127), .B1_f (new_AGEMA_signal_4128), .Z0_t (MCout[5]), .Z0_f (new_AGEMA_signal_5115), .Z1_t (new_AGEMA_signal_5116), .Z1_f (new_AGEMA_signal_5117) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line3_U17 ( .A0_t (MixColumns_line1_S02[6]), .A0_f (new_AGEMA_signal_3967), .A1_t (new_AGEMA_signal_3968), .A1_f (new_AGEMA_signal_3969), .B0_t (MixColumns_line2_S02[6]), .B0_f (new_AGEMA_signal_3019), .B1_t (new_AGEMA_signal_3020), .B1_f (new_AGEMA_signal_3021), .Z0_t (MixColumns_line3_n11), .Z0_f (new_AGEMA_signal_4126), .Z1_t (new_AGEMA_signal_4127), .Z1_f (new_AGEMA_signal_4128) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_U16 ( .A0_t (MixColumns_line3_S02[5]), .A0_f (new_AGEMA_signal_3148), .A1_t (new_AGEMA_signal_3149), .A1_f (new_AGEMA_signal_3150), .B0_t (MixColumns_line3_S13[5]), .B0_f (new_AGEMA_signal_4159), .B1_t (new_AGEMA_signal_4160), .B1_f (new_AGEMA_signal_4161), .Z0_t (MixColumns_line3_n12), .Z0_f (new_AGEMA_signal_4649), .Z1_t (new_AGEMA_signal_4650), .Z1_f (new_AGEMA_signal_4651) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line3_U15 ( .A0_t (MixColumns_line3_n10), .A0_f (new_AGEMA_signal_5118), .A1_t (new_AGEMA_signal_5119), .A1_f (new_AGEMA_signal_5120), .B0_t (MixColumns_line3_n9), .B0_f (new_AGEMA_signal_4129), .B1_t (new_AGEMA_signal_4130), .B1_f (new_AGEMA_signal_4131), .Z0_t (MCout[4]), .Z0_f (new_AGEMA_signal_5274), .Z1_t (new_AGEMA_signal_5275), .Z1_f (new_AGEMA_signal_5276) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line3_U14 ( .A0_t (MixColumns_line1_S02[5]), .A0_f (new_AGEMA_signal_3973), .A1_t (new_AGEMA_signal_3974), .A1_f (new_AGEMA_signal_3975), .B0_t (MixColumns_line2_S02[5]), .B0_f (new_AGEMA_signal_3013), .B1_t (new_AGEMA_signal_3014), .B1_f (new_AGEMA_signal_3015), .Z0_t (MixColumns_line3_n9), .Z0_f (new_AGEMA_signal_4129), .Z1_t (new_AGEMA_signal_4130), .Z1_f (new_AGEMA_signal_4131) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_U13 ( .A0_t (MixColumns_line3_S02[4]), .A0_f (new_AGEMA_signal_4144), .A1_t (new_AGEMA_signal_4145), .A1_f (new_AGEMA_signal_4146), .B0_t (MixColumns_line3_S13[4]), .B0_f (new_AGEMA_signal_4658), .B1_t (new_AGEMA_signal_4659), .B1_f (new_AGEMA_signal_4660), .Z0_t (MixColumns_line3_n10), .Z0_f (new_AGEMA_signal_5118), .Z1_t (new_AGEMA_signal_5119), .Z1_f (new_AGEMA_signal_5120) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line3_U12 ( .A0_t (MixColumns_line3_n8), .A0_f (new_AGEMA_signal_5121), .A1_t (new_AGEMA_signal_5122), .A1_f (new_AGEMA_signal_5123), .B0_t (MixColumns_line3_n7), .B0_f (new_AGEMA_signal_4132), .B1_t (new_AGEMA_signal_4133), .B1_f (new_AGEMA_signal_4134), .Z0_t (MCout[3]), .Z0_f (new_AGEMA_signal_5277), .Z1_t (new_AGEMA_signal_5278), .Z1_f (new_AGEMA_signal_5279) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line3_U11 ( .A0_t (MCin[19]), .A0_f (new_AGEMA_signal_3994), .A1_t (new_AGEMA_signal_3995), .A1_f (new_AGEMA_signal_3996), .B0_t (MCin[11]), .B0_f (new_AGEMA_signal_3007), .B1_t (new_AGEMA_signal_3008), .B1_f (new_AGEMA_signal_3009), .Z0_t (MixColumns_line3_n7), .Z0_f (new_AGEMA_signal_4132), .Z1_t (new_AGEMA_signal_4133), .Z1_f (new_AGEMA_signal_4134) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_U10 ( .A0_t (MixColumns_line3_S02[3]), .A0_f (new_AGEMA_signal_4147), .A1_t (new_AGEMA_signal_4148), .A1_f (new_AGEMA_signal_4149), .B0_t (MixColumns_line3_S13[3]), .B0_f (new_AGEMA_signal_4661), .B1_t (new_AGEMA_signal_4662), .B1_f (new_AGEMA_signal_4663), .Z0_t (MixColumns_line3_n8), .Z0_f (new_AGEMA_signal_5121), .Z1_t (new_AGEMA_signal_5122), .Z1_f (new_AGEMA_signal_5123) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line3_U9 ( .A0_t (MixColumns_line3_n6), .A0_f (new_AGEMA_signal_4652), .A1_t (new_AGEMA_signal_4653), .A1_f (new_AGEMA_signal_4654), .B0_t (MixColumns_line3_n5), .B0_f (new_AGEMA_signal_4135), .B1_t (new_AGEMA_signal_4136), .B1_f (new_AGEMA_signal_4137), .Z0_t (MCout[2]), .Z0_f (new_AGEMA_signal_5124), .Z1_t (new_AGEMA_signal_5125), .Z1_f (new_AGEMA_signal_5126) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line3_U8 ( .A0_t (MCin[18]), .A0_f (new_AGEMA_signal_3979), .A1_t (new_AGEMA_signal_3980), .A1_f (new_AGEMA_signal_3981), .B0_t (MCin[10]), .B0_f (new_AGEMA_signal_3001), .B1_t (new_AGEMA_signal_3002), .B1_f (new_AGEMA_signal_3003), .Z0_t (MixColumns_line3_n5), .Z0_f (new_AGEMA_signal_4135), .Z1_t (new_AGEMA_signal_4136), .Z1_f (new_AGEMA_signal_4137) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_U7 ( .A0_t (MixColumns_line3_S02[2]), .A0_f (new_AGEMA_signal_3121), .A1_t (new_AGEMA_signal_3122), .A1_f (new_AGEMA_signal_3123), .B0_t (MixColumns_line3_S13[2]), .B0_f (new_AGEMA_signal_4162), .B1_t (new_AGEMA_signal_4163), .B1_f (new_AGEMA_signal_4164), .Z0_t (MixColumns_line3_n6), .Z0_f (new_AGEMA_signal_4652), .Z1_t (new_AGEMA_signal_4653), .Z1_f (new_AGEMA_signal_4654) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line3_U6 ( .A0_t (MixColumns_line3_n4), .A0_f (new_AGEMA_signal_5127), .A1_t (new_AGEMA_signal_5128), .A1_f (new_AGEMA_signal_5129), .B0_t (MixColumns_line3_n3), .B0_f (new_AGEMA_signal_4138), .B1_t (new_AGEMA_signal_4139), .B1_f (new_AGEMA_signal_4140), .Z0_t (MCout[1]), .Z0_f (new_AGEMA_signal_5280), .Z1_t (new_AGEMA_signal_5281), .Z1_f (new_AGEMA_signal_5282) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line3_U5 ( .A0_t (MixColumns_line2_S02[2]), .A0_f (new_AGEMA_signal_2995), .A1_t (new_AGEMA_signal_2996), .A1_f (new_AGEMA_signal_2997), .B0_t (MixColumns_line1_S02[2]), .B0_f (new_AGEMA_signal_3982), .B1_t (new_AGEMA_signal_3983), .B1_f (new_AGEMA_signal_3984), .Z0_t (MixColumns_line3_n3), .Z0_f (new_AGEMA_signal_4138), .Z1_t (new_AGEMA_signal_4139), .Z1_f (new_AGEMA_signal_4140) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_U4 ( .A0_t (MixColumns_line3_S02[1]), .A0_f (new_AGEMA_signal_4150), .A1_t (new_AGEMA_signal_4151), .A1_f (new_AGEMA_signal_4152), .B0_t (MixColumns_line3_S13[1]), .B0_f (new_AGEMA_signal_4664), .B1_t (new_AGEMA_signal_4665), .B1_f (new_AGEMA_signal_4666), .Z0_t (MixColumns_line3_n4), .Z0_f (new_AGEMA_signal_5127), .Z1_t (new_AGEMA_signal_5128), .Z1_f (new_AGEMA_signal_5129) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line3_U3 ( .A0_t (MixColumns_line3_n2), .A0_f (new_AGEMA_signal_4655), .A1_t (new_AGEMA_signal_4656), .A1_f (new_AGEMA_signal_4657), .B0_t (MixColumns_line3_n1), .B0_f (new_AGEMA_signal_4141), .B1_t (new_AGEMA_signal_4142), .B1_f (new_AGEMA_signal_4143), .Z0_t (MCout[0]), .Z0_f (new_AGEMA_signal_5130), .Z1_t (new_AGEMA_signal_5131), .Z1_f (new_AGEMA_signal_5132) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) MixColumns_line3_U2 ( .A0_t (MCin[8]), .A0_f (new_AGEMA_signal_2989), .A1_t (new_AGEMA_signal_2990), .A1_f (new_AGEMA_signal_2991), .B0_t (MCin[16]), .B0_f (new_AGEMA_signal_3988), .B1_t (new_AGEMA_signal_3989), .B1_f (new_AGEMA_signal_3990), .Z0_t (MixColumns_line3_n1), .Z0_f (new_AGEMA_signal_4141), .Z1_t (new_AGEMA_signal_4142), .Z1_f (new_AGEMA_signal_4143) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_U1 ( .A0_t (MixColumns_line3_S02[0]), .A0_f (new_AGEMA_signal_3175), .A1_t (new_AGEMA_signal_3176), .A1_f (new_AGEMA_signal_3177), .B0_t (MixColumns_line3_S13[0]), .B0_f (new_AGEMA_signal_4165), .B1_t (new_AGEMA_signal_4166), .B1_f (new_AGEMA_signal_4167), .Z0_t (MixColumns_line3_n2), .Z0_f (new_AGEMA_signal_4655), .Z1_t (new_AGEMA_signal_4656), .Z1_f (new_AGEMA_signal_4657) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_timesTWO_U3 ( .A0_t (MixColumns_line3_S02[0]), .A0_f (new_AGEMA_signal_3175), .A1_t (new_AGEMA_signal_3176), .A1_f (new_AGEMA_signal_3177), .B0_t (MCin[3]), .B0_f (new_AGEMA_signal_3139), .B1_t (new_AGEMA_signal_3140), .B1_f (new_AGEMA_signal_3141), .Z0_t (MixColumns_line3_S02[4]), .Z0_f (new_AGEMA_signal_4144), .Z1_t (new_AGEMA_signal_4145), .Z1_f (new_AGEMA_signal_4146) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_timesTWO_U2 ( .A0_t (MixColumns_line3_S02[0]), .A0_f (new_AGEMA_signal_3175), .A1_t (new_AGEMA_signal_3176), .A1_f (new_AGEMA_signal_3177), .B0_t (MCin[2]), .B0_f (new_AGEMA_signal_3130), .B1_t (new_AGEMA_signal_3131), .B1_f (new_AGEMA_signal_3132), .Z0_t (MixColumns_line3_S02[3]), .Z0_f (new_AGEMA_signal_4147), .Z1_t (new_AGEMA_signal_4148), .Z1_f (new_AGEMA_signal_4149) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_timesTWO_U1 ( .A0_t (MixColumns_line3_S02[0]), .A0_f (new_AGEMA_signal_3175), .A1_t (new_AGEMA_signal_3176), .A1_f (new_AGEMA_signal_3177), .B0_t (MCin[0]), .B0_f (new_AGEMA_signal_3112), .B1_t (new_AGEMA_signal_3113), .B1_f (new_AGEMA_signal_3114), .Z0_t (MixColumns_line3_S02[1]), .Z0_f (new_AGEMA_signal_4150), .Z1_t (new_AGEMA_signal_4151), .Z1_f (new_AGEMA_signal_4152) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_timesTHREE_U8 ( .A0_t (port_out_s0_t[7]), .A0_f (port_out_s0_f[7]), .A1_t (port_out_s1_t[7]), .A1_f (port_out_s1_f[7]), .B0_t (port_out_s0_t[6]), .B0_f (port_out_s0_f[6]), .B1_t (port_out_s1_t[6]), .B1_f (port_out_s1_f[6]), .Z0_t (MixColumns_line3_S13[7]), .Z0_f (new_AGEMA_signal_4153), .Z1_t (new_AGEMA_signal_4154), .Z1_f (new_AGEMA_signal_4155) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_timesTHREE_U7 ( .A0_t (port_out_s0_t[6]), .A0_f (port_out_s0_f[6]), .A1_t (port_out_s1_t[6]), .A1_f (port_out_s1_f[6]), .B0_t (port_out_s0_t[5]), .B0_f (port_out_s0_f[5]), .B1_t (port_out_s1_t[5]), .B1_f (port_out_s1_f[5]), .Z0_t (MixColumns_line3_S13[6]), .Z0_f (new_AGEMA_signal_4156), .Z1_t (new_AGEMA_signal_4157), .Z1_f (new_AGEMA_signal_4158) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_timesTHREE_U6 ( .A0_t (port_out_s0_t[5]), .A0_f (port_out_s0_f[5]), .A1_t (port_out_s1_t[5]), .A1_f (port_out_s1_f[5]), .B0_t (port_out_s0_t[4]), .B0_f (port_out_s0_f[4]), .B1_t (port_out_s1_t[4]), .B1_f (port_out_s1_f[4]), .Z0_t (MixColumns_line3_S13[5]), .Z0_f (new_AGEMA_signal_4159), .Z1_t (new_AGEMA_signal_4160), .Z1_f (new_AGEMA_signal_4161) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_timesTHREE_U5 ( .A0_t (port_out_s0_t[4]), .A0_f (port_out_s0_f[4]), .A1_t (port_out_s1_t[4]), .A1_f (port_out_s1_f[4]), .B0_t (MixColumns_line3_timesTHREE_input2_4_), .B0_f (new_AGEMA_signal_4168), .B1_t (new_AGEMA_signal_4169), .B1_f (new_AGEMA_signal_4170), .Z0_t (MixColumns_line3_S13[4]), .Z0_f (new_AGEMA_signal_4658), .Z1_t (new_AGEMA_signal_4659), .Z1_f (new_AGEMA_signal_4660) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_timesTHREE_U4 ( .A0_t (port_out_s0_t[3]), .A0_f (port_out_s0_f[3]), .A1_t (port_out_s1_t[3]), .A1_f (port_out_s1_f[3]), .B0_t (MixColumns_line3_timesTHREE_input2_3_), .B0_f (new_AGEMA_signal_4171), .B1_t (new_AGEMA_signal_4172), .B1_f (new_AGEMA_signal_4173), .Z0_t (MixColumns_line3_S13[3]), .Z0_f (new_AGEMA_signal_4661), .Z1_t (new_AGEMA_signal_4662), .Z1_f (new_AGEMA_signal_4663) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_timesTHREE_U3 ( .A0_t (port_out_s0_t[2]), .A0_f (port_out_s0_f[2]), .A1_t (port_out_s1_t[2]), .A1_f (port_out_s1_f[2]), .B0_t (port_out_s0_t[1]), .B0_f (port_out_s0_f[1]), .B1_t (port_out_s1_t[1]), .B1_f (port_out_s1_f[1]), .Z0_t (MixColumns_line3_S13[2]), .Z0_f (new_AGEMA_signal_4162), .Z1_t (new_AGEMA_signal_4163), .Z1_f (new_AGEMA_signal_4164) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_timesTHREE_U2 ( .A0_t (port_out_s0_t[1]), .A0_f (port_out_s0_f[1]), .A1_t (port_out_s1_t[1]), .A1_f (port_out_s1_f[1]), .B0_t (MixColumns_line3_timesTHREE_input2_1_), .B0_f (new_AGEMA_signal_4174), .B1_t (new_AGEMA_signal_4175), .B1_f (new_AGEMA_signal_4176), .Z0_t (MixColumns_line3_S13[1]), .Z0_f (new_AGEMA_signal_4664), .Z1_t (new_AGEMA_signal_4665), .Z1_f (new_AGEMA_signal_4666) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_timesTHREE_U1 ( .A0_t (port_out_s0_t[0]), .A0_f (port_out_s0_f[0]), .A1_t (port_out_s1_t[0]), .A1_f (port_out_s1_f[0]), .B0_t (port_out_s0_t[7]), .B0_f (port_out_s0_f[7]), .B1_t (port_out_s1_t[7]), .B1_f (port_out_s1_f[7]), .Z0_t (MixColumns_line3_S13[0]), .Z0_f (new_AGEMA_signal_4165), .Z1_t (new_AGEMA_signal_4166), .Z1_f (new_AGEMA_signal_4167) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_timesTHREE_timesTWO_U3 ( .A0_t (port_out_s0_t[7]), .A0_f (port_out_s0_f[7]), .A1_t (port_out_s1_t[7]), .A1_f (port_out_s1_f[7]), .B0_t (port_out_s0_t[3]), .B0_f (port_out_s0_f[3]), .B1_t (port_out_s1_t[3]), .B1_f (port_out_s1_f[3]), .Z0_t (MixColumns_line3_timesTHREE_input2_4_), .Z0_f (new_AGEMA_signal_4168), .Z1_t (new_AGEMA_signal_4169), .Z1_f (new_AGEMA_signal_4170) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_timesTHREE_timesTWO_U2 ( .A0_t (port_out_s0_t[7]), .A0_f (port_out_s0_f[7]), .A1_t (port_out_s1_t[7]), .A1_f (port_out_s1_f[7]), .B0_t (port_out_s0_t[2]), .B0_f (port_out_s0_f[2]), .B1_t (port_out_s1_t[2]), .B1_f (port_out_s1_f[2]), .Z0_t (MixColumns_line3_timesTHREE_input2_3_), .Z0_f (new_AGEMA_signal_4171), .Z1_t (new_AGEMA_signal_4172), .Z1_f (new_AGEMA_signal_4173) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MixColumns_line3_timesTHREE_timesTWO_U1 ( .A0_t (port_out_s0_t[7]), .A0_f (port_out_s0_f[7]), .A1_t (port_out_s1_t[7]), .A1_f (port_out_s1_f[7]), .B0_t (port_out_s0_t[0]), .B0_f (port_out_s0_f[0]), .B1_t (port_out_s1_t[0]), .B1_f (port_out_s1_f[0]), .Z0_t (MixColumns_line3_timesTHREE_input2_1_), .Z0_f (new_AGEMA_signal_4174), .Z1_t (new_AGEMA_signal_4175), .Z1_f (new_AGEMA_signal_4176) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U53 ( .A0_t (calcRCon_s_current_state_7_), .A0_f (new_AGEMA_signal_4177), .B0_t (enRCon), .B0_f (new_AGEMA_signal_4178), .Z0_t (roundConstant[7]), .Z0_f (new_AGEMA_signal_4179) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U52 ( .A0_t (calcRCon_s_current_state_6_), .A0_f (new_AGEMA_signal_4180), .B0_t (enRCon), .B0_f (new_AGEMA_signal_4178), .Z0_t (roundConstant[6]), .Z0_f (new_AGEMA_signal_4181) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U51 ( .A0_t (calcRCon_s_current_state_5_), .A0_f (new_AGEMA_signal_4182), .B0_t (enRCon), .B0_f (new_AGEMA_signal_4178), .Z0_t (roundConstant[5]), .Z0_f (new_AGEMA_signal_4183) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U50 ( .A0_t (calcRCon_s_current_state_4_), .A0_f (new_AGEMA_signal_4184), .B0_t (enRCon), .B0_f (new_AGEMA_signal_4178), .Z0_t (roundConstant[4]), .Z0_f (new_AGEMA_signal_4185) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U49 ( .A0_t (calcRCon_s_current_state_3_), .A0_f (new_AGEMA_signal_4186), .B0_t (enRCon), .B0_f (new_AGEMA_signal_4178), .Z0_t (roundConstant[3]), .Z0_f (new_AGEMA_signal_4187) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U48 ( .A0_t (calcRCon_s_current_state_2_), .A0_f (new_AGEMA_signal_4188), .B0_t (enRCon), .B0_f (new_AGEMA_signal_4178), .Z0_t (roundConstant[2]), .Z0_f (new_AGEMA_signal_4189) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U47 ( .A0_t (calcRCon_s_current_state_1_), .A0_f (new_AGEMA_signal_4190), .B0_t (enRCon), .B0_f (new_AGEMA_signal_4178), .Z0_t (roundConstant[1]), .Z0_f (new_AGEMA_signal_4191) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U46 ( .A0_t (calcRCon_s_current_state_0_), .A0_f (new_AGEMA_signal_4192), .B0_t (enRCon), .B0_f (new_AGEMA_signal_4178), .Z0_t (roundConstant[0]), .Z0_f (new_AGEMA_signal_4193) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) calcRCon_U44 ( .A0_t (calcRCon_n42), .A0_f (new_AGEMA_signal_4668), .B0_t (calcRCon_n41), .B0_f (new_AGEMA_signal_4667), .Z0_t (notFirst), .Z0_f (new_AGEMA_signal_5133) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U43 ( .A0_t (calcRCon_n40), .A0_f (new_AGEMA_signal_4195), .B0_t (calcRCon_n39), .B0_f (new_AGEMA_signal_4194), .Z0_t (calcRCon_n41), .Z0_f (new_AGEMA_signal_4667) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) calcRCon_U42 ( .A0_t (calcRCon_s_current_state_6_), .A0_f (new_AGEMA_signal_4180), .B0_t (calcRCon_s_current_state_5_), .B0_f (new_AGEMA_signal_4182), .Z0_t (calcRCon_n39), .Z0_f (new_AGEMA_signal_4194) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) calcRCon_U41 ( .A0_t (calcRCon_s_current_state_3_), .A0_f (new_AGEMA_signal_4186), .B0_t (calcRCon_s_current_state_7_), .B0_f (new_AGEMA_signal_4177), .Z0_t (calcRCon_n40), .Z0_f (new_AGEMA_signal_4195) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U40 ( .A0_t (calcRCon_n38), .A0_f (new_AGEMA_signal_4197), .B0_t (calcRCon_n37), .B0_f (new_AGEMA_signal_4196), .Z0_t (calcRCon_n42), .Z0_f (new_AGEMA_signal_4668) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) calcRCon_U39 ( .A0_t (calcRCon_s_current_state_2_), .A0_f (new_AGEMA_signal_4188), .B0_t (calcRCon_s_current_state_0_), .B0_f (new_AGEMA_signal_4192), .Z0_t (calcRCon_n37), .Z0_f (new_AGEMA_signal_4196) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) calcRCon_U38 ( .A0_t (calcRCon_s_current_state_1_), .A0_f (new_AGEMA_signal_4190), .B0_t (calcRCon_s_current_state_4_), .B0_f (new_AGEMA_signal_4184), .Z0_t (calcRCon_n38), .Z0_f (new_AGEMA_signal_4197) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1), .NL(1'b1)) calcRCon_U37 ( .A0_t (calcRCon_n36), .A0_f (new_AGEMA_signal_7254), .B0_t (calcRCon_n35), .B0_f (new_AGEMA_signal_7135), .Z0_t (calcRCon_s_current_state_0_), .Z0_f (new_AGEMA_signal_4192) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) calcRCon_U36 ( .A0_t (calcRCon_n34), .A0_f (new_AGEMA_signal_6303), .B0_t (calcRCon_s_current_state_0_), .B0_f (new_AGEMA_signal_4192), .Z0_t (calcRCon_n35), .Z0_f (new_AGEMA_signal_7135) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U35 ( .A0_t (start_t), .A0_f (start_f), .B0_t (calcRCon_n33), .B0_f (new_AGEMA_signal_7136), .Z0_t (calcRCon_n36), .Z0_f (new_AGEMA_signal_7254) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U34 ( .A0_t (calcRCon_n34), .A0_f (new_AGEMA_signal_6303), .B0_t (calcRCon_s_current_state_7_), .B0_f (new_AGEMA_signal_4177), .Z0_t (calcRCon_n33), .Z0_f (new_AGEMA_signal_7136) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1), .NL(1'b1)) calcRCon_U33 ( .A0_t (calcRCon_n32), .A0_f (new_AGEMA_signal_7255), .B0_t (calcRCon_n31), .B0_f (new_AGEMA_signal_7137), .Z0_t (calcRCon_s_current_state_1_), .Z0_f (new_AGEMA_signal_4190) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) calcRCon_U32 ( .A0_t (calcRCon_n34), .A0_f (new_AGEMA_signal_6303), .B0_t (calcRCon_s_current_state_1_), .B0_f (new_AGEMA_signal_4190), .Z0_t (calcRCon_n31), .Z0_f (new_AGEMA_signal_7137) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) calcRCon_U31 ( .A0_t (calcRCon_n30), .A0_f (new_AGEMA_signal_4198), .B0_t (calcRCon_n29), .B0_f (new_AGEMA_signal_7144), .Z0_t (calcRCon_n32), .Z0_f (new_AGEMA_signal_7255) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) calcRCon_U30 ( .A0_t (calcRCon_s_current_state_0_), .A0_f (new_AGEMA_signal_4192), .B0_t (calcRCon_s_current_state_7_), .B0_f (new_AGEMA_signal_4177), .Z0_t (calcRCon_n30), .Z0_f (new_AGEMA_signal_4198) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b1), .NL(1'b1)) calcRCon_U29 ( .A0_t (start_t), .A0_f (start_f), .B0_t (calcRCon_n28), .B0_f (new_AGEMA_signal_7256), .Z0_t (calcRCon_s_current_state_2_), .Z0_f (new_AGEMA_signal_4188) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U28 ( .A0_t (calcRCon_n27), .A0_f (new_AGEMA_signal_7138), .B0_t (calcRCon_n26), .B0_f (new_AGEMA_signal_6301), .Z0_t (calcRCon_n28), .Z0_f (new_AGEMA_signal_7256) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U27 ( .A0_t (ctrl_n4), .A0_f (new_AGEMA_signal_5778), .B0_t (calcRCon_s_current_state_2_), .B0_f (new_AGEMA_signal_4188), .Z0_t (calcRCon_n26), .Z0_f (new_AGEMA_signal_6301) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U26 ( .A0_t (calcRCon_n34), .A0_f (new_AGEMA_signal_6303), .B0_t (calcRCon_s_current_state_1_), .B0_f (new_AGEMA_signal_4190), .Z0_t (calcRCon_n27), .Z0_f (new_AGEMA_signal_7138) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1), .NL(1'b1)) calcRCon_U25 ( .A0_t (calcRCon_n25), .A0_f (new_AGEMA_signal_7257), .B0_t (calcRCon_n24), .B0_f (new_AGEMA_signal_7139), .Z0_t (calcRCon_s_current_state_3_), .Z0_f (new_AGEMA_signal_4186) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) calcRCon_U24 ( .A0_t (calcRCon_n34), .A0_f (new_AGEMA_signal_6303), .B0_t (calcRCon_s_current_state_3_), .B0_f (new_AGEMA_signal_4186), .Z0_t (calcRCon_n24), .Z0_f (new_AGEMA_signal_7139) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U23 ( .A0_t (calcRCon_n23), .A0_f (new_AGEMA_signal_7140), .B0_t (start_t), .B0_f (start_f), .Z0_t (calcRCon_n25), .Z0_f (new_AGEMA_signal_7257) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U22 ( .A0_t (calcRCon_n34), .A0_f (new_AGEMA_signal_6303), .B0_t (calcRCon_n22), .B0_f (new_AGEMA_signal_4199), .Z0_t (calcRCon_n23), .Z0_f (new_AGEMA_signal_7140) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) calcRCon_U21 ( .A0_t (calcRCon_s_current_state_2_), .A0_f (new_AGEMA_signal_4188), .B0_t (calcRCon_s_current_state_7_), .B0_f (new_AGEMA_signal_4177), .Z0_t (calcRCon_n22), .Z0_f (new_AGEMA_signal_4199) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1), .NL(1'b1)) calcRCon_U20 ( .A0_t (calcRCon_n21), .A0_f (new_AGEMA_signal_7258), .B0_t (calcRCon_n20), .B0_f (new_AGEMA_signal_7141), .Z0_t (calcRCon_s_current_state_4_), .Z0_f (new_AGEMA_signal_4184) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) calcRCon_U19 ( .A0_t (calcRCon_n34), .A0_f (new_AGEMA_signal_6303), .B0_t (calcRCon_s_current_state_4_), .B0_f (new_AGEMA_signal_4184), .Z0_t (calcRCon_n20), .Z0_f (new_AGEMA_signal_7141) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) calcRCon_U18 ( .A0_t (calcRCon_n19), .A0_f (new_AGEMA_signal_4200), .B0_t (calcRCon_n29), .B0_f (new_AGEMA_signal_7144), .Z0_t (calcRCon_n21), .Z0_f (new_AGEMA_signal_7258) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) calcRCon_U17 ( .A0_t (calcRCon_s_current_state_3_), .A0_f (new_AGEMA_signal_4186), .B0_t (calcRCon_s_current_state_7_), .B0_f (new_AGEMA_signal_4177), .Z0_t (calcRCon_n19), .Z0_f (new_AGEMA_signal_4200) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1), .NL(1'b1)) calcRCon_U16 ( .A0_t (calcRCon_n18), .A0_f (new_AGEMA_signal_7259), .B0_t (calcRCon_n17), .B0_f (new_AGEMA_signal_7142), .Z0_t (calcRCon_s_current_state_5_), .Z0_f (new_AGEMA_signal_4182) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) calcRCon_U15 ( .A0_t (calcRCon_s_current_state_5_), .A0_f (new_AGEMA_signal_4182), .B0_t (calcRCon_n34), .B0_f (new_AGEMA_signal_6303), .Z0_t (calcRCon_n17), .Z0_f (new_AGEMA_signal_7142) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) calcRCon_U14 ( .A0_t (calcRCon_s_current_state_4_), .A0_f (new_AGEMA_signal_4184), .B0_t (calcRCon_n29), .B0_f (new_AGEMA_signal_7144), .Z0_t (calcRCon_n18), .Z0_f (new_AGEMA_signal_7259) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b1), .NL(1'b1)) calcRCon_U13 ( .A0_t (calcRCon_n16), .A0_f (new_AGEMA_signal_7260), .B0_t (calcRCon_n15), .B0_f (new_AGEMA_signal_7143), .Z0_t (calcRCon_s_current_state_6_), .Z0_f (new_AGEMA_signal_4180) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) calcRCon_U12 ( .A0_t (calcRCon_s_current_state_6_), .A0_f (new_AGEMA_signal_4180), .B0_t (calcRCon_n34), .B0_f (new_AGEMA_signal_6303), .Z0_t (calcRCon_n15), .Z0_f (new_AGEMA_signal_7143) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) calcRCon_U11 ( .A0_t (calcRCon_s_current_state_5_), .A0_f (new_AGEMA_signal_4182), .B0_t (calcRCon_n29), .B0_f (new_AGEMA_signal_7144), .Z0_t (calcRCon_n16), .Z0_f (new_AGEMA_signal_7260) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U10 ( .A0_t (calcRCon_n34), .A0_f (new_AGEMA_signal_6303), .B0_t (start_t), .B0_f (start_f), .Z0_t (calcRCon_n29), .Z0_f (new_AGEMA_signal_7144) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b1), .NL(1'b1)) calcRCon_U9 ( .A0_t (start_t), .A0_f (start_f), .B0_t (calcRCon_n14), .B0_f (new_AGEMA_signal_7261), .Z0_t (calcRCon_s_current_state_7_), .Z0_f (new_AGEMA_signal_4177) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U8 ( .A0_t (calcRCon_n13), .A0_f (new_AGEMA_signal_7145), .B0_t (calcRCon_n9), .B0_f (new_AGEMA_signal_6302), .Z0_t (calcRCon_n14), .Z0_f (new_AGEMA_signal_7261) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U7 ( .A0_t (ctrl_n4), .A0_f (new_AGEMA_signal_5778), .B0_t (calcRCon_s_current_state_7_), .B0_f (new_AGEMA_signal_4177), .Z0_t (calcRCon_n9), .Z0_f (new_AGEMA_signal_6302) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U6 ( .A0_t (calcRCon_n34), .A0_f (new_AGEMA_signal_6303), .B0_t (calcRCon_s_current_state_6_), .B0_f (new_AGEMA_signal_4180), .Z0_t (calcRCon_n13), .Z0_f (new_AGEMA_signal_7145) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) calcRCon_U5 ( .A0_t (calcRCon_s_current_state_5_), .A0_f (new_AGEMA_signal_4182), .B0_t (calcRCon_s_current_state_4_), .B0_f (new_AGEMA_signal_4184), .Z0_t (calcRCon_n7), .Z0_f (new_AGEMA_signal_4201) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) calcRCon_U4 ( .A0_t (calcRCon_s_current_state_1_), .A0_f (new_AGEMA_signal_4190), .B0_t (calcRCon_s_current_state_2_), .B0_f (new_AGEMA_signal_4188), .Z0_t (calcRCon_n8), .Z0_f (new_AGEMA_signal_4202) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U2 ( .A0_t (ctrl_n4), .A0_f (new_AGEMA_signal_5778), .B0_t (start_t), .B0_f (start_f), .Z0_t (calcRCon_n34), .Z0_f (new_AGEMA_signal_6303) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) calcRCon_U1 ( .A0_t (calcRCon_n8), .A0_f (new_AGEMA_signal_4202), .B0_t (calcRCon_n7), .B0_f (new_AGEMA_signal_4201), .Z0_t (intFinal), .Z0_f (new_AGEMA_signal_4669) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_0_XOR1_U1 ( .A0_t (StateOutXORroundKey[0]), .A0_f (new_AGEMA_signal_2495), .A1_t (new_AGEMA_signal_2496), .A1_f (new_AGEMA_signal_2497), .B0_t (keySBIn[0]), .B0_f (new_AGEMA_signal_3400), .B1_t (new_AGEMA_signal_3401), .B1_f (new_AGEMA_signal_3402), .Z0_t (MUX_SboxIn_mux_inst_0_X), .Z0_f (new_AGEMA_signal_4670), .Z1_t (new_AGEMA_signal_4671), .Z1_f (new_AGEMA_signal_4672) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_0_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (MUX_SboxIn_mux_inst_0_X), .B0_f (new_AGEMA_signal_4670), .B1_t (new_AGEMA_signal_4671), .B1_f (new_AGEMA_signal_4672), .Z0_t (MUX_SboxIn_mux_inst_0_Y), .Z0_f (new_AGEMA_signal_5134), .Z1_t (new_AGEMA_signal_5135), .Z1_f (new_AGEMA_signal_5136) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_0_XOR2_U1 ( .A0_t (MUX_SboxIn_mux_inst_0_Y), .A0_f (new_AGEMA_signal_5134), .A1_t (new_AGEMA_signal_5135), .A1_f (new_AGEMA_signal_5136), .B0_t (StateOutXORroundKey[0]), .B0_f (new_AGEMA_signal_2495), .B1_t (new_AGEMA_signal_2496), .B1_f (new_AGEMA_signal_2497), .Z0_t (SboxIn[0]), .Z0_f (new_AGEMA_signal_5283), .Z1_t (new_AGEMA_signal_5284), .Z1_f (new_AGEMA_signal_5285) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_1_XOR1_U1 ( .A0_t (StateOutXORroundKey[1]), .A0_f (new_AGEMA_signal_2504), .A1_t (new_AGEMA_signal_2505), .A1_f (new_AGEMA_signal_2506), .B0_t (keySBIn[1]), .B0_f (new_AGEMA_signal_3409), .B1_t (new_AGEMA_signal_3410), .B1_f (new_AGEMA_signal_3411), .Z0_t (MUX_SboxIn_mux_inst_1_X), .Z0_f (new_AGEMA_signal_4673), .Z1_t (new_AGEMA_signal_4674), .Z1_f (new_AGEMA_signal_4675) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (MUX_SboxIn_mux_inst_1_X), .B0_f (new_AGEMA_signal_4673), .B1_t (new_AGEMA_signal_4674), .B1_f (new_AGEMA_signal_4675), .Z0_t (MUX_SboxIn_mux_inst_1_Y), .Z0_f (new_AGEMA_signal_5137), .Z1_t (new_AGEMA_signal_5138), .Z1_f (new_AGEMA_signal_5139) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_1_XOR2_U1 ( .A0_t (MUX_SboxIn_mux_inst_1_Y), .A0_f (new_AGEMA_signal_5137), .A1_t (new_AGEMA_signal_5138), .A1_f (new_AGEMA_signal_5139), .B0_t (StateOutXORroundKey[1]), .B0_f (new_AGEMA_signal_2504), .B1_t (new_AGEMA_signal_2505), .B1_f (new_AGEMA_signal_2506), .Z0_t (SboxIn[1]), .Z0_f (new_AGEMA_signal_5286), .Z1_t (new_AGEMA_signal_5287), .Z1_f (new_AGEMA_signal_5288) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_2_XOR1_U1 ( .A0_t (StateOutXORroundKey[2]), .A0_f (new_AGEMA_signal_2513), .A1_t (new_AGEMA_signal_2514), .A1_f (new_AGEMA_signal_2515), .B0_t (keySBIn[2]), .B0_f (new_AGEMA_signal_3418), .B1_t (new_AGEMA_signal_3419), .B1_f (new_AGEMA_signal_3420), .Z0_t (MUX_SboxIn_mux_inst_2_X), .Z0_f (new_AGEMA_signal_4676), .Z1_t (new_AGEMA_signal_4677), .Z1_f (new_AGEMA_signal_4678) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_2_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (MUX_SboxIn_mux_inst_2_X), .B0_f (new_AGEMA_signal_4676), .B1_t (new_AGEMA_signal_4677), .B1_f (new_AGEMA_signal_4678), .Z0_t (MUX_SboxIn_mux_inst_2_Y), .Z0_f (new_AGEMA_signal_5140), .Z1_t (new_AGEMA_signal_5141), .Z1_f (new_AGEMA_signal_5142) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_2_XOR2_U1 ( .A0_t (MUX_SboxIn_mux_inst_2_Y), .A0_f (new_AGEMA_signal_5140), .A1_t (new_AGEMA_signal_5141), .A1_f (new_AGEMA_signal_5142), .B0_t (StateOutXORroundKey[2]), .B0_f (new_AGEMA_signal_2513), .B1_t (new_AGEMA_signal_2514), .B1_f (new_AGEMA_signal_2515), .Z0_t (SboxIn[2]), .Z0_f (new_AGEMA_signal_5289), .Z1_t (new_AGEMA_signal_5290), .Z1_f (new_AGEMA_signal_5291) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_3_XOR1_U1 ( .A0_t (StateOutXORroundKey[3]), .A0_f (new_AGEMA_signal_2522), .A1_t (new_AGEMA_signal_2523), .A1_f (new_AGEMA_signal_2524), .B0_t (keySBIn[3]), .B0_f (new_AGEMA_signal_3427), .B1_t (new_AGEMA_signal_3428), .B1_f (new_AGEMA_signal_3429), .Z0_t (MUX_SboxIn_mux_inst_3_X), .Z0_f (new_AGEMA_signal_4679), .Z1_t (new_AGEMA_signal_4680), .Z1_f (new_AGEMA_signal_4681) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_3_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (MUX_SboxIn_mux_inst_3_X), .B0_f (new_AGEMA_signal_4679), .B1_t (new_AGEMA_signal_4680), .B1_f (new_AGEMA_signal_4681), .Z0_t (MUX_SboxIn_mux_inst_3_Y), .Z0_f (new_AGEMA_signal_5143), .Z1_t (new_AGEMA_signal_5144), .Z1_f (new_AGEMA_signal_5145) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_3_XOR2_U1 ( .A0_t (MUX_SboxIn_mux_inst_3_Y), .A0_f (new_AGEMA_signal_5143), .A1_t (new_AGEMA_signal_5144), .A1_f (new_AGEMA_signal_5145), .B0_t (StateOutXORroundKey[3]), .B0_f (new_AGEMA_signal_2522), .B1_t (new_AGEMA_signal_2523), .B1_f (new_AGEMA_signal_2524), .Z0_t (SboxIn[3]), .Z0_f (new_AGEMA_signal_5292), .Z1_t (new_AGEMA_signal_5293), .Z1_f (new_AGEMA_signal_5294) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_4_XOR1_U1 ( .A0_t (StateOutXORroundKey[4]), .A0_f (new_AGEMA_signal_2531), .A1_t (new_AGEMA_signal_2532), .A1_f (new_AGEMA_signal_2533), .B0_t (keySBIn[4]), .B0_f (new_AGEMA_signal_3436), .B1_t (new_AGEMA_signal_3437), .B1_f (new_AGEMA_signal_3438), .Z0_t (MUX_SboxIn_mux_inst_4_X), .Z0_f (new_AGEMA_signal_4682), .Z1_t (new_AGEMA_signal_4683), .Z1_f (new_AGEMA_signal_4684) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_4_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (MUX_SboxIn_mux_inst_4_X), .B0_f (new_AGEMA_signal_4682), .B1_t (new_AGEMA_signal_4683), .B1_f (new_AGEMA_signal_4684), .Z0_t (MUX_SboxIn_mux_inst_4_Y), .Z0_f (new_AGEMA_signal_5146), .Z1_t (new_AGEMA_signal_5147), .Z1_f (new_AGEMA_signal_5148) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_4_XOR2_U1 ( .A0_t (MUX_SboxIn_mux_inst_4_Y), .A0_f (new_AGEMA_signal_5146), .A1_t (new_AGEMA_signal_5147), .A1_f (new_AGEMA_signal_5148), .B0_t (StateOutXORroundKey[4]), .B0_f (new_AGEMA_signal_2531), .B1_t (new_AGEMA_signal_2532), .B1_f (new_AGEMA_signal_2533), .Z0_t (SboxIn[4]), .Z0_f (new_AGEMA_signal_5295), .Z1_t (new_AGEMA_signal_5296), .Z1_f (new_AGEMA_signal_5297) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_5_XOR1_U1 ( .A0_t (StateOutXORroundKey[5]), .A0_f (new_AGEMA_signal_2540), .A1_t (new_AGEMA_signal_2541), .A1_f (new_AGEMA_signal_2542), .B0_t (keySBIn[5]), .B0_f (new_AGEMA_signal_3445), .B1_t (new_AGEMA_signal_3446), .B1_f (new_AGEMA_signal_3447), .Z0_t (MUX_SboxIn_mux_inst_5_X), .Z0_f (new_AGEMA_signal_4685), .Z1_t (new_AGEMA_signal_4686), .Z1_f (new_AGEMA_signal_4687) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_5_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (MUX_SboxIn_mux_inst_5_X), .B0_f (new_AGEMA_signal_4685), .B1_t (new_AGEMA_signal_4686), .B1_f (new_AGEMA_signal_4687), .Z0_t (MUX_SboxIn_mux_inst_5_Y), .Z0_f (new_AGEMA_signal_5149), .Z1_t (new_AGEMA_signal_5150), .Z1_f (new_AGEMA_signal_5151) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_5_XOR2_U1 ( .A0_t (MUX_SboxIn_mux_inst_5_Y), .A0_f (new_AGEMA_signal_5149), .A1_t (new_AGEMA_signal_5150), .A1_f (new_AGEMA_signal_5151), .B0_t (StateOutXORroundKey[5]), .B0_f (new_AGEMA_signal_2540), .B1_t (new_AGEMA_signal_2541), .B1_f (new_AGEMA_signal_2542), .Z0_t (SboxIn[5]), .Z0_f (new_AGEMA_signal_5298), .Z1_t (new_AGEMA_signal_5299), .Z1_f (new_AGEMA_signal_5300) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_6_XOR1_U1 ( .A0_t (StateOutXORroundKey[6]), .A0_f (new_AGEMA_signal_2549), .A1_t (new_AGEMA_signal_2550), .A1_f (new_AGEMA_signal_2551), .B0_t (keySBIn[6]), .B0_f (new_AGEMA_signal_3454), .B1_t (new_AGEMA_signal_3455), .B1_f (new_AGEMA_signal_3456), .Z0_t (MUX_SboxIn_mux_inst_6_X), .Z0_f (new_AGEMA_signal_4688), .Z1_t (new_AGEMA_signal_4689), .Z1_f (new_AGEMA_signal_4690) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_6_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (MUX_SboxIn_mux_inst_6_X), .B0_f (new_AGEMA_signal_4688), .B1_t (new_AGEMA_signal_4689), .B1_f (new_AGEMA_signal_4690), .Z0_t (MUX_SboxIn_mux_inst_6_Y), .Z0_f (new_AGEMA_signal_5152), .Z1_t (new_AGEMA_signal_5153), .Z1_f (new_AGEMA_signal_5154) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_6_XOR2_U1 ( .A0_t (MUX_SboxIn_mux_inst_6_Y), .A0_f (new_AGEMA_signal_5152), .A1_t (new_AGEMA_signal_5153), .A1_f (new_AGEMA_signal_5154), .B0_t (StateOutXORroundKey[6]), .B0_f (new_AGEMA_signal_2549), .B1_t (new_AGEMA_signal_2550), .B1_f (new_AGEMA_signal_2551), .Z0_t (SboxIn[6]), .Z0_f (new_AGEMA_signal_5301), .Z1_t (new_AGEMA_signal_5302), .Z1_f (new_AGEMA_signal_5303) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_7_XOR1_U1 ( .A0_t (StateOutXORroundKey[7]), .A0_f (new_AGEMA_signal_2558), .A1_t (new_AGEMA_signal_2559), .A1_f (new_AGEMA_signal_2560), .B0_t (keySBIn[7]), .B0_f (new_AGEMA_signal_3463), .B1_t (new_AGEMA_signal_3464), .B1_f (new_AGEMA_signal_3465), .Z0_t (MUX_SboxIn_mux_inst_7_X), .Z0_f (new_AGEMA_signal_4691), .Z1_t (new_AGEMA_signal_4692), .Z1_f (new_AGEMA_signal_4693) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_7_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selMC), .A1_f (new_AGEMA_signal_2573), .B0_t (MUX_SboxIn_mux_inst_7_X), .B0_f (new_AGEMA_signal_4691), .B1_t (new_AGEMA_signal_4692), .B1_f (new_AGEMA_signal_4693), .Z0_t (MUX_SboxIn_mux_inst_7_Y), .Z0_f (new_AGEMA_signal_5155), .Z1_t (new_AGEMA_signal_5156), .Z1_f (new_AGEMA_signal_5157) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_SboxIn_mux_inst_7_XOR2_U1 ( .A0_t (MUX_SboxIn_mux_inst_7_Y), .A0_f (new_AGEMA_signal_5155), .A1_t (new_AGEMA_signal_5156), .A1_f (new_AGEMA_signal_5157), .B0_t (StateOutXORroundKey[7]), .B0_f (new_AGEMA_signal_2558), .B1_t (new_AGEMA_signal_2559), .B1_f (new_AGEMA_signal_2560), .Z0_t (SboxIn[7]), .Z0_f (new_AGEMA_signal_5304), .Z1_t (new_AGEMA_signal_5305), .Z1_f (new_AGEMA_signal_5306) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T1_U1 ( .A0_t (SboxIn[7]), .A0_f (new_AGEMA_signal_5304), .A1_t (new_AGEMA_signal_5305), .A1_f (new_AGEMA_signal_5306), .B0_t (SboxIn[4]), .B0_f (new_AGEMA_signal_5295), .B1_t (new_AGEMA_signal_5296), .B1_f (new_AGEMA_signal_5297), .Z0_t (Inst_bSbox_T1), .Z0_f (new_AGEMA_signal_5431), .Z1_t (new_AGEMA_signal_5432), .Z1_f (new_AGEMA_signal_5433) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T2_U1 ( .A0_t (SboxIn[7]), .A0_f (new_AGEMA_signal_5304), .A1_t (new_AGEMA_signal_5305), .A1_f (new_AGEMA_signal_5306), .B0_t (SboxIn[2]), .B0_f (new_AGEMA_signal_5289), .B1_t (new_AGEMA_signal_5290), .B1_f (new_AGEMA_signal_5291), .Z0_t (Inst_bSbox_T2), .Z0_f (new_AGEMA_signal_5434), .Z1_t (new_AGEMA_signal_5435), .Z1_f (new_AGEMA_signal_5436) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T3_U1 ( .A0_t (SboxIn[7]), .A0_f (new_AGEMA_signal_5304), .A1_t (new_AGEMA_signal_5305), .A1_f (new_AGEMA_signal_5306), .B0_t (SboxIn[1]), .B0_f (new_AGEMA_signal_5286), .B1_t (new_AGEMA_signal_5287), .B1_f (new_AGEMA_signal_5288), .Z0_t (Inst_bSbox_T3), .Z0_f (new_AGEMA_signal_5437), .Z1_t (new_AGEMA_signal_5438), .Z1_f (new_AGEMA_signal_5439) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T4_U1 ( .A0_t (SboxIn[4]), .A0_f (new_AGEMA_signal_5295), .A1_t (new_AGEMA_signal_5296), .A1_f (new_AGEMA_signal_5297), .B0_t (SboxIn[2]), .B0_f (new_AGEMA_signal_5289), .B1_t (new_AGEMA_signal_5290), .B1_f (new_AGEMA_signal_5291), .Z0_t (Inst_bSbox_T4), .Z0_f (new_AGEMA_signal_5440), .Z1_t (new_AGEMA_signal_5441), .Z1_f (new_AGEMA_signal_5442) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T5_U1 ( .A0_t (SboxIn[3]), .A0_f (new_AGEMA_signal_5292), .A1_t (new_AGEMA_signal_5293), .A1_f (new_AGEMA_signal_5294), .B0_t (SboxIn[1]), .B0_f (new_AGEMA_signal_5286), .B1_t (new_AGEMA_signal_5287), .B1_f (new_AGEMA_signal_5288), .Z0_t (Inst_bSbox_T5), .Z0_f (new_AGEMA_signal_5443), .Z1_t (new_AGEMA_signal_5444), .Z1_f (new_AGEMA_signal_5445) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T6_U1 ( .A0_t (Inst_bSbox_T1), .A0_f (new_AGEMA_signal_5431), .A1_t (new_AGEMA_signal_5432), .A1_f (new_AGEMA_signal_5433), .B0_t (Inst_bSbox_T5), .B0_f (new_AGEMA_signal_5443), .B1_t (new_AGEMA_signal_5444), .B1_f (new_AGEMA_signal_5445), .Z0_t (Inst_bSbox_T6), .Z0_f (new_AGEMA_signal_5608), .Z1_t (new_AGEMA_signal_5609), .Z1_f (new_AGEMA_signal_5610) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T7_U1 ( .A0_t (SboxIn[6]), .A0_f (new_AGEMA_signal_5301), .A1_t (new_AGEMA_signal_5302), .A1_f (new_AGEMA_signal_5303), .B0_t (SboxIn[5]), .B0_f (new_AGEMA_signal_5298), .B1_t (new_AGEMA_signal_5299), .B1_f (new_AGEMA_signal_5300), .Z0_t (Inst_bSbox_T7), .Z0_f (new_AGEMA_signal_5446), .Z1_t (new_AGEMA_signal_5447), .Z1_f (new_AGEMA_signal_5448) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T8_U1 ( .A0_t (SboxIn[0]), .A0_f (new_AGEMA_signal_5283), .A1_t (new_AGEMA_signal_5284), .A1_f (new_AGEMA_signal_5285), .B0_t (Inst_bSbox_T6), .B0_f (new_AGEMA_signal_5608), .B1_t (new_AGEMA_signal_5609), .B1_f (new_AGEMA_signal_5610), .Z0_t (Inst_bSbox_T8), .Z0_f (new_AGEMA_signal_5738), .Z1_t (new_AGEMA_signal_5739), .Z1_f (new_AGEMA_signal_5740) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T9_U1 ( .A0_t (SboxIn[0]), .A0_f (new_AGEMA_signal_5283), .A1_t (new_AGEMA_signal_5284), .A1_f (new_AGEMA_signal_5285), .B0_t (Inst_bSbox_T7), .B0_f (new_AGEMA_signal_5446), .B1_t (new_AGEMA_signal_5447), .B1_f (new_AGEMA_signal_5448), .Z0_t (Inst_bSbox_T9), .Z0_f (new_AGEMA_signal_5611), .Z1_t (new_AGEMA_signal_5612), .Z1_f (new_AGEMA_signal_5613) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T10_U1 ( .A0_t (Inst_bSbox_T6), .A0_f (new_AGEMA_signal_5608), .A1_t (new_AGEMA_signal_5609), .A1_f (new_AGEMA_signal_5610), .B0_t (Inst_bSbox_T7), .B0_f (new_AGEMA_signal_5446), .B1_t (new_AGEMA_signal_5447), .B1_f (new_AGEMA_signal_5448), .Z0_t (Inst_bSbox_T10), .Z0_f (new_AGEMA_signal_5741), .Z1_t (new_AGEMA_signal_5742), .Z1_f (new_AGEMA_signal_5743) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T11_U1 ( .A0_t (SboxIn[6]), .A0_f (new_AGEMA_signal_5301), .A1_t (new_AGEMA_signal_5302), .A1_f (new_AGEMA_signal_5303), .B0_t (SboxIn[2]), .B0_f (new_AGEMA_signal_5289), .B1_t (new_AGEMA_signal_5290), .B1_f (new_AGEMA_signal_5291), .Z0_t (Inst_bSbox_T11), .Z0_f (new_AGEMA_signal_5449), .Z1_t (new_AGEMA_signal_5450), .Z1_f (new_AGEMA_signal_5451) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T12_U1 ( .A0_t (SboxIn[5]), .A0_f (new_AGEMA_signal_5298), .A1_t (new_AGEMA_signal_5299), .A1_f (new_AGEMA_signal_5300), .B0_t (SboxIn[2]), .B0_f (new_AGEMA_signal_5289), .B1_t (new_AGEMA_signal_5290), .B1_f (new_AGEMA_signal_5291), .Z0_t (Inst_bSbox_T12), .Z0_f (new_AGEMA_signal_5452), .Z1_t (new_AGEMA_signal_5453), .Z1_f (new_AGEMA_signal_5454) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T13_U1 ( .A0_t (Inst_bSbox_T3), .A0_f (new_AGEMA_signal_5437), .A1_t (new_AGEMA_signal_5438), .A1_f (new_AGEMA_signal_5439), .B0_t (Inst_bSbox_T4), .B0_f (new_AGEMA_signal_5440), .B1_t (new_AGEMA_signal_5441), .B1_f (new_AGEMA_signal_5442), .Z0_t (Inst_bSbox_T13), .Z0_f (new_AGEMA_signal_5614), .Z1_t (new_AGEMA_signal_5615), .Z1_f (new_AGEMA_signal_5616) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T14_U1 ( .A0_t (Inst_bSbox_T6), .A0_f (new_AGEMA_signal_5608), .A1_t (new_AGEMA_signal_5609), .A1_f (new_AGEMA_signal_5610), .B0_t (Inst_bSbox_T11), .B0_f (new_AGEMA_signal_5449), .B1_t (new_AGEMA_signal_5450), .B1_f (new_AGEMA_signal_5451), .Z0_t (Inst_bSbox_T14), .Z0_f (new_AGEMA_signal_5744), .Z1_t (new_AGEMA_signal_5745), .Z1_f (new_AGEMA_signal_5746) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T15_U1 ( .A0_t (Inst_bSbox_T5), .A0_f (new_AGEMA_signal_5443), .A1_t (new_AGEMA_signal_5444), .A1_f (new_AGEMA_signal_5445), .B0_t (Inst_bSbox_T11), .B0_f (new_AGEMA_signal_5449), .B1_t (new_AGEMA_signal_5450), .B1_f (new_AGEMA_signal_5451), .Z0_t (Inst_bSbox_T15), .Z0_f (new_AGEMA_signal_5617), .Z1_t (new_AGEMA_signal_5618), .Z1_f (new_AGEMA_signal_5619) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T16_U1 ( .A0_t (Inst_bSbox_T5), .A0_f (new_AGEMA_signal_5443), .A1_t (new_AGEMA_signal_5444), .A1_f (new_AGEMA_signal_5445), .B0_t (Inst_bSbox_T12), .B0_f (new_AGEMA_signal_5452), .B1_t (new_AGEMA_signal_5453), .B1_f (new_AGEMA_signal_5454), .Z0_t (Inst_bSbox_T16), .Z0_f (new_AGEMA_signal_5620), .Z1_t (new_AGEMA_signal_5621), .Z1_f (new_AGEMA_signal_5622) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T17_U1 ( .A0_t (Inst_bSbox_T9), .A0_f (new_AGEMA_signal_5611), .A1_t (new_AGEMA_signal_5612), .A1_f (new_AGEMA_signal_5613), .B0_t (Inst_bSbox_T16), .B0_f (new_AGEMA_signal_5620), .B1_t (new_AGEMA_signal_5621), .B1_f (new_AGEMA_signal_5622), .Z0_t (Inst_bSbox_T17), .Z0_f (new_AGEMA_signal_5747), .Z1_t (new_AGEMA_signal_5748), .Z1_f (new_AGEMA_signal_5749) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T18_U1 ( .A0_t (SboxIn[4]), .A0_f (new_AGEMA_signal_5295), .A1_t (new_AGEMA_signal_5296), .A1_f (new_AGEMA_signal_5297), .B0_t (SboxIn[0]), .B0_f (new_AGEMA_signal_5283), .B1_t (new_AGEMA_signal_5284), .B1_f (new_AGEMA_signal_5285), .Z0_t (Inst_bSbox_T18), .Z0_f (new_AGEMA_signal_5455), .Z1_t (new_AGEMA_signal_5456), .Z1_f (new_AGEMA_signal_5457) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T19_U1 ( .A0_t (Inst_bSbox_T7), .A0_f (new_AGEMA_signal_5446), .A1_t (new_AGEMA_signal_5447), .A1_f (new_AGEMA_signal_5448), .B0_t (Inst_bSbox_T18), .B0_f (new_AGEMA_signal_5455), .B1_t (new_AGEMA_signal_5456), .B1_f (new_AGEMA_signal_5457), .Z0_t (Inst_bSbox_T19), .Z0_f (new_AGEMA_signal_5623), .Z1_t (new_AGEMA_signal_5624), .Z1_f (new_AGEMA_signal_5625) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T20_U1 ( .A0_t (Inst_bSbox_T1), .A0_f (new_AGEMA_signal_5431), .A1_t (new_AGEMA_signal_5432), .A1_f (new_AGEMA_signal_5433), .B0_t (Inst_bSbox_T19), .B0_f (new_AGEMA_signal_5623), .B1_t (new_AGEMA_signal_5624), .B1_f (new_AGEMA_signal_5625), .Z0_t (Inst_bSbox_T20), .Z0_f (new_AGEMA_signal_5750), .Z1_t (new_AGEMA_signal_5751), .Z1_f (new_AGEMA_signal_5752) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T21_U1 ( .A0_t (SboxIn[1]), .A0_f (new_AGEMA_signal_5286), .A1_t (new_AGEMA_signal_5287), .A1_f (new_AGEMA_signal_5288), .B0_t (SboxIn[0]), .B0_f (new_AGEMA_signal_5283), .B1_t (new_AGEMA_signal_5284), .B1_f (new_AGEMA_signal_5285), .Z0_t (Inst_bSbox_T21), .Z0_f (new_AGEMA_signal_5458), .Z1_t (new_AGEMA_signal_5459), .Z1_f (new_AGEMA_signal_5460) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T22_U1 ( .A0_t (Inst_bSbox_T7), .A0_f (new_AGEMA_signal_5446), .A1_t (new_AGEMA_signal_5447), .A1_f (new_AGEMA_signal_5448), .B0_t (Inst_bSbox_T21), .B0_f (new_AGEMA_signal_5458), .B1_t (new_AGEMA_signal_5459), .B1_f (new_AGEMA_signal_5460), .Z0_t (Inst_bSbox_T22), .Z0_f (new_AGEMA_signal_5626), .Z1_t (new_AGEMA_signal_5627), .Z1_f (new_AGEMA_signal_5628) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T23_U1 ( .A0_t (Inst_bSbox_T2), .A0_f (new_AGEMA_signal_5434), .A1_t (new_AGEMA_signal_5435), .A1_f (new_AGEMA_signal_5436), .B0_t (Inst_bSbox_T22), .B0_f (new_AGEMA_signal_5626), .B1_t (new_AGEMA_signal_5627), .B1_f (new_AGEMA_signal_5628), .Z0_t (Inst_bSbox_T23), .Z0_f (new_AGEMA_signal_5753), .Z1_t (new_AGEMA_signal_5754), .Z1_f (new_AGEMA_signal_5755) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T24_U1 ( .A0_t (Inst_bSbox_T2), .A0_f (new_AGEMA_signal_5434), .A1_t (new_AGEMA_signal_5435), .A1_f (new_AGEMA_signal_5436), .B0_t (Inst_bSbox_T10), .B0_f (new_AGEMA_signal_5741), .B1_t (new_AGEMA_signal_5742), .B1_f (new_AGEMA_signal_5743), .Z0_t (Inst_bSbox_T24), .Z0_f (new_AGEMA_signal_5889), .Z1_t (new_AGEMA_signal_5890), .Z1_f (new_AGEMA_signal_5891) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T25_U1 ( .A0_t (Inst_bSbox_T20), .A0_f (new_AGEMA_signal_5750), .A1_t (new_AGEMA_signal_5751), .A1_f (new_AGEMA_signal_5752), .B0_t (Inst_bSbox_T17), .B0_f (new_AGEMA_signal_5747), .B1_t (new_AGEMA_signal_5748), .B1_f (new_AGEMA_signal_5749), .Z0_t (Inst_bSbox_T25), .Z0_f (new_AGEMA_signal_5892), .Z1_t (new_AGEMA_signal_5893), .Z1_f (new_AGEMA_signal_5894) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T26_U1 ( .A0_t (Inst_bSbox_T3), .A0_f (new_AGEMA_signal_5437), .A1_t (new_AGEMA_signal_5438), .A1_f (new_AGEMA_signal_5439), .B0_t (Inst_bSbox_T16), .B0_f (new_AGEMA_signal_5620), .B1_t (new_AGEMA_signal_5621), .B1_f (new_AGEMA_signal_5622), .Z0_t (Inst_bSbox_T26), .Z0_f (new_AGEMA_signal_5756), .Z1_t (new_AGEMA_signal_5757), .Z1_f (new_AGEMA_signal_5758) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_T27_U1 ( .A0_t (Inst_bSbox_T1), .A0_f (new_AGEMA_signal_5431), .A1_t (new_AGEMA_signal_5432), .A1_f (new_AGEMA_signal_5433), .B0_t (Inst_bSbox_T12), .B0_f (new_AGEMA_signal_5452), .B1_t (new_AGEMA_signal_5453), .B1_f (new_AGEMA_signal_5454), .Z0_t (Inst_bSbox_T27), .Z0_f (new_AGEMA_signal_5629), .Z1_t (new_AGEMA_signal_5630), .Z1_f (new_AGEMA_signal_5631) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M1_U1 ( .A0_t (Inst_bSbox_T13), .A0_f (new_AGEMA_signal_5614), .A1_t (new_AGEMA_signal_5615), .A1_f (new_AGEMA_signal_5616), .B0_t (Inst_bSbox_T6), .B0_f (new_AGEMA_signal_5608), .B1_t (new_AGEMA_signal_5609), .B1_f (new_AGEMA_signal_5610), .Z0_t (Inst_bSbox_M1), .Z0_f (new_AGEMA_signal_5759), .Z1_t (new_AGEMA_signal_5760), .Z1_f (new_AGEMA_signal_5761) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M2_U1 ( .A0_t (Inst_bSbox_T23), .A0_f (new_AGEMA_signal_5753), .A1_t (new_AGEMA_signal_5754), .A1_f (new_AGEMA_signal_5755), .B0_t (Inst_bSbox_T8), .B0_f (new_AGEMA_signal_5738), .B1_t (new_AGEMA_signal_5739), .B1_f (new_AGEMA_signal_5740), .Z0_t (Inst_bSbox_M2), .Z0_f (new_AGEMA_signal_5895), .Z1_t (new_AGEMA_signal_5896), .Z1_f (new_AGEMA_signal_5897) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M3_U1 ( .A0_t (Inst_bSbox_T14), .A0_f (new_AGEMA_signal_5744), .A1_t (new_AGEMA_signal_5745), .A1_f (new_AGEMA_signal_5746), .B0_t (Inst_bSbox_M1), .B0_f (new_AGEMA_signal_5759), .B1_t (new_AGEMA_signal_5760), .B1_f (new_AGEMA_signal_5761), .Z0_t (Inst_bSbox_M3), .Z0_f (new_AGEMA_signal_5898), .Z1_t (new_AGEMA_signal_5899), .Z1_f (new_AGEMA_signal_5900) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M4_U1 ( .A0_t (Inst_bSbox_T19), .A0_f (new_AGEMA_signal_5623), .A1_t (new_AGEMA_signal_5624), .A1_f (new_AGEMA_signal_5625), .B0_t (SboxIn[0]), .B0_f (new_AGEMA_signal_5283), .B1_t (new_AGEMA_signal_5284), .B1_f (new_AGEMA_signal_5285), .Z0_t (Inst_bSbox_M4), .Z0_f (new_AGEMA_signal_5762), .Z1_t (new_AGEMA_signal_5763), .Z1_f (new_AGEMA_signal_5764) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M5_U1 ( .A0_t (Inst_bSbox_M4), .A0_f (new_AGEMA_signal_5762), .A1_t (new_AGEMA_signal_5763), .A1_f (new_AGEMA_signal_5764), .B0_t (Inst_bSbox_M1), .B0_f (new_AGEMA_signal_5759), .B1_t (new_AGEMA_signal_5760), .B1_f (new_AGEMA_signal_5761), .Z0_t (Inst_bSbox_M5), .Z0_f (new_AGEMA_signal_5901), .Z1_t (new_AGEMA_signal_5902), .Z1_f (new_AGEMA_signal_5903) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M6_U1 ( .A0_t (Inst_bSbox_T3), .A0_f (new_AGEMA_signal_5437), .A1_t (new_AGEMA_signal_5438), .A1_f (new_AGEMA_signal_5439), .B0_t (Inst_bSbox_T16), .B0_f (new_AGEMA_signal_5620), .B1_t (new_AGEMA_signal_5621), .B1_f (new_AGEMA_signal_5622), .Z0_t (Inst_bSbox_M6), .Z0_f (new_AGEMA_signal_5765), .Z1_t (new_AGEMA_signal_5766), .Z1_f (new_AGEMA_signal_5767) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M7_U1 ( .A0_t (Inst_bSbox_T22), .A0_f (new_AGEMA_signal_5626), .A1_t (new_AGEMA_signal_5627), .A1_f (new_AGEMA_signal_5628), .B0_t (Inst_bSbox_T9), .B0_f (new_AGEMA_signal_5611), .B1_t (new_AGEMA_signal_5612), .B1_f (new_AGEMA_signal_5613), .Z0_t (Inst_bSbox_M7), .Z0_f (new_AGEMA_signal_5768), .Z1_t (new_AGEMA_signal_5769), .Z1_f (new_AGEMA_signal_5770) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M8_U1 ( .A0_t (Inst_bSbox_T26), .A0_f (new_AGEMA_signal_5756), .A1_t (new_AGEMA_signal_5757), .A1_f (new_AGEMA_signal_5758), .B0_t (Inst_bSbox_M6), .B0_f (new_AGEMA_signal_5765), .B1_t (new_AGEMA_signal_5766), .B1_f (new_AGEMA_signal_5767), .Z0_t (Inst_bSbox_M8), .Z0_f (new_AGEMA_signal_5904), .Z1_t (new_AGEMA_signal_5905), .Z1_f (new_AGEMA_signal_5906) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M9_U1 ( .A0_t (Inst_bSbox_T20), .A0_f (new_AGEMA_signal_5750), .A1_t (new_AGEMA_signal_5751), .A1_f (new_AGEMA_signal_5752), .B0_t (Inst_bSbox_T17), .B0_f (new_AGEMA_signal_5747), .B1_t (new_AGEMA_signal_5748), .B1_f (new_AGEMA_signal_5749), .Z0_t (Inst_bSbox_M9), .Z0_f (new_AGEMA_signal_5907), .Z1_t (new_AGEMA_signal_5908), .Z1_f (new_AGEMA_signal_5909) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M10_U1 ( .A0_t (Inst_bSbox_M9), .A0_f (new_AGEMA_signal_5907), .A1_t (new_AGEMA_signal_5908), .A1_f (new_AGEMA_signal_5909), .B0_t (Inst_bSbox_M6), .B0_f (new_AGEMA_signal_5765), .B1_t (new_AGEMA_signal_5766), .B1_f (new_AGEMA_signal_5767), .Z0_t (Inst_bSbox_M10), .Z0_f (new_AGEMA_signal_6304), .Z1_t (new_AGEMA_signal_6305), .Z1_f (new_AGEMA_signal_6306) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M11_U1 ( .A0_t (Inst_bSbox_T1), .A0_f (new_AGEMA_signal_5431), .A1_t (new_AGEMA_signal_5432), .A1_f (new_AGEMA_signal_5433), .B0_t (Inst_bSbox_T15), .B0_f (new_AGEMA_signal_5617), .B1_t (new_AGEMA_signal_5618), .B1_f (new_AGEMA_signal_5619), .Z0_t (Inst_bSbox_M11), .Z0_f (new_AGEMA_signal_5771), .Z1_t (new_AGEMA_signal_5772), .Z1_f (new_AGEMA_signal_5773) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M12_U1 ( .A0_t (Inst_bSbox_T4), .A0_f (new_AGEMA_signal_5440), .A1_t (new_AGEMA_signal_5441), .A1_f (new_AGEMA_signal_5442), .B0_t (Inst_bSbox_T27), .B0_f (new_AGEMA_signal_5629), .B1_t (new_AGEMA_signal_5630), .B1_f (new_AGEMA_signal_5631), .Z0_t (Inst_bSbox_M12), .Z0_f (new_AGEMA_signal_5774), .Z1_t (new_AGEMA_signal_5775), .Z1_f (new_AGEMA_signal_5776) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M13_U1 ( .A0_t (Inst_bSbox_M12), .A0_f (new_AGEMA_signal_5774), .A1_t (new_AGEMA_signal_5775), .A1_f (new_AGEMA_signal_5776), .B0_t (Inst_bSbox_M11), .B0_f (new_AGEMA_signal_5771), .B1_t (new_AGEMA_signal_5772), .B1_f (new_AGEMA_signal_5773), .Z0_t (Inst_bSbox_M13), .Z0_f (new_AGEMA_signal_5910), .Z1_t (new_AGEMA_signal_5911), .Z1_f (new_AGEMA_signal_5912) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M14_U1 ( .A0_t (Inst_bSbox_T2), .A0_f (new_AGEMA_signal_5434), .A1_t (new_AGEMA_signal_5435), .A1_f (new_AGEMA_signal_5436), .B0_t (Inst_bSbox_T10), .B0_f (new_AGEMA_signal_5741), .B1_t (new_AGEMA_signal_5742), .B1_f (new_AGEMA_signal_5743), .Z0_t (Inst_bSbox_M14), .Z0_f (new_AGEMA_signal_5913), .Z1_t (new_AGEMA_signal_5914), .Z1_f (new_AGEMA_signal_5915) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M15_U1 ( .A0_t (Inst_bSbox_M14), .A0_f (new_AGEMA_signal_5913), .A1_t (new_AGEMA_signal_5914), .A1_f (new_AGEMA_signal_5915), .B0_t (Inst_bSbox_M11), .B0_f (new_AGEMA_signal_5771), .B1_t (new_AGEMA_signal_5772), .B1_f (new_AGEMA_signal_5773), .Z0_t (Inst_bSbox_M15), .Z0_f (new_AGEMA_signal_6307), .Z1_t (new_AGEMA_signal_6308), .Z1_f (new_AGEMA_signal_6309) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M16_U1 ( .A0_t (Inst_bSbox_M3), .A0_f (new_AGEMA_signal_5898), .A1_t (new_AGEMA_signal_5899), .A1_f (new_AGEMA_signal_5900), .B0_t (Inst_bSbox_M2), .B0_f (new_AGEMA_signal_5895), .B1_t (new_AGEMA_signal_5896), .B1_f (new_AGEMA_signal_5897), .Z0_t (Inst_bSbox_M16), .Z0_f (new_AGEMA_signal_6310), .Z1_t (new_AGEMA_signal_6311), .Z1_f (new_AGEMA_signal_6312) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M17_U1 ( .A0_t (Inst_bSbox_M5), .A0_f (new_AGEMA_signal_5901), .A1_t (new_AGEMA_signal_5902), .A1_f (new_AGEMA_signal_5903), .B0_t (Inst_bSbox_T24), .B0_f (new_AGEMA_signal_5889), .B1_t (new_AGEMA_signal_5890), .B1_f (new_AGEMA_signal_5891), .Z0_t (Inst_bSbox_M17), .Z0_f (new_AGEMA_signal_6313), .Z1_t (new_AGEMA_signal_6314), .Z1_f (new_AGEMA_signal_6315) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M18_U1 ( .A0_t (Inst_bSbox_M8), .A0_f (new_AGEMA_signal_5904), .A1_t (new_AGEMA_signal_5905), .A1_f (new_AGEMA_signal_5906), .B0_t (Inst_bSbox_M7), .B0_f (new_AGEMA_signal_5768), .B1_t (new_AGEMA_signal_5769), .B1_f (new_AGEMA_signal_5770), .Z0_t (Inst_bSbox_M18), .Z0_f (new_AGEMA_signal_6316), .Z1_t (new_AGEMA_signal_6317), .Z1_f (new_AGEMA_signal_6318) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M19_U1 ( .A0_t (Inst_bSbox_M10), .A0_f (new_AGEMA_signal_6304), .A1_t (new_AGEMA_signal_6305), .A1_f (new_AGEMA_signal_6306), .B0_t (Inst_bSbox_M15), .B0_f (new_AGEMA_signal_6307), .B1_t (new_AGEMA_signal_6308), .B1_f (new_AGEMA_signal_6309), .Z0_t (Inst_bSbox_M19), .Z0_f (new_AGEMA_signal_7146), .Z1_t (new_AGEMA_signal_7147), .Z1_f (new_AGEMA_signal_7148) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M20_U1 ( .A0_t (Inst_bSbox_M16), .A0_f (new_AGEMA_signal_6310), .A1_t (new_AGEMA_signal_6311), .A1_f (new_AGEMA_signal_6312), .B0_t (Inst_bSbox_M13), .B0_f (new_AGEMA_signal_5910), .B1_t (new_AGEMA_signal_5911), .B1_f (new_AGEMA_signal_5912), .Z0_t (Inst_bSbox_M20), .Z0_f (new_AGEMA_signal_7149), .Z1_t (new_AGEMA_signal_7150), .Z1_f (new_AGEMA_signal_7151) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M21_U1 ( .A0_t (Inst_bSbox_M17), .A0_f (new_AGEMA_signal_6313), .A1_t (new_AGEMA_signal_6314), .A1_f (new_AGEMA_signal_6315), .B0_t (Inst_bSbox_M15), .B0_f (new_AGEMA_signal_6307), .B1_t (new_AGEMA_signal_6308), .B1_f (new_AGEMA_signal_6309), .Z0_t (Inst_bSbox_M21), .Z0_f (new_AGEMA_signal_7152), .Z1_t (new_AGEMA_signal_7153), .Z1_f (new_AGEMA_signal_7154) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M22_U1 ( .A0_t (Inst_bSbox_M18), .A0_f (new_AGEMA_signal_6316), .A1_t (new_AGEMA_signal_6317), .A1_f (new_AGEMA_signal_6318), .B0_t (Inst_bSbox_M13), .B0_f (new_AGEMA_signal_5910), .B1_t (new_AGEMA_signal_5911), .B1_f (new_AGEMA_signal_5912), .Z0_t (Inst_bSbox_M22), .Z0_f (new_AGEMA_signal_7155), .Z1_t (new_AGEMA_signal_7156), .Z1_f (new_AGEMA_signal_7157) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M23_U1 ( .A0_t (Inst_bSbox_M19), .A0_f (new_AGEMA_signal_7146), .A1_t (new_AGEMA_signal_7147), .A1_f (new_AGEMA_signal_7148), .B0_t (Inst_bSbox_T25), .B0_f (new_AGEMA_signal_5892), .B1_t (new_AGEMA_signal_5893), .B1_f (new_AGEMA_signal_5894), .Z0_t (Inst_bSbox_M23), .Z0_f (new_AGEMA_signal_7262), .Z1_t (new_AGEMA_signal_7263), .Z1_f (new_AGEMA_signal_7264) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M24_U1 ( .A0_t (Inst_bSbox_M22), .A0_f (new_AGEMA_signal_7155), .A1_t (new_AGEMA_signal_7156), .A1_f (new_AGEMA_signal_7157), .B0_t (Inst_bSbox_M23), .B0_f (new_AGEMA_signal_7262), .B1_t (new_AGEMA_signal_7263), .B1_f (new_AGEMA_signal_7264), .Z0_t (Inst_bSbox_M24), .Z0_f (new_AGEMA_signal_7301), .Z1_t (new_AGEMA_signal_7302), .Z1_f (new_AGEMA_signal_7303) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M25_U1 ( .A0_t (Inst_bSbox_M22), .A0_f (new_AGEMA_signal_7155), .A1_t (new_AGEMA_signal_7156), .A1_f (new_AGEMA_signal_7157), .B0_t (Inst_bSbox_M20), .B0_f (new_AGEMA_signal_7149), .B1_t (new_AGEMA_signal_7150), .B1_f (new_AGEMA_signal_7151), .Z0_t (Inst_bSbox_M25), .Z0_f (new_AGEMA_signal_7265), .Z1_t (new_AGEMA_signal_7266), .Z1_f (new_AGEMA_signal_7267) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M26_U1 ( .A0_t (Inst_bSbox_M21), .A0_f (new_AGEMA_signal_7152), .A1_t (new_AGEMA_signal_7153), .A1_f (new_AGEMA_signal_7154), .B0_t (Inst_bSbox_M25), .B0_f (new_AGEMA_signal_7265), .B1_t (new_AGEMA_signal_7266), .B1_f (new_AGEMA_signal_7267), .Z0_t (Inst_bSbox_M26), .Z0_f (new_AGEMA_signal_7304), .Z1_t (new_AGEMA_signal_7305), .Z1_f (new_AGEMA_signal_7306) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M27_U1 ( .A0_t (Inst_bSbox_M20), .A0_f (new_AGEMA_signal_7149), .A1_t (new_AGEMA_signal_7150), .A1_f (new_AGEMA_signal_7151), .B0_t (Inst_bSbox_M21), .B0_f (new_AGEMA_signal_7152), .B1_t (new_AGEMA_signal_7153), .B1_f (new_AGEMA_signal_7154), .Z0_t (Inst_bSbox_M27), .Z0_f (new_AGEMA_signal_7268), .Z1_t (new_AGEMA_signal_7269), .Z1_f (new_AGEMA_signal_7270) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M28_U1 ( .A0_t (Inst_bSbox_M23), .A0_f (new_AGEMA_signal_7262), .A1_t (new_AGEMA_signal_7263), .A1_f (new_AGEMA_signal_7264), .B0_t (Inst_bSbox_M25), .B0_f (new_AGEMA_signal_7265), .B1_t (new_AGEMA_signal_7266), .B1_f (new_AGEMA_signal_7267), .Z0_t (Inst_bSbox_M28), .Z0_f (new_AGEMA_signal_7307), .Z1_t (new_AGEMA_signal_7308), .Z1_f (new_AGEMA_signal_7309) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M29_U1 ( .A0_t (Inst_bSbox_M28), .A0_f (new_AGEMA_signal_7307), .A1_t (new_AGEMA_signal_7308), .A1_f (new_AGEMA_signal_7309), .B0_t (Inst_bSbox_M27), .B0_f (new_AGEMA_signal_7268), .B1_t (new_AGEMA_signal_7269), .B1_f (new_AGEMA_signal_7270), .Z0_t (Inst_bSbox_M29), .Z0_f (new_AGEMA_signal_7316), .Z1_t (new_AGEMA_signal_7317), .Z1_f (new_AGEMA_signal_7318) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M30_U1 ( .A0_t (Inst_bSbox_M26), .A0_f (new_AGEMA_signal_7304), .A1_t (new_AGEMA_signal_7305), .A1_f (new_AGEMA_signal_7306), .B0_t (Inst_bSbox_M24), .B0_f (new_AGEMA_signal_7301), .B1_t (new_AGEMA_signal_7302), .B1_f (new_AGEMA_signal_7303), .Z0_t (Inst_bSbox_M30), .Z0_f (new_AGEMA_signal_7319), .Z1_t (new_AGEMA_signal_7320), .Z1_f (new_AGEMA_signal_7321) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M31_U1 ( .A0_t (Inst_bSbox_M20), .A0_f (new_AGEMA_signal_7149), .A1_t (new_AGEMA_signal_7150), .A1_f (new_AGEMA_signal_7151), .B0_t (Inst_bSbox_M23), .B0_f (new_AGEMA_signal_7262), .B1_t (new_AGEMA_signal_7263), .B1_f (new_AGEMA_signal_7264), .Z0_t (Inst_bSbox_M31), .Z0_f (new_AGEMA_signal_7310), .Z1_t (new_AGEMA_signal_7311), .Z1_f (new_AGEMA_signal_7312) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M32_U1 ( .A0_t (Inst_bSbox_M27), .A0_f (new_AGEMA_signal_7268), .A1_t (new_AGEMA_signal_7269), .A1_f (new_AGEMA_signal_7270), .B0_t (Inst_bSbox_M31), .B0_f (new_AGEMA_signal_7310), .B1_t (new_AGEMA_signal_7311), .B1_f (new_AGEMA_signal_7312), .Z0_t (Inst_bSbox_M32), .Z0_f (new_AGEMA_signal_7322), .Z1_t (new_AGEMA_signal_7323), .Z1_f (new_AGEMA_signal_7324) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M33_U1 ( .A0_t (Inst_bSbox_M27), .A0_f (new_AGEMA_signal_7268), .A1_t (new_AGEMA_signal_7269), .A1_f (new_AGEMA_signal_7270), .B0_t (Inst_bSbox_M25), .B0_f (new_AGEMA_signal_7265), .B1_t (new_AGEMA_signal_7266), .B1_f (new_AGEMA_signal_7267), .Z0_t (Inst_bSbox_M33), .Z0_f (new_AGEMA_signal_7313), .Z1_t (new_AGEMA_signal_7314), .Z1_f (new_AGEMA_signal_7315) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M34_U1 ( .A0_t (Inst_bSbox_M21), .A0_f (new_AGEMA_signal_7152), .A1_t (new_AGEMA_signal_7153), .A1_f (new_AGEMA_signal_7154), .B0_t (Inst_bSbox_M22), .B0_f (new_AGEMA_signal_7155), .B1_t (new_AGEMA_signal_7156), .B1_f (new_AGEMA_signal_7157), .Z0_t (Inst_bSbox_M34), .Z0_f (new_AGEMA_signal_7271), .Z1_t (new_AGEMA_signal_7272), .Z1_f (new_AGEMA_signal_7273) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M35_U1 ( .A0_t (Inst_bSbox_M24), .A0_f (new_AGEMA_signal_7301), .A1_t (new_AGEMA_signal_7302), .A1_f (new_AGEMA_signal_7303), .B0_t (Inst_bSbox_M34), .B0_f (new_AGEMA_signal_7271), .B1_t (new_AGEMA_signal_7272), .B1_f (new_AGEMA_signal_7273), .Z0_t (Inst_bSbox_M35), .Z0_f (new_AGEMA_signal_7325), .Z1_t (new_AGEMA_signal_7326), .Z1_f (new_AGEMA_signal_7327) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M36_U1 ( .A0_t (Inst_bSbox_M24), .A0_f (new_AGEMA_signal_7301), .A1_t (new_AGEMA_signal_7302), .A1_f (new_AGEMA_signal_7303), .B0_t (Inst_bSbox_M25), .B0_f (new_AGEMA_signal_7265), .B1_t (new_AGEMA_signal_7266), .B1_f (new_AGEMA_signal_7267), .Z0_t (Inst_bSbox_M36), .Z0_f (new_AGEMA_signal_7328), .Z1_t (new_AGEMA_signal_7329), .Z1_f (new_AGEMA_signal_7330) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M37_U1 ( .A0_t (Inst_bSbox_M21), .A0_f (new_AGEMA_signal_7152), .A1_t (new_AGEMA_signal_7153), .A1_f (new_AGEMA_signal_7154), .B0_t (Inst_bSbox_M29), .B0_f (new_AGEMA_signal_7316), .B1_t (new_AGEMA_signal_7317), .B1_f (new_AGEMA_signal_7318), .Z0_t (Inst_bSbox_M37), .Z0_f (new_AGEMA_signal_7331), .Z1_t (new_AGEMA_signal_7332), .Z1_f (new_AGEMA_signal_7333) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M38_U1 ( .A0_t (Inst_bSbox_M32), .A0_f (new_AGEMA_signal_7322), .A1_t (new_AGEMA_signal_7323), .A1_f (new_AGEMA_signal_7324), .B0_t (Inst_bSbox_M33), .B0_f (new_AGEMA_signal_7313), .B1_t (new_AGEMA_signal_7314), .B1_f (new_AGEMA_signal_7315), .Z0_t (Inst_bSbox_M38), .Z0_f (new_AGEMA_signal_7334), .Z1_t (new_AGEMA_signal_7335), .Z1_f (new_AGEMA_signal_7336) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M39_U1 ( .A0_t (Inst_bSbox_M23), .A0_f (new_AGEMA_signal_7262), .A1_t (new_AGEMA_signal_7263), .A1_f (new_AGEMA_signal_7264), .B0_t (Inst_bSbox_M30), .B0_f (new_AGEMA_signal_7319), .B1_t (new_AGEMA_signal_7320), .B1_f (new_AGEMA_signal_7321), .Z0_t (Inst_bSbox_M39), .Z0_f (new_AGEMA_signal_7337), .Z1_t (new_AGEMA_signal_7338), .Z1_f (new_AGEMA_signal_7339) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M40_U1 ( .A0_t (Inst_bSbox_M35), .A0_f (new_AGEMA_signal_7325), .A1_t (new_AGEMA_signal_7326), .A1_f (new_AGEMA_signal_7327), .B0_t (Inst_bSbox_M36), .B0_f (new_AGEMA_signal_7328), .B1_t (new_AGEMA_signal_7329), .B1_f (new_AGEMA_signal_7330), .Z0_t (Inst_bSbox_M40), .Z0_f (new_AGEMA_signal_7340), .Z1_t (new_AGEMA_signal_7341), .Z1_f (new_AGEMA_signal_7342) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M41_U1 ( .A0_t (Inst_bSbox_M38), .A0_f (new_AGEMA_signal_7334), .A1_t (new_AGEMA_signal_7335), .A1_f (new_AGEMA_signal_7336), .B0_t (Inst_bSbox_M40), .B0_f (new_AGEMA_signal_7340), .B1_t (new_AGEMA_signal_7341), .B1_f (new_AGEMA_signal_7342), .Z0_t (Inst_bSbox_M41), .Z0_f (new_AGEMA_signal_7343), .Z1_t (new_AGEMA_signal_7344), .Z1_f (new_AGEMA_signal_7345) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M42_U1 ( .A0_t (Inst_bSbox_M37), .A0_f (new_AGEMA_signal_7331), .A1_t (new_AGEMA_signal_7332), .A1_f (new_AGEMA_signal_7333), .B0_t (Inst_bSbox_M39), .B0_f (new_AGEMA_signal_7337), .B1_t (new_AGEMA_signal_7338), .B1_f (new_AGEMA_signal_7339), .Z0_t (Inst_bSbox_M42), .Z0_f (new_AGEMA_signal_7346), .Z1_t (new_AGEMA_signal_7347), .Z1_f (new_AGEMA_signal_7348) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M43_U1 ( .A0_t (Inst_bSbox_M37), .A0_f (new_AGEMA_signal_7331), .A1_t (new_AGEMA_signal_7332), .A1_f (new_AGEMA_signal_7333), .B0_t (Inst_bSbox_M38), .B0_f (new_AGEMA_signal_7334), .B1_t (new_AGEMA_signal_7335), .B1_f (new_AGEMA_signal_7336), .Z0_t (Inst_bSbox_M43), .Z0_f (new_AGEMA_signal_7349), .Z1_t (new_AGEMA_signal_7350), .Z1_f (new_AGEMA_signal_7351) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M44_U1 ( .A0_t (Inst_bSbox_M39), .A0_f (new_AGEMA_signal_7337), .A1_t (new_AGEMA_signal_7338), .A1_f (new_AGEMA_signal_7339), .B0_t (Inst_bSbox_M40), .B0_f (new_AGEMA_signal_7340), .B1_t (new_AGEMA_signal_7341), .B1_f (new_AGEMA_signal_7342), .Z0_t (Inst_bSbox_M44), .Z0_f (new_AGEMA_signal_7352), .Z1_t (new_AGEMA_signal_7353), .Z1_f (new_AGEMA_signal_7354) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_M45_U1 ( .A0_t (Inst_bSbox_M42), .A0_f (new_AGEMA_signal_7346), .A1_t (new_AGEMA_signal_7347), .A1_f (new_AGEMA_signal_7348), .B0_t (Inst_bSbox_M41), .B0_f (new_AGEMA_signal_7343), .B1_t (new_AGEMA_signal_7344), .B1_f (new_AGEMA_signal_7345), .Z0_t (Inst_bSbox_M45), .Z0_f (new_AGEMA_signal_7379), .Z1_t (new_AGEMA_signal_7380), .Z1_f (new_AGEMA_signal_7381) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M46_U1 ( .A0_t (Inst_bSbox_M44), .A0_f (new_AGEMA_signal_7352), .A1_t (new_AGEMA_signal_7353), .A1_f (new_AGEMA_signal_7354), .B0_t (Inst_bSbox_T6), .B0_f (new_AGEMA_signal_5608), .B1_t (new_AGEMA_signal_5609), .B1_f (new_AGEMA_signal_5610), .Z0_t (Inst_bSbox_M46), .Z0_f (new_AGEMA_signal_7382), .Z1_t (new_AGEMA_signal_7383), .Z1_f (new_AGEMA_signal_7384) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M47_U1 ( .A0_t (Inst_bSbox_M40), .A0_f (new_AGEMA_signal_7340), .A1_t (new_AGEMA_signal_7341), .A1_f (new_AGEMA_signal_7342), .B0_t (Inst_bSbox_T8), .B0_f (new_AGEMA_signal_5738), .B1_t (new_AGEMA_signal_5739), .B1_f (new_AGEMA_signal_5740), .Z0_t (Inst_bSbox_M47), .Z0_f (new_AGEMA_signal_7355), .Z1_t (new_AGEMA_signal_7356), .Z1_f (new_AGEMA_signal_7357) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M48_U1 ( .A0_t (Inst_bSbox_M39), .A0_f (new_AGEMA_signal_7337), .A1_t (new_AGEMA_signal_7338), .A1_f (new_AGEMA_signal_7339), .B0_t (SboxIn[0]), .B0_f (new_AGEMA_signal_5283), .B1_t (new_AGEMA_signal_5284), .B1_f (new_AGEMA_signal_5285), .Z0_t (Inst_bSbox_M48), .Z0_f (new_AGEMA_signal_7358), .Z1_t (new_AGEMA_signal_7359), .Z1_f (new_AGEMA_signal_7360) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M49_U1 ( .A0_t (Inst_bSbox_M43), .A0_f (new_AGEMA_signal_7349), .A1_t (new_AGEMA_signal_7350), .A1_f (new_AGEMA_signal_7351), .B0_t (Inst_bSbox_T16), .B0_f (new_AGEMA_signal_5620), .B1_t (new_AGEMA_signal_5621), .B1_f (new_AGEMA_signal_5622), .Z0_t (Inst_bSbox_M49), .Z0_f (new_AGEMA_signal_7385), .Z1_t (new_AGEMA_signal_7386), .Z1_f (new_AGEMA_signal_7387) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M50_U1 ( .A0_t (Inst_bSbox_M38), .A0_f (new_AGEMA_signal_7334), .A1_t (new_AGEMA_signal_7335), .A1_f (new_AGEMA_signal_7336), .B0_t (Inst_bSbox_T9), .B0_f (new_AGEMA_signal_5611), .B1_t (new_AGEMA_signal_5612), .B1_f (new_AGEMA_signal_5613), .Z0_t (Inst_bSbox_M50), .Z0_f (new_AGEMA_signal_7361), .Z1_t (new_AGEMA_signal_7362), .Z1_f (new_AGEMA_signal_7363) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M51_U1 ( .A0_t (Inst_bSbox_M37), .A0_f (new_AGEMA_signal_7331), .A1_t (new_AGEMA_signal_7332), .A1_f (new_AGEMA_signal_7333), .B0_t (Inst_bSbox_T17), .B0_f (new_AGEMA_signal_5747), .B1_t (new_AGEMA_signal_5748), .B1_f (new_AGEMA_signal_5749), .Z0_t (Inst_bSbox_M51), .Z0_f (new_AGEMA_signal_7364), .Z1_t (new_AGEMA_signal_7365), .Z1_f (new_AGEMA_signal_7366) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M52_U1 ( .A0_t (Inst_bSbox_M42), .A0_f (new_AGEMA_signal_7346), .A1_t (new_AGEMA_signal_7347), .A1_f (new_AGEMA_signal_7348), .B0_t (Inst_bSbox_T15), .B0_f (new_AGEMA_signal_5617), .B1_t (new_AGEMA_signal_5618), .B1_f (new_AGEMA_signal_5619), .Z0_t (Inst_bSbox_M52), .Z0_f (new_AGEMA_signal_7388), .Z1_t (new_AGEMA_signal_7389), .Z1_f (new_AGEMA_signal_7390) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M53_U1 ( .A0_t (Inst_bSbox_M45), .A0_f (new_AGEMA_signal_7379), .A1_t (new_AGEMA_signal_7380), .A1_f (new_AGEMA_signal_7381), .B0_t (Inst_bSbox_T27), .B0_f (new_AGEMA_signal_5629), .B1_t (new_AGEMA_signal_5630), .B1_f (new_AGEMA_signal_5631), .Z0_t (Inst_bSbox_M53), .Z0_f (new_AGEMA_signal_7415), .Z1_t (new_AGEMA_signal_7416), .Z1_f (new_AGEMA_signal_7417) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M54_U1 ( .A0_t (Inst_bSbox_M41), .A0_f (new_AGEMA_signal_7343), .A1_t (new_AGEMA_signal_7344), .A1_f (new_AGEMA_signal_7345), .B0_t (Inst_bSbox_T10), .B0_f (new_AGEMA_signal_5741), .B1_t (new_AGEMA_signal_5742), .B1_f (new_AGEMA_signal_5743), .Z0_t (Inst_bSbox_M54), .Z0_f (new_AGEMA_signal_7391), .Z1_t (new_AGEMA_signal_7392), .Z1_f (new_AGEMA_signal_7393) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M55_U1 ( .A0_t (Inst_bSbox_M44), .A0_f (new_AGEMA_signal_7352), .A1_t (new_AGEMA_signal_7353), .A1_f (new_AGEMA_signal_7354), .B0_t (Inst_bSbox_T13), .B0_f (new_AGEMA_signal_5614), .B1_t (new_AGEMA_signal_5615), .B1_f (new_AGEMA_signal_5616), .Z0_t (Inst_bSbox_M55), .Z0_f (new_AGEMA_signal_7394), .Z1_t (new_AGEMA_signal_7395), .Z1_f (new_AGEMA_signal_7396) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M56_U1 ( .A0_t (Inst_bSbox_M40), .A0_f (new_AGEMA_signal_7340), .A1_t (new_AGEMA_signal_7341), .A1_f (new_AGEMA_signal_7342), .B0_t (Inst_bSbox_T23), .B0_f (new_AGEMA_signal_5753), .B1_t (new_AGEMA_signal_5754), .B1_f (new_AGEMA_signal_5755), .Z0_t (Inst_bSbox_M56), .Z0_f (new_AGEMA_signal_7367), .Z1_t (new_AGEMA_signal_7368), .Z1_f (new_AGEMA_signal_7369) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M57_U1 ( .A0_t (Inst_bSbox_M39), .A0_f (new_AGEMA_signal_7337), .A1_t (new_AGEMA_signal_7338), .A1_f (new_AGEMA_signal_7339), .B0_t (Inst_bSbox_T19), .B0_f (new_AGEMA_signal_5623), .B1_t (new_AGEMA_signal_5624), .B1_f (new_AGEMA_signal_5625), .Z0_t (Inst_bSbox_M57), .Z0_f (new_AGEMA_signal_7370), .Z1_t (new_AGEMA_signal_7371), .Z1_f (new_AGEMA_signal_7372) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M58_U1 ( .A0_t (Inst_bSbox_M43), .A0_f (new_AGEMA_signal_7349), .A1_t (new_AGEMA_signal_7350), .A1_f (new_AGEMA_signal_7351), .B0_t (Inst_bSbox_T3), .B0_f (new_AGEMA_signal_5437), .B1_t (new_AGEMA_signal_5438), .B1_f (new_AGEMA_signal_5439), .Z0_t (Inst_bSbox_M58), .Z0_f (new_AGEMA_signal_7397), .Z1_t (new_AGEMA_signal_7398), .Z1_f (new_AGEMA_signal_7399) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M59_U1 ( .A0_t (Inst_bSbox_M38), .A0_f (new_AGEMA_signal_7334), .A1_t (new_AGEMA_signal_7335), .A1_f (new_AGEMA_signal_7336), .B0_t (Inst_bSbox_T22), .B0_f (new_AGEMA_signal_5626), .B1_t (new_AGEMA_signal_5627), .B1_f (new_AGEMA_signal_5628), .Z0_t (Inst_bSbox_M59), .Z0_f (new_AGEMA_signal_7373), .Z1_t (new_AGEMA_signal_7374), .Z1_f (new_AGEMA_signal_7375) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M60_U1 ( .A0_t (Inst_bSbox_M37), .A0_f (new_AGEMA_signal_7331), .A1_t (new_AGEMA_signal_7332), .A1_f (new_AGEMA_signal_7333), .B0_t (Inst_bSbox_T20), .B0_f (new_AGEMA_signal_5750), .B1_t (new_AGEMA_signal_5751), .B1_f (new_AGEMA_signal_5752), .Z0_t (Inst_bSbox_M60), .Z0_f (new_AGEMA_signal_7376), .Z1_t (new_AGEMA_signal_7377), .Z1_f (new_AGEMA_signal_7378) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M61_U1 ( .A0_t (Inst_bSbox_M42), .A0_f (new_AGEMA_signal_7346), .A1_t (new_AGEMA_signal_7347), .A1_f (new_AGEMA_signal_7348), .B0_t (Inst_bSbox_T1), .B0_f (new_AGEMA_signal_5431), .B1_t (new_AGEMA_signal_5432), .B1_f (new_AGEMA_signal_5433), .Z0_t (Inst_bSbox_M61), .Z0_f (new_AGEMA_signal_7400), .Z1_t (new_AGEMA_signal_7401), .Z1_f (new_AGEMA_signal_7402) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M62_U1 ( .A0_t (Inst_bSbox_M45), .A0_f (new_AGEMA_signal_7379), .A1_t (new_AGEMA_signal_7380), .A1_f (new_AGEMA_signal_7381), .B0_t (Inst_bSbox_T4), .B0_f (new_AGEMA_signal_5440), .B1_t (new_AGEMA_signal_5441), .B1_f (new_AGEMA_signal_5442), .Z0_t (Inst_bSbox_M62), .Z0_f (new_AGEMA_signal_7418), .Z1_t (new_AGEMA_signal_7419), .Z1_f (new_AGEMA_signal_7420) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_AND_M63_U1 ( .A0_t (Inst_bSbox_M41), .A0_f (new_AGEMA_signal_7343), .A1_t (new_AGEMA_signal_7344), .A1_f (new_AGEMA_signal_7345), .B0_t (Inst_bSbox_T2), .B0_f (new_AGEMA_signal_5434), .B1_t (new_AGEMA_signal_5435), .B1_f (new_AGEMA_signal_5436), .Z0_t (Inst_bSbox_M63), .Z0_f (new_AGEMA_signal_7403), .Z1_t (new_AGEMA_signal_7404), .Z1_f (new_AGEMA_signal_7405) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L0_U1 ( .A0_t (Inst_bSbox_M61), .A0_f (new_AGEMA_signal_7400), .A1_t (new_AGEMA_signal_7401), .A1_f (new_AGEMA_signal_7402), .B0_t (Inst_bSbox_M62), .B0_f (new_AGEMA_signal_7418), .B1_t (new_AGEMA_signal_7419), .B1_f (new_AGEMA_signal_7420), .Z0_t (Inst_bSbox_L0), .Z0_f (new_AGEMA_signal_7445), .Z1_t (new_AGEMA_signal_7446), .Z1_f (new_AGEMA_signal_7447) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L1_U1 ( .A0_t (Inst_bSbox_M50), .A0_f (new_AGEMA_signal_7361), .A1_t (new_AGEMA_signal_7362), .A1_f (new_AGEMA_signal_7363), .B0_t (Inst_bSbox_M56), .B0_f (new_AGEMA_signal_7367), .B1_t (new_AGEMA_signal_7368), .B1_f (new_AGEMA_signal_7369), .Z0_t (Inst_bSbox_L1), .Z0_f (new_AGEMA_signal_7406), .Z1_t (new_AGEMA_signal_7407), .Z1_f (new_AGEMA_signal_7408) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L2_U1 ( .A0_t (Inst_bSbox_M46), .A0_f (new_AGEMA_signal_7382), .A1_t (new_AGEMA_signal_7383), .A1_f (new_AGEMA_signal_7384), .B0_t (Inst_bSbox_M48), .B0_f (new_AGEMA_signal_7358), .B1_t (new_AGEMA_signal_7359), .B1_f (new_AGEMA_signal_7360), .Z0_t (Inst_bSbox_L2), .Z0_f (new_AGEMA_signal_7421), .Z1_t (new_AGEMA_signal_7422), .Z1_f (new_AGEMA_signal_7423) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L3_U1 ( .A0_t (Inst_bSbox_M47), .A0_f (new_AGEMA_signal_7355), .A1_t (new_AGEMA_signal_7356), .A1_f (new_AGEMA_signal_7357), .B0_t (Inst_bSbox_M55), .B0_f (new_AGEMA_signal_7394), .B1_t (new_AGEMA_signal_7395), .B1_f (new_AGEMA_signal_7396), .Z0_t (Inst_bSbox_L3), .Z0_f (new_AGEMA_signal_7424), .Z1_t (new_AGEMA_signal_7425), .Z1_f (new_AGEMA_signal_7426) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L4_U1 ( .A0_t (Inst_bSbox_M54), .A0_f (new_AGEMA_signal_7391), .A1_t (new_AGEMA_signal_7392), .A1_f (new_AGEMA_signal_7393), .B0_t (Inst_bSbox_M58), .B0_f (new_AGEMA_signal_7397), .B1_t (new_AGEMA_signal_7398), .B1_f (new_AGEMA_signal_7399), .Z0_t (Inst_bSbox_L4), .Z0_f (new_AGEMA_signal_7427), .Z1_t (new_AGEMA_signal_7428), .Z1_f (new_AGEMA_signal_7429) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L5_U1 ( .A0_t (Inst_bSbox_M49), .A0_f (new_AGEMA_signal_7385), .A1_t (new_AGEMA_signal_7386), .A1_f (new_AGEMA_signal_7387), .B0_t (Inst_bSbox_M61), .B0_f (new_AGEMA_signal_7400), .B1_t (new_AGEMA_signal_7401), .B1_f (new_AGEMA_signal_7402), .Z0_t (Inst_bSbox_L5), .Z0_f (new_AGEMA_signal_7430), .Z1_t (new_AGEMA_signal_7431), .Z1_f (new_AGEMA_signal_7432) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L6_U1 ( .A0_t (Inst_bSbox_M62), .A0_f (new_AGEMA_signal_7418), .A1_t (new_AGEMA_signal_7419), .A1_f (new_AGEMA_signal_7420), .B0_t (Inst_bSbox_L5), .B0_f (new_AGEMA_signal_7430), .B1_t (new_AGEMA_signal_7431), .B1_f (new_AGEMA_signal_7432), .Z0_t (Inst_bSbox_L6), .Z0_f (new_AGEMA_signal_7448), .Z1_t (new_AGEMA_signal_7449), .Z1_f (new_AGEMA_signal_7450) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L7_U1 ( .A0_t (Inst_bSbox_M46), .A0_f (new_AGEMA_signal_7382), .A1_t (new_AGEMA_signal_7383), .A1_f (new_AGEMA_signal_7384), .B0_t (Inst_bSbox_L3), .B0_f (new_AGEMA_signal_7424), .B1_t (new_AGEMA_signal_7425), .B1_f (new_AGEMA_signal_7426), .Z0_t (Inst_bSbox_L7), .Z0_f (new_AGEMA_signal_7451), .Z1_t (new_AGEMA_signal_7452), .Z1_f (new_AGEMA_signal_7453) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L8_U1 ( .A0_t (Inst_bSbox_M51), .A0_f (new_AGEMA_signal_7364), .A1_t (new_AGEMA_signal_7365), .A1_f (new_AGEMA_signal_7366), .B0_t (Inst_bSbox_M59), .B0_f (new_AGEMA_signal_7373), .B1_t (new_AGEMA_signal_7374), .B1_f (new_AGEMA_signal_7375), .Z0_t (Inst_bSbox_L8), .Z0_f (new_AGEMA_signal_7409), .Z1_t (new_AGEMA_signal_7410), .Z1_f (new_AGEMA_signal_7411) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L9_U1 ( .A0_t (Inst_bSbox_M52), .A0_f (new_AGEMA_signal_7388), .A1_t (new_AGEMA_signal_7389), .A1_f (new_AGEMA_signal_7390), .B0_t (Inst_bSbox_M53), .B0_f (new_AGEMA_signal_7415), .B1_t (new_AGEMA_signal_7416), .B1_f (new_AGEMA_signal_7417), .Z0_t (Inst_bSbox_L9), .Z0_f (new_AGEMA_signal_7454), .Z1_t (new_AGEMA_signal_7455), .Z1_f (new_AGEMA_signal_7456) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L10_U1 ( .A0_t (Inst_bSbox_M53), .A0_f (new_AGEMA_signal_7415), .A1_t (new_AGEMA_signal_7416), .A1_f (new_AGEMA_signal_7417), .B0_t (Inst_bSbox_L4), .B0_f (new_AGEMA_signal_7427), .B1_t (new_AGEMA_signal_7428), .B1_f (new_AGEMA_signal_7429), .Z0_t (Inst_bSbox_L10), .Z0_f (new_AGEMA_signal_7457), .Z1_t (new_AGEMA_signal_7458), .Z1_f (new_AGEMA_signal_7459) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L11_U1 ( .A0_t (Inst_bSbox_M60), .A0_f (new_AGEMA_signal_7376), .A1_t (new_AGEMA_signal_7377), .A1_f (new_AGEMA_signal_7378), .B0_t (Inst_bSbox_L2), .B0_f (new_AGEMA_signal_7421), .B1_t (new_AGEMA_signal_7422), .B1_f (new_AGEMA_signal_7423), .Z0_t (Inst_bSbox_L11), .Z0_f (new_AGEMA_signal_7460), .Z1_t (new_AGEMA_signal_7461), .Z1_f (new_AGEMA_signal_7462) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L12_U1 ( .A0_t (Inst_bSbox_M48), .A0_f (new_AGEMA_signal_7358), .A1_t (new_AGEMA_signal_7359), .A1_f (new_AGEMA_signal_7360), .B0_t (Inst_bSbox_M51), .B0_f (new_AGEMA_signal_7364), .B1_t (new_AGEMA_signal_7365), .B1_f (new_AGEMA_signal_7366), .Z0_t (Inst_bSbox_L12), .Z0_f (new_AGEMA_signal_7412), .Z1_t (new_AGEMA_signal_7413), .Z1_f (new_AGEMA_signal_7414) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L13_U1 ( .A0_t (Inst_bSbox_M50), .A0_f (new_AGEMA_signal_7361), .A1_t (new_AGEMA_signal_7362), .A1_f (new_AGEMA_signal_7363), .B0_t (Inst_bSbox_L0), .B0_f (new_AGEMA_signal_7445), .B1_t (new_AGEMA_signal_7446), .B1_f (new_AGEMA_signal_7447), .Z0_t (Inst_bSbox_L13), .Z0_f (new_AGEMA_signal_7472), .Z1_t (new_AGEMA_signal_7473), .Z1_f (new_AGEMA_signal_7474) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L14_U1 ( .A0_t (Inst_bSbox_M52), .A0_f (new_AGEMA_signal_7388), .A1_t (new_AGEMA_signal_7389), .A1_f (new_AGEMA_signal_7390), .B0_t (Inst_bSbox_M61), .B0_f (new_AGEMA_signal_7400), .B1_t (new_AGEMA_signal_7401), .B1_f (new_AGEMA_signal_7402), .Z0_t (Inst_bSbox_L14), .Z0_f (new_AGEMA_signal_7433), .Z1_t (new_AGEMA_signal_7434), .Z1_f (new_AGEMA_signal_7435) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L15_U1 ( .A0_t (Inst_bSbox_M55), .A0_f (new_AGEMA_signal_7394), .A1_t (new_AGEMA_signal_7395), .A1_f (new_AGEMA_signal_7396), .B0_t (Inst_bSbox_L1), .B0_f (new_AGEMA_signal_7406), .B1_t (new_AGEMA_signal_7407), .B1_f (new_AGEMA_signal_7408), .Z0_t (Inst_bSbox_L15), .Z0_f (new_AGEMA_signal_7436), .Z1_t (new_AGEMA_signal_7437), .Z1_f (new_AGEMA_signal_7438) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L16_U1 ( .A0_t (Inst_bSbox_M56), .A0_f (new_AGEMA_signal_7367), .A1_t (new_AGEMA_signal_7368), .A1_f (new_AGEMA_signal_7369), .B0_t (Inst_bSbox_L0), .B0_f (new_AGEMA_signal_7445), .B1_t (new_AGEMA_signal_7446), .B1_f (new_AGEMA_signal_7447), .Z0_t (Inst_bSbox_L16), .Z0_f (new_AGEMA_signal_7475), .Z1_t (new_AGEMA_signal_7476), .Z1_f (new_AGEMA_signal_7477) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L17_U1 ( .A0_t (Inst_bSbox_M57), .A0_f (new_AGEMA_signal_7370), .A1_t (new_AGEMA_signal_7371), .A1_f (new_AGEMA_signal_7372), .B0_t (Inst_bSbox_L1), .B0_f (new_AGEMA_signal_7406), .B1_t (new_AGEMA_signal_7407), .B1_f (new_AGEMA_signal_7408), .Z0_t (Inst_bSbox_L17), .Z0_f (new_AGEMA_signal_7439), .Z1_t (new_AGEMA_signal_7440), .Z1_f (new_AGEMA_signal_7441) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L18_U1 ( .A0_t (Inst_bSbox_M58), .A0_f (new_AGEMA_signal_7397), .A1_t (new_AGEMA_signal_7398), .A1_f (new_AGEMA_signal_7399), .B0_t (Inst_bSbox_L8), .B0_f (new_AGEMA_signal_7409), .B1_t (new_AGEMA_signal_7410), .B1_f (new_AGEMA_signal_7411), .Z0_t (Inst_bSbox_L18), .Z0_f (new_AGEMA_signal_7442), .Z1_t (new_AGEMA_signal_7443), .Z1_f (new_AGEMA_signal_7444) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L19_U1 ( .A0_t (Inst_bSbox_M63), .A0_f (new_AGEMA_signal_7403), .A1_t (new_AGEMA_signal_7404), .A1_f (new_AGEMA_signal_7405), .B0_t (Inst_bSbox_L4), .B0_f (new_AGEMA_signal_7427), .B1_t (new_AGEMA_signal_7428), .B1_f (new_AGEMA_signal_7429), .Z0_t (Inst_bSbox_L19), .Z0_f (new_AGEMA_signal_7463), .Z1_t (new_AGEMA_signal_7464), .Z1_f (new_AGEMA_signal_7465) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L20_U1 ( .A0_t (Inst_bSbox_L0), .A0_f (new_AGEMA_signal_7445), .A1_t (new_AGEMA_signal_7446), .A1_f (new_AGEMA_signal_7447), .B0_t (Inst_bSbox_L1), .B0_f (new_AGEMA_signal_7406), .B1_t (new_AGEMA_signal_7407), .B1_f (new_AGEMA_signal_7408), .Z0_t (Inst_bSbox_L20), .Z0_f (new_AGEMA_signal_7478), .Z1_t (new_AGEMA_signal_7479), .Z1_f (new_AGEMA_signal_7480) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L21_U1 ( .A0_t (Inst_bSbox_L1), .A0_f (new_AGEMA_signal_7406), .A1_t (new_AGEMA_signal_7407), .A1_f (new_AGEMA_signal_7408), .B0_t (Inst_bSbox_L7), .B0_f (new_AGEMA_signal_7451), .B1_t (new_AGEMA_signal_7452), .B1_f (new_AGEMA_signal_7453), .Z0_t (Inst_bSbox_L21), .Z0_f (new_AGEMA_signal_7481), .Z1_t (new_AGEMA_signal_7482), .Z1_f (new_AGEMA_signal_7483) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L22_U1 ( .A0_t (Inst_bSbox_L3), .A0_f (new_AGEMA_signal_7424), .A1_t (new_AGEMA_signal_7425), .A1_f (new_AGEMA_signal_7426), .B0_t (Inst_bSbox_L12), .B0_f (new_AGEMA_signal_7412), .B1_t (new_AGEMA_signal_7413), .B1_f (new_AGEMA_signal_7414), .Z0_t (Inst_bSbox_L22), .Z0_f (new_AGEMA_signal_7466), .Z1_t (new_AGEMA_signal_7467), .Z1_f (new_AGEMA_signal_7468) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L23_U1 ( .A0_t (Inst_bSbox_L18), .A0_f (new_AGEMA_signal_7442), .A1_t (new_AGEMA_signal_7443), .A1_f (new_AGEMA_signal_7444), .B0_t (Inst_bSbox_L2), .B0_f (new_AGEMA_signal_7421), .B1_t (new_AGEMA_signal_7422), .B1_f (new_AGEMA_signal_7423), .Z0_t (Inst_bSbox_L23), .Z0_f (new_AGEMA_signal_7469), .Z1_t (new_AGEMA_signal_7470), .Z1_f (new_AGEMA_signal_7471) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L24_U1 ( .A0_t (Inst_bSbox_L15), .A0_f (new_AGEMA_signal_7436), .A1_t (new_AGEMA_signal_7437), .A1_f (new_AGEMA_signal_7438), .B0_t (Inst_bSbox_L9), .B0_f (new_AGEMA_signal_7454), .B1_t (new_AGEMA_signal_7455), .B1_f (new_AGEMA_signal_7456), .Z0_t (Inst_bSbox_L24), .Z0_f (new_AGEMA_signal_7484), .Z1_t (new_AGEMA_signal_7485), .Z1_f (new_AGEMA_signal_7486) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L25_U1 ( .A0_t (Inst_bSbox_L6), .A0_f (new_AGEMA_signal_7448), .A1_t (new_AGEMA_signal_7449), .A1_f (new_AGEMA_signal_7450), .B0_t (Inst_bSbox_L10), .B0_f (new_AGEMA_signal_7457), .B1_t (new_AGEMA_signal_7458), .B1_f (new_AGEMA_signal_7459), .Z0_t (Inst_bSbox_L25), .Z0_f (new_AGEMA_signal_7487), .Z1_t (new_AGEMA_signal_7488), .Z1_f (new_AGEMA_signal_7489) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L26_U1 ( .A0_t (Inst_bSbox_L7), .A0_f (new_AGEMA_signal_7451), .A1_t (new_AGEMA_signal_7452), .A1_f (new_AGEMA_signal_7453), .B0_t (Inst_bSbox_L9), .B0_f (new_AGEMA_signal_7454), .B1_t (new_AGEMA_signal_7455), .B1_f (new_AGEMA_signal_7456), .Z0_t (Inst_bSbox_L26), .Z0_f (new_AGEMA_signal_7490), .Z1_t (new_AGEMA_signal_7491), .Z1_f (new_AGEMA_signal_7492) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L27_U1 ( .A0_t (Inst_bSbox_L8), .A0_f (new_AGEMA_signal_7409), .A1_t (new_AGEMA_signal_7410), .A1_f (new_AGEMA_signal_7411), .B0_t (Inst_bSbox_L10), .B0_f (new_AGEMA_signal_7457), .B1_t (new_AGEMA_signal_7458), .B1_f (new_AGEMA_signal_7459), .Z0_t (Inst_bSbox_L27), .Z0_f (new_AGEMA_signal_7493), .Z1_t (new_AGEMA_signal_7494), .Z1_f (new_AGEMA_signal_7495) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L28_U1 ( .A0_t (Inst_bSbox_L11), .A0_f (new_AGEMA_signal_7460), .A1_t (new_AGEMA_signal_7461), .A1_f (new_AGEMA_signal_7462), .B0_t (Inst_bSbox_L14), .B0_f (new_AGEMA_signal_7433), .B1_t (new_AGEMA_signal_7434), .B1_f (new_AGEMA_signal_7435), .Z0_t (Inst_bSbox_L28), .Z0_f (new_AGEMA_signal_7496), .Z1_t (new_AGEMA_signal_7497), .Z1_f (new_AGEMA_signal_7498) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_L29_U1 ( .A0_t (Inst_bSbox_L11), .A0_f (new_AGEMA_signal_7460), .A1_t (new_AGEMA_signal_7461), .A1_f (new_AGEMA_signal_7462), .B0_t (Inst_bSbox_L17), .B0_f (new_AGEMA_signal_7439), .B1_t (new_AGEMA_signal_7440), .B1_f (new_AGEMA_signal_7441), .Z0_t (Inst_bSbox_L29), .Z0_f (new_AGEMA_signal_7499), .Z1_t (new_AGEMA_signal_7500), .Z1_f (new_AGEMA_signal_7501) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_S0_U1 ( .A0_t (Inst_bSbox_L6), .A0_f (new_AGEMA_signal_7448), .A1_t (new_AGEMA_signal_7449), .A1_f (new_AGEMA_signal_7450), .B0_t (Inst_bSbox_L24), .B0_f (new_AGEMA_signal_7484), .B1_t (new_AGEMA_signal_7485), .B1_f (new_AGEMA_signal_7486), .Z0_t (SboxOut[7]), .Z0_f (new_AGEMA_signal_7511), .Z1_t (new_AGEMA_signal_7512), .Z1_f (new_AGEMA_signal_7513) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Inst_bSbox_XOR_S1_U1 ( .A0_t (Inst_bSbox_L16), .A0_f (new_AGEMA_signal_7475), .A1_t (new_AGEMA_signal_7476), .A1_f (new_AGEMA_signal_7477), .B0_t (Inst_bSbox_L26), .B0_f (new_AGEMA_signal_7490), .B1_t (new_AGEMA_signal_7491), .B1_f (new_AGEMA_signal_7492), .Z0_t (SboxOut[6]), .Z0_f (new_AGEMA_signal_7514), .Z1_t (new_AGEMA_signal_7515), .Z1_f (new_AGEMA_signal_7516) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Inst_bSbox_XOR_S2_U1 ( .A0_t (Inst_bSbox_L19), .A0_f (new_AGEMA_signal_7463), .A1_t (new_AGEMA_signal_7464), .A1_f (new_AGEMA_signal_7465), .B0_t (Inst_bSbox_L28), .B0_f (new_AGEMA_signal_7496), .B1_t (new_AGEMA_signal_7497), .B1_f (new_AGEMA_signal_7498), .Z0_t (SboxOut[5]), .Z0_f (new_AGEMA_signal_7517), .Z1_t (new_AGEMA_signal_7518), .Z1_f (new_AGEMA_signal_7519) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_S3_U1 ( .A0_t (Inst_bSbox_L6), .A0_f (new_AGEMA_signal_7448), .A1_t (new_AGEMA_signal_7449), .A1_f (new_AGEMA_signal_7450), .B0_t (Inst_bSbox_L21), .B0_f (new_AGEMA_signal_7481), .B1_t (new_AGEMA_signal_7482), .B1_f (new_AGEMA_signal_7483), .Z0_t (SboxOut[4]), .Z0_f (new_AGEMA_signal_7520), .Z1_t (new_AGEMA_signal_7521), .Z1_f (new_AGEMA_signal_7522) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_S4_U1 ( .A0_t (Inst_bSbox_L20), .A0_f (new_AGEMA_signal_7478), .A1_t (new_AGEMA_signal_7479), .A1_f (new_AGEMA_signal_7480), .B0_t (Inst_bSbox_L22), .B0_f (new_AGEMA_signal_7466), .B1_t (new_AGEMA_signal_7467), .B1_f (new_AGEMA_signal_7468), .Z0_t (SboxOut[3]), .Z0_f (new_AGEMA_signal_7523), .Z1_t (new_AGEMA_signal_7524), .Z1_f (new_AGEMA_signal_7525) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Inst_bSbox_XOR_S5_U1 ( .A0_t (Inst_bSbox_L25), .A0_f (new_AGEMA_signal_7487), .A1_t (new_AGEMA_signal_7488), .A1_f (new_AGEMA_signal_7489), .B0_t (Inst_bSbox_L29), .B0_f (new_AGEMA_signal_7499), .B1_t (new_AGEMA_signal_7500), .B1_f (new_AGEMA_signal_7501), .Z0_t (SboxOut[2]), .Z0_f (new_AGEMA_signal_7526), .Z1_t (new_AGEMA_signal_7527), .Z1_f (new_AGEMA_signal_7528) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Inst_bSbox_XOR_S6_U1 ( .A0_t (Inst_bSbox_L13), .A0_f (new_AGEMA_signal_7472), .A1_t (new_AGEMA_signal_7473), .A1_f (new_AGEMA_signal_7474), .B0_t (Inst_bSbox_L27), .B0_f (new_AGEMA_signal_7493), .B1_t (new_AGEMA_signal_7494), .B1_f (new_AGEMA_signal_7495), .Z0_t (SboxOut[1]), .Z0_f (new_AGEMA_signal_7529), .Z1_t (new_AGEMA_signal_7530), .Z1_f (new_AGEMA_signal_7531) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Inst_bSbox_XOR_S7_U1 ( .A0_t (Inst_bSbox_L6), .A0_f (new_AGEMA_signal_7448), .A1_t (new_AGEMA_signal_7449), .A1_f (new_AGEMA_signal_7450), .B0_t (Inst_bSbox_L23), .B0_f (new_AGEMA_signal_7469), .B1_t (new_AGEMA_signal_7470), .B1_f (new_AGEMA_signal_7471), .Z0_t (SboxOut[0]), .Z0_f (new_AGEMA_signal_7502), .Z1_t (new_AGEMA_signal_7503), .Z1_f (new_AGEMA_signal_7504) ) ;

    /* register cells */
endmodule
