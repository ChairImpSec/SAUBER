/* modified netlist. Source: module LED in file /mnt/c/Users/amirm/Desktop/Papers_in_progress/SAUBER/Design for our FPGA/12-LED_round_based_encryption_PortParallel/4-AGEMA/LED.v */
/* 0 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 1 register stage(s) in total */

module LED_SAUBER_Pipeline_d1 (IN_plaintext_s0_t, IN_key_s0_t, IN_reset_t, IN_reset_f, IN_key_s0_f, IN_key_s1_t, IN_key_s1_f, IN_plaintext_s0_f, IN_plaintext_s1_t, IN_plaintext_s1_f, OUT_ciphertext_s0_t, OUT_done_t, OUT_done_f, OUT_ciphertext_s0_f, OUT_ciphertext_s1_t, OUT_ciphertext_s1_f);
    input [63:0] IN_plaintext_s0_t ;
    input [127:0] IN_key_s0_t ;
    input IN_reset_t ;
    input IN_reset_f ;
    input [127:0] IN_key_s0_f ;
    input [127:0] IN_key_s1_t ;
    input [127:0] IN_key_s1_f ;
    input [63:0] IN_plaintext_s0_f ;
    input [63:0] IN_plaintext_s1_t ;
    input [63:0] IN_plaintext_s1_f ;
    output [63:0] OUT_ciphertext_s0_t ;
    output OUT_done_t ;
    output OUT_done_f ;
    output [63:0] OUT_ciphertext_s0_f ;
    output [63:0] OUT_ciphertext_s1_t ;
    output [63:0] OUT_ciphertext_s1_f ;
    wire n15 ;
    wire n16 ;
    wire n17 ;
    wire n18 ;
    wire n19 ;
    wire n20 ;
    wire LED_128_Instance_n29 ;
    wire LED_128_Instance_n19 ;
    wire LED_128_Instance_n18 ;
    wire LED_128_Instance_n17 ;
    wire LED_128_Instance_n16 ;
    wire LED_128_Instance_n13 ;
    wire LED_128_Instance_n12 ;
    wire LED_128_Instance_n11 ;
    wire LED_128_Instance_n9 ;
    wire LED_128_Instance_n8 ;
    wire LED_128_Instance_n31 ;
    wire LED_128_Instance_n24 ;
    wire LED_128_Instance_ks_0 ;
    wire LED_128_Instance_ks_3_ ;
    wire LED_128_Instance_n23 ;
    wire LED_128_Instance_n22 ;
    wire LED_128_Instance_MUX_state0_mux_inst_0_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_0_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_1_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_1_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_2_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_2_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_3_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_3_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_4_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_4_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_5_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_5_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_6_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_6_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_7_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_7_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_8_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_8_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_9_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_9_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_10_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_10_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_11_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_11_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_12_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_12_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_13_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_13_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_14_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_14_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_15_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_15_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_16_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_16_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_17_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_17_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_18_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_18_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_19_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_19_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_20_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_20_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_21_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_21_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_22_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_22_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_23_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_23_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_24_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_24_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_25_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_25_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_26_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_26_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_27_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_27_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_28_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_28_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_29_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_29_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_30_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_30_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_31_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_31_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_32_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_32_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_33_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_33_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_34_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_34_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_35_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_35_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_36_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_36_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_37_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_37_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_38_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_38_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_39_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_39_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_40_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_40_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_41_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_41_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_42_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_42_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_43_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_43_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_44_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_44_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_45_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_45_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_46_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_46_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_47_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_47_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_48_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_48_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_49_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_49_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_50_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_50_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_51_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_51_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_52_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_52_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_53_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_53_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_54_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_54_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_55_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_55_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_56_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_56_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_57_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_57_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_58_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_58_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_59_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_59_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_60_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_60_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_61_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_61_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_62_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_62_U1_X ;
    wire LED_128_Instance_MUX_state0_mux_inst_63_U1_Y ;
    wire LED_128_Instance_MUX_state0_mux_inst_63_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_0_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_0_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_1_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_1_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_2_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_2_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_3_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_3_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_4_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_4_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_5_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_5_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_6_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_6_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_7_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_7_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_8_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_8_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_9_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_9_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_10_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_10_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_11_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_11_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_12_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_12_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_13_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_13_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_14_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_14_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_15_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_15_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_16_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_16_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_17_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_17_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_18_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_18_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_19_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_19_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_20_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_20_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_21_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_21_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_22_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_22_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_23_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_23_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_24_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_24_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_25_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_25_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_26_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_26_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_27_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_27_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_28_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_28_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_29_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_29_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_30_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_30_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_31_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_31_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_32_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_32_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_33_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_33_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_34_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_34_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_35_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_35_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_36_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_36_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_37_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_37_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_38_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_38_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_39_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_39_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_40_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_40_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_41_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_41_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_42_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_42_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_43_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_43_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_44_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_44_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_45_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_45_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_46_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_46_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_47_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_47_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_48_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_48_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_49_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_49_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_50_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_50_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_51_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_51_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_52_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_52_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_53_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_53_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_54_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_54_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_55_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_55_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_56_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_56_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_57_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_57_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_58_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_58_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_59_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_59_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_60_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_60_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_61_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_61_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_62_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_62_U1_X ;
    wire LED_128_Instance_MUX_state1_mux_inst_63_U1_Y ;
    wire LED_128_Instance_MUX_state1_mux_inst_63_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_0_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_0_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_1_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_1_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_2_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_2_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_3_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_3_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_4_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_4_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_5_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_5_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_6_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_6_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_7_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_7_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_8_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_8_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_9_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_9_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_10_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_10_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_11_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_11_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_12_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_12_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_13_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_13_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_14_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_14_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_15_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_15_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_16_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_16_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_17_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_17_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_18_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_18_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_19_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_19_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_20_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_20_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_21_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_21_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_22_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_22_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_23_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_23_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_24_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_24_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_25_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_25_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_26_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_26_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_27_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_27_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_28_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_28_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_29_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_29_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_30_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_30_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_31_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_31_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_32_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_32_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_33_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_33_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_34_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_34_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_35_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_35_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_36_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_36_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_37_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_37_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_38_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_38_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_39_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_39_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_40_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_40_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_41_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_41_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_42_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_42_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_43_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_43_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_44_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_44_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_45_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_45_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_46_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_46_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_47_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_47_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_48_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_48_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_49_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_49_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_50_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_50_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_51_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_51_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_52_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_52_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_53_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_53_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_54_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_54_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_55_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_55_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_56_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_56_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_57_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_57_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_58_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_58_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_59_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_59_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_60_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_60_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_61_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_61_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_62_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_62_U1_X ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_63_U1_Y ;
    wire LED_128_Instance_MUX_current_roundkey_mux_inst_63_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_0_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_0_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_1_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_1_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_2_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_2_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_3_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_3_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_4_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_4_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_5_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_5_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_6_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_6_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_7_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_7_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_8_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_8_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_9_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_9_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_10_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_10_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_11_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_11_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_12_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_12_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_13_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_13_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_14_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_14_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_15_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_15_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_16_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_16_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_17_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_17_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_18_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_18_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_19_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_19_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_20_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_20_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_21_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_21_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_22_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_22_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_23_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_23_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_24_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_24_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_25_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_25_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_26_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_26_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_27_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_27_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_28_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_28_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_29_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_29_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_30_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_30_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_31_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_31_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_32_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_32_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_33_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_33_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_34_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_34_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_35_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_35_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_36_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_36_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_37_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_37_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_38_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_38_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_39_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_39_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_40_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_40_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_41_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_41_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_42_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_42_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_43_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_43_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_44_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_44_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_45_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_45_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_46_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_46_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_47_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_47_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_48_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_48_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_49_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_49_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_50_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_50_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_51_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_51_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_52_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_52_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_53_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_53_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_54_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_54_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_55_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_55_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_56_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_56_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_57_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_57_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_58_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_58_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_59_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_59_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_60_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_60_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_61_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_61_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_62_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_62_U1_X ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_63_U1_Y ;
    wire LED_128_Instance_MUX_addroundkey_out_mux_inst_63_U1_X ;
    wire LED_128_Instance_SBox_Instance_0_L8 ;
    wire LED_128_Instance_SBox_Instance_0_L7 ;
    wire LED_128_Instance_SBox_Instance_0_T3 ;
    wire LED_128_Instance_SBox_Instance_0_T1 ;
    wire LED_128_Instance_SBox_Instance_0_Q7 ;
    wire LED_128_Instance_SBox_Instance_0_Q6 ;
    wire LED_128_Instance_SBox_Instance_0_L5 ;
    wire LED_128_Instance_SBox_Instance_0_T2 ;
    wire LED_128_Instance_SBox_Instance_0_L4 ;
    wire LED_128_Instance_SBox_Instance_0_Q3 ;
    wire LED_128_Instance_SBox_Instance_0_L3 ;
    wire LED_128_Instance_SBox_Instance_0_Q2 ;
    wire LED_128_Instance_SBox_Instance_0_T0 ;
    wire LED_128_Instance_SBox_Instance_0_L2 ;
    wire LED_128_Instance_SBox_Instance_0_L1 ;
    wire LED_128_Instance_SBox_Instance_0_L0 ;
    wire LED_128_Instance_SBox_Instance_1_L8 ;
    wire LED_128_Instance_SBox_Instance_1_L7 ;
    wire LED_128_Instance_SBox_Instance_1_T3 ;
    wire LED_128_Instance_SBox_Instance_1_T1 ;
    wire LED_128_Instance_SBox_Instance_1_Q7 ;
    wire LED_128_Instance_SBox_Instance_1_Q6 ;
    wire LED_128_Instance_SBox_Instance_1_L5 ;
    wire LED_128_Instance_SBox_Instance_1_T2 ;
    wire LED_128_Instance_SBox_Instance_1_L4 ;
    wire LED_128_Instance_SBox_Instance_1_Q3 ;
    wire LED_128_Instance_SBox_Instance_1_L3 ;
    wire LED_128_Instance_SBox_Instance_1_Q2 ;
    wire LED_128_Instance_SBox_Instance_1_T0 ;
    wire LED_128_Instance_SBox_Instance_1_L2 ;
    wire LED_128_Instance_SBox_Instance_1_L1 ;
    wire LED_128_Instance_SBox_Instance_1_L0 ;
    wire LED_128_Instance_SBox_Instance_2_L8 ;
    wire LED_128_Instance_SBox_Instance_2_L7 ;
    wire LED_128_Instance_SBox_Instance_2_T3 ;
    wire LED_128_Instance_SBox_Instance_2_T1 ;
    wire LED_128_Instance_SBox_Instance_2_Q7 ;
    wire LED_128_Instance_SBox_Instance_2_Q6 ;
    wire LED_128_Instance_SBox_Instance_2_L5 ;
    wire LED_128_Instance_SBox_Instance_2_T2 ;
    wire LED_128_Instance_SBox_Instance_2_L4 ;
    wire LED_128_Instance_SBox_Instance_2_Q3 ;
    wire LED_128_Instance_SBox_Instance_2_L3 ;
    wire LED_128_Instance_SBox_Instance_2_Q2 ;
    wire LED_128_Instance_SBox_Instance_2_T0 ;
    wire LED_128_Instance_SBox_Instance_2_L2 ;
    wire LED_128_Instance_SBox_Instance_2_L1 ;
    wire LED_128_Instance_SBox_Instance_2_L0 ;
    wire LED_128_Instance_SBox_Instance_3_L8 ;
    wire LED_128_Instance_SBox_Instance_3_L7 ;
    wire LED_128_Instance_SBox_Instance_3_T3 ;
    wire LED_128_Instance_SBox_Instance_3_T1 ;
    wire LED_128_Instance_SBox_Instance_3_Q7 ;
    wire LED_128_Instance_SBox_Instance_3_Q6 ;
    wire LED_128_Instance_SBox_Instance_3_L5 ;
    wire LED_128_Instance_SBox_Instance_3_T2 ;
    wire LED_128_Instance_SBox_Instance_3_L4 ;
    wire LED_128_Instance_SBox_Instance_3_Q3 ;
    wire LED_128_Instance_SBox_Instance_3_L3 ;
    wire LED_128_Instance_SBox_Instance_3_Q2 ;
    wire LED_128_Instance_SBox_Instance_3_T0 ;
    wire LED_128_Instance_SBox_Instance_3_L2 ;
    wire LED_128_Instance_SBox_Instance_3_L1 ;
    wire LED_128_Instance_SBox_Instance_3_L0 ;
    wire LED_128_Instance_SBox_Instance_4_L8 ;
    wire LED_128_Instance_SBox_Instance_4_L7 ;
    wire LED_128_Instance_SBox_Instance_4_T3 ;
    wire LED_128_Instance_SBox_Instance_4_T1 ;
    wire LED_128_Instance_SBox_Instance_4_Q7 ;
    wire LED_128_Instance_SBox_Instance_4_Q6 ;
    wire LED_128_Instance_SBox_Instance_4_L5 ;
    wire LED_128_Instance_SBox_Instance_4_T2 ;
    wire LED_128_Instance_SBox_Instance_4_L4 ;
    wire LED_128_Instance_SBox_Instance_4_Q3 ;
    wire LED_128_Instance_SBox_Instance_4_L3 ;
    wire LED_128_Instance_SBox_Instance_4_Q2 ;
    wire LED_128_Instance_SBox_Instance_4_T0 ;
    wire LED_128_Instance_SBox_Instance_4_L2 ;
    wire LED_128_Instance_SBox_Instance_4_L1 ;
    wire LED_128_Instance_SBox_Instance_4_L0 ;
    wire LED_128_Instance_SBox_Instance_5_L8 ;
    wire LED_128_Instance_SBox_Instance_5_L7 ;
    wire LED_128_Instance_SBox_Instance_5_T3 ;
    wire LED_128_Instance_SBox_Instance_5_T1 ;
    wire LED_128_Instance_SBox_Instance_5_Q7 ;
    wire LED_128_Instance_SBox_Instance_5_Q6 ;
    wire LED_128_Instance_SBox_Instance_5_L5 ;
    wire LED_128_Instance_SBox_Instance_5_T2 ;
    wire LED_128_Instance_SBox_Instance_5_L4 ;
    wire LED_128_Instance_SBox_Instance_5_Q3 ;
    wire LED_128_Instance_SBox_Instance_5_L3 ;
    wire LED_128_Instance_SBox_Instance_5_Q2 ;
    wire LED_128_Instance_SBox_Instance_5_T0 ;
    wire LED_128_Instance_SBox_Instance_5_L2 ;
    wire LED_128_Instance_SBox_Instance_5_L1 ;
    wire LED_128_Instance_SBox_Instance_5_L0 ;
    wire LED_128_Instance_SBox_Instance_6_L8 ;
    wire LED_128_Instance_SBox_Instance_6_L7 ;
    wire LED_128_Instance_SBox_Instance_6_T3 ;
    wire LED_128_Instance_SBox_Instance_6_T1 ;
    wire LED_128_Instance_SBox_Instance_6_Q7 ;
    wire LED_128_Instance_SBox_Instance_6_Q6 ;
    wire LED_128_Instance_SBox_Instance_6_L5 ;
    wire LED_128_Instance_SBox_Instance_6_T2 ;
    wire LED_128_Instance_SBox_Instance_6_L4 ;
    wire LED_128_Instance_SBox_Instance_6_Q3 ;
    wire LED_128_Instance_SBox_Instance_6_L3 ;
    wire LED_128_Instance_SBox_Instance_6_Q2 ;
    wire LED_128_Instance_SBox_Instance_6_T0 ;
    wire LED_128_Instance_SBox_Instance_6_L2 ;
    wire LED_128_Instance_SBox_Instance_6_L1 ;
    wire LED_128_Instance_SBox_Instance_6_L0 ;
    wire LED_128_Instance_SBox_Instance_7_L8 ;
    wire LED_128_Instance_SBox_Instance_7_L7 ;
    wire LED_128_Instance_SBox_Instance_7_T3 ;
    wire LED_128_Instance_SBox_Instance_7_T1 ;
    wire LED_128_Instance_SBox_Instance_7_Q7 ;
    wire LED_128_Instance_SBox_Instance_7_Q6 ;
    wire LED_128_Instance_SBox_Instance_7_L5 ;
    wire LED_128_Instance_SBox_Instance_7_T2 ;
    wire LED_128_Instance_SBox_Instance_7_L4 ;
    wire LED_128_Instance_SBox_Instance_7_Q3 ;
    wire LED_128_Instance_SBox_Instance_7_L3 ;
    wire LED_128_Instance_SBox_Instance_7_Q2 ;
    wire LED_128_Instance_SBox_Instance_7_T0 ;
    wire LED_128_Instance_SBox_Instance_7_L2 ;
    wire LED_128_Instance_SBox_Instance_7_L1 ;
    wire LED_128_Instance_SBox_Instance_7_L0 ;
    wire LED_128_Instance_SBox_Instance_8_L8 ;
    wire LED_128_Instance_SBox_Instance_8_L7 ;
    wire LED_128_Instance_SBox_Instance_8_T3 ;
    wire LED_128_Instance_SBox_Instance_8_T1 ;
    wire LED_128_Instance_SBox_Instance_8_Q7 ;
    wire LED_128_Instance_SBox_Instance_8_Q6 ;
    wire LED_128_Instance_SBox_Instance_8_L5 ;
    wire LED_128_Instance_SBox_Instance_8_T2 ;
    wire LED_128_Instance_SBox_Instance_8_L4 ;
    wire LED_128_Instance_SBox_Instance_8_Q3 ;
    wire LED_128_Instance_SBox_Instance_8_L3 ;
    wire LED_128_Instance_SBox_Instance_8_Q2 ;
    wire LED_128_Instance_SBox_Instance_8_T0 ;
    wire LED_128_Instance_SBox_Instance_8_L2 ;
    wire LED_128_Instance_SBox_Instance_8_L1 ;
    wire LED_128_Instance_SBox_Instance_8_L0 ;
    wire LED_128_Instance_SBox_Instance_9_L8 ;
    wire LED_128_Instance_SBox_Instance_9_L7 ;
    wire LED_128_Instance_SBox_Instance_9_T3 ;
    wire LED_128_Instance_SBox_Instance_9_T1 ;
    wire LED_128_Instance_SBox_Instance_9_Q7 ;
    wire LED_128_Instance_SBox_Instance_9_Q6 ;
    wire LED_128_Instance_SBox_Instance_9_L5 ;
    wire LED_128_Instance_SBox_Instance_9_T2 ;
    wire LED_128_Instance_SBox_Instance_9_L4 ;
    wire LED_128_Instance_SBox_Instance_9_Q3 ;
    wire LED_128_Instance_SBox_Instance_9_L3 ;
    wire LED_128_Instance_SBox_Instance_9_Q2 ;
    wire LED_128_Instance_SBox_Instance_9_T0 ;
    wire LED_128_Instance_SBox_Instance_9_L2 ;
    wire LED_128_Instance_SBox_Instance_9_L1 ;
    wire LED_128_Instance_SBox_Instance_9_L0 ;
    wire LED_128_Instance_SBox_Instance_10_L8 ;
    wire LED_128_Instance_SBox_Instance_10_L7 ;
    wire LED_128_Instance_SBox_Instance_10_T3 ;
    wire LED_128_Instance_SBox_Instance_10_T1 ;
    wire LED_128_Instance_SBox_Instance_10_Q7 ;
    wire LED_128_Instance_SBox_Instance_10_Q6 ;
    wire LED_128_Instance_SBox_Instance_10_L5 ;
    wire LED_128_Instance_SBox_Instance_10_T2 ;
    wire LED_128_Instance_SBox_Instance_10_L4 ;
    wire LED_128_Instance_SBox_Instance_10_Q3 ;
    wire LED_128_Instance_SBox_Instance_10_L3 ;
    wire LED_128_Instance_SBox_Instance_10_Q2 ;
    wire LED_128_Instance_SBox_Instance_10_T0 ;
    wire LED_128_Instance_SBox_Instance_10_L2 ;
    wire LED_128_Instance_SBox_Instance_10_L1 ;
    wire LED_128_Instance_SBox_Instance_10_L0 ;
    wire LED_128_Instance_SBox_Instance_11_L8 ;
    wire LED_128_Instance_SBox_Instance_11_L7 ;
    wire LED_128_Instance_SBox_Instance_11_T3 ;
    wire LED_128_Instance_SBox_Instance_11_T1 ;
    wire LED_128_Instance_SBox_Instance_11_Q7 ;
    wire LED_128_Instance_SBox_Instance_11_Q6 ;
    wire LED_128_Instance_SBox_Instance_11_L5 ;
    wire LED_128_Instance_SBox_Instance_11_T2 ;
    wire LED_128_Instance_SBox_Instance_11_L4 ;
    wire LED_128_Instance_SBox_Instance_11_Q3 ;
    wire LED_128_Instance_SBox_Instance_11_L3 ;
    wire LED_128_Instance_SBox_Instance_11_Q2 ;
    wire LED_128_Instance_SBox_Instance_11_T0 ;
    wire LED_128_Instance_SBox_Instance_11_L2 ;
    wire LED_128_Instance_SBox_Instance_11_L1 ;
    wire LED_128_Instance_SBox_Instance_11_L0 ;
    wire LED_128_Instance_SBox_Instance_12_L8 ;
    wire LED_128_Instance_SBox_Instance_12_L7 ;
    wire LED_128_Instance_SBox_Instance_12_T3 ;
    wire LED_128_Instance_SBox_Instance_12_T1 ;
    wire LED_128_Instance_SBox_Instance_12_Q7 ;
    wire LED_128_Instance_SBox_Instance_12_Q6 ;
    wire LED_128_Instance_SBox_Instance_12_L5 ;
    wire LED_128_Instance_SBox_Instance_12_T2 ;
    wire LED_128_Instance_SBox_Instance_12_L4 ;
    wire LED_128_Instance_SBox_Instance_12_Q3 ;
    wire LED_128_Instance_SBox_Instance_12_L3 ;
    wire LED_128_Instance_SBox_Instance_12_Q2 ;
    wire LED_128_Instance_SBox_Instance_12_T0 ;
    wire LED_128_Instance_SBox_Instance_12_L2 ;
    wire LED_128_Instance_SBox_Instance_12_L1 ;
    wire LED_128_Instance_SBox_Instance_12_L0 ;
    wire LED_128_Instance_SBox_Instance_13_L8 ;
    wire LED_128_Instance_SBox_Instance_13_L7 ;
    wire LED_128_Instance_SBox_Instance_13_T3 ;
    wire LED_128_Instance_SBox_Instance_13_T1 ;
    wire LED_128_Instance_SBox_Instance_13_Q7 ;
    wire LED_128_Instance_SBox_Instance_13_Q6 ;
    wire LED_128_Instance_SBox_Instance_13_L5 ;
    wire LED_128_Instance_SBox_Instance_13_T2 ;
    wire LED_128_Instance_SBox_Instance_13_L4 ;
    wire LED_128_Instance_SBox_Instance_13_Q3 ;
    wire LED_128_Instance_SBox_Instance_13_L3 ;
    wire LED_128_Instance_SBox_Instance_13_Q2 ;
    wire LED_128_Instance_SBox_Instance_13_T0 ;
    wire LED_128_Instance_SBox_Instance_13_L2 ;
    wire LED_128_Instance_SBox_Instance_13_L1 ;
    wire LED_128_Instance_SBox_Instance_13_L0 ;
    wire LED_128_Instance_SBox_Instance_14_L8 ;
    wire LED_128_Instance_SBox_Instance_14_L7 ;
    wire LED_128_Instance_SBox_Instance_14_T3 ;
    wire LED_128_Instance_SBox_Instance_14_T1 ;
    wire LED_128_Instance_SBox_Instance_14_Q7 ;
    wire LED_128_Instance_SBox_Instance_14_Q6 ;
    wire LED_128_Instance_SBox_Instance_14_L5 ;
    wire LED_128_Instance_SBox_Instance_14_T2 ;
    wire LED_128_Instance_SBox_Instance_14_L4 ;
    wire LED_128_Instance_SBox_Instance_14_Q3 ;
    wire LED_128_Instance_SBox_Instance_14_L3 ;
    wire LED_128_Instance_SBox_Instance_14_Q2 ;
    wire LED_128_Instance_SBox_Instance_14_T0 ;
    wire LED_128_Instance_SBox_Instance_14_L2 ;
    wire LED_128_Instance_SBox_Instance_14_L1 ;
    wire LED_128_Instance_SBox_Instance_14_L0 ;
    wire LED_128_Instance_SBox_Instance_15_L8 ;
    wire LED_128_Instance_SBox_Instance_15_L7 ;
    wire LED_128_Instance_SBox_Instance_15_T3 ;
    wire LED_128_Instance_SBox_Instance_15_T1 ;
    wire LED_128_Instance_SBox_Instance_15_Q7 ;
    wire LED_128_Instance_SBox_Instance_15_Q6 ;
    wire LED_128_Instance_SBox_Instance_15_L5 ;
    wire LED_128_Instance_SBox_Instance_15_T2 ;
    wire LED_128_Instance_SBox_Instance_15_L4 ;
    wire LED_128_Instance_SBox_Instance_15_Q3 ;
    wire LED_128_Instance_SBox_Instance_15_L3 ;
    wire LED_128_Instance_SBox_Instance_15_Q2 ;
    wire LED_128_Instance_SBox_Instance_15_T0 ;
    wire LED_128_Instance_SBox_Instance_15_L2 ;
    wire LED_128_Instance_SBox_Instance_15_L1 ;
    wire LED_128_Instance_SBox_Instance_15_L0 ;
    wire LED_128_Instance_MCS_Instance_0_n42 ;
    wire LED_128_Instance_MCS_Instance_0_n41 ;
    wire LED_128_Instance_MCS_Instance_0_n40 ;
    wire LED_128_Instance_MCS_Instance_0_n39 ;
    wire LED_128_Instance_MCS_Instance_0_n38 ;
    wire LED_128_Instance_MCS_Instance_0_n37 ;
    wire LED_128_Instance_MCS_Instance_0_n36 ;
    wire LED_128_Instance_MCS_Instance_0_n35 ;
    wire LED_128_Instance_MCS_Instance_0_n34 ;
    wire LED_128_Instance_MCS_Instance_0_n33 ;
    wire LED_128_Instance_MCS_Instance_0_n32 ;
    wire LED_128_Instance_MCS_Instance_0_n31 ;
    wire LED_128_Instance_MCS_Instance_0_n30 ;
    wire LED_128_Instance_MCS_Instance_0_n29 ;
    wire LED_128_Instance_MCS_Instance_0_n28 ;
    wire LED_128_Instance_MCS_Instance_0_n27 ;
    wire LED_128_Instance_MCS_Instance_0_n26 ;
    wire LED_128_Instance_MCS_Instance_0_n25 ;
    wire LED_128_Instance_MCS_Instance_0_n24 ;
    wire LED_128_Instance_MCS_Instance_0_n23 ;
    wire LED_128_Instance_MCS_Instance_0_n22 ;
    wire LED_128_Instance_MCS_Instance_0_n21 ;
    wire LED_128_Instance_MCS_Instance_0_n20 ;
    wire LED_128_Instance_MCS_Instance_0_n19 ;
    wire LED_128_Instance_MCS_Instance_0_n18 ;
    wire LED_128_Instance_MCS_Instance_0_n17 ;
    wire LED_128_Instance_MCS_Instance_0_n16 ;
    wire LED_128_Instance_MCS_Instance_0_n15 ;
    wire LED_128_Instance_MCS_Instance_0_n14 ;
    wire LED_128_Instance_MCS_Instance_0_n13 ;
    wire LED_128_Instance_MCS_Instance_0_n12 ;
    wire LED_128_Instance_MCS_Instance_0_n11 ;
    wire LED_128_Instance_MCS_Instance_0_n10 ;
    wire LED_128_Instance_MCS_Instance_0_n9 ;
    wire LED_128_Instance_MCS_Instance_0_n8 ;
    wire LED_128_Instance_MCS_Instance_0_n7 ;
    wire LED_128_Instance_MCS_Instance_0_n6 ;
    wire LED_128_Instance_MCS_Instance_0_n5 ;
    wire LED_128_Instance_MCS_Instance_0_n4 ;
    wire LED_128_Instance_MCS_Instance_0_n3 ;
    wire LED_128_Instance_MCS_Instance_0_n2 ;
    wire LED_128_Instance_MCS_Instance_0_n1 ;
    wire LED_128_Instance_MCS_Instance_1_n42 ;
    wire LED_128_Instance_MCS_Instance_1_n41 ;
    wire LED_128_Instance_MCS_Instance_1_n40 ;
    wire LED_128_Instance_MCS_Instance_1_n39 ;
    wire LED_128_Instance_MCS_Instance_1_n38 ;
    wire LED_128_Instance_MCS_Instance_1_n37 ;
    wire LED_128_Instance_MCS_Instance_1_n36 ;
    wire LED_128_Instance_MCS_Instance_1_n35 ;
    wire LED_128_Instance_MCS_Instance_1_n34 ;
    wire LED_128_Instance_MCS_Instance_1_n33 ;
    wire LED_128_Instance_MCS_Instance_1_n32 ;
    wire LED_128_Instance_MCS_Instance_1_n31 ;
    wire LED_128_Instance_MCS_Instance_1_n30 ;
    wire LED_128_Instance_MCS_Instance_1_n29 ;
    wire LED_128_Instance_MCS_Instance_1_n28 ;
    wire LED_128_Instance_MCS_Instance_1_n27 ;
    wire LED_128_Instance_MCS_Instance_1_n26 ;
    wire LED_128_Instance_MCS_Instance_1_n25 ;
    wire LED_128_Instance_MCS_Instance_1_n24 ;
    wire LED_128_Instance_MCS_Instance_1_n23 ;
    wire LED_128_Instance_MCS_Instance_1_n22 ;
    wire LED_128_Instance_MCS_Instance_1_n21 ;
    wire LED_128_Instance_MCS_Instance_1_n20 ;
    wire LED_128_Instance_MCS_Instance_1_n19 ;
    wire LED_128_Instance_MCS_Instance_1_n18 ;
    wire LED_128_Instance_MCS_Instance_1_n17 ;
    wire LED_128_Instance_MCS_Instance_1_n16 ;
    wire LED_128_Instance_MCS_Instance_1_n15 ;
    wire LED_128_Instance_MCS_Instance_1_n14 ;
    wire LED_128_Instance_MCS_Instance_1_n13 ;
    wire LED_128_Instance_MCS_Instance_1_n12 ;
    wire LED_128_Instance_MCS_Instance_1_n11 ;
    wire LED_128_Instance_MCS_Instance_1_n10 ;
    wire LED_128_Instance_MCS_Instance_1_n9 ;
    wire LED_128_Instance_MCS_Instance_1_n8 ;
    wire LED_128_Instance_MCS_Instance_1_n7 ;
    wire LED_128_Instance_MCS_Instance_1_n6 ;
    wire LED_128_Instance_MCS_Instance_1_n5 ;
    wire LED_128_Instance_MCS_Instance_1_n4 ;
    wire LED_128_Instance_MCS_Instance_1_n3 ;
    wire LED_128_Instance_MCS_Instance_1_n2 ;
    wire LED_128_Instance_MCS_Instance_1_n1 ;
    wire LED_128_Instance_MCS_Instance_2_n42 ;
    wire LED_128_Instance_MCS_Instance_2_n41 ;
    wire LED_128_Instance_MCS_Instance_2_n40 ;
    wire LED_128_Instance_MCS_Instance_2_n39 ;
    wire LED_128_Instance_MCS_Instance_2_n38 ;
    wire LED_128_Instance_MCS_Instance_2_n37 ;
    wire LED_128_Instance_MCS_Instance_2_n36 ;
    wire LED_128_Instance_MCS_Instance_2_n35 ;
    wire LED_128_Instance_MCS_Instance_2_n34 ;
    wire LED_128_Instance_MCS_Instance_2_n33 ;
    wire LED_128_Instance_MCS_Instance_2_n32 ;
    wire LED_128_Instance_MCS_Instance_2_n31 ;
    wire LED_128_Instance_MCS_Instance_2_n30 ;
    wire LED_128_Instance_MCS_Instance_2_n29 ;
    wire LED_128_Instance_MCS_Instance_2_n28 ;
    wire LED_128_Instance_MCS_Instance_2_n27 ;
    wire LED_128_Instance_MCS_Instance_2_n26 ;
    wire LED_128_Instance_MCS_Instance_2_n25 ;
    wire LED_128_Instance_MCS_Instance_2_n24 ;
    wire LED_128_Instance_MCS_Instance_2_n23 ;
    wire LED_128_Instance_MCS_Instance_2_n22 ;
    wire LED_128_Instance_MCS_Instance_2_n21 ;
    wire LED_128_Instance_MCS_Instance_2_n20 ;
    wire LED_128_Instance_MCS_Instance_2_n19 ;
    wire LED_128_Instance_MCS_Instance_2_n18 ;
    wire LED_128_Instance_MCS_Instance_2_n17 ;
    wire LED_128_Instance_MCS_Instance_2_n16 ;
    wire LED_128_Instance_MCS_Instance_2_n15 ;
    wire LED_128_Instance_MCS_Instance_2_n14 ;
    wire LED_128_Instance_MCS_Instance_2_n13 ;
    wire LED_128_Instance_MCS_Instance_2_n12 ;
    wire LED_128_Instance_MCS_Instance_2_n11 ;
    wire LED_128_Instance_MCS_Instance_2_n10 ;
    wire LED_128_Instance_MCS_Instance_2_n9 ;
    wire LED_128_Instance_MCS_Instance_2_n8 ;
    wire LED_128_Instance_MCS_Instance_2_n7 ;
    wire LED_128_Instance_MCS_Instance_2_n6 ;
    wire LED_128_Instance_MCS_Instance_2_n5 ;
    wire LED_128_Instance_MCS_Instance_2_n4 ;
    wire LED_128_Instance_MCS_Instance_2_n3 ;
    wire LED_128_Instance_MCS_Instance_2_n2 ;
    wire LED_128_Instance_MCS_Instance_2_n1 ;
    wire LED_128_Instance_MCS_Instance_3_n42 ;
    wire LED_128_Instance_MCS_Instance_3_n41 ;
    wire LED_128_Instance_MCS_Instance_3_n40 ;
    wire LED_128_Instance_MCS_Instance_3_n39 ;
    wire LED_128_Instance_MCS_Instance_3_n38 ;
    wire LED_128_Instance_MCS_Instance_3_n37 ;
    wire LED_128_Instance_MCS_Instance_3_n36 ;
    wire LED_128_Instance_MCS_Instance_3_n35 ;
    wire LED_128_Instance_MCS_Instance_3_n34 ;
    wire LED_128_Instance_MCS_Instance_3_n33 ;
    wire LED_128_Instance_MCS_Instance_3_n32 ;
    wire LED_128_Instance_MCS_Instance_3_n31 ;
    wire LED_128_Instance_MCS_Instance_3_n30 ;
    wire LED_128_Instance_MCS_Instance_3_n29 ;
    wire LED_128_Instance_MCS_Instance_3_n28 ;
    wire LED_128_Instance_MCS_Instance_3_n27 ;
    wire LED_128_Instance_MCS_Instance_3_n26 ;
    wire LED_128_Instance_MCS_Instance_3_n25 ;
    wire LED_128_Instance_MCS_Instance_3_n24 ;
    wire LED_128_Instance_MCS_Instance_3_n23 ;
    wire LED_128_Instance_MCS_Instance_3_n22 ;
    wire LED_128_Instance_MCS_Instance_3_n21 ;
    wire LED_128_Instance_MCS_Instance_3_n20 ;
    wire LED_128_Instance_MCS_Instance_3_n19 ;
    wire LED_128_Instance_MCS_Instance_3_n18 ;
    wire LED_128_Instance_MCS_Instance_3_n17 ;
    wire LED_128_Instance_MCS_Instance_3_n16 ;
    wire LED_128_Instance_MCS_Instance_3_n15 ;
    wire LED_128_Instance_MCS_Instance_3_n14 ;
    wire LED_128_Instance_MCS_Instance_3_n13 ;
    wire LED_128_Instance_MCS_Instance_3_n12 ;
    wire LED_128_Instance_MCS_Instance_3_n11 ;
    wire LED_128_Instance_MCS_Instance_3_n10 ;
    wire LED_128_Instance_MCS_Instance_3_n9 ;
    wire LED_128_Instance_MCS_Instance_3_n8 ;
    wire LED_128_Instance_MCS_Instance_3_n7 ;
    wire LED_128_Instance_MCS_Instance_3_n6 ;
    wire LED_128_Instance_MCS_Instance_3_n5 ;
    wire LED_128_Instance_MCS_Instance_3_n4 ;
    wire LED_128_Instance_MCS_Instance_3_n3 ;
    wire LED_128_Instance_MCS_Instance_3_n2 ;
    wire LED_128_Instance_MCS_Instance_3_n1 ;
    wire LED_128_Instance_ks_reg_2__Q ;
    wire [5:0] roundconstant ;
    wire [63:0] LED_128_Instance_subcells_out ;
    wire [63:0] LED_128_Instance_addconst_out ;
    wire [63:0] LED_128_Instance_addroundkey_tmp ;
    wire [63:0] LED_128_Instance_current_roundkey ;
    wire [63:0] LED_128_Instance_state0 ;
    wire [54:3] LED_128_Instance_addroundkey_out ;
    wire [63:0] LED_128_Instance_mixcolumns_out ;
    wire new_AGEMA_signal_1877 ;
    wire new_AGEMA_signal_1878 ;
    wire new_AGEMA_signal_1879 ;
    wire new_AGEMA_signal_1880 ;
    wire new_AGEMA_signal_1882 ;
    wire new_AGEMA_signal_1883 ;
    wire new_AGEMA_signal_1884 ;
    wire new_AGEMA_signal_1885 ;
    wire new_AGEMA_signal_1886 ;
    wire new_AGEMA_signal_1887 ;
    wire new_AGEMA_signal_1888 ;
    wire new_AGEMA_signal_1889 ;
    wire new_AGEMA_signal_1890 ;
    wire new_AGEMA_signal_1891 ;
    wire new_AGEMA_signal_1892 ;
    wire new_AGEMA_signal_1893 ;
    wire new_AGEMA_signal_1900 ;
    wire new_AGEMA_signal_1901 ;
    wire new_AGEMA_signal_1902 ;
    wire new_AGEMA_signal_1909 ;
    wire new_AGEMA_signal_1910 ;
    wire new_AGEMA_signal_1911 ;
    wire new_AGEMA_signal_1918 ;
    wire new_AGEMA_signal_1919 ;
    wire new_AGEMA_signal_1920 ;
    wire new_AGEMA_signal_1927 ;
    wire new_AGEMA_signal_1928 ;
    wire new_AGEMA_signal_1929 ;
    wire new_AGEMA_signal_1936 ;
    wire new_AGEMA_signal_1937 ;
    wire new_AGEMA_signal_1938 ;
    wire new_AGEMA_signal_1945 ;
    wire new_AGEMA_signal_1946 ;
    wire new_AGEMA_signal_1947 ;
    wire new_AGEMA_signal_1954 ;
    wire new_AGEMA_signal_1955 ;
    wire new_AGEMA_signal_1956 ;
    wire new_AGEMA_signal_1963 ;
    wire new_AGEMA_signal_1964 ;
    wire new_AGEMA_signal_1965 ;
    wire new_AGEMA_signal_1972 ;
    wire new_AGEMA_signal_1973 ;
    wire new_AGEMA_signal_1974 ;
    wire new_AGEMA_signal_1981 ;
    wire new_AGEMA_signal_1982 ;
    wire new_AGEMA_signal_1983 ;
    wire new_AGEMA_signal_1990 ;
    wire new_AGEMA_signal_1991 ;
    wire new_AGEMA_signal_1992 ;
    wire new_AGEMA_signal_1999 ;
    wire new_AGEMA_signal_2000 ;
    wire new_AGEMA_signal_2001 ;
    wire new_AGEMA_signal_2008 ;
    wire new_AGEMA_signal_2009 ;
    wire new_AGEMA_signal_2010 ;
    wire new_AGEMA_signal_2017 ;
    wire new_AGEMA_signal_2018 ;
    wire new_AGEMA_signal_2019 ;
    wire new_AGEMA_signal_2026 ;
    wire new_AGEMA_signal_2027 ;
    wire new_AGEMA_signal_2028 ;
    wire new_AGEMA_signal_2035 ;
    wire new_AGEMA_signal_2036 ;
    wire new_AGEMA_signal_2037 ;
    wire new_AGEMA_signal_2044 ;
    wire new_AGEMA_signal_2045 ;
    wire new_AGEMA_signal_2046 ;
    wire new_AGEMA_signal_2053 ;
    wire new_AGEMA_signal_2054 ;
    wire new_AGEMA_signal_2055 ;
    wire new_AGEMA_signal_2062 ;
    wire new_AGEMA_signal_2063 ;
    wire new_AGEMA_signal_2064 ;
    wire new_AGEMA_signal_2071 ;
    wire new_AGEMA_signal_2072 ;
    wire new_AGEMA_signal_2073 ;
    wire new_AGEMA_signal_2080 ;
    wire new_AGEMA_signal_2081 ;
    wire new_AGEMA_signal_2082 ;
    wire new_AGEMA_signal_2089 ;
    wire new_AGEMA_signal_2090 ;
    wire new_AGEMA_signal_2091 ;
    wire new_AGEMA_signal_2098 ;
    wire new_AGEMA_signal_2099 ;
    wire new_AGEMA_signal_2100 ;
    wire new_AGEMA_signal_2107 ;
    wire new_AGEMA_signal_2108 ;
    wire new_AGEMA_signal_2109 ;
    wire new_AGEMA_signal_2116 ;
    wire new_AGEMA_signal_2117 ;
    wire new_AGEMA_signal_2118 ;
    wire new_AGEMA_signal_2125 ;
    wire new_AGEMA_signal_2126 ;
    wire new_AGEMA_signal_2127 ;
    wire new_AGEMA_signal_2134 ;
    wire new_AGEMA_signal_2135 ;
    wire new_AGEMA_signal_2136 ;
    wire new_AGEMA_signal_2143 ;
    wire new_AGEMA_signal_2144 ;
    wire new_AGEMA_signal_2145 ;
    wire new_AGEMA_signal_2152 ;
    wire new_AGEMA_signal_2153 ;
    wire new_AGEMA_signal_2154 ;
    wire new_AGEMA_signal_2161 ;
    wire new_AGEMA_signal_2162 ;
    wire new_AGEMA_signal_2163 ;
    wire new_AGEMA_signal_2170 ;
    wire new_AGEMA_signal_2171 ;
    wire new_AGEMA_signal_2172 ;
    wire new_AGEMA_signal_2179 ;
    wire new_AGEMA_signal_2180 ;
    wire new_AGEMA_signal_2181 ;
    wire new_AGEMA_signal_2188 ;
    wire new_AGEMA_signal_2189 ;
    wire new_AGEMA_signal_2190 ;
    wire new_AGEMA_signal_2197 ;
    wire new_AGEMA_signal_2198 ;
    wire new_AGEMA_signal_2199 ;
    wire new_AGEMA_signal_2206 ;
    wire new_AGEMA_signal_2207 ;
    wire new_AGEMA_signal_2208 ;
    wire new_AGEMA_signal_2215 ;
    wire new_AGEMA_signal_2216 ;
    wire new_AGEMA_signal_2217 ;
    wire new_AGEMA_signal_2224 ;
    wire new_AGEMA_signal_2225 ;
    wire new_AGEMA_signal_2226 ;
    wire new_AGEMA_signal_2233 ;
    wire new_AGEMA_signal_2234 ;
    wire new_AGEMA_signal_2235 ;
    wire new_AGEMA_signal_2242 ;
    wire new_AGEMA_signal_2243 ;
    wire new_AGEMA_signal_2244 ;
    wire new_AGEMA_signal_2251 ;
    wire new_AGEMA_signal_2252 ;
    wire new_AGEMA_signal_2253 ;
    wire new_AGEMA_signal_2260 ;
    wire new_AGEMA_signal_2261 ;
    wire new_AGEMA_signal_2262 ;
    wire new_AGEMA_signal_2269 ;
    wire new_AGEMA_signal_2270 ;
    wire new_AGEMA_signal_2271 ;
    wire new_AGEMA_signal_2278 ;
    wire new_AGEMA_signal_2279 ;
    wire new_AGEMA_signal_2280 ;
    wire new_AGEMA_signal_2287 ;
    wire new_AGEMA_signal_2288 ;
    wire new_AGEMA_signal_2289 ;
    wire new_AGEMA_signal_2296 ;
    wire new_AGEMA_signal_2297 ;
    wire new_AGEMA_signal_2298 ;
    wire new_AGEMA_signal_2305 ;
    wire new_AGEMA_signal_2306 ;
    wire new_AGEMA_signal_2307 ;
    wire new_AGEMA_signal_2314 ;
    wire new_AGEMA_signal_2315 ;
    wire new_AGEMA_signal_2316 ;
    wire new_AGEMA_signal_2323 ;
    wire new_AGEMA_signal_2324 ;
    wire new_AGEMA_signal_2325 ;
    wire new_AGEMA_signal_2332 ;
    wire new_AGEMA_signal_2333 ;
    wire new_AGEMA_signal_2334 ;
    wire new_AGEMA_signal_2341 ;
    wire new_AGEMA_signal_2342 ;
    wire new_AGEMA_signal_2343 ;
    wire new_AGEMA_signal_2350 ;
    wire new_AGEMA_signal_2351 ;
    wire new_AGEMA_signal_2352 ;
    wire new_AGEMA_signal_2359 ;
    wire new_AGEMA_signal_2360 ;
    wire new_AGEMA_signal_2361 ;
    wire new_AGEMA_signal_2368 ;
    wire new_AGEMA_signal_2369 ;
    wire new_AGEMA_signal_2370 ;
    wire new_AGEMA_signal_2377 ;
    wire new_AGEMA_signal_2378 ;
    wire new_AGEMA_signal_2379 ;
    wire new_AGEMA_signal_2386 ;
    wire new_AGEMA_signal_2387 ;
    wire new_AGEMA_signal_2388 ;
    wire new_AGEMA_signal_2395 ;
    wire new_AGEMA_signal_2396 ;
    wire new_AGEMA_signal_2397 ;
    wire new_AGEMA_signal_2404 ;
    wire new_AGEMA_signal_2405 ;
    wire new_AGEMA_signal_2406 ;
    wire new_AGEMA_signal_2413 ;
    wire new_AGEMA_signal_2414 ;
    wire new_AGEMA_signal_2415 ;
    wire new_AGEMA_signal_2422 ;
    wire new_AGEMA_signal_2423 ;
    wire new_AGEMA_signal_2424 ;
    wire new_AGEMA_signal_2431 ;
    wire new_AGEMA_signal_2432 ;
    wire new_AGEMA_signal_2433 ;
    wire new_AGEMA_signal_2440 ;
    wire new_AGEMA_signal_2441 ;
    wire new_AGEMA_signal_2442 ;
    wire new_AGEMA_signal_2449 ;
    wire new_AGEMA_signal_2450 ;
    wire new_AGEMA_signal_2451 ;
    wire new_AGEMA_signal_2458 ;
    wire new_AGEMA_signal_2459 ;
    wire new_AGEMA_signal_2460 ;
    wire new_AGEMA_signal_2467 ;
    wire new_AGEMA_signal_2468 ;
    wire new_AGEMA_signal_2469 ;
    wire new_AGEMA_signal_2470 ;
    wire new_AGEMA_signal_2471 ;
    wire new_AGEMA_signal_2472 ;
    wire new_AGEMA_signal_2473 ;
    wire new_AGEMA_signal_2474 ;
    wire new_AGEMA_signal_2475 ;
    wire new_AGEMA_signal_2476 ;
    wire new_AGEMA_signal_2477 ;
    wire new_AGEMA_signal_2478 ;
    wire new_AGEMA_signal_2479 ;
    wire new_AGEMA_signal_2480 ;
    wire new_AGEMA_signal_2481 ;
    wire new_AGEMA_signal_2482 ;
    wire new_AGEMA_signal_2483 ;
    wire new_AGEMA_signal_2484 ;
    wire new_AGEMA_signal_2485 ;
    wire new_AGEMA_signal_2486 ;
    wire new_AGEMA_signal_2487 ;
    wire new_AGEMA_signal_2488 ;
    wire new_AGEMA_signal_2489 ;
    wire new_AGEMA_signal_2490 ;
    wire new_AGEMA_signal_2491 ;
    wire new_AGEMA_signal_2492 ;
    wire new_AGEMA_signal_2493 ;
    wire new_AGEMA_signal_2494 ;
    wire new_AGEMA_signal_2495 ;
    wire new_AGEMA_signal_2496 ;
    wire new_AGEMA_signal_2497 ;
    wire new_AGEMA_signal_2498 ;
    wire new_AGEMA_signal_2499 ;
    wire new_AGEMA_signal_2500 ;
    wire new_AGEMA_signal_2501 ;
    wire new_AGEMA_signal_2502 ;
    wire new_AGEMA_signal_2503 ;
    wire new_AGEMA_signal_2504 ;
    wire new_AGEMA_signal_2505 ;
    wire new_AGEMA_signal_2506 ;
    wire new_AGEMA_signal_2507 ;
    wire new_AGEMA_signal_2508 ;
    wire new_AGEMA_signal_2509 ;
    wire new_AGEMA_signal_2510 ;
    wire new_AGEMA_signal_2511 ;
    wire new_AGEMA_signal_2512 ;
    wire new_AGEMA_signal_2513 ;
    wire new_AGEMA_signal_2514 ;
    wire new_AGEMA_signal_2515 ;
    wire new_AGEMA_signal_2516 ;
    wire new_AGEMA_signal_2517 ;
    wire new_AGEMA_signal_2518 ;
    wire new_AGEMA_signal_2519 ;
    wire new_AGEMA_signal_2520 ;
    wire new_AGEMA_signal_2521 ;
    wire new_AGEMA_signal_2522 ;
    wire new_AGEMA_signal_2523 ;
    wire new_AGEMA_signal_2524 ;
    wire new_AGEMA_signal_2525 ;
    wire new_AGEMA_signal_2526 ;
    wire new_AGEMA_signal_2527 ;
    wire new_AGEMA_signal_2528 ;
    wire new_AGEMA_signal_2529 ;
    wire new_AGEMA_signal_2530 ;
    wire new_AGEMA_signal_2531 ;
    wire new_AGEMA_signal_2532 ;
    wire new_AGEMA_signal_2533 ;
    wire new_AGEMA_signal_2534 ;
    wire new_AGEMA_signal_2535 ;
    wire new_AGEMA_signal_2536 ;
    wire new_AGEMA_signal_2537 ;
    wire new_AGEMA_signal_2538 ;
    wire new_AGEMA_signal_2539 ;
    wire new_AGEMA_signal_2540 ;
    wire new_AGEMA_signal_2541 ;
    wire new_AGEMA_signal_2542 ;
    wire new_AGEMA_signal_2543 ;
    wire new_AGEMA_signal_2544 ;
    wire new_AGEMA_signal_2545 ;
    wire new_AGEMA_signal_2546 ;
    wire new_AGEMA_signal_2547 ;
    wire new_AGEMA_signal_2548 ;
    wire new_AGEMA_signal_2549 ;
    wire new_AGEMA_signal_2550 ;
    wire new_AGEMA_signal_2551 ;
    wire new_AGEMA_signal_2552 ;
    wire new_AGEMA_signal_2553 ;
    wire new_AGEMA_signal_2554 ;
    wire new_AGEMA_signal_2555 ;
    wire new_AGEMA_signal_2556 ;
    wire new_AGEMA_signal_2557 ;
    wire new_AGEMA_signal_2558 ;
    wire new_AGEMA_signal_2559 ;
    wire new_AGEMA_signal_2560 ;
    wire new_AGEMA_signal_2561 ;
    wire new_AGEMA_signal_2562 ;
    wire new_AGEMA_signal_2563 ;
    wire new_AGEMA_signal_2564 ;
    wire new_AGEMA_signal_2565 ;
    wire new_AGEMA_signal_2566 ;
    wire new_AGEMA_signal_2567 ;
    wire new_AGEMA_signal_2568 ;
    wire new_AGEMA_signal_2569 ;
    wire new_AGEMA_signal_2570 ;
    wire new_AGEMA_signal_2571 ;
    wire new_AGEMA_signal_2572 ;
    wire new_AGEMA_signal_2573 ;
    wire new_AGEMA_signal_2574 ;
    wire new_AGEMA_signal_2575 ;
    wire new_AGEMA_signal_2576 ;
    wire new_AGEMA_signal_2577 ;
    wire new_AGEMA_signal_2578 ;
    wire new_AGEMA_signal_2579 ;
    wire new_AGEMA_signal_2580 ;
    wire new_AGEMA_signal_2581 ;
    wire new_AGEMA_signal_2582 ;
    wire new_AGEMA_signal_2583 ;
    wire new_AGEMA_signal_2584 ;
    wire new_AGEMA_signal_2585 ;
    wire new_AGEMA_signal_2586 ;
    wire new_AGEMA_signal_2587 ;
    wire new_AGEMA_signal_2588 ;
    wire new_AGEMA_signal_2589 ;
    wire new_AGEMA_signal_2590 ;
    wire new_AGEMA_signal_2591 ;
    wire new_AGEMA_signal_2592 ;
    wire new_AGEMA_signal_2593 ;
    wire new_AGEMA_signal_2594 ;
    wire new_AGEMA_signal_2595 ;
    wire new_AGEMA_signal_2596 ;
    wire new_AGEMA_signal_2597 ;
    wire new_AGEMA_signal_2598 ;
    wire new_AGEMA_signal_2599 ;
    wire new_AGEMA_signal_2600 ;
    wire new_AGEMA_signal_2601 ;
    wire new_AGEMA_signal_2602 ;
    wire new_AGEMA_signal_2603 ;
    wire new_AGEMA_signal_2604 ;
    wire new_AGEMA_signal_2605 ;
    wire new_AGEMA_signal_2606 ;
    wire new_AGEMA_signal_2607 ;
    wire new_AGEMA_signal_2608 ;
    wire new_AGEMA_signal_2609 ;
    wire new_AGEMA_signal_2610 ;
    wire new_AGEMA_signal_2611 ;
    wire new_AGEMA_signal_2612 ;
    wire new_AGEMA_signal_2613 ;
    wire new_AGEMA_signal_2614 ;
    wire new_AGEMA_signal_2615 ;
    wire new_AGEMA_signal_2616 ;
    wire new_AGEMA_signal_2617 ;
    wire new_AGEMA_signal_2618 ;
    wire new_AGEMA_signal_2619 ;
    wire new_AGEMA_signal_2620 ;
    wire new_AGEMA_signal_2621 ;
    wire new_AGEMA_signal_2622 ;
    wire new_AGEMA_signal_2623 ;
    wire new_AGEMA_signal_2624 ;
    wire new_AGEMA_signal_2625 ;
    wire new_AGEMA_signal_2626 ;
    wire new_AGEMA_signal_2627 ;
    wire new_AGEMA_signal_2628 ;
    wire new_AGEMA_signal_2629 ;
    wire new_AGEMA_signal_2630 ;
    wire new_AGEMA_signal_2631 ;
    wire new_AGEMA_signal_2632 ;
    wire new_AGEMA_signal_2633 ;
    wire new_AGEMA_signal_2634 ;
    wire new_AGEMA_signal_2635 ;
    wire new_AGEMA_signal_2636 ;
    wire new_AGEMA_signal_2637 ;
    wire new_AGEMA_signal_2638 ;
    wire new_AGEMA_signal_2639 ;
    wire new_AGEMA_signal_2640 ;
    wire new_AGEMA_signal_2641 ;
    wire new_AGEMA_signal_2642 ;
    wire new_AGEMA_signal_2643 ;
    wire new_AGEMA_signal_2644 ;
    wire new_AGEMA_signal_2645 ;
    wire new_AGEMA_signal_2646 ;
    wire new_AGEMA_signal_2647 ;
    wire new_AGEMA_signal_2648 ;
    wire new_AGEMA_signal_2649 ;
    wire new_AGEMA_signal_2650 ;
    wire new_AGEMA_signal_2651 ;
    wire new_AGEMA_signal_2652 ;
    wire new_AGEMA_signal_2653 ;
    wire new_AGEMA_signal_2654 ;
    wire new_AGEMA_signal_2655 ;
    wire new_AGEMA_signal_2656 ;
    wire new_AGEMA_signal_2657 ;
    wire new_AGEMA_signal_2658 ;
    wire new_AGEMA_signal_2659 ;
    wire new_AGEMA_signal_2660 ;
    wire new_AGEMA_signal_2661 ;
    wire new_AGEMA_signal_2662 ;
    wire new_AGEMA_signal_2663 ;
    wire new_AGEMA_signal_2664 ;
    wire new_AGEMA_signal_2665 ;
    wire new_AGEMA_signal_2666 ;
    wire new_AGEMA_signal_2667 ;
    wire new_AGEMA_signal_2668 ;
    wire new_AGEMA_signal_2669 ;
    wire new_AGEMA_signal_2670 ;
    wire new_AGEMA_signal_2671 ;
    wire new_AGEMA_signal_2672 ;
    wire new_AGEMA_signal_2673 ;
    wire new_AGEMA_signal_2674 ;
    wire new_AGEMA_signal_2675 ;
    wire new_AGEMA_signal_2676 ;
    wire new_AGEMA_signal_2677 ;
    wire new_AGEMA_signal_2678 ;
    wire new_AGEMA_signal_2679 ;
    wire new_AGEMA_signal_2680 ;
    wire new_AGEMA_signal_2681 ;
    wire new_AGEMA_signal_2682 ;
    wire new_AGEMA_signal_2683 ;
    wire new_AGEMA_signal_2684 ;
    wire new_AGEMA_signal_2685 ;
    wire new_AGEMA_signal_2686 ;
    wire new_AGEMA_signal_2687 ;
    wire new_AGEMA_signal_2688 ;
    wire new_AGEMA_signal_2689 ;
    wire new_AGEMA_signal_2690 ;
    wire new_AGEMA_signal_2691 ;
    wire new_AGEMA_signal_2692 ;
    wire new_AGEMA_signal_2693 ;
    wire new_AGEMA_signal_2694 ;
    wire new_AGEMA_signal_2695 ;
    wire new_AGEMA_signal_2696 ;
    wire new_AGEMA_signal_2697 ;
    wire new_AGEMA_signal_2698 ;
    wire new_AGEMA_signal_2699 ;
    wire new_AGEMA_signal_2700 ;
    wire new_AGEMA_signal_2701 ;
    wire new_AGEMA_signal_2702 ;
    wire new_AGEMA_signal_2703 ;
    wire new_AGEMA_signal_2704 ;
    wire new_AGEMA_signal_2705 ;
    wire new_AGEMA_signal_2706 ;
    wire new_AGEMA_signal_2707 ;
    wire new_AGEMA_signal_2708 ;
    wire new_AGEMA_signal_2709 ;
    wire new_AGEMA_signal_2710 ;
    wire new_AGEMA_signal_2711 ;
    wire new_AGEMA_signal_2712 ;
    wire new_AGEMA_signal_2713 ;
    wire new_AGEMA_signal_2714 ;
    wire new_AGEMA_signal_2715 ;
    wire new_AGEMA_signal_2716 ;
    wire new_AGEMA_signal_2717 ;
    wire new_AGEMA_signal_2718 ;
    wire new_AGEMA_signal_2719 ;
    wire new_AGEMA_signal_2720 ;
    wire new_AGEMA_signal_2721 ;
    wire new_AGEMA_signal_2722 ;
    wire new_AGEMA_signal_2723 ;
    wire new_AGEMA_signal_2724 ;
    wire new_AGEMA_signal_2725 ;
    wire new_AGEMA_signal_2726 ;
    wire new_AGEMA_signal_2727 ;
    wire new_AGEMA_signal_2728 ;
    wire new_AGEMA_signal_2729 ;
    wire new_AGEMA_signal_2730 ;
    wire new_AGEMA_signal_2731 ;
    wire new_AGEMA_signal_2732 ;
    wire new_AGEMA_signal_2733 ;
    wire new_AGEMA_signal_2734 ;
    wire new_AGEMA_signal_2735 ;
    wire new_AGEMA_signal_2736 ;
    wire new_AGEMA_signal_2737 ;
    wire new_AGEMA_signal_2738 ;
    wire new_AGEMA_signal_2739 ;
    wire new_AGEMA_signal_2740 ;
    wire new_AGEMA_signal_2741 ;
    wire new_AGEMA_signal_2742 ;
    wire new_AGEMA_signal_2743 ;
    wire new_AGEMA_signal_2744 ;
    wire new_AGEMA_signal_2745 ;
    wire new_AGEMA_signal_2746 ;
    wire new_AGEMA_signal_2747 ;
    wire new_AGEMA_signal_2748 ;
    wire new_AGEMA_signal_2749 ;
    wire new_AGEMA_signal_2750 ;
    wire new_AGEMA_signal_2751 ;
    wire new_AGEMA_signal_2752 ;
    wire new_AGEMA_signal_2753 ;
    wire new_AGEMA_signal_2754 ;
    wire new_AGEMA_signal_2755 ;
    wire new_AGEMA_signal_2756 ;
    wire new_AGEMA_signal_2757 ;
    wire new_AGEMA_signal_2758 ;
    wire new_AGEMA_signal_2759 ;
    wire new_AGEMA_signal_2760 ;
    wire new_AGEMA_signal_2761 ;
    wire new_AGEMA_signal_2762 ;
    wire new_AGEMA_signal_2763 ;
    wire new_AGEMA_signal_2764 ;
    wire new_AGEMA_signal_2765 ;
    wire new_AGEMA_signal_2766 ;
    wire new_AGEMA_signal_2767 ;
    wire new_AGEMA_signal_2768 ;
    wire new_AGEMA_signal_2769 ;
    wire new_AGEMA_signal_2770 ;
    wire new_AGEMA_signal_2771 ;
    wire new_AGEMA_signal_2772 ;
    wire new_AGEMA_signal_2773 ;
    wire new_AGEMA_signal_2774 ;
    wire new_AGEMA_signal_2775 ;
    wire new_AGEMA_signal_2776 ;
    wire new_AGEMA_signal_2777 ;
    wire new_AGEMA_signal_2778 ;
    wire new_AGEMA_signal_2779 ;
    wire new_AGEMA_signal_2780 ;
    wire new_AGEMA_signal_2781 ;
    wire new_AGEMA_signal_2782 ;
    wire new_AGEMA_signal_2783 ;
    wire new_AGEMA_signal_2784 ;
    wire new_AGEMA_signal_2785 ;
    wire new_AGEMA_signal_2786 ;
    wire new_AGEMA_signal_2787 ;
    wire new_AGEMA_signal_2788 ;
    wire new_AGEMA_signal_2789 ;
    wire new_AGEMA_signal_2790 ;
    wire new_AGEMA_signal_2791 ;
    wire new_AGEMA_signal_2792 ;
    wire new_AGEMA_signal_2793 ;
    wire new_AGEMA_signal_2794 ;
    wire new_AGEMA_signal_2795 ;
    wire new_AGEMA_signal_2796 ;
    wire new_AGEMA_signal_2797 ;
    wire new_AGEMA_signal_2798 ;
    wire new_AGEMA_signal_2799 ;
    wire new_AGEMA_signal_2800 ;
    wire new_AGEMA_signal_2801 ;
    wire new_AGEMA_signal_2802 ;
    wire new_AGEMA_signal_2803 ;
    wire new_AGEMA_signal_2804 ;
    wire new_AGEMA_signal_2805 ;
    wire new_AGEMA_signal_2806 ;
    wire new_AGEMA_signal_2807 ;
    wire new_AGEMA_signal_2808 ;
    wire new_AGEMA_signal_2809 ;
    wire new_AGEMA_signal_2810 ;
    wire new_AGEMA_signal_2811 ;
    wire new_AGEMA_signal_2812 ;
    wire new_AGEMA_signal_2813 ;
    wire new_AGEMA_signal_2814 ;
    wire new_AGEMA_signal_2815 ;
    wire new_AGEMA_signal_2816 ;
    wire new_AGEMA_signal_2817 ;
    wire new_AGEMA_signal_2818 ;
    wire new_AGEMA_signal_2819 ;
    wire new_AGEMA_signal_2820 ;
    wire new_AGEMA_signal_2821 ;
    wire new_AGEMA_signal_2822 ;
    wire new_AGEMA_signal_2823 ;
    wire new_AGEMA_signal_2824 ;
    wire new_AGEMA_signal_2825 ;
    wire new_AGEMA_signal_2826 ;
    wire new_AGEMA_signal_2827 ;
    wire new_AGEMA_signal_2828 ;
    wire new_AGEMA_signal_2829 ;
    wire new_AGEMA_signal_2830 ;
    wire new_AGEMA_signal_2831 ;
    wire new_AGEMA_signal_2832 ;
    wire new_AGEMA_signal_2833 ;
    wire new_AGEMA_signal_2834 ;
    wire new_AGEMA_signal_2835 ;
    wire new_AGEMA_signal_2836 ;
    wire new_AGEMA_signal_2837 ;
    wire new_AGEMA_signal_2838 ;
    wire new_AGEMA_signal_2839 ;
    wire new_AGEMA_signal_2840 ;
    wire new_AGEMA_signal_2841 ;
    wire new_AGEMA_signal_2842 ;
    wire new_AGEMA_signal_2843 ;
    wire new_AGEMA_signal_2844 ;
    wire new_AGEMA_signal_2845 ;
    wire new_AGEMA_signal_2846 ;
    wire new_AGEMA_signal_2847 ;
    wire new_AGEMA_signal_2848 ;
    wire new_AGEMA_signal_2849 ;
    wire new_AGEMA_signal_2850 ;
    wire new_AGEMA_signal_2851 ;
    wire new_AGEMA_signal_2852 ;
    wire new_AGEMA_signal_2853 ;
    wire new_AGEMA_signal_2854 ;
    wire new_AGEMA_signal_2855 ;
    wire new_AGEMA_signal_2856 ;
    wire new_AGEMA_signal_2857 ;
    wire new_AGEMA_signal_2858 ;
    wire new_AGEMA_signal_2859 ;
    wire new_AGEMA_signal_2860 ;
    wire new_AGEMA_signal_2861 ;
    wire new_AGEMA_signal_2862 ;
    wire new_AGEMA_signal_2863 ;
    wire new_AGEMA_signal_2864 ;
    wire new_AGEMA_signal_2865 ;
    wire new_AGEMA_signal_2867 ;
    wire new_AGEMA_signal_2871 ;
    wire new_AGEMA_signal_2872 ;
    wire new_AGEMA_signal_2873 ;
    wire new_AGEMA_signal_2877 ;
    wire new_AGEMA_signal_2878 ;
    wire new_AGEMA_signal_2879 ;
    wire new_AGEMA_signal_2883 ;
    wire new_AGEMA_signal_2884 ;
    wire new_AGEMA_signal_2885 ;
    wire new_AGEMA_signal_2889 ;
    wire new_AGEMA_signal_2890 ;
    wire new_AGEMA_signal_2891 ;
    wire new_AGEMA_signal_2895 ;
    wire new_AGEMA_signal_2896 ;
    wire new_AGEMA_signal_2897 ;
    wire new_AGEMA_signal_2901 ;
    wire new_AGEMA_signal_2902 ;
    wire new_AGEMA_signal_2903 ;
    wire new_AGEMA_signal_2907 ;
    wire new_AGEMA_signal_2908 ;
    wire new_AGEMA_signal_2909 ;
    wire new_AGEMA_signal_2913 ;
    wire new_AGEMA_signal_2914 ;
    wire new_AGEMA_signal_2915 ;
    wire new_AGEMA_signal_2919 ;
    wire new_AGEMA_signal_2920 ;
    wire new_AGEMA_signal_2921 ;
    wire new_AGEMA_signal_2925 ;
    wire new_AGEMA_signal_2926 ;
    wire new_AGEMA_signal_2927 ;
    wire new_AGEMA_signal_2931 ;
    wire new_AGEMA_signal_2932 ;
    wire new_AGEMA_signal_2933 ;
    wire new_AGEMA_signal_2937 ;
    wire new_AGEMA_signal_2938 ;
    wire new_AGEMA_signal_2939 ;
    wire new_AGEMA_signal_2943 ;
    wire new_AGEMA_signal_2944 ;
    wire new_AGEMA_signal_2945 ;
    wire new_AGEMA_signal_2949 ;
    wire new_AGEMA_signal_2950 ;
    wire new_AGEMA_signal_2951 ;
    wire new_AGEMA_signal_2955 ;
    wire new_AGEMA_signal_2956 ;
    wire new_AGEMA_signal_2957 ;
    wire new_AGEMA_signal_2961 ;
    wire new_AGEMA_signal_2962 ;
    wire new_AGEMA_signal_2963 ;
    wire new_AGEMA_signal_2967 ;
    wire new_AGEMA_signal_2968 ;
    wire new_AGEMA_signal_2969 ;
    wire new_AGEMA_signal_2973 ;
    wire new_AGEMA_signal_2974 ;
    wire new_AGEMA_signal_2975 ;
    wire new_AGEMA_signal_2979 ;
    wire new_AGEMA_signal_2980 ;
    wire new_AGEMA_signal_2981 ;
    wire new_AGEMA_signal_2985 ;
    wire new_AGEMA_signal_2986 ;
    wire new_AGEMA_signal_2987 ;
    wire new_AGEMA_signal_2991 ;
    wire new_AGEMA_signal_2992 ;
    wire new_AGEMA_signal_2993 ;
    wire new_AGEMA_signal_2997 ;
    wire new_AGEMA_signal_2998 ;
    wire new_AGEMA_signal_2999 ;
    wire new_AGEMA_signal_3003 ;
    wire new_AGEMA_signal_3004 ;
    wire new_AGEMA_signal_3005 ;
    wire new_AGEMA_signal_3009 ;
    wire new_AGEMA_signal_3010 ;
    wire new_AGEMA_signal_3011 ;
    wire new_AGEMA_signal_3015 ;
    wire new_AGEMA_signal_3016 ;
    wire new_AGEMA_signal_3017 ;
    wire new_AGEMA_signal_3021 ;
    wire new_AGEMA_signal_3022 ;
    wire new_AGEMA_signal_3023 ;
    wire new_AGEMA_signal_3027 ;
    wire new_AGEMA_signal_3028 ;
    wire new_AGEMA_signal_3029 ;
    wire new_AGEMA_signal_3033 ;
    wire new_AGEMA_signal_3034 ;
    wire new_AGEMA_signal_3035 ;
    wire new_AGEMA_signal_3039 ;
    wire new_AGEMA_signal_3040 ;
    wire new_AGEMA_signal_3041 ;
    wire new_AGEMA_signal_3045 ;
    wire new_AGEMA_signal_3046 ;
    wire new_AGEMA_signal_3047 ;
    wire new_AGEMA_signal_3051 ;
    wire new_AGEMA_signal_3052 ;
    wire new_AGEMA_signal_3053 ;
    wire new_AGEMA_signal_3057 ;
    wire new_AGEMA_signal_3058 ;
    wire new_AGEMA_signal_3059 ;
    wire new_AGEMA_signal_3063 ;
    wire new_AGEMA_signal_3064 ;
    wire new_AGEMA_signal_3065 ;
    wire new_AGEMA_signal_3069 ;
    wire new_AGEMA_signal_3070 ;
    wire new_AGEMA_signal_3071 ;
    wire new_AGEMA_signal_3075 ;
    wire new_AGEMA_signal_3076 ;
    wire new_AGEMA_signal_3077 ;
    wire new_AGEMA_signal_3081 ;
    wire new_AGEMA_signal_3082 ;
    wire new_AGEMA_signal_3083 ;
    wire new_AGEMA_signal_3087 ;
    wire new_AGEMA_signal_3088 ;
    wire new_AGEMA_signal_3089 ;
    wire new_AGEMA_signal_3093 ;
    wire new_AGEMA_signal_3094 ;
    wire new_AGEMA_signal_3095 ;
    wire new_AGEMA_signal_3099 ;
    wire new_AGEMA_signal_3100 ;
    wire new_AGEMA_signal_3101 ;
    wire new_AGEMA_signal_3105 ;
    wire new_AGEMA_signal_3106 ;
    wire new_AGEMA_signal_3107 ;
    wire new_AGEMA_signal_3111 ;
    wire new_AGEMA_signal_3112 ;
    wire new_AGEMA_signal_3113 ;
    wire new_AGEMA_signal_3117 ;
    wire new_AGEMA_signal_3118 ;
    wire new_AGEMA_signal_3119 ;
    wire new_AGEMA_signal_3123 ;
    wire new_AGEMA_signal_3124 ;
    wire new_AGEMA_signal_3125 ;
    wire new_AGEMA_signal_3129 ;
    wire new_AGEMA_signal_3130 ;
    wire new_AGEMA_signal_3131 ;
    wire new_AGEMA_signal_3135 ;
    wire new_AGEMA_signal_3136 ;
    wire new_AGEMA_signal_3137 ;
    wire new_AGEMA_signal_3141 ;
    wire new_AGEMA_signal_3142 ;
    wire new_AGEMA_signal_3143 ;
    wire new_AGEMA_signal_3147 ;
    wire new_AGEMA_signal_3148 ;
    wire new_AGEMA_signal_3149 ;
    wire new_AGEMA_signal_3153 ;
    wire new_AGEMA_signal_3154 ;
    wire new_AGEMA_signal_3155 ;
    wire new_AGEMA_signal_3159 ;
    wire new_AGEMA_signal_3160 ;
    wire new_AGEMA_signal_3161 ;
    wire new_AGEMA_signal_3165 ;
    wire new_AGEMA_signal_3166 ;
    wire new_AGEMA_signal_3167 ;
    wire new_AGEMA_signal_3171 ;
    wire new_AGEMA_signal_3172 ;
    wire new_AGEMA_signal_3173 ;
    wire new_AGEMA_signal_3177 ;
    wire new_AGEMA_signal_3178 ;
    wire new_AGEMA_signal_3179 ;
    wire new_AGEMA_signal_3183 ;
    wire new_AGEMA_signal_3184 ;
    wire new_AGEMA_signal_3185 ;
    wire new_AGEMA_signal_3189 ;
    wire new_AGEMA_signal_3190 ;
    wire new_AGEMA_signal_3191 ;
    wire new_AGEMA_signal_3195 ;
    wire new_AGEMA_signal_3196 ;
    wire new_AGEMA_signal_3197 ;
    wire new_AGEMA_signal_3201 ;
    wire new_AGEMA_signal_3202 ;
    wire new_AGEMA_signal_3203 ;
    wire new_AGEMA_signal_3207 ;
    wire new_AGEMA_signal_3208 ;
    wire new_AGEMA_signal_3209 ;
    wire new_AGEMA_signal_3213 ;
    wire new_AGEMA_signal_3214 ;
    wire new_AGEMA_signal_3215 ;
    wire new_AGEMA_signal_3219 ;
    wire new_AGEMA_signal_3220 ;
    wire new_AGEMA_signal_3221 ;
    wire new_AGEMA_signal_3225 ;
    wire new_AGEMA_signal_3226 ;
    wire new_AGEMA_signal_3227 ;
    wire new_AGEMA_signal_3231 ;
    wire new_AGEMA_signal_3232 ;
    wire new_AGEMA_signal_3233 ;
    wire new_AGEMA_signal_3237 ;
    wire new_AGEMA_signal_3238 ;
    wire new_AGEMA_signal_3239 ;
    wire new_AGEMA_signal_3243 ;
    wire new_AGEMA_signal_3244 ;
    wire new_AGEMA_signal_3245 ;
    wire new_AGEMA_signal_3249 ;
    wire new_AGEMA_signal_3250 ;
    wire new_AGEMA_signal_3251 ;
    wire new_AGEMA_signal_3252 ;
    wire new_AGEMA_signal_3253 ;
    wire new_AGEMA_signal_3254 ;
    wire new_AGEMA_signal_3255 ;
    wire new_AGEMA_signal_3256 ;
    wire new_AGEMA_signal_3257 ;
    wire new_AGEMA_signal_3258 ;
    wire new_AGEMA_signal_3259 ;
    wire new_AGEMA_signal_3260 ;
    wire new_AGEMA_signal_3261 ;
    wire new_AGEMA_signal_3262 ;
    wire new_AGEMA_signal_3263 ;
    wire new_AGEMA_signal_3264 ;
    wire new_AGEMA_signal_3265 ;
    wire new_AGEMA_signal_3266 ;
    wire new_AGEMA_signal_3267 ;
    wire new_AGEMA_signal_3268 ;
    wire new_AGEMA_signal_3269 ;
    wire new_AGEMA_signal_3270 ;
    wire new_AGEMA_signal_3271 ;
    wire new_AGEMA_signal_3272 ;
    wire new_AGEMA_signal_3273 ;
    wire new_AGEMA_signal_3274 ;
    wire new_AGEMA_signal_3275 ;
    wire new_AGEMA_signal_3276 ;
    wire new_AGEMA_signal_3277 ;
    wire new_AGEMA_signal_3278 ;
    wire new_AGEMA_signal_3279 ;
    wire new_AGEMA_signal_3280 ;
    wire new_AGEMA_signal_3281 ;
    wire new_AGEMA_signal_3282 ;
    wire new_AGEMA_signal_3283 ;
    wire new_AGEMA_signal_3284 ;
    wire new_AGEMA_signal_3285 ;
    wire new_AGEMA_signal_3286 ;
    wire new_AGEMA_signal_3287 ;
    wire new_AGEMA_signal_3288 ;
    wire new_AGEMA_signal_3289 ;
    wire new_AGEMA_signal_3290 ;
    wire new_AGEMA_signal_3291 ;
    wire new_AGEMA_signal_3292 ;
    wire new_AGEMA_signal_3293 ;
    wire new_AGEMA_signal_3294 ;
    wire new_AGEMA_signal_3295 ;
    wire new_AGEMA_signal_3296 ;
    wire new_AGEMA_signal_3297 ;
    wire new_AGEMA_signal_3298 ;
    wire new_AGEMA_signal_3299 ;
    wire new_AGEMA_signal_3300 ;
    wire new_AGEMA_signal_3301 ;
    wire new_AGEMA_signal_3302 ;
    wire new_AGEMA_signal_3303 ;
    wire new_AGEMA_signal_3304 ;
    wire new_AGEMA_signal_3305 ;
    wire new_AGEMA_signal_3306 ;
    wire new_AGEMA_signal_3307 ;
    wire new_AGEMA_signal_3308 ;
    wire new_AGEMA_signal_3309 ;
    wire new_AGEMA_signal_3310 ;
    wire new_AGEMA_signal_3311 ;
    wire new_AGEMA_signal_3312 ;
    wire new_AGEMA_signal_3313 ;
    wire new_AGEMA_signal_3314 ;
    wire new_AGEMA_signal_3315 ;
    wire new_AGEMA_signal_3316 ;
    wire new_AGEMA_signal_3317 ;
    wire new_AGEMA_signal_3318 ;
    wire new_AGEMA_signal_3319 ;
    wire new_AGEMA_signal_3320 ;
    wire new_AGEMA_signal_3321 ;
    wire new_AGEMA_signal_3322 ;
    wire new_AGEMA_signal_3323 ;
    wire new_AGEMA_signal_3324 ;
    wire new_AGEMA_signal_3325 ;
    wire new_AGEMA_signal_3326 ;
    wire new_AGEMA_signal_3327 ;
    wire new_AGEMA_signal_3328 ;
    wire new_AGEMA_signal_3329 ;
    wire new_AGEMA_signal_3330 ;
    wire new_AGEMA_signal_3331 ;
    wire new_AGEMA_signal_3332 ;
    wire new_AGEMA_signal_3333 ;
    wire new_AGEMA_signal_3334 ;
    wire new_AGEMA_signal_3335 ;
    wire new_AGEMA_signal_3336 ;
    wire new_AGEMA_signal_3337 ;
    wire new_AGEMA_signal_3338 ;
    wire new_AGEMA_signal_3339 ;
    wire new_AGEMA_signal_3340 ;
    wire new_AGEMA_signal_3341 ;
    wire new_AGEMA_signal_3342 ;
    wire new_AGEMA_signal_3343 ;
    wire new_AGEMA_signal_3344 ;
    wire new_AGEMA_signal_3345 ;
    wire new_AGEMA_signal_3346 ;
    wire new_AGEMA_signal_3347 ;
    wire new_AGEMA_signal_3348 ;
    wire new_AGEMA_signal_3349 ;
    wire new_AGEMA_signal_3350 ;
    wire new_AGEMA_signal_3351 ;
    wire new_AGEMA_signal_3352 ;
    wire new_AGEMA_signal_3353 ;
    wire new_AGEMA_signal_3354 ;
    wire new_AGEMA_signal_3355 ;
    wire new_AGEMA_signal_3356 ;
    wire new_AGEMA_signal_3357 ;
    wire new_AGEMA_signal_3358 ;
    wire new_AGEMA_signal_3359 ;
    wire new_AGEMA_signal_3360 ;
    wire new_AGEMA_signal_3361 ;
    wire new_AGEMA_signal_3362 ;
    wire new_AGEMA_signal_3363 ;
    wire new_AGEMA_signal_3364 ;
    wire new_AGEMA_signal_3365 ;
    wire new_AGEMA_signal_3366 ;
    wire new_AGEMA_signal_3367 ;
    wire new_AGEMA_signal_3368 ;
    wire new_AGEMA_signal_3369 ;
    wire new_AGEMA_signal_3370 ;
    wire new_AGEMA_signal_3371 ;
    wire new_AGEMA_signal_3372 ;
    wire new_AGEMA_signal_3373 ;
    wire new_AGEMA_signal_3374 ;
    wire new_AGEMA_signal_3375 ;
    wire new_AGEMA_signal_3376 ;
    wire new_AGEMA_signal_3377 ;
    wire new_AGEMA_signal_3378 ;
    wire new_AGEMA_signal_3379 ;
    wire new_AGEMA_signal_3380 ;
    wire new_AGEMA_signal_3381 ;
    wire new_AGEMA_signal_3382 ;
    wire new_AGEMA_signal_3383 ;
    wire new_AGEMA_signal_3384 ;
    wire new_AGEMA_signal_3385 ;
    wire new_AGEMA_signal_3386 ;
    wire new_AGEMA_signal_3387 ;
    wire new_AGEMA_signal_3388 ;
    wire new_AGEMA_signal_3389 ;
    wire new_AGEMA_signal_3390 ;
    wire new_AGEMA_signal_3391 ;
    wire new_AGEMA_signal_3392 ;
    wire new_AGEMA_signal_3393 ;
    wire new_AGEMA_signal_3394 ;
    wire new_AGEMA_signal_3395 ;
    wire new_AGEMA_signal_3396 ;
    wire new_AGEMA_signal_3397 ;
    wire new_AGEMA_signal_3398 ;
    wire new_AGEMA_signal_3399 ;
    wire new_AGEMA_signal_3400 ;
    wire new_AGEMA_signal_3401 ;
    wire new_AGEMA_signal_3402 ;
    wire new_AGEMA_signal_3403 ;
    wire new_AGEMA_signal_3404 ;
    wire new_AGEMA_signal_3405 ;
    wire new_AGEMA_signal_3406 ;
    wire new_AGEMA_signal_3407 ;
    wire new_AGEMA_signal_3408 ;
    wire new_AGEMA_signal_3409 ;
    wire new_AGEMA_signal_3410 ;
    wire new_AGEMA_signal_3411 ;
    wire new_AGEMA_signal_3412 ;
    wire new_AGEMA_signal_3413 ;
    wire new_AGEMA_signal_3414 ;
    wire new_AGEMA_signal_3415 ;
    wire new_AGEMA_signal_3416 ;
    wire new_AGEMA_signal_3417 ;
    wire new_AGEMA_signal_3418 ;
    wire new_AGEMA_signal_3419 ;
    wire new_AGEMA_signal_3420 ;
    wire new_AGEMA_signal_3421 ;
    wire new_AGEMA_signal_3422 ;
    wire new_AGEMA_signal_3423 ;
    wire new_AGEMA_signal_3424 ;
    wire new_AGEMA_signal_3425 ;
    wire new_AGEMA_signal_3426 ;
    wire new_AGEMA_signal_3427 ;
    wire new_AGEMA_signal_3428 ;
    wire new_AGEMA_signal_3429 ;
    wire new_AGEMA_signal_3430 ;
    wire new_AGEMA_signal_3431 ;
    wire new_AGEMA_signal_3432 ;
    wire new_AGEMA_signal_3433 ;
    wire new_AGEMA_signal_3434 ;
    wire new_AGEMA_signal_3435 ;
    wire new_AGEMA_signal_3436 ;
    wire new_AGEMA_signal_3437 ;
    wire new_AGEMA_signal_3438 ;
    wire new_AGEMA_signal_3439 ;
    wire new_AGEMA_signal_3440 ;
    wire new_AGEMA_signal_3441 ;
    wire new_AGEMA_signal_3442 ;
    wire new_AGEMA_signal_3443 ;
    wire new_AGEMA_signal_3444 ;
    wire new_AGEMA_signal_3445 ;
    wire new_AGEMA_signal_3446 ;
    wire new_AGEMA_signal_3447 ;
    wire new_AGEMA_signal_3448 ;
    wire new_AGEMA_signal_3449 ;
    wire new_AGEMA_signal_3450 ;
    wire new_AGEMA_signal_3451 ;
    wire new_AGEMA_signal_3452 ;
    wire new_AGEMA_signal_3453 ;
    wire new_AGEMA_signal_3454 ;
    wire new_AGEMA_signal_3455 ;
    wire new_AGEMA_signal_3456 ;
    wire new_AGEMA_signal_3457 ;
    wire new_AGEMA_signal_3458 ;
    wire new_AGEMA_signal_3459 ;
    wire new_AGEMA_signal_3460 ;
    wire new_AGEMA_signal_3461 ;
    wire new_AGEMA_signal_3462 ;
    wire new_AGEMA_signal_3463 ;
    wire new_AGEMA_signal_3464 ;
    wire new_AGEMA_signal_3465 ;
    wire new_AGEMA_signal_3466 ;
    wire new_AGEMA_signal_3467 ;
    wire new_AGEMA_signal_3468 ;
    wire new_AGEMA_signal_3469 ;
    wire new_AGEMA_signal_3470 ;
    wire new_AGEMA_signal_3471 ;
    wire new_AGEMA_signal_3472 ;
    wire new_AGEMA_signal_3473 ;
    wire new_AGEMA_signal_3474 ;
    wire new_AGEMA_signal_3475 ;
    wire new_AGEMA_signal_3476 ;
    wire new_AGEMA_signal_3477 ;
    wire new_AGEMA_signal_3478 ;
    wire new_AGEMA_signal_3479 ;
    wire new_AGEMA_signal_3480 ;
    wire new_AGEMA_signal_3481 ;
    wire new_AGEMA_signal_3482 ;
    wire new_AGEMA_signal_3483 ;
    wire new_AGEMA_signal_3484 ;
    wire new_AGEMA_signal_3485 ;
    wire new_AGEMA_signal_3486 ;
    wire new_AGEMA_signal_3487 ;
    wire new_AGEMA_signal_3488 ;
    wire new_AGEMA_signal_3489 ;
    wire new_AGEMA_signal_3490 ;
    wire new_AGEMA_signal_3491 ;
    wire new_AGEMA_signal_3492 ;
    wire new_AGEMA_signal_3493 ;
    wire new_AGEMA_signal_3494 ;
    wire new_AGEMA_signal_3495 ;
    wire new_AGEMA_signal_3496 ;
    wire new_AGEMA_signal_3497 ;
    wire new_AGEMA_signal_3498 ;
    wire new_AGEMA_signal_3499 ;
    wire new_AGEMA_signal_3500 ;
    wire new_AGEMA_signal_3501 ;
    wire new_AGEMA_signal_3502 ;
    wire new_AGEMA_signal_3503 ;
    wire new_AGEMA_signal_3504 ;
    wire new_AGEMA_signal_3505 ;
    wire new_AGEMA_signal_3506 ;
    wire new_AGEMA_signal_3507 ;
    wire new_AGEMA_signal_3508 ;
    wire new_AGEMA_signal_3509 ;
    wire new_AGEMA_signal_3510 ;
    wire new_AGEMA_signal_3511 ;
    wire new_AGEMA_signal_3512 ;
    wire new_AGEMA_signal_3513 ;
    wire new_AGEMA_signal_3514 ;
    wire new_AGEMA_signal_3515 ;
    wire new_AGEMA_signal_3516 ;
    wire new_AGEMA_signal_3517 ;
    wire new_AGEMA_signal_3518 ;
    wire new_AGEMA_signal_3519 ;
    wire new_AGEMA_signal_3520 ;
    wire new_AGEMA_signal_3521 ;
    wire new_AGEMA_signal_3522 ;
    wire new_AGEMA_signal_3523 ;
    wire new_AGEMA_signal_3524 ;
    wire new_AGEMA_signal_3525 ;
    wire new_AGEMA_signal_3526 ;
    wire new_AGEMA_signal_3527 ;
    wire new_AGEMA_signal_3528 ;
    wire new_AGEMA_signal_3529 ;
    wire new_AGEMA_signal_3530 ;
    wire new_AGEMA_signal_3531 ;
    wire new_AGEMA_signal_3532 ;
    wire new_AGEMA_signal_3533 ;
    wire new_AGEMA_signal_3534 ;
    wire new_AGEMA_signal_3535 ;
    wire new_AGEMA_signal_3536 ;
    wire new_AGEMA_signal_3537 ;
    wire new_AGEMA_signal_3538 ;
    wire new_AGEMA_signal_3539 ;
    wire new_AGEMA_signal_3540 ;
    wire new_AGEMA_signal_3541 ;
    wire new_AGEMA_signal_3542 ;
    wire new_AGEMA_signal_3543 ;
    wire new_AGEMA_signal_3544 ;
    wire new_AGEMA_signal_3545 ;
    wire new_AGEMA_signal_3546 ;
    wire new_AGEMA_signal_3547 ;
    wire new_AGEMA_signal_3548 ;
    wire new_AGEMA_signal_3549 ;
    wire new_AGEMA_signal_3550 ;
    wire new_AGEMA_signal_3551 ;
    wire new_AGEMA_signal_3552 ;
    wire new_AGEMA_signal_3553 ;
    wire new_AGEMA_signal_3554 ;
    wire new_AGEMA_signal_3555 ;
    wire new_AGEMA_signal_3556 ;
    wire new_AGEMA_signal_3557 ;
    wire new_AGEMA_signal_3558 ;
    wire new_AGEMA_signal_3559 ;
    wire new_AGEMA_signal_3560 ;
    wire new_AGEMA_signal_3561 ;
    wire new_AGEMA_signal_3562 ;
    wire new_AGEMA_signal_3563 ;
    wire new_AGEMA_signal_3564 ;
    wire new_AGEMA_signal_3565 ;
    wire new_AGEMA_signal_3566 ;
    wire new_AGEMA_signal_3567 ;
    wire new_AGEMA_signal_3568 ;
    wire new_AGEMA_signal_3569 ;
    wire new_AGEMA_signal_3570 ;
    wire new_AGEMA_signal_3571 ;
    wire new_AGEMA_signal_3572 ;
    wire new_AGEMA_signal_3573 ;
    wire new_AGEMA_signal_3574 ;
    wire new_AGEMA_signal_3575 ;
    wire new_AGEMA_signal_3576 ;
    wire new_AGEMA_signal_3577 ;
    wire new_AGEMA_signal_3578 ;
    wire new_AGEMA_signal_3579 ;
    wire new_AGEMA_signal_3580 ;
    wire new_AGEMA_signal_3581 ;
    wire new_AGEMA_signal_3582 ;
    wire new_AGEMA_signal_3583 ;
    wire new_AGEMA_signal_3584 ;
    wire new_AGEMA_signal_3585 ;
    wire new_AGEMA_signal_3586 ;
    wire new_AGEMA_signal_3587 ;
    wire new_AGEMA_signal_3588 ;
    wire new_AGEMA_signal_3589 ;
    wire new_AGEMA_signal_3590 ;
    wire new_AGEMA_signal_3591 ;
    wire new_AGEMA_signal_3592 ;
    wire new_AGEMA_signal_3593 ;
    wire new_AGEMA_signal_3594 ;
    wire new_AGEMA_signal_3595 ;
    wire new_AGEMA_signal_3596 ;
    wire new_AGEMA_signal_3597 ;
    wire new_AGEMA_signal_3598 ;
    wire new_AGEMA_signal_3599 ;
    wire new_AGEMA_signal_3600 ;
    wire new_AGEMA_signal_3601 ;
    wire new_AGEMA_signal_3602 ;
    wire new_AGEMA_signal_3603 ;
    wire new_AGEMA_signal_3604 ;
    wire new_AGEMA_signal_3605 ;
    wire new_AGEMA_signal_3606 ;
    wire new_AGEMA_signal_3607 ;
    wire new_AGEMA_signal_3608 ;
    wire new_AGEMA_signal_3609 ;
    wire new_AGEMA_signal_3610 ;
    wire new_AGEMA_signal_3611 ;
    wire new_AGEMA_signal_3612 ;
    wire new_AGEMA_signal_3613 ;
    wire new_AGEMA_signal_3614 ;
    wire new_AGEMA_signal_3615 ;
    wire new_AGEMA_signal_3616 ;
    wire new_AGEMA_signal_3617 ;
    wire new_AGEMA_signal_3618 ;
    wire new_AGEMA_signal_3619 ;
    wire new_AGEMA_signal_3620 ;
    wire new_AGEMA_signal_3621 ;
    wire new_AGEMA_signal_3622 ;
    wire new_AGEMA_signal_3623 ;
    wire new_AGEMA_signal_3624 ;
    wire new_AGEMA_signal_3625 ;
    wire new_AGEMA_signal_3626 ;
    wire new_AGEMA_signal_3627 ;
    wire new_AGEMA_signal_3628 ;
    wire new_AGEMA_signal_3629 ;
    wire new_AGEMA_signal_3630 ;
    wire new_AGEMA_signal_3631 ;
    wire new_AGEMA_signal_3632 ;
    wire new_AGEMA_signal_3633 ;
    wire new_AGEMA_signal_3634 ;
    wire new_AGEMA_signal_3635 ;
    wire new_AGEMA_signal_3636 ;
    wire new_AGEMA_signal_3637 ;
    wire new_AGEMA_signal_3638 ;
    wire new_AGEMA_signal_3639 ;
    wire new_AGEMA_signal_3640 ;
    wire new_AGEMA_signal_3641 ;
    wire new_AGEMA_signal_3642 ;
    wire new_AGEMA_signal_3643 ;
    wire new_AGEMA_signal_3644 ;
    wire new_AGEMA_signal_3645 ;
    wire new_AGEMA_signal_3646 ;
    wire new_AGEMA_signal_3647 ;
    wire new_AGEMA_signal_3648 ;
    wire new_AGEMA_signal_3649 ;
    wire new_AGEMA_signal_3650 ;
    wire new_AGEMA_signal_3651 ;
    wire new_AGEMA_signal_3652 ;
    wire new_AGEMA_signal_3653 ;
    wire new_AGEMA_signal_3654 ;
    wire new_AGEMA_signal_3655 ;
    wire new_AGEMA_signal_3656 ;
    wire new_AGEMA_signal_3657 ;
    wire new_AGEMA_signal_3658 ;
    wire new_AGEMA_signal_3659 ;
    wire new_AGEMA_signal_3660 ;
    wire new_AGEMA_signal_3661 ;
    wire new_AGEMA_signal_3662 ;
    wire new_AGEMA_signal_3663 ;
    wire new_AGEMA_signal_3664 ;
    wire new_AGEMA_signal_3665 ;
    wire new_AGEMA_signal_3666 ;
    wire new_AGEMA_signal_3667 ;
    wire new_AGEMA_signal_3668 ;
    wire new_AGEMA_signal_3669 ;
    wire new_AGEMA_signal_3670 ;
    wire new_AGEMA_signal_3671 ;
    wire new_AGEMA_signal_3672 ;
    wire new_AGEMA_signal_3673 ;
    wire new_AGEMA_signal_3674 ;
    wire new_AGEMA_signal_3675 ;
    wire new_AGEMA_signal_3676 ;
    wire new_AGEMA_signal_3677 ;
    wire new_AGEMA_signal_3678 ;
    wire new_AGEMA_signal_3679 ;
    wire new_AGEMA_signal_3680 ;
    wire new_AGEMA_signal_3681 ;
    wire new_AGEMA_signal_3682 ;
    wire new_AGEMA_signal_3683 ;
    wire new_AGEMA_signal_3684 ;
    wire new_AGEMA_signal_3685 ;
    wire new_AGEMA_signal_3686 ;
    wire new_AGEMA_signal_3687 ;
    wire new_AGEMA_signal_3688 ;
    wire new_AGEMA_signal_3689 ;
    wire new_AGEMA_signal_3690 ;
    wire new_AGEMA_signal_3691 ;
    wire new_AGEMA_signal_3692 ;
    wire new_AGEMA_signal_3693 ;
    wire new_AGEMA_signal_3694 ;
    wire new_AGEMA_signal_3695 ;
    wire new_AGEMA_signal_3696 ;
    wire new_AGEMA_signal_3697 ;
    wire new_AGEMA_signal_3698 ;
    wire new_AGEMA_signal_3699 ;
    wire new_AGEMA_signal_3700 ;
    wire new_AGEMA_signal_3701 ;
    wire new_AGEMA_signal_3702 ;
    wire new_AGEMA_signal_3703 ;
    wire new_AGEMA_signal_3704 ;
    wire new_AGEMA_signal_3705 ;
    wire new_AGEMA_signal_3706 ;
    wire new_AGEMA_signal_3707 ;
    wire new_AGEMA_signal_3708 ;
    wire new_AGEMA_signal_3709 ;
    wire new_AGEMA_signal_3710 ;
    wire new_AGEMA_signal_3711 ;
    wire new_AGEMA_signal_3712 ;
    wire new_AGEMA_signal_3713 ;
    wire new_AGEMA_signal_3714 ;
    wire new_AGEMA_signal_3715 ;
    wire new_AGEMA_signal_3716 ;
    wire new_AGEMA_signal_3717 ;
    wire new_AGEMA_signal_3718 ;
    wire new_AGEMA_signal_3719 ;
    wire new_AGEMA_signal_3720 ;
    wire new_AGEMA_signal_3721 ;
    wire new_AGEMA_signal_3722 ;
    wire new_AGEMA_signal_3723 ;
    wire new_AGEMA_signal_3724 ;
    wire new_AGEMA_signal_3725 ;
    wire new_AGEMA_signal_3726 ;
    wire new_AGEMA_signal_3727 ;
    wire new_AGEMA_signal_3728 ;
    wire new_AGEMA_signal_3729 ;
    wire new_AGEMA_signal_3730 ;
    wire new_AGEMA_signal_3731 ;
    wire new_AGEMA_signal_3732 ;
    wire new_AGEMA_signal_3733 ;
    wire new_AGEMA_signal_3734 ;
    wire new_AGEMA_signal_3735 ;
    wire new_AGEMA_signal_3736 ;
    wire new_AGEMA_signal_3737 ;
    wire new_AGEMA_signal_3738 ;
    wire new_AGEMA_signal_3739 ;
    wire new_AGEMA_signal_3740 ;
    wire new_AGEMA_signal_3741 ;
    wire new_AGEMA_signal_3742 ;
    wire new_AGEMA_signal_3743 ;
    wire new_AGEMA_signal_3744 ;
    wire new_AGEMA_signal_3745 ;
    wire new_AGEMA_signal_3746 ;
    wire new_AGEMA_signal_3747 ;
    wire new_AGEMA_signal_3748 ;
    wire new_AGEMA_signal_3749 ;
    wire new_AGEMA_signal_3750 ;
    wire new_AGEMA_signal_3751 ;
    wire new_AGEMA_signal_3752 ;
    wire new_AGEMA_signal_3753 ;
    wire new_AGEMA_signal_3754 ;
    wire new_AGEMA_signal_3755 ;
    wire new_AGEMA_signal_3756 ;
    wire new_AGEMA_signal_3757 ;
    wire new_AGEMA_signal_3758 ;
    wire new_AGEMA_signal_3759 ;
    wire new_AGEMA_signal_3760 ;
    wire new_AGEMA_signal_3761 ;
    wire new_AGEMA_signal_3762 ;
    wire new_AGEMA_signal_3763 ;
    wire new_AGEMA_signal_3764 ;
    wire new_AGEMA_signal_3765 ;
    wire new_AGEMA_signal_3766 ;
    wire new_AGEMA_signal_3767 ;
    wire new_AGEMA_signal_3768 ;
    wire new_AGEMA_signal_3769 ;
    wire new_AGEMA_signal_3770 ;
    wire new_AGEMA_signal_3771 ;
    wire new_AGEMA_signal_3772 ;
    wire new_AGEMA_signal_3773 ;
    wire new_AGEMA_signal_3774 ;
    wire new_AGEMA_signal_3775 ;
    wire new_AGEMA_signal_3776 ;
    wire new_AGEMA_signal_3777 ;
    wire new_AGEMA_signal_3778 ;
    wire new_AGEMA_signal_3779 ;
    wire new_AGEMA_signal_3780 ;
    wire new_AGEMA_signal_3781 ;
    wire new_AGEMA_signal_3782 ;
    wire new_AGEMA_signal_3783 ;
    wire new_AGEMA_signal_3784 ;
    wire new_AGEMA_signal_3785 ;
    wire new_AGEMA_signal_3786 ;
    wire new_AGEMA_signal_3787 ;
    wire new_AGEMA_signal_3788 ;
    wire new_AGEMA_signal_3789 ;
    wire new_AGEMA_signal_3790 ;
    wire new_AGEMA_signal_3791 ;
    wire new_AGEMA_signal_3792 ;
    wire new_AGEMA_signal_3793 ;
    wire new_AGEMA_signal_3794 ;
    wire new_AGEMA_signal_3795 ;
    wire new_AGEMA_signal_3796 ;
    wire new_AGEMA_signal_3797 ;
    wire new_AGEMA_signal_3798 ;
    wire new_AGEMA_signal_3799 ;
    wire new_AGEMA_signal_3800 ;
    wire new_AGEMA_signal_3801 ;
    wire new_AGEMA_signal_3802 ;
    wire new_AGEMA_signal_3803 ;
    wire new_AGEMA_signal_3804 ;
    wire new_AGEMA_signal_3805 ;
    wire new_AGEMA_signal_3806 ;
    wire new_AGEMA_signal_3807 ;
    wire new_AGEMA_signal_3808 ;
    wire new_AGEMA_signal_3809 ;
    wire new_AGEMA_signal_3810 ;
    wire new_AGEMA_signal_3811 ;
    wire new_AGEMA_signal_3812 ;
    wire new_AGEMA_signal_3813 ;
    wire new_AGEMA_signal_3814 ;
    wire new_AGEMA_signal_3815 ;
    wire new_AGEMA_signal_3816 ;
    wire new_AGEMA_signal_3817 ;
    wire new_AGEMA_signal_3818 ;
    wire new_AGEMA_signal_3819 ;
    wire new_AGEMA_signal_3820 ;
    wire new_AGEMA_signal_3821 ;
    wire new_AGEMA_signal_3822 ;
    wire new_AGEMA_signal_3823 ;
    wire new_AGEMA_signal_3824 ;
    wire new_AGEMA_signal_3825 ;
    wire new_AGEMA_signal_3826 ;
    wire new_AGEMA_signal_3827 ;
    wire new_AGEMA_signal_3828 ;
    wire new_AGEMA_signal_3829 ;
    wire new_AGEMA_signal_3830 ;
    wire new_AGEMA_signal_3831 ;
    wire new_AGEMA_signal_3832 ;
    wire new_AGEMA_signal_3833 ;
    wire new_AGEMA_signal_3834 ;
    wire new_AGEMA_signal_3835 ;
    wire new_AGEMA_signal_3836 ;
    wire new_AGEMA_signal_3837 ;
    wire new_AGEMA_signal_3838 ;
    wire new_AGEMA_signal_3839 ;
    wire new_AGEMA_signal_3840 ;
    wire new_AGEMA_signal_3841 ;
    wire new_AGEMA_signal_3842 ;
    wire new_AGEMA_signal_3843 ;
    wire new_AGEMA_signal_3844 ;
    wire new_AGEMA_signal_3845 ;
    wire new_AGEMA_signal_3846 ;
    wire new_AGEMA_signal_3847 ;
    wire new_AGEMA_signal_3848 ;
    wire new_AGEMA_signal_3849 ;
    wire new_AGEMA_signal_3850 ;
    wire new_AGEMA_signal_3851 ;
    wire new_AGEMA_signal_3852 ;
    wire new_AGEMA_signal_3853 ;
    wire new_AGEMA_signal_3854 ;
    wire new_AGEMA_signal_3855 ;
    wire new_AGEMA_signal_3856 ;
    wire new_AGEMA_signal_3857 ;
    wire new_AGEMA_signal_3858 ;
    wire new_AGEMA_signal_3859 ;
    wire new_AGEMA_signal_3860 ;
    wire new_AGEMA_signal_3861 ;
    wire new_AGEMA_signal_3862 ;
    wire new_AGEMA_signal_3863 ;
    wire new_AGEMA_signal_3864 ;
    wire new_AGEMA_signal_3865 ;
    wire new_AGEMA_signal_3866 ;
    wire new_AGEMA_signal_3867 ;
    wire new_AGEMA_signal_3868 ;
    wire new_AGEMA_signal_3869 ;
    wire new_AGEMA_signal_3870 ;
    wire new_AGEMA_signal_3871 ;
    wire new_AGEMA_signal_3872 ;
    wire new_AGEMA_signal_3873 ;
    wire new_AGEMA_signal_3874 ;
    wire new_AGEMA_signal_3875 ;
    wire new_AGEMA_signal_3876 ;
    wire new_AGEMA_signal_3877 ;
    wire new_AGEMA_signal_3878 ;
    wire new_AGEMA_signal_3879 ;
    wire new_AGEMA_signal_3880 ;
    wire new_AGEMA_signal_3881 ;
    wire new_AGEMA_signal_3882 ;
    wire new_AGEMA_signal_3883 ;
    wire new_AGEMA_signal_3884 ;
    wire new_AGEMA_signal_3885 ;
    wire new_AGEMA_signal_3886 ;
    wire new_AGEMA_signal_3887 ;
    wire new_AGEMA_signal_3888 ;
    wire new_AGEMA_signal_3889 ;
    wire new_AGEMA_signal_3890 ;
    wire new_AGEMA_signal_3891 ;
    wire new_AGEMA_signal_3892 ;
    wire new_AGEMA_signal_3893 ;
    wire new_AGEMA_signal_3894 ;
    wire new_AGEMA_signal_3895 ;
    wire new_AGEMA_signal_3896 ;
    wire new_AGEMA_signal_3897 ;
    wire new_AGEMA_signal_3898 ;
    wire new_AGEMA_signal_3899 ;
    wire new_AGEMA_signal_3900 ;
    wire new_AGEMA_signal_3901 ;
    wire new_AGEMA_signal_3902 ;
    wire new_AGEMA_signal_3903 ;
    wire new_AGEMA_signal_3904 ;
    wire new_AGEMA_signal_3905 ;
    wire new_AGEMA_signal_3906 ;
    wire new_AGEMA_signal_3907 ;
    wire new_AGEMA_signal_3908 ;
    wire new_AGEMA_signal_3909 ;
    wire new_AGEMA_signal_3910 ;
    wire new_AGEMA_signal_3911 ;
    wire new_AGEMA_signal_3912 ;
    wire new_AGEMA_signal_3913 ;
    wire new_AGEMA_signal_3914 ;
    wire new_AGEMA_signal_3915 ;
    wire new_AGEMA_signal_3916 ;
    wire new_AGEMA_signal_3917 ;
    wire new_AGEMA_signal_3918 ;
    wire new_AGEMA_signal_3919 ;
    wire new_AGEMA_signal_3920 ;
    wire new_AGEMA_signal_3921 ;
    wire new_AGEMA_signal_3922 ;
    wire new_AGEMA_signal_3923 ;
    wire new_AGEMA_signal_3924 ;
    wire new_AGEMA_signal_3925 ;
    wire new_AGEMA_signal_3926 ;
    wire new_AGEMA_signal_3927 ;
    wire new_AGEMA_signal_3928 ;
    wire new_AGEMA_signal_3929 ;
    wire new_AGEMA_signal_3930 ;
    wire new_AGEMA_signal_3931 ;
    wire new_AGEMA_signal_3932 ;
    wire new_AGEMA_signal_3933 ;
    wire new_AGEMA_signal_3934 ;
    wire new_AGEMA_signal_3935 ;
    wire new_AGEMA_signal_3936 ;
    wire new_AGEMA_signal_3937 ;
    wire new_AGEMA_signal_3938 ;
    wire new_AGEMA_signal_3939 ;
    wire new_AGEMA_signal_3940 ;
    wire new_AGEMA_signal_3941 ;
    wire new_AGEMA_signal_3942 ;
    wire new_AGEMA_signal_3943 ;
    wire new_AGEMA_signal_3944 ;
    wire new_AGEMA_signal_3945 ;
    wire new_AGEMA_signal_3946 ;
    wire new_AGEMA_signal_3947 ;
    wire new_AGEMA_signal_3948 ;
    wire new_AGEMA_signal_3949 ;
    wire new_AGEMA_signal_3950 ;
    wire new_AGEMA_signal_3951 ;
    wire new_AGEMA_signal_3952 ;
    wire new_AGEMA_signal_3953 ;
    wire new_AGEMA_signal_3954 ;
    wire new_AGEMA_signal_3955 ;
    wire new_AGEMA_signal_3956 ;
    wire new_AGEMA_signal_3957 ;
    wire new_AGEMA_signal_3958 ;
    wire new_AGEMA_signal_3959 ;
    wire new_AGEMA_signal_3960 ;
    wire new_AGEMA_signal_3961 ;
    wire new_AGEMA_signal_3962 ;
    wire new_AGEMA_signal_3963 ;
    wire new_AGEMA_signal_3964 ;
    wire new_AGEMA_signal_3965 ;
    wire new_AGEMA_signal_3966 ;
    wire new_AGEMA_signal_3967 ;
    wire new_AGEMA_signal_3968 ;
    wire new_AGEMA_signal_3969 ;
    wire new_AGEMA_signal_3970 ;
    wire new_AGEMA_signal_3971 ;
    wire new_AGEMA_signal_3972 ;
    wire new_AGEMA_signal_3973 ;
    wire new_AGEMA_signal_3974 ;
    wire new_AGEMA_signal_3975 ;
    wire new_AGEMA_signal_3976 ;
    wire new_AGEMA_signal_3977 ;
    wire new_AGEMA_signal_3978 ;
    wire new_AGEMA_signal_3979 ;
    wire new_AGEMA_signal_3980 ;
    wire new_AGEMA_signal_3981 ;
    wire new_AGEMA_signal_3982 ;
    wire new_AGEMA_signal_3983 ;
    wire new_AGEMA_signal_3984 ;
    wire new_AGEMA_signal_3985 ;
    wire new_AGEMA_signal_3986 ;
    wire new_AGEMA_signal_3987 ;
    wire new_AGEMA_signal_3988 ;
    wire new_AGEMA_signal_3989 ;
    wire new_AGEMA_signal_3990 ;
    wire new_AGEMA_signal_3991 ;
    wire new_AGEMA_signal_3992 ;
    wire new_AGEMA_signal_3993 ;
    wire new_AGEMA_signal_3994 ;
    wire new_AGEMA_signal_3995 ;
    wire new_AGEMA_signal_3996 ;
    wire new_AGEMA_signal_3997 ;
    wire new_AGEMA_signal_3998 ;
    wire new_AGEMA_signal_3999 ;
    wire new_AGEMA_signal_4000 ;
    wire new_AGEMA_signal_4001 ;
    wire new_AGEMA_signal_4002 ;
    wire new_AGEMA_signal_4003 ;
    wire new_AGEMA_signal_4004 ;
    wire new_AGEMA_signal_4005 ;
    wire new_AGEMA_signal_4006 ;
    wire new_AGEMA_signal_4007 ;
    wire new_AGEMA_signal_4008 ;
    wire new_AGEMA_signal_4009 ;
    wire new_AGEMA_signal_4010 ;
    wire new_AGEMA_signal_4011 ;
    wire new_AGEMA_signal_4012 ;
    wire new_AGEMA_signal_4013 ;
    wire new_AGEMA_signal_4014 ;
    wire new_AGEMA_signal_4015 ;
    wire new_AGEMA_signal_4016 ;
    wire new_AGEMA_signal_4017 ;
    wire new_AGEMA_signal_4018 ;
    wire new_AGEMA_signal_4019 ;
    wire new_AGEMA_signal_4020 ;
    wire new_AGEMA_signal_4021 ;
    wire new_AGEMA_signal_4022 ;
    wire new_AGEMA_signal_4023 ;
    wire new_AGEMA_signal_4024 ;
    wire new_AGEMA_signal_4025 ;
    wire new_AGEMA_signal_4026 ;
    wire new_AGEMA_signal_4027 ;
    wire new_AGEMA_signal_4028 ;
    wire new_AGEMA_signal_4029 ;
    wire new_AGEMA_signal_4030 ;
    wire new_AGEMA_signal_4031 ;
    wire new_AGEMA_signal_4032 ;
    wire new_AGEMA_signal_4033 ;
    wire new_AGEMA_signal_4034 ;
    wire new_AGEMA_signal_4035 ;
    wire new_AGEMA_signal_4036 ;
    wire new_AGEMA_signal_4037 ;
    wire new_AGEMA_signal_4038 ;
    wire new_AGEMA_signal_4039 ;
    wire new_AGEMA_signal_4040 ;
    wire new_AGEMA_signal_4041 ;
    wire new_AGEMA_signal_4042 ;
    wire new_AGEMA_signal_4043 ;
    wire new_AGEMA_signal_4044 ;
    wire new_AGEMA_signal_4045 ;
    wire new_AGEMA_signal_4046 ;
    wire new_AGEMA_signal_4047 ;
    wire new_AGEMA_signal_4048 ;
    wire new_AGEMA_signal_4049 ;
    wire new_AGEMA_signal_4050 ;
    wire new_AGEMA_signal_4051 ;
    wire new_AGEMA_signal_4052 ;
    wire new_AGEMA_signal_4053 ;
    wire new_AGEMA_signal_4054 ;
    wire new_AGEMA_signal_4055 ;
    wire new_AGEMA_signal_4056 ;
    wire new_AGEMA_signal_4057 ;
    wire new_AGEMA_signal_4058 ;
    wire new_AGEMA_signal_4059 ;
    wire new_AGEMA_signal_4060 ;
    wire new_AGEMA_signal_4061 ;
    wire new_AGEMA_signal_4062 ;
    wire new_AGEMA_signal_4063 ;
    wire new_AGEMA_signal_4064 ;
    wire new_AGEMA_signal_4065 ;
    wire new_AGEMA_signal_4066 ;
    wire new_AGEMA_signal_4067 ;
    wire new_AGEMA_signal_4068 ;
    wire new_AGEMA_signal_4069 ;
    wire new_AGEMA_signal_4070 ;
    wire new_AGEMA_signal_4071 ;
    wire new_AGEMA_signal_4072 ;
    wire new_AGEMA_signal_4073 ;
    wire new_AGEMA_signal_4074 ;
    wire new_AGEMA_signal_4075 ;
    wire new_AGEMA_signal_4076 ;
    wire new_AGEMA_signal_4077 ;
    wire new_AGEMA_signal_4078 ;
    wire new_AGEMA_signal_4079 ;
    wire new_AGEMA_signal_4080 ;
    wire new_AGEMA_signal_4081 ;
    wire new_AGEMA_signal_4082 ;
    wire new_AGEMA_signal_4083 ;
    wire new_AGEMA_signal_4084 ;
    wire new_AGEMA_signal_4085 ;
    wire new_AGEMA_signal_4086 ;
    wire new_AGEMA_signal_4087 ;
    wire new_AGEMA_signal_4088 ;
    wire new_AGEMA_signal_4089 ;
    wire new_AGEMA_signal_4090 ;
    wire new_AGEMA_signal_4091 ;
    wire new_AGEMA_signal_4092 ;
    wire new_AGEMA_signal_4093 ;
    wire new_AGEMA_signal_4094 ;
    wire new_AGEMA_signal_4095 ;
    wire new_AGEMA_signal_4096 ;
    wire new_AGEMA_signal_4097 ;
    wire new_AGEMA_signal_4098 ;
    wire new_AGEMA_signal_4099 ;
    wire new_AGEMA_signal_4100 ;
    wire new_AGEMA_signal_4101 ;
    wire new_AGEMA_signal_4102 ;
    wire new_AGEMA_signal_4103 ;
    wire new_AGEMA_signal_4104 ;
    wire new_AGEMA_signal_4105 ;
    wire new_AGEMA_signal_4106 ;
    wire new_AGEMA_signal_4107 ;
    wire new_AGEMA_signal_4108 ;
    wire new_AGEMA_signal_4109 ;
    wire new_AGEMA_signal_4110 ;
    wire new_AGEMA_signal_4111 ;
    wire new_AGEMA_signal_4112 ;
    wire new_AGEMA_signal_4113 ;
    wire new_AGEMA_signal_4114 ;
    wire new_AGEMA_signal_4115 ;
    wire new_AGEMA_signal_4116 ;
    wire new_AGEMA_signal_4117 ;
    wire new_AGEMA_signal_4118 ;
    wire new_AGEMA_signal_4119 ;
    wire new_AGEMA_signal_4120 ;
    wire new_AGEMA_signal_4121 ;
    wire new_AGEMA_signal_4122 ;
    wire new_AGEMA_signal_4123 ;
    wire new_AGEMA_signal_4124 ;
    wire new_AGEMA_signal_4125 ;
    wire new_AGEMA_signal_4126 ;
    wire new_AGEMA_signal_4127 ;
    wire new_AGEMA_signal_4128 ;
    wire new_AGEMA_signal_4129 ;
    wire new_AGEMA_signal_4130 ;
    wire new_AGEMA_signal_4131 ;
    wire new_AGEMA_signal_4132 ;
    wire new_AGEMA_signal_4133 ;
    wire new_AGEMA_signal_4134 ;
    wire new_AGEMA_signal_4135 ;
    wire new_AGEMA_signal_4136 ;
    wire new_AGEMA_signal_4137 ;
    wire new_AGEMA_signal_4138 ;
    wire new_AGEMA_signal_4139 ;
    wire new_AGEMA_signal_4140 ;
    wire new_AGEMA_signal_4141 ;
    wire new_AGEMA_signal_4142 ;
    wire new_AGEMA_signal_4143 ;
    wire new_AGEMA_signal_4144 ;
    wire new_AGEMA_signal_4145 ;
    wire new_AGEMA_signal_4146 ;
    wire new_AGEMA_signal_4147 ;
    wire new_AGEMA_signal_4148 ;
    wire new_AGEMA_signal_4149 ;
    wire new_AGEMA_signal_4150 ;
    wire new_AGEMA_signal_4151 ;
    wire new_AGEMA_signal_4152 ;
    wire new_AGEMA_signal_4153 ;
    wire new_AGEMA_signal_4154 ;
    wire new_AGEMA_signal_4155 ;
    wire new_AGEMA_signal_4156 ;
    wire new_AGEMA_signal_4157 ;
    wire new_AGEMA_signal_4158 ;
    wire new_AGEMA_signal_4159 ;
    wire new_AGEMA_signal_4160 ;
    wire new_AGEMA_signal_4161 ;
    wire new_AGEMA_signal_4162 ;
    wire new_AGEMA_signal_4163 ;
    wire new_AGEMA_signal_4164 ;
    wire new_AGEMA_signal_4165 ;
    wire new_AGEMA_signal_4166 ;
    wire new_AGEMA_signal_4167 ;
    wire new_AGEMA_signal_4168 ;
    wire new_AGEMA_signal_4169 ;
    wire new_AGEMA_signal_4170 ;
    wire new_AGEMA_signal_4171 ;
    wire new_AGEMA_signal_4172 ;
    wire new_AGEMA_signal_4173 ;
    wire new_AGEMA_signal_4174 ;
    wire new_AGEMA_signal_4175 ;
    wire new_AGEMA_signal_4176 ;
    wire new_AGEMA_signal_4177 ;
    wire new_AGEMA_signal_4178 ;
    wire new_AGEMA_signal_4179 ;
    wire new_AGEMA_signal_4180 ;
    wire new_AGEMA_signal_4181 ;
    wire new_AGEMA_signal_4182 ;
    wire new_AGEMA_signal_4183 ;
    wire new_AGEMA_signal_4184 ;
    wire new_AGEMA_signal_4185 ;
    wire new_AGEMA_signal_4186 ;
    wire new_AGEMA_signal_4187 ;
    wire new_AGEMA_signal_4188 ;
    wire new_AGEMA_signal_4189 ;
    wire new_AGEMA_signal_4190 ;
    wire new_AGEMA_signal_4191 ;
    wire new_AGEMA_signal_4192 ;
    wire new_AGEMA_signal_4193 ;
    wire new_AGEMA_signal_4194 ;
    wire new_AGEMA_signal_4195 ;
    wire new_AGEMA_signal_4196 ;
    wire new_AGEMA_signal_4197 ;
    wire new_AGEMA_signal_4198 ;
    wire new_AGEMA_signal_4199 ;
    wire new_AGEMA_signal_4200 ;
    wire new_AGEMA_signal_4201 ;
    wire new_AGEMA_signal_4202 ;
    wire new_AGEMA_signal_4203 ;
    wire new_AGEMA_signal_4204 ;
    wire new_AGEMA_signal_4205 ;
    wire new_AGEMA_signal_4206 ;
    wire new_AGEMA_signal_4207 ;
    wire new_AGEMA_signal_4208 ;
    wire new_AGEMA_signal_4209 ;
    wire new_AGEMA_signal_4210 ;
    wire new_AGEMA_signal_4211 ;
    wire new_AGEMA_signal_4212 ;
    wire new_AGEMA_signal_4213 ;
    wire new_AGEMA_signal_4214 ;
    wire new_AGEMA_signal_4215 ;
    wire new_AGEMA_signal_4216 ;
    wire new_AGEMA_signal_4217 ;
    wire new_AGEMA_signal_4218 ;
    wire new_AGEMA_signal_4219 ;
    wire new_AGEMA_signal_4220 ;
    wire new_AGEMA_signal_4221 ;
    wire new_AGEMA_signal_4222 ;
    wire new_AGEMA_signal_4223 ;
    wire new_AGEMA_signal_4224 ;
    wire new_AGEMA_signal_4225 ;
    wire new_AGEMA_signal_4226 ;
    wire new_AGEMA_signal_4227 ;
    wire new_AGEMA_signal_4228 ;
    wire new_AGEMA_signal_4229 ;
    wire new_AGEMA_signal_4230 ;
    wire new_AGEMA_signal_4231 ;
    wire new_AGEMA_signal_4232 ;
    wire new_AGEMA_signal_4233 ;
    wire new_AGEMA_signal_4234 ;
    wire new_AGEMA_signal_4235 ;
    wire new_AGEMA_signal_4236 ;
    wire new_AGEMA_signal_4237 ;
    wire new_AGEMA_signal_4238 ;
    wire new_AGEMA_signal_4239 ;
    wire new_AGEMA_signal_4240 ;
    wire new_AGEMA_signal_4241 ;
    wire new_AGEMA_signal_4242 ;
    wire new_AGEMA_signal_4243 ;
    wire new_AGEMA_signal_4244 ;
    wire new_AGEMA_signal_4245 ;
    wire new_AGEMA_signal_4246 ;
    wire new_AGEMA_signal_4247 ;
    wire new_AGEMA_signal_4248 ;
    wire new_AGEMA_signal_4249 ;
    wire new_AGEMA_signal_4250 ;
    wire new_AGEMA_signal_4251 ;
    wire new_AGEMA_signal_4252 ;
    wire new_AGEMA_signal_4253 ;
    wire new_AGEMA_signal_4254 ;
    wire new_AGEMA_signal_4255 ;
    wire new_AGEMA_signal_4256 ;
    wire new_AGEMA_signal_4257 ;
    wire new_AGEMA_signal_4258 ;
    wire new_AGEMA_signal_4259 ;
    wire new_AGEMA_signal_4260 ;
    wire new_AGEMA_signal_4261 ;
    wire new_AGEMA_signal_4262 ;
    wire new_AGEMA_signal_4263 ;
    wire new_AGEMA_signal_4264 ;
    wire new_AGEMA_signal_4265 ;
    wire new_AGEMA_signal_4266 ;
    wire new_AGEMA_signal_4267 ;
    wire new_AGEMA_signal_4268 ;
    wire new_AGEMA_signal_4269 ;
    wire new_AGEMA_signal_4270 ;
    wire new_AGEMA_signal_4271 ;
    wire new_AGEMA_signal_4272 ;
    wire new_AGEMA_signal_4273 ;
    wire new_AGEMA_signal_4274 ;
    wire new_AGEMA_signal_4275 ;
    wire new_AGEMA_signal_4276 ;
    wire new_AGEMA_signal_4277 ;
    wire new_AGEMA_signal_4278 ;
    wire new_AGEMA_signal_4279 ;
    wire new_AGEMA_signal_4280 ;
    wire new_AGEMA_signal_4281 ;
    wire new_AGEMA_signal_4282 ;
    wire new_AGEMA_signal_4283 ;
    wire new_AGEMA_signal_4284 ;
    wire new_AGEMA_signal_4285 ;
    wire new_AGEMA_signal_4286 ;
    wire new_AGEMA_signal_4287 ;
    wire new_AGEMA_signal_4288 ;
    wire new_AGEMA_signal_4289 ;
    wire new_AGEMA_signal_4290 ;
    wire new_AGEMA_signal_4291 ;
    wire new_AGEMA_signal_4292 ;
    wire new_AGEMA_signal_4293 ;
    wire new_AGEMA_signal_4294 ;
    wire new_AGEMA_signal_4295 ;
    wire new_AGEMA_signal_4296 ;
    wire new_AGEMA_signal_4297 ;
    wire new_AGEMA_signal_4298 ;
    wire new_AGEMA_signal_4299 ;
    wire new_AGEMA_signal_4300 ;
    wire new_AGEMA_signal_4301 ;
    wire new_AGEMA_signal_4302 ;
    wire new_AGEMA_signal_4303 ;
    wire new_AGEMA_signal_4304 ;
    wire new_AGEMA_signal_4305 ;
    wire new_AGEMA_signal_4306 ;
    wire new_AGEMA_signal_4307 ;
    wire new_AGEMA_signal_4308 ;
    wire new_AGEMA_signal_4309 ;
    wire new_AGEMA_signal_4310 ;
    wire new_AGEMA_signal_4311 ;
    wire new_AGEMA_signal_4312 ;
    wire new_AGEMA_signal_4313 ;
    wire new_AGEMA_signal_4314 ;
    wire new_AGEMA_signal_4315 ;
    wire new_AGEMA_signal_4316 ;
    wire new_AGEMA_signal_4317 ;
    wire new_AGEMA_signal_4318 ;
    wire new_AGEMA_signal_4319 ;
    wire new_AGEMA_signal_4320 ;
    wire new_AGEMA_signal_4321 ;
    wire new_AGEMA_signal_4322 ;
    wire new_AGEMA_signal_4323 ;
    wire new_AGEMA_signal_4324 ;
    wire new_AGEMA_signal_4325 ;
    wire new_AGEMA_signal_4326 ;
    wire new_AGEMA_signal_4327 ;
    wire new_AGEMA_signal_4328 ;
    wire new_AGEMA_signal_4329 ;
    wire new_AGEMA_signal_4330 ;
    wire new_AGEMA_signal_4331 ;
    wire new_AGEMA_signal_4332 ;
    wire new_AGEMA_signal_4333 ;
    wire new_AGEMA_signal_4334 ;
    wire new_AGEMA_signal_4335 ;
    wire new_AGEMA_signal_4336 ;
    wire new_AGEMA_signal_4337 ;
    wire new_AGEMA_signal_4338 ;
    wire new_AGEMA_signal_4339 ;
    wire new_AGEMA_signal_4340 ;
    wire new_AGEMA_signal_4341 ;
    wire new_AGEMA_signal_4342 ;
    wire new_AGEMA_signal_4343 ;
    wire new_AGEMA_signal_4344 ;
    wire new_AGEMA_signal_4345 ;
    wire new_AGEMA_signal_4346 ;
    wire new_AGEMA_signal_4347 ;
    wire new_AGEMA_signal_4348 ;
    wire new_AGEMA_signal_4349 ;
    wire new_AGEMA_signal_4350 ;
    wire new_AGEMA_signal_4351 ;
    wire new_AGEMA_signal_4352 ;
    wire new_AGEMA_signal_4353 ;
    wire new_AGEMA_signal_4354 ;
    wire new_AGEMA_signal_4355 ;
    wire new_AGEMA_signal_4356 ;
    wire new_AGEMA_signal_4357 ;
    wire new_AGEMA_signal_4358 ;
    wire new_AGEMA_signal_4359 ;
    wire new_AGEMA_signal_4360 ;
    wire new_AGEMA_signal_4361 ;
    wire new_AGEMA_signal_4362 ;
    wire new_AGEMA_signal_4363 ;
    wire new_AGEMA_signal_4364 ;
    wire new_AGEMA_signal_4365 ;
    wire new_AGEMA_signal_4366 ;
    wire new_AGEMA_signal_4367 ;
    wire new_AGEMA_signal_4368 ;
    wire new_AGEMA_signal_4369 ;
    wire new_AGEMA_signal_4370 ;
    wire new_AGEMA_signal_4371 ;
    wire new_AGEMA_signal_4372 ;
    wire new_AGEMA_signal_4373 ;
    wire new_AGEMA_signal_4374 ;
    wire new_AGEMA_signal_4375 ;
    wire new_AGEMA_signal_4376 ;
    wire new_AGEMA_signal_4377 ;
    wire new_AGEMA_signal_4378 ;
    wire new_AGEMA_signal_4379 ;
    wire new_AGEMA_signal_4380 ;
    wire new_AGEMA_signal_4381 ;
    wire new_AGEMA_signal_4382 ;
    wire new_AGEMA_signal_4383 ;
    wire new_AGEMA_signal_4384 ;
    wire new_AGEMA_signal_4385 ;
    wire new_AGEMA_signal_4386 ;
    wire new_AGEMA_signal_4387 ;
    wire new_AGEMA_signal_4388 ;
    wire new_AGEMA_signal_4389 ;
    wire new_AGEMA_signal_4390 ;
    wire new_AGEMA_signal_4391 ;
    wire new_AGEMA_signal_4392 ;
    wire new_AGEMA_signal_4393 ;
    wire new_AGEMA_signal_4394 ;
    wire new_AGEMA_signal_4395 ;
    wire new_AGEMA_signal_4396 ;
    wire new_AGEMA_signal_4397 ;
    wire new_AGEMA_signal_4398 ;
    wire new_AGEMA_signal_4399 ;
    wire new_AGEMA_signal_4400 ;
    wire new_AGEMA_signal_4401 ;
    wire new_AGEMA_signal_4402 ;
    wire new_AGEMA_signal_4403 ;
    wire new_AGEMA_signal_4404 ;
    wire new_AGEMA_signal_4405 ;
    wire new_AGEMA_signal_4406 ;
    wire new_AGEMA_signal_4407 ;
    wire new_AGEMA_signal_4408 ;
    wire new_AGEMA_signal_4409 ;
    wire new_AGEMA_signal_4410 ;
    wire new_AGEMA_signal_4411 ;
    wire new_AGEMA_signal_4412 ;
    wire new_AGEMA_signal_4413 ;
    wire new_AGEMA_signal_4414 ;
    wire new_AGEMA_signal_4415 ;
    wire new_AGEMA_signal_4416 ;
    wire new_AGEMA_signal_4417 ;
    wire new_AGEMA_signal_4418 ;
    wire new_AGEMA_signal_4419 ;
    wire new_AGEMA_signal_4420 ;
    wire new_AGEMA_signal_4421 ;
    wire new_AGEMA_signal_4422 ;
    wire new_AGEMA_signal_4423 ;
    wire new_AGEMA_signal_4424 ;
    wire new_AGEMA_signal_4425 ;
    wire new_AGEMA_signal_4426 ;
    wire new_AGEMA_signal_4427 ;
    wire new_AGEMA_signal_4428 ;
    wire new_AGEMA_signal_4429 ;
    wire new_AGEMA_signal_4430 ;
    wire new_AGEMA_signal_4431 ;
    wire new_AGEMA_signal_4432 ;
    wire new_AGEMA_signal_4433 ;
    wire new_AGEMA_signal_4434 ;
    wire new_AGEMA_signal_4435 ;
    wire new_AGEMA_signal_4436 ;
    wire new_AGEMA_signal_4437 ;
    wire new_AGEMA_signal_4438 ;
    wire new_AGEMA_signal_4439 ;
    wire new_AGEMA_signal_4440 ;
    wire new_AGEMA_signal_4441 ;
    wire new_AGEMA_signal_4442 ;
    wire new_AGEMA_signal_4443 ;
    wire new_AGEMA_signal_4444 ;
    wire new_AGEMA_signal_4445 ;
    wire new_AGEMA_signal_4446 ;
    wire new_AGEMA_signal_4447 ;
    wire new_AGEMA_signal_4448 ;
    wire new_AGEMA_signal_4449 ;
    wire new_AGEMA_signal_4450 ;
    wire new_AGEMA_signal_4451 ;
    wire new_AGEMA_signal_4452 ;
    wire new_AGEMA_signal_4453 ;
    wire new_AGEMA_signal_4454 ;
    wire new_AGEMA_signal_4455 ;
    wire new_AGEMA_signal_4456 ;
    wire new_AGEMA_signal_4457 ;
    wire new_AGEMA_signal_4458 ;
    wire new_AGEMA_signal_4459 ;
    wire new_AGEMA_signal_4460 ;
    wire new_AGEMA_signal_4461 ;
    wire new_AGEMA_signal_4462 ;
    wire new_AGEMA_signal_4463 ;
    wire new_AGEMA_signal_4464 ;
    wire new_AGEMA_signal_4465 ;
    wire new_AGEMA_signal_4466 ;
    wire new_AGEMA_signal_4467 ;
    wire new_AGEMA_signal_4468 ;
    wire new_AGEMA_signal_4469 ;
    wire new_AGEMA_signal_4470 ;
    wire new_AGEMA_signal_4471 ;
    wire new_AGEMA_signal_4472 ;
    wire new_AGEMA_signal_4473 ;
    wire new_AGEMA_signal_4474 ;
    wire new_AGEMA_signal_4475 ;
    wire new_AGEMA_signal_4476 ;
    wire new_AGEMA_signal_4477 ;
    wire new_AGEMA_signal_4478 ;
    wire new_AGEMA_signal_4479 ;
    wire new_AGEMA_signal_4480 ;
    wire new_AGEMA_signal_4481 ;
    wire new_AGEMA_signal_4482 ;
    wire new_AGEMA_signal_4483 ;
    wire new_AGEMA_signal_4484 ;
    wire new_AGEMA_signal_4485 ;
    wire new_AGEMA_signal_4486 ;
    wire new_AGEMA_signal_4487 ;
    wire new_AGEMA_signal_4488 ;
    wire new_AGEMA_signal_4489 ;
    wire new_AGEMA_signal_4490 ;
    wire new_AGEMA_signal_4491 ;
    wire new_AGEMA_signal_4492 ;
    wire new_AGEMA_signal_4493 ;
    wire new_AGEMA_signal_4494 ;
    wire new_AGEMA_signal_4495 ;
    wire new_AGEMA_signal_4496 ;
    wire new_AGEMA_signal_4497 ;
    wire new_AGEMA_signal_4498 ;
    wire new_AGEMA_signal_4499 ;
    wire new_AGEMA_signal_4500 ;
    wire new_AGEMA_signal_4501 ;
    wire new_AGEMA_signal_4502 ;
    wire new_AGEMA_signal_4503 ;
    wire new_AGEMA_signal_4504 ;
    wire new_AGEMA_signal_4505 ;
    wire new_AGEMA_signal_4506 ;
    wire new_AGEMA_signal_4507 ;
    wire new_AGEMA_signal_4508 ;
    wire new_AGEMA_signal_4509 ;
    wire new_AGEMA_signal_4510 ;
    wire new_AGEMA_signal_4511 ;
    wire new_AGEMA_signal_4512 ;
    wire new_AGEMA_signal_4513 ;
    wire new_AGEMA_signal_4514 ;
    wire new_AGEMA_signal_4515 ;
    wire new_AGEMA_signal_4516 ;
    wire new_AGEMA_signal_4517 ;
    wire new_AGEMA_signal_4518 ;
    wire new_AGEMA_signal_4519 ;
    wire new_AGEMA_signal_4520 ;
    wire new_AGEMA_signal_4521 ;
    wire new_AGEMA_signal_4522 ;
    wire new_AGEMA_signal_4523 ;
    wire new_AGEMA_signal_4524 ;
    wire new_AGEMA_signal_4525 ;
    wire new_AGEMA_signal_4526 ;
    wire new_AGEMA_signal_4527 ;
    wire new_AGEMA_signal_4528 ;
    wire new_AGEMA_signal_4529 ;
    wire new_AGEMA_signal_4530 ;
    wire new_AGEMA_signal_4531 ;
    wire new_AGEMA_signal_4532 ;
    wire new_AGEMA_signal_4533 ;
    wire new_AGEMA_signal_4534 ;
    wire new_AGEMA_signal_4535 ;
    wire new_AGEMA_signal_4536 ;
    wire new_AGEMA_signal_4537 ;
    wire new_AGEMA_signal_4538 ;
    wire new_AGEMA_signal_4539 ;
    wire new_AGEMA_signal_4540 ;
    wire new_AGEMA_signal_4541 ;
    wire new_AGEMA_signal_4542 ;
    wire new_AGEMA_signal_4543 ;
    wire new_AGEMA_signal_4544 ;
    wire new_AGEMA_signal_4545 ;
    wire new_AGEMA_signal_4546 ;
    wire new_AGEMA_signal_4547 ;
    wire new_AGEMA_signal_4548 ;
    wire new_AGEMA_signal_4549 ;
    wire new_AGEMA_signal_4550 ;
    wire new_AGEMA_signal_4551 ;
    wire new_AGEMA_signal_4552 ;
    wire new_AGEMA_signal_4553 ;
    wire new_AGEMA_signal_4554 ;
    wire new_AGEMA_signal_4555 ;
    wire new_AGEMA_signal_4556 ;
    wire new_AGEMA_signal_4557 ;
    wire new_AGEMA_signal_4558 ;
    wire new_AGEMA_signal_4559 ;
    wire new_AGEMA_signal_4560 ;
    wire new_AGEMA_signal_4561 ;
    wire new_AGEMA_signal_4562 ;
    wire new_AGEMA_signal_4563 ;
    wire new_AGEMA_signal_4564 ;
    wire new_AGEMA_signal_4565 ;
    wire new_AGEMA_signal_4566 ;
    wire new_AGEMA_signal_4567 ;
    wire new_AGEMA_signal_4568 ;
    wire new_AGEMA_signal_4569 ;
    wire new_AGEMA_signal_4570 ;
    wire new_AGEMA_signal_4571 ;
    wire new_AGEMA_signal_4572 ;
    wire new_AGEMA_signal_4573 ;
    wire new_AGEMA_signal_4574 ;
    wire new_AGEMA_signal_4575 ;
    wire new_AGEMA_signal_4576 ;
    wire new_AGEMA_signal_4577 ;
    wire new_AGEMA_signal_4578 ;
    wire new_AGEMA_signal_4579 ;
    wire new_AGEMA_signal_4580 ;
    wire new_AGEMA_signal_4581 ;
    wire new_AGEMA_signal_4582 ;
    wire new_AGEMA_signal_4583 ;
    wire new_AGEMA_signal_4584 ;
    wire new_AGEMA_signal_4585 ;
    wire new_AGEMA_signal_4586 ;
    wire new_AGEMA_signal_4587 ;
    wire new_AGEMA_signal_4588 ;
    wire new_AGEMA_signal_4589 ;
    wire new_AGEMA_signal_4590 ;
    wire new_AGEMA_signal_4591 ;
    wire new_AGEMA_signal_4592 ;
    wire new_AGEMA_signal_4593 ;
    wire new_AGEMA_signal_4594 ;
    wire new_AGEMA_signal_4595 ;
    wire new_AGEMA_signal_4596 ;
    wire new_AGEMA_signal_4597 ;
    wire new_AGEMA_signal_4598 ;
    wire new_AGEMA_signal_4599 ;
    wire new_AGEMA_signal_4600 ;
    wire new_AGEMA_signal_4601 ;
    wire new_AGEMA_signal_4602 ;
    wire new_AGEMA_signal_4603 ;
    wire new_AGEMA_signal_4604 ;
    wire new_AGEMA_signal_4605 ;
    wire new_AGEMA_signal_4606 ;
    wire new_AGEMA_signal_4607 ;
    wire new_AGEMA_signal_4608 ;
    wire new_AGEMA_signal_4609 ;
    wire new_AGEMA_signal_4610 ;
    wire new_AGEMA_signal_4611 ;
    wire new_AGEMA_signal_4612 ;
    wire new_AGEMA_signal_4613 ;
    wire new_AGEMA_signal_4614 ;
    wire new_AGEMA_signal_4615 ;
    wire new_AGEMA_signal_4616 ;
    wire new_AGEMA_signal_4617 ;
    wire new_AGEMA_signal_4618 ;
    wire new_AGEMA_signal_4619 ;
    wire new_AGEMA_signal_4620 ;
    wire new_AGEMA_signal_4621 ;
    wire new_AGEMA_signal_4622 ;
    wire new_AGEMA_signal_4623 ;
    wire new_AGEMA_signal_4624 ;
    wire new_AGEMA_signal_4625 ;
    wire new_AGEMA_signal_4626 ;
    wire new_AGEMA_signal_4627 ;
    wire new_AGEMA_signal_4628 ;
    wire new_AGEMA_signal_4629 ;
    wire new_AGEMA_signal_4630 ;
    wire new_AGEMA_signal_4631 ;
    wire new_AGEMA_signal_4632 ;
    wire new_AGEMA_signal_4633 ;
    wire new_AGEMA_signal_4634 ;
    wire new_AGEMA_signal_4635 ;
    wire new_AGEMA_signal_4636 ;
    wire new_AGEMA_signal_4637 ;
    wire new_AGEMA_signal_4638 ;
    wire new_AGEMA_signal_4639 ;
    wire new_AGEMA_signal_4640 ;
    wire new_AGEMA_signal_4641 ;
    wire new_AGEMA_signal_4642 ;
    wire new_AGEMA_signal_4643 ;
    wire new_AGEMA_signal_4644 ;
    wire new_AGEMA_signal_4645 ;
    wire new_AGEMA_signal_4646 ;
    wire new_AGEMA_signal_4647 ;
    wire new_AGEMA_signal_4648 ;
    wire new_AGEMA_signal_4649 ;
    wire new_AGEMA_signal_4650 ;
    wire new_AGEMA_signal_4651 ;
    wire new_AGEMA_signal_4652 ;
    wire new_AGEMA_signal_4653 ;
    wire new_AGEMA_signal_4654 ;
    wire new_AGEMA_signal_4655 ;
    wire new_AGEMA_signal_4656 ;
    wire new_AGEMA_signal_4657 ;
    wire new_AGEMA_signal_4658 ;
    wire new_AGEMA_signal_4659 ;
    wire new_AGEMA_signal_4660 ;
    wire new_AGEMA_signal_4661 ;
    wire new_AGEMA_signal_4662 ;
    wire new_AGEMA_signal_4663 ;
    wire new_AGEMA_signal_4664 ;
    wire new_AGEMA_signal_4665 ;
    wire new_AGEMA_signal_4666 ;
    wire new_AGEMA_signal_4667 ;
    wire new_AGEMA_signal_4668 ;
    wire new_AGEMA_signal_4669 ;
    wire new_AGEMA_signal_4670 ;
    wire new_AGEMA_signal_4671 ;
    wire new_AGEMA_signal_4672 ;
    wire new_AGEMA_signal_4673 ;
    wire new_AGEMA_signal_4674 ;
    wire new_AGEMA_signal_4675 ;
    wire new_AGEMA_signal_4676 ;
    wire new_AGEMA_signal_4677 ;
    wire new_AGEMA_signal_4678 ;
    wire new_AGEMA_signal_4679 ;
    wire new_AGEMA_signal_4680 ;
    wire new_AGEMA_signal_4681 ;
    wire new_AGEMA_signal_4682 ;
    wire new_AGEMA_signal_4683 ;
    wire new_AGEMA_signal_4684 ;
    wire new_AGEMA_signal_4685 ;
    wire new_AGEMA_signal_4686 ;
    wire new_AGEMA_signal_4687 ;
    wire new_AGEMA_signal_4688 ;
    wire new_AGEMA_signal_4689 ;
    wire new_AGEMA_signal_4690 ;
    wire new_AGEMA_signal_4691 ;
    wire new_AGEMA_signal_4692 ;
    wire new_AGEMA_signal_4693 ;
    wire new_AGEMA_signal_4694 ;
    wire new_AGEMA_signal_4695 ;
    wire new_AGEMA_signal_4696 ;
    wire new_AGEMA_signal_4697 ;
    wire new_AGEMA_signal_4698 ;
    wire new_AGEMA_signal_4699 ;
    wire new_AGEMA_signal_4700 ;
    wire new_AGEMA_signal_4701 ;
    wire new_AGEMA_signal_4702 ;
    wire new_AGEMA_signal_4703 ;
    wire new_AGEMA_signal_4704 ;
    wire new_AGEMA_signal_4705 ;
    wire new_AGEMA_signal_4706 ;
    wire new_AGEMA_signal_4707 ;
    wire new_AGEMA_signal_4708 ;
    wire new_AGEMA_signal_4709 ;
    wire new_AGEMA_signal_4710 ;
    wire new_AGEMA_signal_4711 ;
    wire new_AGEMA_signal_4712 ;
    wire new_AGEMA_signal_4713 ;
    wire new_AGEMA_signal_4714 ;
    wire new_AGEMA_signal_4715 ;
    wire new_AGEMA_signal_4716 ;
    wire new_AGEMA_signal_4717 ;
    wire new_AGEMA_signal_4718 ;
    wire new_AGEMA_signal_4719 ;
    wire new_AGEMA_signal_4720 ;
    wire new_AGEMA_signal_4721 ;
    wire new_AGEMA_signal_4722 ;
    wire new_AGEMA_signal_4723 ;
    wire new_AGEMA_signal_4724 ;
    wire new_AGEMA_signal_4725 ;
    wire new_AGEMA_signal_4726 ;
    wire new_AGEMA_signal_4727 ;
    wire new_AGEMA_signal_4728 ;
    wire new_AGEMA_signal_4729 ;
    wire new_AGEMA_signal_4730 ;
    wire new_AGEMA_signal_4731 ;
    wire new_AGEMA_signal_4732 ;
    wire new_AGEMA_signal_4733 ;
    wire new_AGEMA_signal_4734 ;
    wire new_AGEMA_signal_4735 ;
    wire new_AGEMA_signal_4736 ;
    wire new_AGEMA_signal_4737 ;
    wire new_AGEMA_signal_4738 ;
    wire new_AGEMA_signal_4739 ;
    wire new_AGEMA_signal_4740 ;
    wire new_AGEMA_signal_4741 ;
    wire new_AGEMA_signal_4742 ;
    wire new_AGEMA_signal_4743 ;
    wire new_AGEMA_signal_4744 ;
    wire new_AGEMA_signal_4745 ;
    wire new_AGEMA_signal_4746 ;
    wire new_AGEMA_signal_4747 ;
    wire new_AGEMA_signal_4748 ;
    wire new_AGEMA_signal_4749 ;
    wire new_AGEMA_signal_4750 ;
    wire new_AGEMA_signal_4751 ;
    wire new_AGEMA_signal_4752 ;
    wire new_AGEMA_signal_4753 ;
    wire new_AGEMA_signal_4754 ;
    wire new_AGEMA_signal_4755 ;
    wire new_AGEMA_signal_4756 ;
    wire new_AGEMA_signal_4757 ;
    wire new_AGEMA_signal_4758 ;
    wire new_AGEMA_signal_4759 ;
    wire new_AGEMA_signal_4760 ;
    wire new_AGEMA_signal_4761 ;
    wire new_AGEMA_signal_4762 ;
    wire new_AGEMA_signal_4763 ;
    wire new_AGEMA_signal_4764 ;
    wire new_AGEMA_signal_4765 ;
    wire new_AGEMA_signal_4766 ;
    wire new_AGEMA_signal_4767 ;
    wire new_AGEMA_signal_4768 ;
    wire new_AGEMA_signal_4769 ;
    wire new_AGEMA_signal_4770 ;
    wire new_AGEMA_signal_4771 ;
    wire new_AGEMA_signal_4772 ;
    wire new_AGEMA_signal_4773 ;
    wire new_AGEMA_signal_4774 ;
    wire new_AGEMA_signal_4775 ;
    wire new_AGEMA_signal_4776 ;
    wire new_AGEMA_signal_4777 ;
    wire new_AGEMA_signal_4778 ;
    wire new_AGEMA_signal_4779 ;
    wire new_AGEMA_signal_4780 ;
    wire new_AGEMA_signal_4781 ;
    wire new_AGEMA_signal_4782 ;
    wire new_AGEMA_signal_4783 ;
    wire new_AGEMA_signal_4784 ;
    wire new_AGEMA_signal_4785 ;
    wire new_AGEMA_signal_4786 ;
    wire new_AGEMA_signal_4787 ;
    wire new_AGEMA_signal_4788 ;
    wire new_AGEMA_signal_4789 ;
    wire new_AGEMA_signal_4790 ;
    wire new_AGEMA_signal_4791 ;
    wire new_AGEMA_signal_4792 ;
    wire new_AGEMA_signal_4793 ;
    wire new_AGEMA_signal_4794 ;
    wire new_AGEMA_signal_4795 ;
    wire new_AGEMA_signal_4796 ;
    wire new_AGEMA_signal_4797 ;
    wire new_AGEMA_signal_4798 ;
    wire new_AGEMA_signal_4799 ;
    wire new_AGEMA_signal_4800 ;
    wire new_AGEMA_signal_4801 ;
    wire new_AGEMA_signal_4802 ;
    wire new_AGEMA_signal_4803 ;
    wire new_AGEMA_signal_4804 ;
    wire new_AGEMA_signal_4805 ;
    wire new_AGEMA_signal_4806 ;
    wire new_AGEMA_signal_4807 ;
    wire new_AGEMA_signal_4808 ;
    wire new_AGEMA_signal_4809 ;
    wire new_AGEMA_signal_4810 ;
    wire new_AGEMA_signal_4811 ;
    wire new_AGEMA_signal_4812 ;
    wire new_AGEMA_signal_4813 ;
    wire new_AGEMA_signal_4814 ;
    wire new_AGEMA_signal_4815 ;
    wire new_AGEMA_signal_4816 ;
    wire new_AGEMA_signal_4817 ;
    wire new_AGEMA_signal_4818 ;
    wire new_AGEMA_signal_4819 ;
    wire new_AGEMA_signal_4820 ;
    wire new_AGEMA_signal_4821 ;
    wire new_AGEMA_signal_4822 ;
    wire new_AGEMA_signal_4823 ;
    wire new_AGEMA_signal_4824 ;
    wire new_AGEMA_signal_4825 ;
    wire new_AGEMA_signal_4826 ;
    wire new_AGEMA_signal_4827 ;
    wire new_AGEMA_signal_4828 ;
    wire new_AGEMA_signal_4829 ;
    wire new_AGEMA_signal_4830 ;
    wire new_AGEMA_signal_4831 ;
    wire new_AGEMA_signal_4832 ;
    wire new_AGEMA_signal_4833 ;
    wire new_AGEMA_signal_4834 ;
    wire new_AGEMA_signal_4835 ;
    wire new_AGEMA_signal_4836 ;
    wire new_AGEMA_signal_4837 ;
    wire new_AGEMA_signal_4838 ;
    wire new_AGEMA_signal_4839 ;
    wire new_AGEMA_signal_4840 ;
    wire new_AGEMA_signal_4841 ;
    wire new_AGEMA_signal_4842 ;
    wire new_AGEMA_signal_4843 ;
    wire new_AGEMA_signal_4844 ;
    wire new_AGEMA_signal_4845 ;
    wire new_AGEMA_signal_4846 ;
    wire new_AGEMA_signal_4847 ;
    wire new_AGEMA_signal_4848 ;
    wire new_AGEMA_signal_4849 ;
    wire new_AGEMA_signal_4850 ;
    wire new_AGEMA_signal_4851 ;
    wire new_AGEMA_signal_4852 ;
    wire new_AGEMA_signal_4853 ;
    wire new_AGEMA_signal_4854 ;
    wire new_AGEMA_signal_4855 ;
    wire new_AGEMA_signal_4856 ;
    wire new_AGEMA_signal_4857 ;
    wire new_AGEMA_signal_4858 ;
    wire new_AGEMA_signal_4859 ;
    wire new_AGEMA_signal_4860 ;
    wire new_AGEMA_signal_4861 ;
    wire new_AGEMA_signal_4862 ;
    wire new_AGEMA_signal_4863 ;
    wire new_AGEMA_signal_4864 ;
    wire new_AGEMA_signal_4865 ;
    wire new_AGEMA_signal_4866 ;
    wire new_AGEMA_signal_4867 ;
    wire new_AGEMA_signal_4868 ;
    wire new_AGEMA_signal_4869 ;
    wire new_AGEMA_signal_4870 ;
    wire new_AGEMA_signal_4871 ;
    wire new_AGEMA_signal_4872 ;
    wire new_AGEMA_signal_4873 ;
    wire new_AGEMA_signal_4874 ;
    wire new_AGEMA_signal_4875 ;
    wire new_AGEMA_signal_4876 ;
    wire new_AGEMA_signal_4877 ;
    wire new_AGEMA_signal_4878 ;
    wire new_AGEMA_signal_4879 ;
    wire new_AGEMA_signal_4880 ;
    wire new_AGEMA_signal_4881 ;
    wire new_AGEMA_signal_4882 ;
    wire new_AGEMA_signal_4883 ;
    wire new_AGEMA_signal_4884 ;
    wire new_AGEMA_signal_4885 ;
    wire new_AGEMA_signal_4886 ;
    wire new_AGEMA_signal_4887 ;
    wire new_AGEMA_signal_4888 ;
    wire new_AGEMA_signal_4889 ;
    wire new_AGEMA_signal_4890 ;
    wire new_AGEMA_signal_4891 ;
    wire new_AGEMA_signal_4892 ;
    wire new_AGEMA_signal_4893 ;
    wire new_AGEMA_signal_4894 ;
    wire new_AGEMA_signal_4895 ;
    wire new_AGEMA_signal_4896 ;
    wire new_AGEMA_signal_4897 ;
    wire new_AGEMA_signal_4898 ;
    wire new_AGEMA_signal_4899 ;
    wire new_AGEMA_signal_4900 ;
    wire new_AGEMA_signal_4901 ;
    wire new_AGEMA_signal_4902 ;
    wire new_AGEMA_signal_4903 ;
    wire new_AGEMA_signal_4904 ;
    wire new_AGEMA_signal_4905 ;
    wire new_AGEMA_signal_4906 ;
    wire new_AGEMA_signal_4907 ;
    wire new_AGEMA_signal_4908 ;
    wire new_AGEMA_signal_4909 ;
    wire new_AGEMA_signal_4910 ;
    wire new_AGEMA_signal_4911 ;
    wire new_AGEMA_signal_4912 ;
    wire new_AGEMA_signal_4913 ;
    wire new_AGEMA_signal_4914 ;
    wire new_AGEMA_signal_4915 ;
    wire new_AGEMA_signal_4916 ;
    wire new_AGEMA_signal_4917 ;
    wire new_AGEMA_signal_4918 ;
    wire new_AGEMA_signal_4919 ;
    wire new_AGEMA_signal_4920 ;
    wire new_AGEMA_signal_4921 ;
    wire new_AGEMA_signal_4922 ;
    wire new_AGEMA_signal_4923 ;
    wire new_AGEMA_signal_4924 ;
    wire new_AGEMA_signal_4925 ;
    wire new_AGEMA_signal_4926 ;
    wire new_AGEMA_signal_4927 ;
    wire new_AGEMA_signal_4928 ;
    wire new_AGEMA_signal_4929 ;
    wire new_AGEMA_signal_4930 ;
    wire new_AGEMA_signal_4931 ;
    wire new_AGEMA_signal_4932 ;
    wire new_AGEMA_signal_4933 ;
    wire new_AGEMA_signal_4934 ;
    wire new_AGEMA_signal_4935 ;
    wire new_AGEMA_signal_4936 ;
    wire new_AGEMA_signal_4937 ;
    wire new_AGEMA_signal_4938 ;
    wire new_AGEMA_signal_4939 ;
    wire new_AGEMA_signal_4940 ;
    wire new_AGEMA_signal_4941 ;
    wire new_AGEMA_signal_4942 ;
    wire new_AGEMA_signal_4943 ;
    wire new_AGEMA_signal_4944 ;
    wire new_AGEMA_signal_4945 ;
    wire new_AGEMA_signal_4946 ;
    wire new_AGEMA_signal_4947 ;
    wire new_AGEMA_signal_4948 ;
    wire new_AGEMA_signal_4949 ;
    wire new_AGEMA_signal_4950 ;
    wire new_AGEMA_signal_4951 ;
    wire new_AGEMA_signal_4952 ;
    wire new_AGEMA_signal_4953 ;
    wire new_AGEMA_signal_4954 ;
    wire new_AGEMA_signal_4955 ;
    wire new_AGEMA_signal_4956 ;
    wire new_AGEMA_signal_4957 ;
    wire new_AGEMA_signal_4958 ;
    wire new_AGEMA_signal_4959 ;
    wire new_AGEMA_signal_4960 ;
    wire new_AGEMA_signal_4961 ;
    wire new_AGEMA_signal_4962 ;
    wire new_AGEMA_signal_4963 ;
    wire new_AGEMA_signal_4964 ;
    wire new_AGEMA_signal_4965 ;
    wire new_AGEMA_signal_4966 ;
    wire new_AGEMA_signal_4967 ;
    wire new_AGEMA_signal_4968 ;
    wire new_AGEMA_signal_4969 ;
    wire new_AGEMA_signal_4970 ;
    wire new_AGEMA_signal_4971 ;
    wire new_AGEMA_signal_4972 ;
    wire new_AGEMA_signal_4973 ;
    wire new_AGEMA_signal_4974 ;
    wire new_AGEMA_signal_4975 ;
    wire new_AGEMA_signal_4976 ;
    wire new_AGEMA_signal_4977 ;
    wire new_AGEMA_signal_4978 ;
    wire new_AGEMA_signal_4979 ;
    wire new_AGEMA_signal_4980 ;
    wire new_AGEMA_signal_4981 ;
    wire new_AGEMA_signal_4982 ;
    wire new_AGEMA_signal_4983 ;
    wire new_AGEMA_signal_4984 ;
    wire new_AGEMA_signal_4985 ;
    wire new_AGEMA_signal_4986 ;
    wire new_AGEMA_signal_4987 ;
    wire new_AGEMA_signal_4988 ;
    wire new_AGEMA_signal_4989 ;
    wire new_AGEMA_signal_4990 ;
    wire new_AGEMA_signal_4991 ;
    wire new_AGEMA_signal_4992 ;
    wire new_AGEMA_signal_4993 ;
    wire new_AGEMA_signal_4994 ;
    wire new_AGEMA_signal_4995 ;
    wire new_AGEMA_signal_4996 ;
    wire new_AGEMA_signal_4997 ;
    wire new_AGEMA_signal_4998 ;
    wire new_AGEMA_signal_4999 ;
    wire new_AGEMA_signal_5000 ;
    wire new_AGEMA_signal_5001 ;
    wire new_AGEMA_signal_5002 ;
    wire new_AGEMA_signal_5003 ;
    wire new_AGEMA_signal_5004 ;
    wire new_AGEMA_signal_5005 ;
    wire new_AGEMA_signal_5006 ;
    wire new_AGEMA_signal_5007 ;
    wire new_AGEMA_signal_5008 ;
    wire new_AGEMA_signal_5009 ;
    wire new_AGEMA_signal_5010 ;
    wire new_AGEMA_signal_5011 ;
    wire new_AGEMA_signal_5012 ;
    wire new_AGEMA_signal_5013 ;
    wire new_AGEMA_signal_5014 ;
    wire new_AGEMA_signal_5015 ;
    wire new_AGEMA_signal_5016 ;
    wire new_AGEMA_signal_5017 ;
    wire new_AGEMA_signal_5018 ;
    wire new_AGEMA_signal_5019 ;
    wire new_AGEMA_signal_5020 ;
    wire new_AGEMA_signal_5021 ;
    wire new_AGEMA_signal_5022 ;
    wire new_AGEMA_signal_5023 ;
    wire new_AGEMA_signal_5024 ;
    wire new_AGEMA_signal_5025 ;
    wire new_AGEMA_signal_5026 ;
    wire new_AGEMA_signal_5027 ;
    wire new_AGEMA_signal_5028 ;
    wire new_AGEMA_signal_5029 ;
    wire new_AGEMA_signal_5030 ;
    wire new_AGEMA_signal_5031 ;
    wire new_AGEMA_signal_5032 ;
    wire new_AGEMA_signal_5033 ;
    wire new_AGEMA_signal_5034 ;
    wire new_AGEMA_signal_5035 ;
    wire new_AGEMA_signal_5036 ;
    wire new_AGEMA_signal_5037 ;
    wire new_AGEMA_signal_5038 ;
    wire new_AGEMA_signal_5039 ;
    wire new_AGEMA_signal_5040 ;
    wire new_AGEMA_signal_5041 ;
    wire new_AGEMA_signal_5042 ;
    wire new_AGEMA_signal_5043 ;
    wire new_AGEMA_signal_5044 ;
    wire new_AGEMA_signal_5045 ;
    wire new_AGEMA_signal_5046 ;
    wire new_AGEMA_signal_5047 ;
    wire new_AGEMA_signal_5048 ;
    wire new_AGEMA_signal_5049 ;
    wire new_AGEMA_signal_5050 ;
    wire new_AGEMA_signal_5051 ;
    wire new_AGEMA_signal_5052 ;
    wire new_AGEMA_signal_5053 ;
    wire new_AGEMA_signal_5054 ;
    wire new_AGEMA_signal_5055 ;
    wire new_AGEMA_signal_5056 ;
    wire new_AGEMA_signal_5057 ;
    wire new_AGEMA_signal_5058 ;
    wire new_AGEMA_signal_5059 ;
    wire new_AGEMA_signal_5060 ;
    wire new_AGEMA_signal_5061 ;
    wire new_AGEMA_signal_5062 ;
    wire new_AGEMA_signal_5063 ;
    wire new_AGEMA_signal_5064 ;
    wire new_AGEMA_signal_5065 ;
    wire new_AGEMA_signal_5066 ;
    wire new_AGEMA_signal_5067 ;
    wire new_AGEMA_signal_5068 ;
    wire new_AGEMA_signal_5069 ;
    wire new_AGEMA_signal_5070 ;
    wire new_AGEMA_signal_5071 ;
    wire new_AGEMA_signal_5072 ;
    wire new_AGEMA_signal_5073 ;
    wire new_AGEMA_signal_5074 ;
    wire new_AGEMA_signal_5075 ;
    wire new_AGEMA_signal_5076 ;
    wire new_AGEMA_signal_5077 ;
    wire new_AGEMA_signal_5078 ;
    wire new_AGEMA_signal_5079 ;
    wire new_AGEMA_signal_5080 ;
    wire new_AGEMA_signal_5081 ;
    wire new_AGEMA_signal_5082 ;
    wire new_AGEMA_signal_5083 ;
    wire new_AGEMA_signal_5084 ;
    wire new_AGEMA_signal_5085 ;
    wire new_AGEMA_signal_5086 ;
    wire new_AGEMA_signal_5087 ;
    wire new_AGEMA_signal_5088 ;
    wire new_AGEMA_signal_5089 ;
    wire new_AGEMA_signal_5090 ;
    wire new_AGEMA_signal_5091 ;
    wire new_AGEMA_signal_5092 ;
    wire new_AGEMA_signal_5093 ;
    wire new_AGEMA_signal_5094 ;
    wire new_AGEMA_signal_5095 ;
    wire new_AGEMA_signal_5096 ;
    wire new_AGEMA_signal_5097 ;
    wire new_AGEMA_signal_5098 ;
    wire new_AGEMA_signal_5099 ;
    wire new_AGEMA_signal_5100 ;
    wire new_AGEMA_signal_5101 ;
    wire new_AGEMA_signal_5102 ;
    wire new_AGEMA_signal_5103 ;
    wire new_AGEMA_signal_5104 ;
    wire new_AGEMA_signal_5105 ;
    wire new_AGEMA_signal_5106 ;
    wire new_AGEMA_signal_5107 ;
    wire new_AGEMA_signal_5108 ;
    wire new_AGEMA_signal_5109 ;
    wire new_AGEMA_signal_5110 ;
    wire new_AGEMA_signal_5111 ;
    wire new_AGEMA_signal_5112 ;
    wire new_AGEMA_signal_5113 ;
    wire new_AGEMA_signal_5114 ;
    wire new_AGEMA_signal_5115 ;
    wire new_AGEMA_signal_5116 ;
    wire new_AGEMA_signal_5117 ;
    wire new_AGEMA_signal_5118 ;
    wire new_AGEMA_signal_5119 ;
    wire new_AGEMA_signal_5120 ;
    wire new_AGEMA_signal_5121 ;
    wire new_AGEMA_signal_5122 ;
    wire new_AGEMA_signal_5123 ;
    wire new_AGEMA_signal_5124 ;
    wire new_AGEMA_signal_5125 ;
    wire new_AGEMA_signal_5126 ;
    wire new_AGEMA_signal_5127 ;
    wire new_AGEMA_signal_5128 ;
    wire new_AGEMA_signal_5129 ;
    wire new_AGEMA_signal_5130 ;
    wire new_AGEMA_signal_5131 ;
    wire new_AGEMA_signal_5132 ;
    wire new_AGEMA_signal_5133 ;
    wire new_AGEMA_signal_5134 ;
    wire new_AGEMA_signal_5135 ;
    wire new_AGEMA_signal_5136 ;
    wire new_AGEMA_signal_5137 ;
    wire new_AGEMA_signal_5138 ;
    wire new_AGEMA_signal_5139 ;
    wire new_AGEMA_signal_5140 ;
    wire new_AGEMA_signal_5141 ;
    wire new_AGEMA_signal_5142 ;
    wire new_AGEMA_signal_5143 ;
    wire new_AGEMA_signal_5144 ;
    wire new_AGEMA_signal_5145 ;
    wire new_AGEMA_signal_5146 ;
    wire new_AGEMA_signal_5147 ;
    wire new_AGEMA_signal_5148 ;
    wire new_AGEMA_signal_5149 ;
    wire new_AGEMA_signal_5150 ;
    wire new_AGEMA_signal_5151 ;
    wire new_AGEMA_signal_5152 ;
    wire new_AGEMA_signal_5153 ;
    wire new_AGEMA_signal_5154 ;
    wire new_AGEMA_signal_5155 ;
    wire new_AGEMA_signal_5156 ;
    wire new_AGEMA_signal_5157 ;
    wire new_AGEMA_signal_5158 ;
    wire new_AGEMA_signal_5159 ;
    wire new_AGEMA_signal_5160 ;
    wire new_AGEMA_signal_5161 ;
    wire new_AGEMA_signal_5162 ;
    wire new_AGEMA_signal_5163 ;
    wire new_AGEMA_signal_5164 ;
    wire new_AGEMA_signal_5165 ;
    wire new_AGEMA_signal_5166 ;
    wire new_AGEMA_signal_5167 ;
    wire new_AGEMA_signal_5168 ;
    wire new_AGEMA_signal_5169 ;
    wire new_AGEMA_signal_5170 ;
    wire new_AGEMA_signal_5171 ;
    wire new_AGEMA_signal_5172 ;
    wire new_AGEMA_signal_5173 ;
    wire new_AGEMA_signal_5174 ;
    wire new_AGEMA_signal_5175 ;
    wire new_AGEMA_signal_5176 ;
    wire new_AGEMA_signal_5177 ;
    wire new_AGEMA_signal_5178 ;
    wire new_AGEMA_signal_5179 ;
    wire new_AGEMA_signal_5180 ;
    wire new_AGEMA_signal_5181 ;
    wire new_AGEMA_signal_5182 ;
    wire new_AGEMA_signal_5183 ;
    wire new_AGEMA_signal_5184 ;
    wire new_AGEMA_signal_5185 ;
    wire new_AGEMA_signal_5186 ;
    wire new_AGEMA_signal_5187 ;
    wire new_AGEMA_signal_5188 ;
    wire new_AGEMA_signal_5189 ;
    wire new_AGEMA_signal_5190 ;
    wire new_AGEMA_signal_5191 ;
    wire new_AGEMA_signal_5192 ;
    wire new_AGEMA_signal_5193 ;
    wire new_AGEMA_signal_5194 ;
    wire new_AGEMA_signal_5195 ;
    wire new_AGEMA_signal_5196 ;
    wire new_AGEMA_signal_5197 ;
    wire new_AGEMA_signal_5198 ;
    wire new_AGEMA_signal_5199 ;
    wire new_AGEMA_signal_5200 ;
    wire new_AGEMA_signal_5201 ;
    wire new_AGEMA_signal_5202 ;
    wire new_AGEMA_signal_5203 ;
    wire new_AGEMA_signal_5204 ;
    wire new_AGEMA_signal_5205 ;
    wire new_AGEMA_signal_5206 ;
    wire new_AGEMA_signal_5207 ;
    wire new_AGEMA_signal_5208 ;
    wire new_AGEMA_signal_5209 ;
    wire new_AGEMA_signal_5210 ;
    wire new_AGEMA_signal_5211 ;
    wire new_AGEMA_signal_5212 ;
    wire new_AGEMA_signal_5213 ;
    wire new_AGEMA_signal_5214 ;
    wire new_AGEMA_signal_5215 ;
    wire new_AGEMA_signal_5216 ;
    wire new_AGEMA_signal_5217 ;
    wire new_AGEMA_signal_5218 ;
    wire new_AGEMA_signal_5219 ;
    wire new_AGEMA_signal_5220 ;
    wire new_AGEMA_signal_5221 ;
    wire new_AGEMA_signal_5222 ;
    wire new_AGEMA_signal_5223 ;
    wire new_AGEMA_signal_5224 ;
    wire new_AGEMA_signal_5225 ;
    wire new_AGEMA_signal_5226 ;
    wire new_AGEMA_signal_5227 ;
    wire new_AGEMA_signal_5228 ;
    wire new_AGEMA_signal_5229 ;
    wire new_AGEMA_signal_5230 ;
    wire new_AGEMA_signal_5231 ;
    wire new_AGEMA_signal_5232 ;
    wire new_AGEMA_signal_5233 ;
    wire new_AGEMA_signal_5234 ;
    wire new_AGEMA_signal_5235 ;
    wire new_AGEMA_signal_5236 ;
    wire new_AGEMA_signal_5237 ;
    wire new_AGEMA_signal_5238 ;
    wire new_AGEMA_signal_5239 ;
    wire new_AGEMA_signal_5240 ;
    wire new_AGEMA_signal_5241 ;
    wire new_AGEMA_signal_5242 ;
    wire new_AGEMA_signal_5243 ;
    wire new_AGEMA_signal_5244 ;
    wire new_AGEMA_signal_5245 ;
    wire new_AGEMA_signal_5246 ;
    wire new_AGEMA_signal_5247 ;
    wire new_AGEMA_signal_5248 ;
    wire new_AGEMA_signal_5249 ;
    wire new_AGEMA_signal_5250 ;
    wire new_AGEMA_signal_5251 ;
    wire new_AGEMA_signal_5252 ;
    wire new_AGEMA_signal_5253 ;
    wire new_AGEMA_signal_5254 ;
    wire new_AGEMA_signal_5255 ;
    wire new_AGEMA_signal_5256 ;
    wire new_AGEMA_signal_5257 ;
    wire new_AGEMA_signal_5258 ;
    wire new_AGEMA_signal_5259 ;
    wire new_AGEMA_signal_5260 ;
    wire new_AGEMA_signal_5261 ;
    wire new_AGEMA_signal_5262 ;
    wire new_AGEMA_signal_5263 ;
    wire new_AGEMA_signal_5264 ;
    wire new_AGEMA_signal_5265 ;
    wire new_AGEMA_signal_5266 ;
    wire new_AGEMA_signal_5267 ;
    wire new_AGEMA_signal_5268 ;
    wire new_AGEMA_signal_5269 ;
    wire new_AGEMA_signal_5270 ;
    wire new_AGEMA_signal_5271 ;
    wire new_AGEMA_signal_5272 ;
    wire new_AGEMA_signal_5273 ;
    wire new_AGEMA_signal_5274 ;
    wire new_AGEMA_signal_5275 ;
    wire new_AGEMA_signal_5276 ;
    wire new_AGEMA_signal_5277 ;
    wire new_AGEMA_signal_5278 ;
    wire new_AGEMA_signal_5279 ;
    wire new_AGEMA_signal_5280 ;
    wire new_AGEMA_signal_5281 ;
    wire new_AGEMA_signal_5282 ;
    wire new_AGEMA_signal_5283 ;
    wire new_AGEMA_signal_5284 ;
    wire new_AGEMA_signal_5285 ;
    wire new_AGEMA_signal_5286 ;
    wire new_AGEMA_signal_5287 ;
    wire new_AGEMA_signal_5288 ;
    wire new_AGEMA_signal_5289 ;
    wire new_AGEMA_signal_5290 ;
    wire new_AGEMA_signal_5291 ;
    wire new_AGEMA_signal_5292 ;
    wire new_AGEMA_signal_5293 ;
    wire new_AGEMA_signal_5294 ;
    wire new_AGEMA_signal_5295 ;
    wire new_AGEMA_signal_5296 ;
    wire new_AGEMA_signal_5297 ;
    wire new_AGEMA_signal_5298 ;
    wire new_AGEMA_signal_5299 ;
    wire new_AGEMA_signal_5300 ;
    wire new_AGEMA_signal_5301 ;
    wire new_AGEMA_signal_5302 ;
    wire new_AGEMA_signal_5303 ;
    wire new_AGEMA_signal_5304 ;
    wire new_AGEMA_signal_5305 ;
    wire new_AGEMA_signal_5306 ;
    wire new_AGEMA_signal_5307 ;
    wire new_AGEMA_signal_5308 ;
    wire new_AGEMA_signal_5309 ;
    wire new_AGEMA_signal_5310 ;
    wire new_AGEMA_signal_5311 ;
    wire new_AGEMA_signal_5312 ;
    wire new_AGEMA_signal_5313 ;
    wire new_AGEMA_signal_5314 ;
    wire new_AGEMA_signal_5315 ;
    wire new_AGEMA_signal_5316 ;
    wire new_AGEMA_signal_5317 ;
    wire new_AGEMA_signal_5318 ;
    wire new_AGEMA_signal_5319 ;
    wire new_AGEMA_signal_5320 ;
    wire new_AGEMA_signal_5321 ;
    wire new_AGEMA_signal_5322 ;
    wire new_AGEMA_signal_5323 ;
    wire new_AGEMA_signal_5324 ;
    wire new_AGEMA_signal_5325 ;
    wire new_AGEMA_signal_5326 ;
    wire new_AGEMA_signal_5327 ;
    wire new_AGEMA_signal_5328 ;
    wire new_AGEMA_signal_5329 ;
    wire new_AGEMA_signal_5330 ;
    wire new_AGEMA_signal_5331 ;
    wire new_AGEMA_signal_5332 ;
    wire new_AGEMA_signal_5333 ;
    wire new_AGEMA_signal_5334 ;
    wire new_AGEMA_signal_5335 ;
    wire new_AGEMA_signal_5336 ;
    wire new_AGEMA_signal_5337 ;
    wire new_AGEMA_signal_5338 ;
    wire new_AGEMA_signal_5339 ;
    wire new_AGEMA_signal_5340 ;
    wire new_AGEMA_signal_5341 ;
    wire new_AGEMA_signal_5342 ;
    wire new_AGEMA_signal_5343 ;
    wire new_AGEMA_signal_5344 ;
    wire new_AGEMA_signal_5345 ;
    wire new_AGEMA_signal_5346 ;
    wire new_AGEMA_signal_5347 ;
    wire new_AGEMA_signal_5348 ;
    wire new_AGEMA_signal_5349 ;
    wire new_AGEMA_signal_5350 ;
    wire new_AGEMA_signal_5351 ;
    wire new_AGEMA_signal_5352 ;
    wire new_AGEMA_signal_5353 ;
    wire new_AGEMA_signal_5354 ;
    wire new_AGEMA_signal_5355 ;
    wire new_AGEMA_signal_5356 ;
    wire new_AGEMA_signal_5357 ;
    wire new_AGEMA_signal_5358 ;
    wire new_AGEMA_signal_5359 ;
    wire new_AGEMA_signal_5360 ;
    wire new_AGEMA_signal_5361 ;
    wire new_AGEMA_signal_5362 ;
    wire new_AGEMA_signal_5363 ;
    wire new_AGEMA_signal_5364 ;
    wire new_AGEMA_signal_5365 ;
    wire new_AGEMA_signal_5366 ;
    wire new_AGEMA_signal_5367 ;
    wire new_AGEMA_signal_5368 ;
    wire new_AGEMA_signal_5369 ;
    wire new_AGEMA_signal_5370 ;
    wire new_AGEMA_signal_5371 ;
    wire new_AGEMA_signal_5372 ;
    wire new_AGEMA_signal_5373 ;
    wire new_AGEMA_signal_5374 ;
    wire new_AGEMA_signal_5375 ;
    wire new_AGEMA_signal_5376 ;
    wire new_AGEMA_signal_5377 ;
    wire new_AGEMA_signal_5378 ;
    wire new_AGEMA_signal_5379 ;
    wire new_AGEMA_signal_5380 ;
    wire new_AGEMA_signal_5381 ;
    wire new_AGEMA_signal_5382 ;
    wire new_AGEMA_signal_5383 ;
    wire new_AGEMA_signal_5384 ;
    wire new_AGEMA_signal_5385 ;
    wire new_AGEMA_signal_5386 ;
    wire new_AGEMA_signal_5387 ;
    wire new_AGEMA_signal_5388 ;
    wire new_AGEMA_signal_5389 ;
    wire new_AGEMA_signal_5390 ;
    wire new_AGEMA_signal_5391 ;
    wire new_AGEMA_signal_5392 ;
    wire new_AGEMA_signal_5393 ;
    wire new_AGEMA_signal_5394 ;
    wire new_AGEMA_signal_5395 ;
    wire new_AGEMA_signal_5396 ;
    wire new_AGEMA_signal_5397 ;
    wire new_AGEMA_signal_5398 ;
    wire new_AGEMA_signal_5399 ;
    wire new_AGEMA_signal_5400 ;
    wire new_AGEMA_signal_5401 ;
    wire new_AGEMA_signal_5402 ;
    wire new_AGEMA_signal_5403 ;
    wire new_AGEMA_signal_5404 ;
    wire new_AGEMA_signal_5405 ;
    wire new_AGEMA_signal_5406 ;
    wire new_AGEMA_signal_5407 ;
    wire new_AGEMA_signal_5408 ;
    wire new_AGEMA_signal_5409 ;
    wire new_AGEMA_signal_5410 ;
    wire new_AGEMA_signal_5411 ;
    wire new_AGEMA_signal_5412 ;
    wire new_AGEMA_signal_5413 ;
    wire new_AGEMA_signal_5414 ;
    wire new_AGEMA_signal_5415 ;
    wire new_AGEMA_signal_5416 ;
    wire new_AGEMA_signal_5417 ;
    wire new_AGEMA_signal_5418 ;
    wire new_AGEMA_signal_5419 ;
    wire new_AGEMA_signal_5420 ;
    wire new_AGEMA_signal_5421 ;
    wire new_AGEMA_signal_5422 ;
    wire new_AGEMA_signal_5423 ;
    wire new_AGEMA_signal_5424 ;
    wire new_AGEMA_signal_5425 ;
    wire new_AGEMA_signal_5426 ;
    wire new_AGEMA_signal_5427 ;
    wire new_AGEMA_signal_5428 ;
    wire new_AGEMA_signal_5429 ;
    wire new_AGEMA_signal_5430 ;
    wire new_AGEMA_signal_5431 ;
    wire new_AGEMA_signal_5432 ;
    wire new_AGEMA_signal_5433 ;
    wire new_AGEMA_signal_5434 ;
    wire new_AGEMA_signal_5435 ;
    wire new_AGEMA_signal_5436 ;
    wire new_AGEMA_signal_5437 ;
    wire new_AGEMA_signal_5438 ;
    wire new_AGEMA_signal_5439 ;
    wire new_AGEMA_signal_5440 ;
    wire new_AGEMA_signal_5441 ;
    wire new_AGEMA_signal_5442 ;
    wire new_AGEMA_signal_5443 ;
    wire new_AGEMA_signal_5444 ;
    wire new_AGEMA_signal_5445 ;
    wire new_AGEMA_signal_5446 ;
    wire new_AGEMA_signal_5447 ;
    wire new_AGEMA_signal_5448 ;
    wire new_AGEMA_signal_5449 ;
    wire new_AGEMA_signal_5450 ;
    wire new_AGEMA_signal_5451 ;
    wire new_AGEMA_signal_5452 ;
    wire new_AGEMA_signal_5453 ;
    wire new_AGEMA_signal_5454 ;
    wire new_AGEMA_signal_5455 ;
    wire new_AGEMA_signal_5456 ;
    wire new_AGEMA_signal_5457 ;
    wire new_AGEMA_signal_5458 ;
    wire new_AGEMA_signal_5459 ;
    wire new_AGEMA_signal_5460 ;
    wire new_AGEMA_signal_5461 ;
    wire new_AGEMA_signal_5462 ;
    wire new_AGEMA_signal_5463 ;
    wire new_AGEMA_signal_5464 ;
    wire new_AGEMA_signal_5465 ;
    wire new_AGEMA_signal_5466 ;
    wire new_AGEMA_signal_5467 ;
    wire new_AGEMA_signal_5468 ;
    wire new_AGEMA_signal_5469 ;
    wire new_AGEMA_signal_5470 ;
    wire new_AGEMA_signal_5471 ;
    wire new_AGEMA_signal_5472 ;
    wire new_AGEMA_signal_5473 ;
    wire new_AGEMA_signal_5474 ;
    wire new_AGEMA_signal_5475 ;
    wire new_AGEMA_signal_5476 ;
    wire new_AGEMA_signal_5477 ;
    wire new_AGEMA_signal_5478 ;
    wire new_AGEMA_signal_5479 ;
    wire new_AGEMA_signal_5480 ;
    wire new_AGEMA_signal_5481 ;
    wire new_AGEMA_signal_5482 ;
    wire new_AGEMA_signal_5483 ;
    wire new_AGEMA_signal_5484 ;
    wire new_AGEMA_signal_5485 ;
    wire new_AGEMA_signal_5486 ;
    wire new_AGEMA_signal_5487 ;
    wire new_AGEMA_signal_5488 ;
    wire new_AGEMA_signal_5489 ;
    wire new_AGEMA_signal_5490 ;
    wire new_AGEMA_signal_5491 ;
    wire new_AGEMA_signal_5492 ;
    wire new_AGEMA_signal_5493 ;
    wire new_AGEMA_signal_5494 ;
    wire new_AGEMA_signal_5495 ;
    wire new_AGEMA_signal_5496 ;
    wire new_AGEMA_signal_5497 ;
    wire new_AGEMA_signal_5498 ;
    wire new_AGEMA_signal_5499 ;
    wire new_AGEMA_signal_5500 ;
    wire new_AGEMA_signal_5501 ;
    wire new_AGEMA_signal_5502 ;
    wire new_AGEMA_signal_5503 ;
    wire new_AGEMA_signal_5504 ;
    wire new_AGEMA_signal_5505 ;
    wire new_AGEMA_signal_5506 ;
    wire new_AGEMA_signal_5507 ;
    wire new_AGEMA_signal_5508 ;
    wire new_AGEMA_signal_5509 ;
    wire new_AGEMA_signal_5510 ;
    wire new_AGEMA_signal_5511 ;
    wire new_AGEMA_signal_5512 ;
    wire new_AGEMA_signal_5513 ;
    wire new_AGEMA_signal_5514 ;
    wire new_AGEMA_signal_5515 ;
    wire new_AGEMA_signal_5516 ;
    wire new_AGEMA_signal_5517 ;
    wire new_AGEMA_signal_5518 ;
    wire new_AGEMA_signal_5519 ;
    wire new_AGEMA_signal_5520 ;
    wire new_AGEMA_signal_5521 ;
    wire new_AGEMA_signal_5522 ;
    wire new_AGEMA_signal_5523 ;
    wire new_AGEMA_signal_5524 ;
    wire new_AGEMA_signal_5525 ;
    wire new_AGEMA_signal_5526 ;
    wire new_AGEMA_signal_5527 ;
    wire new_AGEMA_signal_5528 ;
    wire new_AGEMA_signal_5529 ;
    wire new_AGEMA_signal_5530 ;
    wire new_AGEMA_signal_5531 ;
    wire new_AGEMA_signal_5532 ;
    wire new_AGEMA_signal_5533 ;
    wire new_AGEMA_signal_5534 ;
    wire new_AGEMA_signal_5535 ;
    wire new_AGEMA_signal_5536 ;
    wire new_AGEMA_signal_5537 ;
    wire new_AGEMA_signal_5538 ;
    wire new_AGEMA_signal_5539 ;
    wire new_AGEMA_signal_5540 ;
    wire new_AGEMA_signal_5541 ;
    wire new_AGEMA_signal_5542 ;
    wire new_AGEMA_signal_5543 ;
    wire new_AGEMA_signal_5544 ;
    wire new_AGEMA_signal_5545 ;
    wire new_AGEMA_signal_5546 ;
    wire new_AGEMA_signal_5547 ;
    wire new_AGEMA_signal_5548 ;
    wire new_AGEMA_signal_5549 ;
    wire new_AGEMA_signal_5550 ;
    wire new_AGEMA_signal_5551 ;
    wire new_AGEMA_signal_5552 ;
    wire new_AGEMA_signal_5553 ;
    wire new_AGEMA_signal_5554 ;
    wire new_AGEMA_signal_5555 ;
    wire new_AGEMA_signal_5556 ;
    wire new_AGEMA_signal_5557 ;
    wire new_AGEMA_signal_5558 ;
    wire new_AGEMA_signal_5559 ;
    wire new_AGEMA_signal_5560 ;
    wire new_AGEMA_signal_5561 ;
    wire new_AGEMA_signal_5562 ;
    wire new_AGEMA_signal_5563 ;
    wire new_AGEMA_signal_5564 ;
    wire new_AGEMA_signal_5565 ;
    wire new_AGEMA_signal_5566 ;
    wire new_AGEMA_signal_5567 ;
    wire new_AGEMA_signal_5568 ;
    wire new_AGEMA_signal_5569 ;
    wire new_AGEMA_signal_5570 ;
    wire new_AGEMA_signal_5571 ;
    wire new_AGEMA_signal_5572 ;
    wire new_AGEMA_signal_5573 ;
    wire new_AGEMA_signal_5574 ;
    wire new_AGEMA_signal_5575 ;
    wire new_AGEMA_signal_5576 ;
    wire new_AGEMA_signal_5577 ;
    wire new_AGEMA_signal_5578 ;
    wire new_AGEMA_signal_5579 ;
    wire new_AGEMA_signal_5580 ;
    wire new_AGEMA_signal_5581 ;
    wire new_AGEMA_signal_5582 ;
    wire new_AGEMA_signal_5583 ;
    wire new_AGEMA_signal_5584 ;
    wire new_AGEMA_signal_5585 ;
    wire new_AGEMA_signal_5586 ;
    wire new_AGEMA_signal_5587 ;
    wire new_AGEMA_signal_5588 ;
    wire new_AGEMA_signal_5589 ;
    wire new_AGEMA_signal_5590 ;
    wire new_AGEMA_signal_5591 ;
    wire new_AGEMA_signal_5592 ;
    wire new_AGEMA_signal_5593 ;
    wire new_AGEMA_signal_5594 ;
    wire new_AGEMA_signal_5595 ;
    wire new_AGEMA_signal_5596 ;
    wire new_AGEMA_signal_5597 ;
    wire new_AGEMA_signal_5598 ;
    wire new_AGEMA_signal_5599 ;
    wire new_AGEMA_signal_5600 ;
    wire new_AGEMA_signal_5601 ;
    wire new_AGEMA_signal_5602 ;
    wire new_AGEMA_signal_5603 ;
    wire new_AGEMA_signal_5604 ;
    wire new_AGEMA_signal_5605 ;
    wire new_AGEMA_signal_5606 ;
    wire new_AGEMA_signal_5607 ;
    wire new_AGEMA_signal_5608 ;
    wire new_AGEMA_signal_5609 ;
    wire new_AGEMA_signal_5610 ;
    wire new_AGEMA_signal_5611 ;
    wire new_AGEMA_signal_5612 ;
    wire new_AGEMA_signal_5613 ;
    wire new_AGEMA_signal_5614 ;
    wire new_AGEMA_signal_5615 ;
    wire new_AGEMA_signal_5616 ;
    wire new_AGEMA_signal_5617 ;
    wire new_AGEMA_signal_5618 ;
    wire new_AGEMA_signal_5619 ;
    wire new_AGEMA_signal_5620 ;
    wire new_AGEMA_signal_5621 ;
    wire new_AGEMA_signal_5622 ;
    wire new_AGEMA_signal_5623 ;
    wire new_AGEMA_signal_5624 ;
    wire new_AGEMA_signal_5625 ;
    wire new_AGEMA_signal_5626 ;
    wire new_AGEMA_signal_5627 ;
    wire new_AGEMA_signal_5628 ;
    wire new_AGEMA_signal_5629 ;
    wire new_AGEMA_signal_5630 ;
    wire new_AGEMA_signal_5631 ;
    wire new_AGEMA_signal_5632 ;
    wire new_AGEMA_signal_5633 ;
    wire new_AGEMA_signal_5634 ;
    wire new_AGEMA_signal_5635 ;
    wire new_AGEMA_signal_5636 ;
    wire new_AGEMA_signal_5637 ;
    wire new_AGEMA_signal_5638 ;
    wire new_AGEMA_signal_5639 ;
    wire new_AGEMA_signal_5640 ;
    wire new_AGEMA_signal_5641 ;
    wire new_AGEMA_signal_5642 ;
    wire new_AGEMA_signal_5643 ;
    wire new_AGEMA_signal_5644 ;
    wire new_AGEMA_signal_5645 ;
    wire new_AGEMA_signal_5646 ;
    wire new_AGEMA_signal_5647 ;
    wire new_AGEMA_signal_5648 ;
    wire new_AGEMA_signal_5649 ;
    wire new_AGEMA_signal_5650 ;
    wire new_AGEMA_signal_5651 ;
    wire new_AGEMA_signal_5652 ;
    wire new_AGEMA_signal_5653 ;
    wire new_AGEMA_signal_5654 ;
    wire new_AGEMA_signal_5655 ;
    wire new_AGEMA_signal_5656 ;
    wire new_AGEMA_signal_5657 ;
    wire new_AGEMA_signal_5658 ;
    wire new_AGEMA_signal_5659 ;
    wire new_AGEMA_signal_5660 ;
    wire new_AGEMA_signal_5661 ;
    wire new_AGEMA_signal_5662 ;
    wire new_AGEMA_signal_5663 ;
    wire new_AGEMA_signal_5664 ;
    wire new_AGEMA_signal_5665 ;
    wire new_AGEMA_signal_5666 ;
    wire new_AGEMA_signal_5667 ;
    wire new_AGEMA_signal_5668 ;
    wire new_AGEMA_signal_5669 ;
    wire new_AGEMA_signal_5670 ;
    wire new_AGEMA_signal_5671 ;
    wire new_AGEMA_signal_5672 ;
    wire new_AGEMA_signal_5673 ;
    wire new_AGEMA_signal_5674 ;
    wire new_AGEMA_signal_5675 ;
    wire new_AGEMA_signal_5676 ;
    wire new_AGEMA_signal_5677 ;
    wire new_AGEMA_signal_5678 ;
    wire new_AGEMA_signal_5679 ;
    wire new_AGEMA_signal_5680 ;
    wire new_AGEMA_signal_5681 ;
    wire new_AGEMA_signal_5682 ;
    wire new_AGEMA_signal_5683 ;
    wire new_AGEMA_signal_5684 ;
    wire new_AGEMA_signal_5685 ;
    wire new_AGEMA_signal_5686 ;
    wire new_AGEMA_signal_5687 ;
    wire new_AGEMA_signal_5688 ;
    wire new_AGEMA_signal_5689 ;
    wire new_AGEMA_signal_5690 ;
    wire new_AGEMA_signal_5691 ;
    wire new_AGEMA_signal_5692 ;
    wire new_AGEMA_signal_5693 ;
    wire new_AGEMA_signal_5694 ;
    wire new_AGEMA_signal_5695 ;
    wire new_AGEMA_signal_5696 ;
    wire new_AGEMA_signal_5697 ;
    wire new_AGEMA_signal_5698 ;
    wire new_AGEMA_signal_5699 ;
    wire new_AGEMA_signal_5700 ;
    wire new_AGEMA_signal_5701 ;
    wire new_AGEMA_signal_5702 ;
    wire new_AGEMA_signal_5703 ;
    wire new_AGEMA_signal_5704 ;
    wire new_AGEMA_signal_5705 ;
    wire new_AGEMA_signal_5706 ;
    wire new_AGEMA_signal_5707 ;
    wire new_AGEMA_signal_5708 ;
    wire new_AGEMA_signal_5709 ;
    wire new_AGEMA_signal_5710 ;
    wire new_AGEMA_signal_5711 ;
    wire new_AGEMA_signal_5712 ;
    wire new_AGEMA_signal_5713 ;
    wire new_AGEMA_signal_5714 ;
    wire new_AGEMA_signal_5715 ;
    wire new_AGEMA_signal_5716 ;
    wire new_AGEMA_signal_5717 ;
    wire new_AGEMA_signal_5718 ;
    wire new_AGEMA_signal_5719 ;
    wire new_AGEMA_signal_5720 ;
    wire new_AGEMA_signal_5721 ;
    wire new_AGEMA_signal_5722 ;
    wire new_AGEMA_signal_5723 ;
    wire new_AGEMA_signal_5724 ;
    wire new_AGEMA_signal_5725 ;
    wire new_AGEMA_signal_5726 ;
    wire new_AGEMA_signal_5727 ;
    wire new_AGEMA_signal_5728 ;
    wire new_AGEMA_signal_5729 ;
    wire new_AGEMA_signal_5730 ;
    wire new_AGEMA_signal_5731 ;
    wire new_AGEMA_signal_5732 ;
    wire new_AGEMA_signal_5733 ;
    wire new_AGEMA_signal_5734 ;
    wire new_AGEMA_signal_5735 ;
    wire new_AGEMA_signal_5736 ;
    wire new_AGEMA_signal_5737 ;
    wire new_AGEMA_signal_5738 ;
    wire new_AGEMA_signal_5739 ;
    wire new_AGEMA_signal_5740 ;
    wire new_AGEMA_signal_5741 ;
    wire new_AGEMA_signal_5742 ;
    wire new_AGEMA_signal_5743 ;
    wire new_AGEMA_signal_5744 ;
    wire new_AGEMA_signal_5745 ;
    wire new_AGEMA_signal_5746 ;
    wire new_AGEMA_signal_5747 ;
    wire new_AGEMA_signal_5748 ;
    wire new_AGEMA_signal_5749 ;
    wire new_AGEMA_signal_5750 ;
    wire new_AGEMA_signal_5751 ;
    wire new_AGEMA_signal_5752 ;
    wire new_AGEMA_signal_5753 ;
    wire new_AGEMA_signal_5754 ;
    wire new_AGEMA_signal_5755 ;
    wire new_AGEMA_signal_5756 ;
    wire new_AGEMA_signal_5757 ;
    wire new_AGEMA_signal_5758 ;
    wire new_AGEMA_signal_5759 ;
    wire new_AGEMA_signal_5760 ;
    wire new_AGEMA_signal_5761 ;
    wire new_AGEMA_signal_5762 ;
    wire new_AGEMA_signal_5763 ;
    wire new_AGEMA_signal_5764 ;
    wire new_AGEMA_signal_5765 ;
    wire new_AGEMA_signal_5766 ;
    wire new_AGEMA_signal_5767 ;
    wire new_AGEMA_signal_5768 ;
    wire new_AGEMA_signal_5769 ;
    wire new_AGEMA_signal_5770 ;
    wire new_AGEMA_signal_5771 ;
    wire new_AGEMA_signal_5772 ;
    wire new_AGEMA_signal_5773 ;
    wire new_AGEMA_signal_5774 ;
    wire new_AGEMA_signal_5775 ;
    wire new_AGEMA_signal_5776 ;
    wire new_AGEMA_signal_5777 ;
    wire new_AGEMA_signal_5778 ;
    wire new_AGEMA_signal_5779 ;
    wire new_AGEMA_signal_5780 ;
    wire new_AGEMA_signal_5781 ;
    wire new_AGEMA_signal_5782 ;
    wire new_AGEMA_signal_5783 ;
    wire new_AGEMA_signal_5784 ;
    wire new_AGEMA_signal_5785 ;
    wire new_AGEMA_signal_5786 ;
    wire new_AGEMA_signal_5787 ;
    wire new_AGEMA_signal_5788 ;
    wire new_AGEMA_signal_5789 ;
    wire new_AGEMA_signal_5790 ;
    wire new_AGEMA_signal_5791 ;
    wire new_AGEMA_signal_5792 ;
    wire new_AGEMA_signal_5793 ;
    wire new_AGEMA_signal_5794 ;
    wire new_AGEMA_signal_5795 ;
    wire new_AGEMA_signal_5799 ;
    wire new_AGEMA_signal_5800 ;
    wire new_AGEMA_signal_5801 ;
    wire new_AGEMA_signal_5805 ;
    wire new_AGEMA_signal_5806 ;
    wire new_AGEMA_signal_5807 ;
    wire new_AGEMA_signal_5811 ;
    wire new_AGEMA_signal_5812 ;
    wire new_AGEMA_signal_5813 ;
    wire new_AGEMA_signal_5817 ;
    wire new_AGEMA_signal_5818 ;
    wire new_AGEMA_signal_5819 ;
    wire new_AGEMA_signal_5820 ;
    wire new_AGEMA_signal_5821 ;
    wire new_AGEMA_signal_5822 ;
    wire new_AGEMA_signal_5823 ;
    wire new_AGEMA_signal_5824 ;
    wire new_AGEMA_signal_5825 ;
    wire new_AGEMA_signal_5826 ;
    wire new_AGEMA_signal_5827 ;
    wire new_AGEMA_signal_5828 ;
    wire new_AGEMA_signal_5829 ;
    wire new_AGEMA_signal_5830 ;
    wire new_AGEMA_signal_5831 ;
    wire new_AGEMA_signal_5832 ;
    wire new_AGEMA_signal_5833 ;
    wire new_AGEMA_signal_5834 ;
    wire new_AGEMA_signal_5835 ;
    wire new_AGEMA_signal_5836 ;
    wire new_AGEMA_signal_5837 ;
    wire new_AGEMA_signal_5838 ;
    wire new_AGEMA_signal_5839 ;
    wire new_AGEMA_signal_5840 ;
    wire new_AGEMA_signal_5841 ;
    wire new_AGEMA_signal_5842 ;
    wire new_AGEMA_signal_5843 ;
    wire new_AGEMA_signal_5844 ;
    wire new_AGEMA_signal_5845 ;
    wire new_AGEMA_signal_5846 ;
    wire new_AGEMA_signal_5847 ;
    wire new_AGEMA_signal_5848 ;
    wire new_AGEMA_signal_5849 ;
    wire new_AGEMA_signal_5850 ;
    wire new_AGEMA_signal_5851 ;
    wire new_AGEMA_signal_5852 ;
    wire new_AGEMA_signal_5853 ;
    wire new_AGEMA_signal_5854 ;
    wire new_AGEMA_signal_5855 ;
    wire new_AGEMA_signal_5856 ;
    wire new_AGEMA_signal_5857 ;
    wire new_AGEMA_signal_5858 ;
    wire new_AGEMA_signal_5859 ;
    wire new_AGEMA_signal_5860 ;
    wire new_AGEMA_signal_5861 ;
    wire new_AGEMA_signal_5862 ;
    wire new_AGEMA_signal_5863 ;
    wire new_AGEMA_signal_5864 ;
    wire new_AGEMA_signal_5865 ;
    wire new_AGEMA_signal_5866 ;
    wire new_AGEMA_signal_5867 ;
    wire new_AGEMA_signal_5868 ;
    wire new_AGEMA_signal_5869 ;
    wire new_AGEMA_signal_5870 ;
    wire new_AGEMA_signal_5871 ;
    wire new_AGEMA_signal_5872 ;
    wire new_AGEMA_signal_5873 ;
    wire new_AGEMA_signal_5874 ;
    wire new_AGEMA_signal_5875 ;
    wire new_AGEMA_signal_5876 ;
    wire new_AGEMA_signal_5877 ;
    wire new_AGEMA_signal_5878 ;
    wire new_AGEMA_signal_5879 ;
    wire new_AGEMA_signal_5880 ;
    wire new_AGEMA_signal_5881 ;
    wire new_AGEMA_signal_5882 ;
    wire new_AGEMA_signal_5883 ;
    wire new_AGEMA_signal_5884 ;
    wire new_AGEMA_signal_5885 ;
    wire new_AGEMA_signal_5886 ;
    wire new_AGEMA_signal_5887 ;
    wire new_AGEMA_signal_5888 ;
    wire new_AGEMA_signal_5889 ;
    wire new_AGEMA_signal_5890 ;
    wire new_AGEMA_signal_5891 ;
    wire new_AGEMA_signal_5892 ;
    wire new_AGEMA_signal_5893 ;
    wire new_AGEMA_signal_5894 ;
    wire new_AGEMA_signal_5895 ;
    wire new_AGEMA_signal_5896 ;
    wire new_AGEMA_signal_5897 ;
    wire new_AGEMA_signal_5898 ;
    wire new_AGEMA_signal_5899 ;
    wire new_AGEMA_signal_5900 ;
    wire new_AGEMA_signal_5901 ;
    wire new_AGEMA_signal_5902 ;
    wire new_AGEMA_signal_5903 ;
    wire new_AGEMA_signal_5904 ;
    wire new_AGEMA_signal_5905 ;
    wire new_AGEMA_signal_5906 ;
    wire new_AGEMA_signal_5907 ;
    wire new_AGEMA_signal_5908 ;
    wire new_AGEMA_signal_5909 ;
    wire new_AGEMA_signal_5910 ;
    wire new_AGEMA_signal_5911 ;
    wire new_AGEMA_signal_5912 ;
    wire new_AGEMA_signal_5913 ;
    wire new_AGEMA_signal_5914 ;
    wire new_AGEMA_signal_5915 ;
    wire new_AGEMA_signal_5916 ;
    wire new_AGEMA_signal_5917 ;
    wire new_AGEMA_signal_5918 ;
    wire new_AGEMA_signal_5919 ;
    wire new_AGEMA_signal_5920 ;
    wire new_AGEMA_signal_5921 ;
    wire new_AGEMA_signal_5922 ;
    wire new_AGEMA_signal_5923 ;
    wire new_AGEMA_signal_5924 ;
    wire new_AGEMA_signal_5925 ;
    wire new_AGEMA_signal_5926 ;
    wire new_AGEMA_signal_5927 ;
    wire new_AGEMA_signal_5928 ;
    wire new_AGEMA_signal_5929 ;
    wire new_AGEMA_signal_5930 ;
    wire new_AGEMA_signal_5931 ;
    wire new_AGEMA_signal_5932 ;
    wire new_AGEMA_signal_5933 ;
    wire new_AGEMA_signal_5934 ;
    wire new_AGEMA_signal_5935 ;
    wire new_AGEMA_signal_5936 ;
    wire new_AGEMA_signal_5937 ;
    wire new_AGEMA_signal_5938 ;
    wire new_AGEMA_signal_5939 ;
    wire new_AGEMA_signal_5940 ;
    wire new_AGEMA_signal_5941 ;
    wire new_AGEMA_signal_5942 ;
    wire new_AGEMA_signal_5943 ;
    wire new_AGEMA_signal_5944 ;
    wire new_AGEMA_signal_5945 ;
    wire new_AGEMA_signal_5946 ;
    wire new_AGEMA_signal_5947 ;
    wire new_AGEMA_signal_5948 ;
    wire new_AGEMA_signal_5949 ;
    wire new_AGEMA_signal_5950 ;
    wire new_AGEMA_signal_5951 ;
    wire new_AGEMA_signal_5952 ;
    wire new_AGEMA_signal_5953 ;
    wire new_AGEMA_signal_5954 ;
    wire new_AGEMA_signal_5955 ;
    wire new_AGEMA_signal_5956 ;
    wire new_AGEMA_signal_5957 ;
    wire new_AGEMA_signal_5958 ;
    wire new_AGEMA_signal_5959 ;
    wire new_AGEMA_signal_5960 ;
    wire new_AGEMA_signal_5961 ;
    wire new_AGEMA_signal_5962 ;
    wire new_AGEMA_signal_5963 ;
    wire new_AGEMA_signal_5964 ;
    wire new_AGEMA_signal_5965 ;
    wire new_AGEMA_signal_5966 ;
    wire new_AGEMA_signal_5967 ;
    wire new_AGEMA_signal_5968 ;
    wire new_AGEMA_signal_5969 ;
    wire new_AGEMA_signal_5970 ;
    wire new_AGEMA_signal_5971 ;
    wire new_AGEMA_signal_5972 ;
    wire new_AGEMA_signal_5973 ;
    wire new_AGEMA_signal_5974 ;
    wire new_AGEMA_signal_5975 ;
    wire new_AGEMA_signal_5976 ;
    wire new_AGEMA_signal_5977 ;
    wire new_AGEMA_signal_5978 ;
    wire new_AGEMA_signal_5979 ;
    wire new_AGEMA_signal_5980 ;
    wire new_AGEMA_signal_5981 ;
    wire new_AGEMA_signal_5982 ;
    wire new_AGEMA_signal_5983 ;
    wire new_AGEMA_signal_5984 ;
    wire new_AGEMA_signal_5985 ;
    wire new_AGEMA_signal_5986 ;
    wire new_AGEMA_signal_5987 ;
    wire new_AGEMA_signal_5988 ;
    wire new_AGEMA_signal_5989 ;
    wire new_AGEMA_signal_5990 ;
    wire new_AGEMA_signal_5991 ;
    wire new_AGEMA_signal_5992 ;
    wire new_AGEMA_signal_5993 ;
    wire new_AGEMA_signal_5994 ;
    wire new_AGEMA_signal_5995 ;
    wire new_AGEMA_signal_5996 ;
    wire new_AGEMA_signal_5997 ;
    wire new_AGEMA_signal_5998 ;
    wire new_AGEMA_signal_5999 ;
    wire new_AGEMA_signal_6000 ;
    wire new_AGEMA_signal_6001 ;
    wire new_AGEMA_signal_6002 ;
    wire new_AGEMA_signal_6006 ;
    wire new_AGEMA_signal_6007 ;
    wire new_AGEMA_signal_6008 ;
    wire new_AGEMA_signal_6012 ;
    wire new_AGEMA_signal_6013 ;
    wire new_AGEMA_signal_6014 ;
    wire new_AGEMA_signal_6018 ;
    wire new_AGEMA_signal_6019 ;
    wire new_AGEMA_signal_6020 ;
    wire new_AGEMA_signal_6021 ;
    wire new_AGEMA_signal_6022 ;
    wire new_AGEMA_signal_6023 ;
    wire new_AGEMA_signal_6027 ;
    wire new_AGEMA_signal_6028 ;
    wire new_AGEMA_signal_6029 ;
    wire new_AGEMA_signal_6033 ;
    wire new_AGEMA_signal_6034 ;
    wire new_AGEMA_signal_6035 ;
    wire new_AGEMA_signal_6039 ;
    wire new_AGEMA_signal_6040 ;
    wire new_AGEMA_signal_6041 ;
    wire new_AGEMA_signal_6042 ;
    wire new_AGEMA_signal_6043 ;
    wire new_AGEMA_signal_6044 ;
    wire new_AGEMA_signal_6048 ;
    wire new_AGEMA_signal_6049 ;
    wire new_AGEMA_signal_6050 ;
    wire new_AGEMA_signal_6054 ;
    wire new_AGEMA_signal_6055 ;
    wire new_AGEMA_signal_6056 ;
    wire new_AGEMA_signal_6060 ;
    wire new_AGEMA_signal_6061 ;
    wire new_AGEMA_signal_6062 ;
    wire new_AGEMA_signal_6063 ;
    wire new_AGEMA_signal_6064 ;
    wire new_AGEMA_signal_6065 ;
    wire new_AGEMA_signal_6066 ;
    wire new_AGEMA_signal_6067 ;
    wire new_AGEMA_signal_6068 ;
    wire new_AGEMA_signal_6069 ;
    wire new_AGEMA_signal_6070 ;
    wire new_AGEMA_signal_6071 ;
    wire new_AGEMA_signal_6072 ;
    wire new_AGEMA_signal_6073 ;
    wire new_AGEMA_signal_6074 ;
    wire new_AGEMA_signal_6075 ;
    wire new_AGEMA_signal_6076 ;
    wire new_AGEMA_signal_6077 ;
    wire new_AGEMA_signal_6078 ;
    wire new_AGEMA_signal_6079 ;
    wire new_AGEMA_signal_6080 ;
    wire new_AGEMA_signal_6081 ;
    wire new_AGEMA_signal_6082 ;
    wire new_AGEMA_signal_6083 ;
    wire new_AGEMA_signal_6084 ;
    wire new_AGEMA_signal_6085 ;
    wire new_AGEMA_signal_6086 ;
    wire new_AGEMA_signal_6087 ;
    wire new_AGEMA_signal_6088 ;
    wire new_AGEMA_signal_6089 ;
    wire new_AGEMA_signal_6090 ;
    wire new_AGEMA_signal_6091 ;
    wire new_AGEMA_signal_6092 ;
    wire new_AGEMA_signal_6093 ;
    wire new_AGEMA_signal_6094 ;
    wire new_AGEMA_signal_6095 ;
    wire new_AGEMA_signal_6096 ;
    wire new_AGEMA_signal_6097 ;
    wire new_AGEMA_signal_6098 ;
    wire new_AGEMA_signal_6099 ;
    wire new_AGEMA_signal_6100 ;
    wire new_AGEMA_signal_6101 ;
    wire new_AGEMA_signal_6102 ;
    wire new_AGEMA_signal_6103 ;
    wire new_AGEMA_signal_6104 ;
    wire new_AGEMA_signal_6105 ;
    wire new_AGEMA_signal_6106 ;
    wire new_AGEMA_signal_6107 ;
    wire new_AGEMA_signal_6108 ;
    wire new_AGEMA_signal_6109 ;
    wire new_AGEMA_signal_6110 ;
    wire new_AGEMA_signal_6111 ;
    wire new_AGEMA_signal_6112 ;
    wire new_AGEMA_signal_6113 ;
    wire new_AGEMA_signal_6114 ;
    wire new_AGEMA_signal_6115 ;
    wire new_AGEMA_signal_6116 ;
    wire new_AGEMA_signal_6117 ;
    wire new_AGEMA_signal_6118 ;
    wire new_AGEMA_signal_6119 ;
    wire new_AGEMA_signal_6120 ;
    wire new_AGEMA_signal_6121 ;
    wire new_AGEMA_signal_6122 ;
    wire new_AGEMA_signal_6123 ;
    wire new_AGEMA_signal_6124 ;
    wire new_AGEMA_signal_6125 ;
    wire new_AGEMA_signal_6126 ;
    wire new_AGEMA_signal_6127 ;
    wire new_AGEMA_signal_6128 ;
    wire new_AGEMA_signal_6129 ;
    wire new_AGEMA_signal_6130 ;
    wire new_AGEMA_signal_6131 ;
    wire new_AGEMA_signal_6132 ;
    wire new_AGEMA_signal_6133 ;
    wire new_AGEMA_signal_6134 ;
    wire new_AGEMA_signal_6135 ;
    wire new_AGEMA_signal_6136 ;
    wire new_AGEMA_signal_6137 ;
    wire new_AGEMA_signal_6138 ;
    wire new_AGEMA_signal_6139 ;
    wire new_AGEMA_signal_6140 ;
    wire new_AGEMA_signal_6141 ;
    wire new_AGEMA_signal_6142 ;
    wire new_AGEMA_signal_6143 ;
    wire new_AGEMA_signal_6144 ;
    wire new_AGEMA_signal_6145 ;
    wire new_AGEMA_signal_6146 ;
    wire new_AGEMA_signal_6147 ;
    wire new_AGEMA_signal_6148 ;
    wire new_AGEMA_signal_6149 ;
    wire new_AGEMA_signal_6150 ;
    wire new_AGEMA_signal_6151 ;
    wire new_AGEMA_signal_6152 ;
    wire new_AGEMA_signal_6153 ;
    wire new_AGEMA_signal_6154 ;
    wire new_AGEMA_signal_6155 ;
    wire new_AGEMA_signal_6159 ;
    wire new_AGEMA_signal_6160 ;
    wire new_AGEMA_signal_6161 ;
    wire new_AGEMA_signal_6165 ;
    wire new_AGEMA_signal_6166 ;
    wire new_AGEMA_signal_6167 ;
    wire new_AGEMA_signal_6168 ;
    wire new_AGEMA_signal_6169 ;
    wire new_AGEMA_signal_6170 ;
    wire new_AGEMA_signal_6174 ;
    wire new_AGEMA_signal_6175 ;
    wire new_AGEMA_signal_6176 ;
    wire new_AGEMA_signal_6177 ;
    wire new_AGEMA_signal_6178 ;
    wire new_AGEMA_signal_6179 ;
    wire new_AGEMA_signal_6180 ;
    wire new_AGEMA_signal_6181 ;
    wire new_AGEMA_signal_6182 ;
    wire new_AGEMA_signal_6186 ;
    wire new_AGEMA_signal_6187 ;
    wire new_AGEMA_signal_6188 ;
    wire new_AGEMA_signal_6189 ;
    wire new_AGEMA_signal_6190 ;
    wire new_AGEMA_signal_6191 ;
    wire new_AGEMA_signal_6192 ;
    wire new_AGEMA_signal_6193 ;
    wire new_AGEMA_signal_6194 ;
    wire new_AGEMA_signal_6195 ;
    wire new_AGEMA_signal_6196 ;
    wire new_AGEMA_signal_6197 ;
    wire new_AGEMA_signal_6198 ;
    wire new_AGEMA_signal_6199 ;
    wire new_AGEMA_signal_6200 ;
    wire new_AGEMA_signal_6204 ;
    wire new_AGEMA_signal_6205 ;
    wire new_AGEMA_signal_6206 ;
    wire new_AGEMA_signal_6210 ;
    wire new_AGEMA_signal_6211 ;
    wire new_AGEMA_signal_6212 ;
    wire new_AGEMA_signal_6213 ;
    wire new_AGEMA_signal_6214 ;
    wire new_AGEMA_signal_6215 ;
    wire new_AGEMA_signal_6219 ;
    wire new_AGEMA_signal_6220 ;
    wire new_AGEMA_signal_6221 ;
    wire new_AGEMA_signal_6225 ;
    wire new_AGEMA_signal_6226 ;
    wire new_AGEMA_signal_6227 ;
    wire new_AGEMA_signal_6231 ;
    wire new_AGEMA_signal_6232 ;
    wire new_AGEMA_signal_6233 ;
    wire new_AGEMA_signal_6237 ;
    wire new_AGEMA_signal_6238 ;
    wire new_AGEMA_signal_6239 ;
    wire new_AGEMA_signal_6243 ;
    wire new_AGEMA_signal_6244 ;
    wire new_AGEMA_signal_6245 ;
    wire new_AGEMA_signal_6249 ;
    wire new_AGEMA_signal_6250 ;
    wire new_AGEMA_signal_6251 ;
    wire new_AGEMA_signal_6255 ;
    wire new_AGEMA_signal_6256 ;
    wire new_AGEMA_signal_6257 ;
    wire new_AGEMA_signal_6261 ;
    wire new_AGEMA_signal_6262 ;
    wire new_AGEMA_signal_6263 ;
    wire new_AGEMA_signal_6267 ;
    wire new_AGEMA_signal_6268 ;
    wire new_AGEMA_signal_6269 ;
    wire new_AGEMA_signal_6273 ;
    wire new_AGEMA_signal_6274 ;
    wire new_AGEMA_signal_6275 ;
    wire new_AGEMA_signal_6279 ;
    wire new_AGEMA_signal_6280 ;
    wire new_AGEMA_signal_6281 ;
    wire new_AGEMA_signal_6285 ;
    wire new_AGEMA_signal_6286 ;
    wire new_AGEMA_signal_6287 ;
    wire new_AGEMA_signal_6288 ;
    wire new_AGEMA_signal_6289 ;
    wire new_AGEMA_signal_6290 ;
    wire new_AGEMA_signal_6294 ;
    wire new_AGEMA_signal_6295 ;
    wire new_AGEMA_signal_6296 ;
    wire new_AGEMA_signal_6300 ;
    wire new_AGEMA_signal_6301 ;
    wire new_AGEMA_signal_6302 ;
    wire new_AGEMA_signal_6306 ;
    wire new_AGEMA_signal_6307 ;
    wire new_AGEMA_signal_6308 ;
    wire new_AGEMA_signal_6309 ;
    wire new_AGEMA_signal_6310 ;
    wire new_AGEMA_signal_6311 ;
    wire new_AGEMA_signal_6312 ;
    wire new_AGEMA_signal_6313 ;
    wire new_AGEMA_signal_6314 ;
    wire new_AGEMA_signal_6315 ;
    wire new_AGEMA_signal_6316 ;
    wire new_AGEMA_signal_6317 ;
    wire new_AGEMA_signal_6318 ;
    wire new_AGEMA_signal_6319 ;
    wire new_AGEMA_signal_6320 ;
    wire new_AGEMA_signal_6321 ;
    wire new_AGEMA_signal_6322 ;
    wire new_AGEMA_signal_6323 ;
    wire new_AGEMA_signal_6324 ;
    wire new_AGEMA_signal_6325 ;
    wire new_AGEMA_signal_6326 ;
    wire new_AGEMA_signal_6327 ;
    wire new_AGEMA_signal_6328 ;
    wire new_AGEMA_signal_6329 ;
    wire new_AGEMA_signal_6330 ;
    wire new_AGEMA_signal_6331 ;
    wire new_AGEMA_signal_6332 ;
    wire new_AGEMA_signal_6333 ;
    wire new_AGEMA_signal_6334 ;
    wire new_AGEMA_signal_6335 ;
    wire new_AGEMA_signal_6336 ;
    wire new_AGEMA_signal_6337 ;
    wire new_AGEMA_signal_6338 ;
    wire new_AGEMA_signal_6339 ;
    wire new_AGEMA_signal_6340 ;
    wire new_AGEMA_signal_6341 ;
    wire new_AGEMA_signal_6342 ;
    wire new_AGEMA_signal_6343 ;
    wire new_AGEMA_signal_6344 ;
    wire new_AGEMA_signal_6345 ;
    wire new_AGEMA_signal_6346 ;
    wire new_AGEMA_signal_6347 ;
    wire new_AGEMA_signal_6351 ;
    wire new_AGEMA_signal_6352 ;
    wire new_AGEMA_signal_6353 ;
    wire new_AGEMA_signal_6357 ;
    wire new_AGEMA_signal_6358 ;
    wire new_AGEMA_signal_6359 ;
    wire new_AGEMA_signal_6360 ;
    wire new_AGEMA_signal_6361 ;
    wire new_AGEMA_signal_6362 ;
    wire new_AGEMA_signal_6366 ;
    wire new_AGEMA_signal_6367 ;
    wire new_AGEMA_signal_6368 ;
    wire new_AGEMA_signal_6372 ;
    wire new_AGEMA_signal_6373 ;
    wire new_AGEMA_signal_6374 ;
    wire new_AGEMA_signal_6375 ;
    wire new_AGEMA_signal_6376 ;
    wire new_AGEMA_signal_6377 ;
    wire new_AGEMA_signal_6381 ;
    wire new_AGEMA_signal_6382 ;
    wire new_AGEMA_signal_6383 ;
    wire new_AGEMA_signal_6387 ;
    wire new_AGEMA_signal_6388 ;
    wire new_AGEMA_signal_6389 ;
    wire new_AGEMA_signal_6390 ;
    wire new_AGEMA_signal_6391 ;
    wire new_AGEMA_signal_6392 ;
    wire new_AGEMA_signal_6393 ;
    wire new_AGEMA_signal_6394 ;
    wire new_AGEMA_signal_6395 ;
    wire new_AGEMA_signal_6399 ;
    wire new_AGEMA_signal_6400 ;
    wire new_AGEMA_signal_6401 ;
    wire new_AGEMA_signal_6405 ;
    wire new_AGEMA_signal_6406 ;
    wire new_AGEMA_signal_6407 ;
    wire new_AGEMA_signal_6408 ;
    wire new_AGEMA_signal_6409 ;
    wire new_AGEMA_signal_6410 ;
    wire new_AGEMA_signal_6411 ;
    wire new_AGEMA_signal_6412 ;
    wire new_AGEMA_signal_6413 ;
    wire new_AGEMA_signal_6417 ;
    wire new_AGEMA_signal_6418 ;
    wire new_AGEMA_signal_6419 ;
    wire new_AGEMA_signal_6420 ;
    wire new_AGEMA_signal_6421 ;
    wire new_AGEMA_signal_6422 ;
    wire new_AGEMA_signal_6423 ;
    wire new_AGEMA_signal_6424 ;
    wire new_AGEMA_signal_6425 ;
    wire new_AGEMA_signal_6429 ;
    wire new_AGEMA_signal_6430 ;
    wire new_AGEMA_signal_6431 ;
    wire new_AGEMA_signal_6432 ;
    wire new_AGEMA_signal_6433 ;
    wire new_AGEMA_signal_6434 ;
    wire new_AGEMA_signal_6438 ;
    wire new_AGEMA_signal_6439 ;
    wire new_AGEMA_signal_6440 ;
    wire new_AGEMA_signal_6444 ;
    wire new_AGEMA_signal_6445 ;
    wire new_AGEMA_signal_6446 ;
    wire new_AGEMA_signal_6447 ;
    wire new_AGEMA_signal_6448 ;
    wire new_AGEMA_signal_6449 ;
    wire new_AGEMA_signal_6450 ;
    wire new_AGEMA_signal_6451 ;
    wire new_AGEMA_signal_6452 ;
    wire new_AGEMA_signal_6456 ;
    wire new_AGEMA_signal_6457 ;
    wire new_AGEMA_signal_6458 ;
    wire new_AGEMA_signal_6462 ;
    wire new_AGEMA_signal_6463 ;
    wire new_AGEMA_signal_6464 ;
    wire new_AGEMA_signal_6468 ;
    wire new_AGEMA_signal_6469 ;
    wire new_AGEMA_signal_6470 ;
    wire new_AGEMA_signal_6474 ;
    wire new_AGEMA_signal_6475 ;
    wire new_AGEMA_signal_6476 ;
    wire new_AGEMA_signal_6477 ;
    wire new_AGEMA_signal_6478 ;
    wire new_AGEMA_signal_6479 ;
    wire new_AGEMA_signal_6480 ;
    wire new_AGEMA_signal_6481 ;
    wire new_AGEMA_signal_6482 ;
    wire new_AGEMA_signal_6486 ;
    wire new_AGEMA_signal_6487 ;
    wire new_AGEMA_signal_6488 ;
    wire new_AGEMA_signal_6492 ;
    wire new_AGEMA_signal_6493 ;
    wire new_AGEMA_signal_6494 ;
    wire new_AGEMA_signal_6495 ;
    wire new_AGEMA_signal_6496 ;
    wire new_AGEMA_signal_6497 ;
    wire new_AGEMA_signal_6501 ;
    wire new_AGEMA_signal_6502 ;
    wire new_AGEMA_signal_6503 ;
    wire new_AGEMA_signal_6504 ;
    wire new_AGEMA_signal_6505 ;
    wire new_AGEMA_signal_6506 ;
    wire new_AGEMA_signal_6510 ;
    wire new_AGEMA_signal_6511 ;
    wire new_AGEMA_signal_6512 ;
    wire new_AGEMA_signal_6516 ;
    wire new_AGEMA_signal_6517 ;
    wire new_AGEMA_signal_6518 ;
    wire new_AGEMA_signal_6519 ;
    wire new_AGEMA_signal_6520 ;
    wire new_AGEMA_signal_6521 ;
    wire new_AGEMA_signal_6522 ;
    wire new_AGEMA_signal_6523 ;
    wire new_AGEMA_signal_6524 ;
    wire new_AGEMA_signal_6525 ;
    wire new_AGEMA_signal_6526 ;
    wire new_AGEMA_signal_6527 ;
    wire new_AGEMA_signal_6528 ;
    wire new_AGEMA_signal_6529 ;
    wire new_AGEMA_signal_6530 ;
    wire new_AGEMA_signal_6531 ;
    wire new_AGEMA_signal_6532 ;
    wire new_AGEMA_signal_6533 ;
    wire new_AGEMA_signal_6534 ;
    wire new_AGEMA_signal_6535 ;
    wire new_AGEMA_signal_6536 ;
    wire new_AGEMA_signal_6537 ;
    wire new_AGEMA_signal_6538 ;
    wire new_AGEMA_signal_6539 ;
    wire new_AGEMA_signal_6540 ;
    wire new_AGEMA_signal_6541 ;
    wire new_AGEMA_signal_6542 ;
    wire new_AGEMA_signal_6543 ;
    wire new_AGEMA_signal_6544 ;
    wire new_AGEMA_signal_6545 ;
    wire new_AGEMA_signal_6546 ;
    wire new_AGEMA_signal_6547 ;
    wire new_AGEMA_signal_6548 ;
    wire new_AGEMA_signal_6549 ;
    wire new_AGEMA_signal_6550 ;
    wire new_AGEMA_signal_6551 ;
    wire new_AGEMA_signal_6555 ;
    wire new_AGEMA_signal_6556 ;
    wire new_AGEMA_signal_6557 ;
    wire new_AGEMA_signal_6561 ;
    wire new_AGEMA_signal_6562 ;
    wire new_AGEMA_signal_6563 ;
    wire new_AGEMA_signal_6567 ;
    wire new_AGEMA_signal_6568 ;
    wire new_AGEMA_signal_6569 ;
    wire new_AGEMA_signal_6570 ;
    wire new_AGEMA_signal_6571 ;
    wire new_AGEMA_signal_6572 ;
    wire new_AGEMA_signal_6576 ;
    wire new_AGEMA_signal_6577 ;
    wire new_AGEMA_signal_6578 ;
    wire new_AGEMA_signal_6579 ;
    wire new_AGEMA_signal_6580 ;
    wire new_AGEMA_signal_6581 ;
    wire new_AGEMA_signal_6582 ;
    wire new_AGEMA_signal_6583 ;
    wire new_AGEMA_signal_6584 ;
    wire new_AGEMA_signal_6588 ;
    wire new_AGEMA_signal_6589 ;
    wire new_AGEMA_signal_6590 ;
    wire new_AGEMA_signal_6591 ;
    wire new_AGEMA_signal_6592 ;
    wire new_AGEMA_signal_6593 ;
    wire new_AGEMA_signal_6597 ;
    wire new_AGEMA_signal_6598 ;
    wire new_AGEMA_signal_6599 ;
    wire new_AGEMA_signal_6600 ;
    wire new_AGEMA_signal_6601 ;
    wire new_AGEMA_signal_6602 ;
    wire new_AGEMA_signal_6603 ;
    wire new_AGEMA_signal_6604 ;
    wire new_AGEMA_signal_6605 ;
    wire new_AGEMA_signal_6606 ;
    wire new_AGEMA_signal_6607 ;
    wire new_AGEMA_signal_6608 ;
    wire new_AGEMA_signal_6609 ;
    wire new_AGEMA_signal_6610 ;
    wire new_AGEMA_signal_6611 ;
    wire new_AGEMA_signal_6612 ;
    wire new_AGEMA_signal_6613 ;
    wire new_AGEMA_signal_6614 ;
    wire new_AGEMA_signal_6615 ;
    wire new_AGEMA_signal_6616 ;
    wire new_AGEMA_signal_6617 ;
    wire new_AGEMA_signal_6621 ;
    wire new_AGEMA_signal_6622 ;
    wire new_AGEMA_signal_6623 ;
    wire new_AGEMA_signal_6627 ;
    wire new_AGEMA_signal_6628 ;
    wire new_AGEMA_signal_6629 ;
    wire new_AGEMA_signal_6630 ;
    wire new_AGEMA_signal_6631 ;
    wire new_AGEMA_signal_6632 ;
    wire new_AGEMA_signal_6633 ;
    wire new_AGEMA_signal_6634 ;
    wire new_AGEMA_signal_6635 ;
    wire new_AGEMA_signal_6636 ;
    wire new_AGEMA_signal_6637 ;
    wire new_AGEMA_signal_6638 ;
    wire new_AGEMA_signal_6639 ;
    wire new_AGEMA_signal_6640 ;
    wire new_AGEMA_signal_6641 ;
    wire new_AGEMA_signal_6642 ;
    wire new_AGEMA_signal_6643 ;
    wire new_AGEMA_signal_6644 ;
    wire new_AGEMA_signal_6645 ;
    wire new_AGEMA_signal_6646 ;
    wire new_AGEMA_signal_6647 ;
    wire new_AGEMA_signal_6648 ;
    wire new_AGEMA_signal_6649 ;
    wire new_AGEMA_signal_6650 ;
    wire new_AGEMA_signal_6651 ;
    wire new_AGEMA_signal_6652 ;
    wire new_AGEMA_signal_6653 ;
    wire new_AGEMA_signal_6657 ;
    wire new_AGEMA_signal_6658 ;
    wire new_AGEMA_signal_6659 ;
    wire new_AGEMA_signal_6660 ;
    wire new_AGEMA_signal_6661 ;
    wire new_AGEMA_signal_6662 ;
    wire new_AGEMA_signal_6663 ;
    wire new_AGEMA_signal_6664 ;
    wire new_AGEMA_signal_6665 ;
    wire new_AGEMA_signal_6666 ;
    wire new_AGEMA_signal_6667 ;
    wire new_AGEMA_signal_6668 ;
    wire new_AGEMA_signal_6669 ;
    wire new_AGEMA_signal_6670 ;
    wire new_AGEMA_signal_6671 ;

    /* cells in depth 0 */
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) U16 ( .A0_t (roundconstant[5]), .A0_f (new_AGEMA_signal_1877), .B0_t (roundconstant[1]), .B0_f (new_AGEMA_signal_1878), .Z0_t (n15), .Z0_f (new_AGEMA_signal_1879) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) U17 ( .A0_t (roundconstant[0]), .A0_f (new_AGEMA_signal_1888), .B0_t (n15), .B0_f (new_AGEMA_signal_1879), .Z0_t (n16), .Z0_f (new_AGEMA_signal_2470) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) U18 ( .A0_t (roundconstant[2]), .A0_f (new_AGEMA_signal_1887), .B0_t (n16), .B0_f (new_AGEMA_signal_2470), .Z0_t (n17), .Z0_f (new_AGEMA_signal_2474) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) U19 ( .A0_t (roundconstant[3]), .A0_f (new_AGEMA_signal_1880), .B0_t (n17), .B0_f (new_AGEMA_signal_2474), .Z0_t (n18), .Z0_f (new_AGEMA_signal_2478) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) U20 ( .A0_t (roundconstant[4]), .A0_f (new_AGEMA_signal_1882), .B0_t (n18), .B0_f (new_AGEMA_signal_2478), .Z0_t (n19), .Z0_f (new_AGEMA_signal_2673) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) U21 ( .A0_t (OUT_done_t), .A0_f (OUT_done_f), .B0_t (n19), .B0_f (new_AGEMA_signal_2673), .Z0_t (n20), .Z0_f (new_AGEMA_signal_2867) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) U22 ( .A0_t (IN_reset_t), .A0_f (IN_reset_f), .B0_t (n20), .B0_f (new_AGEMA_signal_2867), .Z0_t (OUT_done_t), .Z0_f (OUT_done_f) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) LED_128_Instance_U31 ( .A0_t (roundconstant[3]), .A0_f (new_AGEMA_signal_1880), .B0_t (IN_reset_t), .B0_f (IN_reset_f), .Z0_t (roundconstant[4]), .Z0_f (new_AGEMA_signal_1882) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) LED_128_Instance_U30 ( .A0_t (IN_reset_t), .A0_f (IN_reset_f), .B0_t (LED_128_Instance_n24), .B0_f (new_AGEMA_signal_1883), .Z0_t (LED_128_Instance_ks_reg_2__Q), .Z0_f (new_AGEMA_signal_1884) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) LED_128_Instance_U29 ( .A0_t (IN_reset_t), .A0_f (IN_reset_f), .B0_t (LED_128_Instance_ks_0), .B0_f (new_AGEMA_signal_1885), .Z0_t (LED_128_Instance_n24), .Z0_f (new_AGEMA_signal_1883) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) LED_128_Instance_U28 ( .A0_t (IN_reset_t), .A0_f (IN_reset_f), .B0_t (LED_128_Instance_ks_3_), .B0_f (new_AGEMA_signal_1886), .Z0_t (LED_128_Instance_ks_0), .Z0_f (new_AGEMA_signal_1885) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) LED_128_Instance_U27 ( .A0_t (roundconstant[4]), .A0_f (new_AGEMA_signal_1882), .B0_t (IN_reset_t), .B0_f (IN_reset_f), .Z0_t (roundconstant[5]), .Z0_f (new_AGEMA_signal_1877) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) LED_128_Instance_U26 ( .A0_t (roundconstant[2]), .A0_f (new_AGEMA_signal_1887), .B0_t (IN_reset_t), .B0_f (IN_reset_f), .Z0_t (roundconstant[3]), .Z0_f (new_AGEMA_signal_1880) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) LED_128_Instance_U25 ( .A0_t (roundconstant[1]), .A0_f (new_AGEMA_signal_1878), .B0_t (IN_reset_t), .B0_f (IN_reset_f), .Z0_t (roundconstant[2]), .Z0_f (new_AGEMA_signal_1887) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) LED_128_Instance_U24 ( .A0_t (roundconstant[0]), .A0_f (new_AGEMA_signal_1888), .B0_t (IN_reset_t), .B0_f (IN_reset_f), .Z0_t (roundconstant[1]), .Z0_f (new_AGEMA_signal_1878) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) LED_128_Instance_U23 ( .A0_t (IN_reset_t), .A0_f (IN_reset_f), .B0_t (LED_128_Instance_ks_reg_2__Q), .B0_f (new_AGEMA_signal_1884), .Z0_t (LED_128_Instance_ks_3_), .Z0_f (new_AGEMA_signal_1886) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b1), .NL(1'b1)) LED_128_Instance_U22 ( .A0_t (LED_128_Instance_n29), .A0_f (new_AGEMA_signal_1889), .B0_t (IN_reset_t), .B0_f (IN_reset_f), .Z0_t (roundconstant[0]), .Z0_f (new_AGEMA_signal_1888) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) LED_128_Instance_U20 ( .A0_t (roundconstant[5]), .A0_f (new_AGEMA_signal_1877), .B0_t (roundconstant[4]), .B0_f (new_AGEMA_signal_1882), .Z0_t (LED_128_Instance_n29), .Z0_f (new_AGEMA_signal_1889) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) LED_128_Instance_U17 ( .A0_t (roundconstant[0]), .A0_f (new_AGEMA_signal_1888), .B0_t (LED_128_Instance_n19), .B0_f (new_AGEMA_signal_2475), .Z0_t (LED_128_Instance_n22), .Z0_f (new_AGEMA_signal_2479) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) LED_128_Instance_U16 ( .A0_t (roundconstant[5]), .A0_f (new_AGEMA_signal_1877), .B0_t (LED_128_Instance_n18), .B0_f (new_AGEMA_signal_2471), .Z0_t (LED_128_Instance_n19), .Z0_f (new_AGEMA_signal_2475) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) LED_128_Instance_U15 ( .A0_t (LED_128_Instance_n17), .A0_f (new_AGEMA_signal_1891), .B0_t (LED_128_Instance_n16), .B0_f (new_AGEMA_signal_1890), .Z0_t (LED_128_Instance_n18), .Z0_f (new_AGEMA_signal_2471) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) LED_128_Instance_U14 ( .A0_t (roundconstant[2]), .A0_f (new_AGEMA_signal_1887), .B0_t (roundconstant[1]), .B0_f (new_AGEMA_signal_1878), .Z0_t (LED_128_Instance_n16), .Z0_f (new_AGEMA_signal_1890) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) LED_128_Instance_U13 ( .A0_t (roundconstant[4]), .A0_f (new_AGEMA_signal_1882), .B0_t (roundconstant[3]), .B0_f (new_AGEMA_signal_1880), .Z0_t (LED_128_Instance_n17), .Z0_f (new_AGEMA_signal_1891) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) LED_128_Instance_U11 ( .A0_t (LED_128_Instance_n31), .A0_f (new_AGEMA_signal_2477), .B0_t (LED_128_Instance_n13), .B0_f (new_AGEMA_signal_2476), .Z0_t (LED_128_Instance_n23), .Z0_f (new_AGEMA_signal_2480) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) LED_128_Instance_U10 ( .A0_t (LED_128_Instance_ks_0), .A0_f (new_AGEMA_signal_1885), .B0_t (LED_128_Instance_n12), .B0_f (new_AGEMA_signal_2472), .Z0_t (LED_128_Instance_n13), .Z0_f (new_AGEMA_signal_2476) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) LED_128_Instance_U9 ( .A0_t (LED_128_Instance_ks_3_), .A0_f (new_AGEMA_signal_1886), .B0_t (LED_128_Instance_n11), .B0_f (new_AGEMA_signal_1892), .Z0_t (LED_128_Instance_n12), .Z0_f (new_AGEMA_signal_2472) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) LED_128_Instance_U8 ( .A0_t (LED_128_Instance_n24), .A0_f (new_AGEMA_signal_1883), .B0_t (LED_128_Instance_ks_reg_2__Q), .B0_f (new_AGEMA_signal_1884), .Z0_t (LED_128_Instance_n11), .Z0_f (new_AGEMA_signal_1892) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) LED_128_Instance_U6 ( .A0_t (LED_128_Instance_ks_0), .A0_f (new_AGEMA_signal_1885), .B0_t (LED_128_Instance_n9), .B0_f (new_AGEMA_signal_2473), .Z0_t (LED_128_Instance_n31), .Z0_f (new_AGEMA_signal_2477) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) LED_128_Instance_U5 ( .A0_t (LED_128_Instance_ks_3_), .A0_f (new_AGEMA_signal_1886), .B0_t (LED_128_Instance_n8), .B0_f (new_AGEMA_signal_1893), .Z0_t (LED_128_Instance_n9), .Z0_f (new_AGEMA_signal_2473) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) LED_128_Instance_U4 ( .A0_t (LED_128_Instance_n24), .A0_f (new_AGEMA_signal_1883), .B0_t (LED_128_Instance_ks_reg_2__Q), .B0_f (new_AGEMA_signal_1884), .Z0_t (LED_128_Instance_n8), .Z0_f (new_AGEMA_signal_1893) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_0_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[0]), .A0_f (new_AGEMA_signal_5019), .A1_t (new_AGEMA_signal_5020), .A1_f (new_AGEMA_signal_5021), .B0_t (LED_128_Instance_addconst_out[0]), .B0_f (new_AGEMA_signal_3636), .B1_t (new_AGEMA_signal_3637), .B1_f (new_AGEMA_signal_3638), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_0_U1_X), .Z0_f (new_AGEMA_signal_5127), .Z1_t (new_AGEMA_signal_5128), .Z1_f (new_AGEMA_signal_5129) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_0_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n22), .A1_f (new_AGEMA_signal_2479), .B0_t (LED_128_Instance_MUX_state0_mux_inst_0_U1_X), .B0_f (new_AGEMA_signal_5127), .B1_t (new_AGEMA_signal_5128), .B1_f (new_AGEMA_signal_5129), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_0_U1_Y), .Z0_f (new_AGEMA_signal_5280), .Z1_t (new_AGEMA_signal_5281), .Z1_f (new_AGEMA_signal_5282) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_0_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_0_U1_Y), .A0_f (new_AGEMA_signal_5280), .A1_t (new_AGEMA_signal_5281), .A1_f (new_AGEMA_signal_5282), .B0_t (LED_128_Instance_mixcolumns_out[0]), .B0_f (new_AGEMA_signal_5019), .B1_t (new_AGEMA_signal_5020), .B1_f (new_AGEMA_signal_5021), .Z0_t (LED_128_Instance_state0[0]), .Z0_f (new_AGEMA_signal_5454), .Z1_t (new_AGEMA_signal_5455), .Z1_f (new_AGEMA_signal_5456) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_1_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[1]), .A0_f (new_AGEMA_signal_5319), .A1_t (new_AGEMA_signal_5320), .A1_f (new_AGEMA_signal_5321), .B0_t (LED_128_Instance_addconst_out[1]), .B0_f (new_AGEMA_signal_3639), .B1_t (new_AGEMA_signal_3640), .B1_f (new_AGEMA_signal_3641), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_1_U1_X), .Z0_f (new_AGEMA_signal_5457), .Z1_t (new_AGEMA_signal_5458), .Z1_f (new_AGEMA_signal_5459) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_1_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n22), .A1_f (new_AGEMA_signal_2479), .B0_t (LED_128_Instance_MUX_state0_mux_inst_1_U1_X), .B0_f (new_AGEMA_signal_5457), .B1_t (new_AGEMA_signal_5458), .B1_f (new_AGEMA_signal_5459), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_1_U1_Y), .Z0_f (new_AGEMA_signal_5643), .Z1_t (new_AGEMA_signal_5644), .Z1_f (new_AGEMA_signal_5645) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_1_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_1_U1_Y), .A0_f (new_AGEMA_signal_5643), .A1_t (new_AGEMA_signal_5644), .A1_f (new_AGEMA_signal_5645), .B0_t (LED_128_Instance_mixcolumns_out[1]), .B0_f (new_AGEMA_signal_5319), .B1_t (new_AGEMA_signal_5320), .B1_f (new_AGEMA_signal_5321), .Z0_t (LED_128_Instance_state0[1]), .Z0_f (new_AGEMA_signal_5847), .Z1_t (new_AGEMA_signal_5848), .Z1_f (new_AGEMA_signal_5849) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_2_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[2]), .A0_f (new_AGEMA_signal_5010), .A1_t (new_AGEMA_signal_5011), .A1_f (new_AGEMA_signal_5012), .B0_t (LED_128_Instance_addconst_out[2]), .B0_f (new_AGEMA_signal_3642), .B1_t (new_AGEMA_signal_3643), .B1_f (new_AGEMA_signal_3644), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_2_U1_X), .Z0_f (new_AGEMA_signal_5130), .Z1_t (new_AGEMA_signal_5131), .Z1_f (new_AGEMA_signal_5132) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_2_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n22), .A1_f (new_AGEMA_signal_2479), .B0_t (LED_128_Instance_MUX_state0_mux_inst_2_U1_X), .B0_f (new_AGEMA_signal_5130), .B1_t (new_AGEMA_signal_5131), .B1_f (new_AGEMA_signal_5132), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_2_U1_Y), .Z0_f (new_AGEMA_signal_5283), .Z1_t (new_AGEMA_signal_5284), .Z1_f (new_AGEMA_signal_5285) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_2_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_2_U1_Y), .A0_f (new_AGEMA_signal_5283), .A1_t (new_AGEMA_signal_5284), .A1_f (new_AGEMA_signal_5285), .B0_t (LED_128_Instance_mixcolumns_out[2]), .B0_f (new_AGEMA_signal_5010), .B1_t (new_AGEMA_signal_5011), .B1_f (new_AGEMA_signal_5012), .Z0_t (LED_128_Instance_state0[2]), .Z0_f (new_AGEMA_signal_5460), .Z1_t (new_AGEMA_signal_5461), .Z1_f (new_AGEMA_signal_5462) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_3_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[3]), .A0_f (new_AGEMA_signal_5349), .A1_t (new_AGEMA_signal_5350), .A1_f (new_AGEMA_signal_5351), .B0_t (LED_128_Instance_addroundkey_out[3]), .B0_f (new_AGEMA_signal_3645), .B1_t (new_AGEMA_signal_3646), .B1_f (new_AGEMA_signal_3647), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_3_U1_X), .Z0_f (new_AGEMA_signal_5463), .Z1_t (new_AGEMA_signal_5464), .Z1_f (new_AGEMA_signal_5465) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_3_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n22), .A1_f (new_AGEMA_signal_2479), .B0_t (LED_128_Instance_MUX_state0_mux_inst_3_U1_X), .B0_f (new_AGEMA_signal_5463), .B1_t (new_AGEMA_signal_5464), .B1_f (new_AGEMA_signal_5465), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_3_U1_Y), .Z0_f (new_AGEMA_signal_5646), .Z1_t (new_AGEMA_signal_5647), .Z1_f (new_AGEMA_signal_5648) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_3_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_3_U1_Y), .A0_f (new_AGEMA_signal_5646), .A1_t (new_AGEMA_signal_5647), .A1_f (new_AGEMA_signal_5648), .B0_t (LED_128_Instance_mixcolumns_out[3]), .B0_f (new_AGEMA_signal_5349), .B1_t (new_AGEMA_signal_5350), .B1_f (new_AGEMA_signal_5351), .Z0_t (LED_128_Instance_state0[3]), .Z0_f (new_AGEMA_signal_5850), .Z1_t (new_AGEMA_signal_5851), .Z1_f (new_AGEMA_signal_5852) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_4_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[4]), .A0_f (new_AGEMA_signal_5208), .A1_t (new_AGEMA_signal_5209), .A1_f (new_AGEMA_signal_5210), .B0_t (LED_128_Instance_addroundkey_out[4]), .B0_f (new_AGEMA_signal_3648), .B1_t (new_AGEMA_signal_3649), .B1_f (new_AGEMA_signal_3650), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_4_U1_X), .Z0_f (new_AGEMA_signal_5286), .Z1_t (new_AGEMA_signal_5287), .Z1_f (new_AGEMA_signal_5288) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_4_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n22), .A1_f (new_AGEMA_signal_2479), .B0_t (LED_128_Instance_MUX_state0_mux_inst_4_U1_X), .B0_f (new_AGEMA_signal_5286), .B1_t (new_AGEMA_signal_5287), .B1_f (new_AGEMA_signal_5288), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_4_U1_Y), .Z0_f (new_AGEMA_signal_5466), .Z1_t (new_AGEMA_signal_5467), .Z1_f (new_AGEMA_signal_5468) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_4_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_4_U1_Y), .A0_f (new_AGEMA_signal_5466), .A1_t (new_AGEMA_signal_5467), .A1_f (new_AGEMA_signal_5468), .B0_t (LED_128_Instance_mixcolumns_out[4]), .B0_f (new_AGEMA_signal_5208), .B1_t (new_AGEMA_signal_5209), .B1_f (new_AGEMA_signal_5210), .Z0_t (LED_128_Instance_state0[4]), .Z0_f (new_AGEMA_signal_5649), .Z1_t (new_AGEMA_signal_5650), .Z1_f (new_AGEMA_signal_5651) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_5_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[5]), .A0_f (new_AGEMA_signal_5358), .A1_t (new_AGEMA_signal_5359), .A1_f (new_AGEMA_signal_5360), .B0_t (LED_128_Instance_addroundkey_out[5]), .B0_f (new_AGEMA_signal_3651), .B1_t (new_AGEMA_signal_3652), .B1_f (new_AGEMA_signal_3653), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_5_U1_X), .Z0_f (new_AGEMA_signal_5469), .Z1_t (new_AGEMA_signal_5470), .Z1_f (new_AGEMA_signal_5471) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_5_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n22), .A1_f (new_AGEMA_signal_2479), .B0_t (LED_128_Instance_MUX_state0_mux_inst_5_U1_X), .B0_f (new_AGEMA_signal_5469), .B1_t (new_AGEMA_signal_5470), .B1_f (new_AGEMA_signal_5471), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_5_U1_Y), .Z0_f (new_AGEMA_signal_5652), .Z1_t (new_AGEMA_signal_5653), .Z1_f (new_AGEMA_signal_5654) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_5_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_5_U1_Y), .A0_f (new_AGEMA_signal_5652), .A1_t (new_AGEMA_signal_5653), .A1_f (new_AGEMA_signal_5654), .B0_t (LED_128_Instance_mixcolumns_out[5]), .B0_f (new_AGEMA_signal_5358), .B1_t (new_AGEMA_signal_5359), .B1_f (new_AGEMA_signal_5360), .Z0_t (LED_128_Instance_state0[5]), .Z0_f (new_AGEMA_signal_5853), .Z1_t (new_AGEMA_signal_5854), .Z1_f (new_AGEMA_signal_5855) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_6_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[6]), .A0_f (new_AGEMA_signal_5196), .A1_t (new_AGEMA_signal_5197), .A1_f (new_AGEMA_signal_5198), .B0_t (LED_128_Instance_addroundkey_out[6]), .B0_f (new_AGEMA_signal_3654), .B1_t (new_AGEMA_signal_3655), .B1_f (new_AGEMA_signal_3656), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_6_U1_X), .Z0_f (new_AGEMA_signal_5289), .Z1_t (new_AGEMA_signal_5290), .Z1_f (new_AGEMA_signal_5291) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_6_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n22), .A1_f (new_AGEMA_signal_2479), .B0_t (LED_128_Instance_MUX_state0_mux_inst_6_U1_X), .B0_f (new_AGEMA_signal_5289), .B1_t (new_AGEMA_signal_5290), .B1_f (new_AGEMA_signal_5291), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_6_U1_Y), .Z0_f (new_AGEMA_signal_5472), .Z1_t (new_AGEMA_signal_5473), .Z1_f (new_AGEMA_signal_5474) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_6_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_6_U1_Y), .A0_f (new_AGEMA_signal_5472), .A1_t (new_AGEMA_signal_5473), .A1_f (new_AGEMA_signal_5474), .B0_t (LED_128_Instance_mixcolumns_out[6]), .B0_f (new_AGEMA_signal_5196), .B1_t (new_AGEMA_signal_5197), .B1_f (new_AGEMA_signal_5198), .Z0_t (LED_128_Instance_state0[6]), .Z0_f (new_AGEMA_signal_5655), .Z1_t (new_AGEMA_signal_5656), .Z1_f (new_AGEMA_signal_5657) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_7_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[7]), .A0_f (new_AGEMA_signal_5202), .A1_t (new_AGEMA_signal_5203), .A1_f (new_AGEMA_signal_5204), .B0_t (LED_128_Instance_addconst_out[7]), .B0_f (new_AGEMA_signal_3657), .B1_t (new_AGEMA_signal_3658), .B1_f (new_AGEMA_signal_3659), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_7_U1_X), .Z0_f (new_AGEMA_signal_5292), .Z1_t (new_AGEMA_signal_5293), .Z1_f (new_AGEMA_signal_5294) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_7_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n22), .A1_f (new_AGEMA_signal_2479), .B0_t (LED_128_Instance_MUX_state0_mux_inst_7_U1_X), .B0_f (new_AGEMA_signal_5292), .B1_t (new_AGEMA_signal_5293), .B1_f (new_AGEMA_signal_5294), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_7_U1_Y), .Z0_f (new_AGEMA_signal_5475), .Z1_t (new_AGEMA_signal_5476), .Z1_f (new_AGEMA_signal_5477) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_7_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_7_U1_Y), .A0_f (new_AGEMA_signal_5475), .A1_t (new_AGEMA_signal_5476), .A1_f (new_AGEMA_signal_5477), .B0_t (LED_128_Instance_mixcolumns_out[7]), .B0_f (new_AGEMA_signal_5202), .B1_t (new_AGEMA_signal_5203), .B1_f (new_AGEMA_signal_5204), .Z0_t (LED_128_Instance_state0[7]), .Z0_f (new_AGEMA_signal_5658), .Z1_t (new_AGEMA_signal_5659), .Z1_f (new_AGEMA_signal_5660) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_8_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[8]), .A0_f (new_AGEMA_signal_5088), .A1_t (new_AGEMA_signal_5089), .A1_f (new_AGEMA_signal_5090), .B0_t (LED_128_Instance_addconst_out[8]), .B0_f (new_AGEMA_signal_3660), .B1_t (new_AGEMA_signal_3661), .B1_f (new_AGEMA_signal_3662), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_8_U1_X), .Z0_f (new_AGEMA_signal_5133), .Z1_t (new_AGEMA_signal_5134), .Z1_f (new_AGEMA_signal_5135) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_8_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n22), .A1_f (new_AGEMA_signal_2479), .B0_t (LED_128_Instance_MUX_state0_mux_inst_8_U1_X), .B0_f (new_AGEMA_signal_5133), .B1_t (new_AGEMA_signal_5134), .B1_f (new_AGEMA_signal_5135), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_8_U1_Y), .Z0_f (new_AGEMA_signal_5295), .Z1_t (new_AGEMA_signal_5296), .Z1_f (new_AGEMA_signal_5297) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_8_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_8_U1_Y), .A0_f (new_AGEMA_signal_5295), .A1_t (new_AGEMA_signal_5296), .A1_f (new_AGEMA_signal_5297), .B0_t (LED_128_Instance_mixcolumns_out[8]), .B0_f (new_AGEMA_signal_5088), .B1_t (new_AGEMA_signal_5089), .B1_f (new_AGEMA_signal_5090), .Z0_t (LED_128_Instance_state0[8]), .Z0_f (new_AGEMA_signal_5478), .Z1_t (new_AGEMA_signal_5479), .Z1_f (new_AGEMA_signal_5480) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_9_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[9]), .A0_f (new_AGEMA_signal_5388), .A1_t (new_AGEMA_signal_5389), .A1_f (new_AGEMA_signal_5390), .B0_t (LED_128_Instance_addconst_out[9]), .B0_f (new_AGEMA_signal_3663), .B1_t (new_AGEMA_signal_3664), .B1_f (new_AGEMA_signal_3665), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_9_U1_X), .Z0_f (new_AGEMA_signal_5481), .Z1_t (new_AGEMA_signal_5482), .Z1_f (new_AGEMA_signal_5483) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_9_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n22), .A1_f (new_AGEMA_signal_2479), .B0_t (LED_128_Instance_MUX_state0_mux_inst_9_U1_X), .B0_f (new_AGEMA_signal_5481), .B1_t (new_AGEMA_signal_5482), .B1_f (new_AGEMA_signal_5483), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_9_U1_Y), .Z0_f (new_AGEMA_signal_5661), .Z1_t (new_AGEMA_signal_5662), .Z1_f (new_AGEMA_signal_5663) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_9_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_9_U1_Y), .A0_f (new_AGEMA_signal_5661), .A1_t (new_AGEMA_signal_5662), .A1_f (new_AGEMA_signal_5663), .B0_t (LED_128_Instance_mixcolumns_out[9]), .B0_f (new_AGEMA_signal_5388), .B1_t (new_AGEMA_signal_5389), .B1_f (new_AGEMA_signal_5390), .Z0_t (LED_128_Instance_state0[9]), .Z0_f (new_AGEMA_signal_5856), .Z1_t (new_AGEMA_signal_5857), .Z1_f (new_AGEMA_signal_5858) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_10_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[10]), .A0_f (new_AGEMA_signal_5235), .A1_t (new_AGEMA_signal_5236), .A1_f (new_AGEMA_signal_5237), .B0_t (LED_128_Instance_addconst_out[10]), .B0_f (new_AGEMA_signal_3666), .B1_t (new_AGEMA_signal_3667), .B1_f (new_AGEMA_signal_3668), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_10_U1_X), .Z0_f (new_AGEMA_signal_5298), .Z1_t (new_AGEMA_signal_5299), .Z1_f (new_AGEMA_signal_5300) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_10_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n22), .A1_f (new_AGEMA_signal_2479), .B0_t (LED_128_Instance_MUX_state0_mux_inst_10_U1_X), .B0_f (new_AGEMA_signal_5298), .B1_t (new_AGEMA_signal_5299), .B1_f (new_AGEMA_signal_5300), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_10_U1_Y), .Z0_f (new_AGEMA_signal_5484), .Z1_t (new_AGEMA_signal_5485), .Z1_f (new_AGEMA_signal_5486) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_10_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_10_U1_Y), .A0_f (new_AGEMA_signal_5484), .A1_t (new_AGEMA_signal_5485), .A1_f (new_AGEMA_signal_5486), .B0_t (LED_128_Instance_mixcolumns_out[10]), .B0_f (new_AGEMA_signal_5235), .B1_t (new_AGEMA_signal_5236), .B1_f (new_AGEMA_signal_5237), .Z0_t (LED_128_Instance_state0[10]), .Z0_f (new_AGEMA_signal_5664), .Z1_t (new_AGEMA_signal_5665), .Z1_f (new_AGEMA_signal_5666) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_11_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[11]), .A0_f (new_AGEMA_signal_5241), .A1_t (new_AGEMA_signal_5242), .A1_f (new_AGEMA_signal_5243), .B0_t (LED_128_Instance_addconst_out[11]), .B0_f (new_AGEMA_signal_3669), .B1_t (new_AGEMA_signal_3670), .B1_f (new_AGEMA_signal_3671), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_11_U1_X), .Z0_f (new_AGEMA_signal_5301), .Z1_t (new_AGEMA_signal_5302), .Z1_f (new_AGEMA_signal_5303) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_11_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n22), .A1_f (new_AGEMA_signal_2479), .B0_t (LED_128_Instance_MUX_state0_mux_inst_11_U1_X), .B0_f (new_AGEMA_signal_5301), .B1_t (new_AGEMA_signal_5302), .B1_f (new_AGEMA_signal_5303), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_11_U1_Y), .Z0_f (new_AGEMA_signal_5487), .Z1_t (new_AGEMA_signal_5488), .Z1_f (new_AGEMA_signal_5489) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_11_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_11_U1_Y), .A0_f (new_AGEMA_signal_5487), .A1_t (new_AGEMA_signal_5488), .A1_f (new_AGEMA_signal_5489), .B0_t (LED_128_Instance_mixcolumns_out[11]), .B0_f (new_AGEMA_signal_5241), .B1_t (new_AGEMA_signal_5242), .B1_f (new_AGEMA_signal_5243), .Z0_t (LED_128_Instance_state0[11]), .Z0_f (new_AGEMA_signal_5667), .Z1_t (new_AGEMA_signal_5668), .Z1_f (new_AGEMA_signal_5669) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_12_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[12]), .A0_f (new_AGEMA_signal_5274), .A1_t (new_AGEMA_signal_5275), .A1_f (new_AGEMA_signal_5276), .B0_t (LED_128_Instance_addconst_out[12]), .B0_f (new_AGEMA_signal_3672), .B1_t (new_AGEMA_signal_3673), .B1_f (new_AGEMA_signal_3674), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_12_U1_X), .Z0_f (new_AGEMA_signal_5304), .Z1_t (new_AGEMA_signal_5305), .Z1_f (new_AGEMA_signal_5306) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_12_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n22), .A1_f (new_AGEMA_signal_2479), .B0_t (LED_128_Instance_MUX_state0_mux_inst_12_U1_X), .B0_f (new_AGEMA_signal_5304), .B1_t (new_AGEMA_signal_5305), .B1_f (new_AGEMA_signal_5306), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_12_U1_Y), .Z0_f (new_AGEMA_signal_5490), .Z1_t (new_AGEMA_signal_5491), .Z1_f (new_AGEMA_signal_5492) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_12_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_12_U1_Y), .A0_f (new_AGEMA_signal_5490), .A1_t (new_AGEMA_signal_5491), .A1_f (new_AGEMA_signal_5492), .B0_t (LED_128_Instance_mixcolumns_out[12]), .B0_f (new_AGEMA_signal_5274), .B1_t (new_AGEMA_signal_5275), .B1_f (new_AGEMA_signal_5276), .Z0_t (LED_128_Instance_state0[12]), .Z0_f (new_AGEMA_signal_5670), .Z1_t (new_AGEMA_signal_5671), .Z1_f (new_AGEMA_signal_5672) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_13_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[13]), .A0_f (new_AGEMA_signal_5619), .A1_t (new_AGEMA_signal_5620), .A1_f (new_AGEMA_signal_5621), .B0_t (LED_128_Instance_addconst_out[13]), .B0_f (new_AGEMA_signal_3675), .B1_t (new_AGEMA_signal_3676), .B1_f (new_AGEMA_signal_3677), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_13_U1_X), .Z0_f (new_AGEMA_signal_5673), .Z1_t (new_AGEMA_signal_5674), .Z1_f (new_AGEMA_signal_5675) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_13_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n22), .A1_f (new_AGEMA_signal_2479), .B0_t (LED_128_Instance_MUX_state0_mux_inst_13_U1_X), .B0_f (new_AGEMA_signal_5673), .B1_t (new_AGEMA_signal_5674), .B1_f (new_AGEMA_signal_5675), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_13_U1_Y), .Z0_f (new_AGEMA_signal_5859), .Z1_t (new_AGEMA_signal_5860), .Z1_f (new_AGEMA_signal_5861) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_13_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_13_U1_Y), .A0_f (new_AGEMA_signal_5859), .A1_t (new_AGEMA_signal_5860), .A1_f (new_AGEMA_signal_5861), .B0_t (LED_128_Instance_mixcolumns_out[13]), .B0_f (new_AGEMA_signal_5619), .B1_t (new_AGEMA_signal_5620), .B1_f (new_AGEMA_signal_5621), .Z0_t (LED_128_Instance_state0[13]), .Z0_f (new_AGEMA_signal_6066), .Z1_t (new_AGEMA_signal_6067), .Z1_f (new_AGEMA_signal_6068) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_14_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[14]), .A0_f (new_AGEMA_signal_5112), .A1_t (new_AGEMA_signal_5113), .A1_f (new_AGEMA_signal_5114), .B0_t (LED_128_Instance_addconst_out[14]), .B0_f (new_AGEMA_signal_3678), .B1_t (new_AGEMA_signal_3679), .B1_f (new_AGEMA_signal_3680), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_14_U1_X), .Z0_f (new_AGEMA_signal_5136), .Z1_t (new_AGEMA_signal_5137), .Z1_f (new_AGEMA_signal_5138) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_14_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n22), .A1_f (new_AGEMA_signal_2479), .B0_t (LED_128_Instance_MUX_state0_mux_inst_14_U1_X), .B0_f (new_AGEMA_signal_5136), .B1_t (new_AGEMA_signal_5137), .B1_f (new_AGEMA_signal_5138), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_14_U1_Y), .Z0_f (new_AGEMA_signal_5307), .Z1_t (new_AGEMA_signal_5308), .Z1_f (new_AGEMA_signal_5309) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_14_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_14_U1_Y), .A0_f (new_AGEMA_signal_5307), .A1_t (new_AGEMA_signal_5308), .A1_f (new_AGEMA_signal_5309), .B0_t (LED_128_Instance_mixcolumns_out[14]), .B0_f (new_AGEMA_signal_5112), .B1_t (new_AGEMA_signal_5113), .B1_f (new_AGEMA_signal_5114), .Z0_t (LED_128_Instance_state0[14]), .Z0_f (new_AGEMA_signal_5493), .Z1_t (new_AGEMA_signal_5494), .Z1_f (new_AGEMA_signal_5495) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_15_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[15]), .A0_f (new_AGEMA_signal_5268), .A1_t (new_AGEMA_signal_5269), .A1_f (new_AGEMA_signal_5270), .B0_t (LED_128_Instance_addconst_out[15]), .B0_f (new_AGEMA_signal_3681), .B1_t (new_AGEMA_signal_3682), .B1_f (new_AGEMA_signal_3683), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_15_U1_X), .Z0_f (new_AGEMA_signal_5310), .Z1_t (new_AGEMA_signal_5311), .Z1_f (new_AGEMA_signal_5312) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_15_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n22), .A1_f (new_AGEMA_signal_2479), .B0_t (LED_128_Instance_MUX_state0_mux_inst_15_U1_X), .B0_f (new_AGEMA_signal_5310), .B1_t (new_AGEMA_signal_5311), .B1_f (new_AGEMA_signal_5312), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_15_U1_Y), .Z0_f (new_AGEMA_signal_5496), .Z1_t (new_AGEMA_signal_5497), .Z1_f (new_AGEMA_signal_5498) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_15_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_15_U1_Y), .A0_f (new_AGEMA_signal_5496), .A1_t (new_AGEMA_signal_5497), .A1_f (new_AGEMA_signal_5498), .B0_t (LED_128_Instance_mixcolumns_out[15]), .B0_f (new_AGEMA_signal_5268), .B1_t (new_AGEMA_signal_5269), .B1_f (new_AGEMA_signal_5270), .Z0_t (LED_128_Instance_state0[15]), .Z0_f (new_AGEMA_signal_5676), .Z1_t (new_AGEMA_signal_5677), .Z1_f (new_AGEMA_signal_5678) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_16_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[16]), .A0_f (new_AGEMA_signal_5574), .A1_t (new_AGEMA_signal_5575), .A1_f (new_AGEMA_signal_5576), .B0_t (LED_128_Instance_addroundkey_out[16]), .B0_f (new_AGEMA_signal_3684), .B1_t (new_AGEMA_signal_3685), .B1_f (new_AGEMA_signal_3686), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_16_U1_X), .Z0_f (new_AGEMA_signal_5679), .Z1_t (new_AGEMA_signal_5680), .Z1_f (new_AGEMA_signal_5681) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_16_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n22), .A1_f (new_AGEMA_signal_2479), .B0_t (LED_128_Instance_MUX_state0_mux_inst_16_U1_X), .B0_f (new_AGEMA_signal_5679), .B1_t (new_AGEMA_signal_5680), .B1_f (new_AGEMA_signal_5681), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_16_U1_Y), .Z0_f (new_AGEMA_signal_5862), .Z1_t (new_AGEMA_signal_5863), .Z1_f (new_AGEMA_signal_5864) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_16_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_16_U1_Y), .A0_f (new_AGEMA_signal_5862), .A1_t (new_AGEMA_signal_5863), .A1_f (new_AGEMA_signal_5864), .B0_t (LED_128_Instance_mixcolumns_out[16]), .B0_f (new_AGEMA_signal_5574), .B1_t (new_AGEMA_signal_5575), .B1_f (new_AGEMA_signal_5576), .Z0_t (LED_128_Instance_state0[16]), .Z0_f (new_AGEMA_signal_6069), .Z1_t (new_AGEMA_signal_6070), .Z1_f (new_AGEMA_signal_6071) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_17_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[17]), .A0_f (new_AGEMA_signal_5346), .A1_t (new_AGEMA_signal_5347), .A1_f (new_AGEMA_signal_5348), .B0_t (LED_128_Instance_addconst_out[17]), .B0_f (new_AGEMA_signal_3687), .B1_t (new_AGEMA_signal_3688), .B1_f (new_AGEMA_signal_3689), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_17_U1_X), .Z0_f (new_AGEMA_signal_5499), .Z1_t (new_AGEMA_signal_5500), .Z1_f (new_AGEMA_signal_5501) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_17_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n22), .A1_f (new_AGEMA_signal_2479), .B0_t (LED_128_Instance_MUX_state0_mux_inst_17_U1_X), .B0_f (new_AGEMA_signal_5499), .B1_t (new_AGEMA_signal_5500), .B1_f (new_AGEMA_signal_5501), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_17_U1_Y), .Z0_f (new_AGEMA_signal_5682), .Z1_t (new_AGEMA_signal_5683), .Z1_f (new_AGEMA_signal_5684) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_17_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_17_U1_Y), .A0_f (new_AGEMA_signal_5682), .A1_t (new_AGEMA_signal_5683), .A1_f (new_AGEMA_signal_5684), .B0_t (LED_128_Instance_mixcolumns_out[17]), .B0_f (new_AGEMA_signal_5346), .B1_t (new_AGEMA_signal_5347), .B1_f (new_AGEMA_signal_5348), .Z0_t (LED_128_Instance_state0[17]), .Z0_f (new_AGEMA_signal_5865), .Z1_t (new_AGEMA_signal_5866), .Z1_f (new_AGEMA_signal_5867) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_18_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[18]), .A0_f (new_AGEMA_signal_5559), .A1_t (new_AGEMA_signal_5560), .A1_f (new_AGEMA_signal_5561), .B0_t (LED_128_Instance_addconst_out[18]), .B0_f (new_AGEMA_signal_3690), .B1_t (new_AGEMA_signal_3691), .B1_f (new_AGEMA_signal_3692), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_18_U1_X), .Z0_f (new_AGEMA_signal_5685), .Z1_t (new_AGEMA_signal_5686), .Z1_f (new_AGEMA_signal_5687) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_18_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n22), .A1_f (new_AGEMA_signal_2479), .B0_t (LED_128_Instance_MUX_state0_mux_inst_18_U1_X), .B0_f (new_AGEMA_signal_5685), .B1_t (new_AGEMA_signal_5686), .B1_f (new_AGEMA_signal_5687), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_18_U1_Y), .Z0_f (new_AGEMA_signal_5868), .Z1_t (new_AGEMA_signal_5869), .Z1_f (new_AGEMA_signal_5870) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_18_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_18_U1_Y), .A0_f (new_AGEMA_signal_5868), .A1_t (new_AGEMA_signal_5869), .A1_f (new_AGEMA_signal_5870), .B0_t (LED_128_Instance_mixcolumns_out[18]), .B0_f (new_AGEMA_signal_5559), .B1_t (new_AGEMA_signal_5560), .B1_f (new_AGEMA_signal_5561), .Z0_t (LED_128_Instance_state0[18]), .Z0_f (new_AGEMA_signal_6072), .Z1_t (new_AGEMA_signal_6073), .Z1_f (new_AGEMA_signal_6074) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_19_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[19]), .A0_f (new_AGEMA_signal_5556), .A1_t (new_AGEMA_signal_5557), .A1_f (new_AGEMA_signal_5558), .B0_t (LED_128_Instance_addroundkey_out[19]), .B0_f (new_AGEMA_signal_3693), .B1_t (new_AGEMA_signal_3694), .B1_f (new_AGEMA_signal_3695), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_19_U1_X), .Z0_f (new_AGEMA_signal_5688), .Z1_t (new_AGEMA_signal_5689), .Z1_f (new_AGEMA_signal_5690) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_19_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n22), .A1_f (new_AGEMA_signal_2479), .B0_t (LED_128_Instance_MUX_state0_mux_inst_19_U1_X), .B0_f (new_AGEMA_signal_5688), .B1_t (new_AGEMA_signal_5689), .B1_f (new_AGEMA_signal_5690), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_19_U1_Y), .Z0_f (new_AGEMA_signal_5871), .Z1_t (new_AGEMA_signal_5872), .Z1_f (new_AGEMA_signal_5873) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_19_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_19_U1_Y), .A0_f (new_AGEMA_signal_5871), .A1_t (new_AGEMA_signal_5872), .A1_f (new_AGEMA_signal_5873), .B0_t (LED_128_Instance_mixcolumns_out[19]), .B0_f (new_AGEMA_signal_5556), .B1_t (new_AGEMA_signal_5557), .B1_f (new_AGEMA_signal_5558), .Z0_t (LED_128_Instance_state0[19]), .Z0_f (new_AGEMA_signal_6075), .Z1_t (new_AGEMA_signal_6076), .Z1_f (new_AGEMA_signal_6077) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_20_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[20]), .A0_f (new_AGEMA_signal_5382), .A1_t (new_AGEMA_signal_5383), .A1_f (new_AGEMA_signal_5384), .B0_t (LED_128_Instance_addroundkey_out[20]), .B0_f (new_AGEMA_signal_3696), .B1_t (new_AGEMA_signal_3697), .B1_f (new_AGEMA_signal_3698), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_20_U1_X), .Z0_f (new_AGEMA_signal_5502), .Z1_t (new_AGEMA_signal_5503), .Z1_f (new_AGEMA_signal_5504) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_20_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n22), .A1_f (new_AGEMA_signal_2479), .B0_t (LED_128_Instance_MUX_state0_mux_inst_20_U1_X), .B0_f (new_AGEMA_signal_5502), .B1_t (new_AGEMA_signal_5503), .B1_f (new_AGEMA_signal_5504), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_20_U1_Y), .Z0_f (new_AGEMA_signal_5691), .Z1_t (new_AGEMA_signal_5692), .Z1_f (new_AGEMA_signal_5693) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_20_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_20_U1_Y), .A0_f (new_AGEMA_signal_5691), .A1_t (new_AGEMA_signal_5692), .A1_f (new_AGEMA_signal_5693), .B0_t (LED_128_Instance_mixcolumns_out[20]), .B0_f (new_AGEMA_signal_5382), .B1_t (new_AGEMA_signal_5383), .B1_f (new_AGEMA_signal_5384), .Z0_t (LED_128_Instance_state0[20]), .Z0_f (new_AGEMA_signal_5874), .Z1_t (new_AGEMA_signal_5875), .Z1_f (new_AGEMA_signal_5876) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_21_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[21]), .A0_f (new_AGEMA_signal_5199), .A1_t (new_AGEMA_signal_5200), .A1_f (new_AGEMA_signal_5201), .B0_t (LED_128_Instance_addroundkey_out[21]), .B0_f (new_AGEMA_signal_3699), .B1_t (new_AGEMA_signal_3700), .B1_f (new_AGEMA_signal_3701), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_21_U1_X), .Z0_f (new_AGEMA_signal_5313), .Z1_t (new_AGEMA_signal_5314), .Z1_f (new_AGEMA_signal_5315) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_21_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n22), .A1_f (new_AGEMA_signal_2479), .B0_t (LED_128_Instance_MUX_state0_mux_inst_21_U1_X), .B0_f (new_AGEMA_signal_5313), .B1_t (new_AGEMA_signal_5314), .B1_f (new_AGEMA_signal_5315), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_21_U1_Y), .Z0_f (new_AGEMA_signal_5505), .Z1_t (new_AGEMA_signal_5506), .Z1_f (new_AGEMA_signal_5507) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_21_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_21_U1_Y), .A0_f (new_AGEMA_signal_5505), .A1_t (new_AGEMA_signal_5506), .A1_f (new_AGEMA_signal_5507), .B0_t (LED_128_Instance_mixcolumns_out[21]), .B0_f (new_AGEMA_signal_5199), .B1_t (new_AGEMA_signal_5200), .B1_f (new_AGEMA_signal_5201), .Z0_t (LED_128_Instance_state0[21]), .Z0_f (new_AGEMA_signal_5694), .Z1_t (new_AGEMA_signal_5695), .Z1_f (new_AGEMA_signal_5696) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_22_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[22]), .A0_f (new_AGEMA_signal_5580), .A1_t (new_AGEMA_signal_5581), .A1_f (new_AGEMA_signal_5582), .B0_t (LED_128_Instance_addroundkey_out[22]), .B0_f (new_AGEMA_signal_3702), .B1_t (new_AGEMA_signal_3703), .B1_f (new_AGEMA_signal_3704), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_22_U1_X), .Z0_f (new_AGEMA_signal_5697), .Z1_t (new_AGEMA_signal_5698), .Z1_f (new_AGEMA_signal_5699) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_22_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n22), .A1_f (new_AGEMA_signal_2479), .B0_t (LED_128_Instance_MUX_state0_mux_inst_22_U1_X), .B0_f (new_AGEMA_signal_5697), .B1_t (new_AGEMA_signal_5698), .B1_f (new_AGEMA_signal_5699), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_22_U1_Y), .Z0_f (new_AGEMA_signal_5877), .Z1_t (new_AGEMA_signal_5878), .Z1_f (new_AGEMA_signal_5879) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_22_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_22_U1_Y), .A0_f (new_AGEMA_signal_5877), .A1_t (new_AGEMA_signal_5878), .A1_f (new_AGEMA_signal_5879), .B0_t (LED_128_Instance_mixcolumns_out[22]), .B0_f (new_AGEMA_signal_5580), .B1_t (new_AGEMA_signal_5581), .B1_f (new_AGEMA_signal_5582), .Z0_t (LED_128_Instance_state0[22]), .Z0_f (new_AGEMA_signal_6078), .Z1_t (new_AGEMA_signal_6079), .Z1_f (new_AGEMA_signal_6080) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_23_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[23]), .A0_f (new_AGEMA_signal_5577), .A1_t (new_AGEMA_signal_5578), .A1_f (new_AGEMA_signal_5579), .B0_t (LED_128_Instance_addconst_out[23]), .B0_f (new_AGEMA_signal_3705), .B1_t (new_AGEMA_signal_3706), .B1_f (new_AGEMA_signal_3707), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_23_U1_X), .Z0_f (new_AGEMA_signal_5700), .Z1_t (new_AGEMA_signal_5701), .Z1_f (new_AGEMA_signal_5702) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_23_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n22), .A1_f (new_AGEMA_signal_2479), .B0_t (LED_128_Instance_MUX_state0_mux_inst_23_U1_X), .B0_f (new_AGEMA_signal_5700), .B1_t (new_AGEMA_signal_5701), .B1_f (new_AGEMA_signal_5702), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_23_U1_Y), .Z0_f (new_AGEMA_signal_5880), .Z1_t (new_AGEMA_signal_5881), .Z1_f (new_AGEMA_signal_5882) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_23_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_23_U1_Y), .A0_f (new_AGEMA_signal_5880), .A1_t (new_AGEMA_signal_5881), .A1_f (new_AGEMA_signal_5882), .B0_t (LED_128_Instance_mixcolumns_out[23]), .B0_f (new_AGEMA_signal_5577), .B1_t (new_AGEMA_signal_5578), .B1_f (new_AGEMA_signal_5579), .Z0_t (LED_128_Instance_state0[23]), .Z0_f (new_AGEMA_signal_6081), .Z1_t (new_AGEMA_signal_6082), .Z1_f (new_AGEMA_signal_6083) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_24_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[24]), .A0_f (new_AGEMA_signal_5418), .A1_t (new_AGEMA_signal_5419), .A1_f (new_AGEMA_signal_5420), .B0_t (LED_128_Instance_addconst_out[24]), .B0_f (new_AGEMA_signal_3708), .B1_t (new_AGEMA_signal_3709), .B1_f (new_AGEMA_signal_3710), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_24_U1_X), .Z0_f (new_AGEMA_signal_5508), .Z1_t (new_AGEMA_signal_5509), .Z1_f (new_AGEMA_signal_5510) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_24_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n22), .A1_f (new_AGEMA_signal_2479), .B0_t (LED_128_Instance_MUX_state0_mux_inst_24_U1_X), .B0_f (new_AGEMA_signal_5508), .B1_t (new_AGEMA_signal_5509), .B1_f (new_AGEMA_signal_5510), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_24_U1_Y), .Z0_f (new_AGEMA_signal_5703), .Z1_t (new_AGEMA_signal_5704), .Z1_f (new_AGEMA_signal_5705) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_24_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_24_U1_Y), .A0_f (new_AGEMA_signal_5703), .A1_t (new_AGEMA_signal_5704), .A1_f (new_AGEMA_signal_5705), .B0_t (LED_128_Instance_mixcolumns_out[24]), .B0_f (new_AGEMA_signal_5418), .B1_t (new_AGEMA_signal_5419), .B1_f (new_AGEMA_signal_5420), .Z0_t (LED_128_Instance_state0[24]), .Z0_f (new_AGEMA_signal_5883), .Z1_t (new_AGEMA_signal_5884), .Z1_f (new_AGEMA_signal_5885) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_25_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[25]), .A0_f (new_AGEMA_signal_5415), .A1_t (new_AGEMA_signal_5416), .A1_f (new_AGEMA_signal_5417), .B0_t (LED_128_Instance_addconst_out[25]), .B0_f (new_AGEMA_signal_3711), .B1_t (new_AGEMA_signal_3712), .B1_f (new_AGEMA_signal_3713), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_25_U1_X), .Z0_f (new_AGEMA_signal_5511), .Z1_t (new_AGEMA_signal_5512), .Z1_f (new_AGEMA_signal_5513) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_25_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n22), .A1_f (new_AGEMA_signal_2479), .B0_t (LED_128_Instance_MUX_state0_mux_inst_25_U1_X), .B0_f (new_AGEMA_signal_5511), .B1_t (new_AGEMA_signal_5512), .B1_f (new_AGEMA_signal_5513), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_25_U1_Y), .Z0_f (new_AGEMA_signal_5706), .Z1_t (new_AGEMA_signal_5707), .Z1_f (new_AGEMA_signal_5708) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_25_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_25_U1_Y), .A0_f (new_AGEMA_signal_5706), .A1_t (new_AGEMA_signal_5707), .A1_f (new_AGEMA_signal_5708), .B0_t (LED_128_Instance_mixcolumns_out[25]), .B0_f (new_AGEMA_signal_5415), .B1_t (new_AGEMA_signal_5416), .B1_f (new_AGEMA_signal_5417), .Z0_t (LED_128_Instance_state0[25]), .Z0_f (new_AGEMA_signal_5886), .Z1_t (new_AGEMA_signal_5887), .Z1_f (new_AGEMA_signal_5888) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_26_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[26]), .A0_f (new_AGEMA_signal_5601), .A1_t (new_AGEMA_signal_5602), .A1_f (new_AGEMA_signal_5603), .B0_t (LED_128_Instance_addconst_out[26]), .B0_f (new_AGEMA_signal_3714), .B1_t (new_AGEMA_signal_3715), .B1_f (new_AGEMA_signal_3716), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_26_U1_X), .Z0_f (new_AGEMA_signal_5709), .Z1_t (new_AGEMA_signal_5710), .Z1_f (new_AGEMA_signal_5711) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_26_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n22), .A1_f (new_AGEMA_signal_2479), .B0_t (LED_128_Instance_MUX_state0_mux_inst_26_U1_X), .B0_f (new_AGEMA_signal_5709), .B1_t (new_AGEMA_signal_5710), .B1_f (new_AGEMA_signal_5711), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_26_U1_Y), .Z0_f (new_AGEMA_signal_5889), .Z1_t (new_AGEMA_signal_5890), .Z1_f (new_AGEMA_signal_5891) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_26_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_26_U1_Y), .A0_f (new_AGEMA_signal_5889), .A1_t (new_AGEMA_signal_5890), .A1_f (new_AGEMA_signal_5891), .B0_t (LED_128_Instance_mixcolumns_out[26]), .B0_f (new_AGEMA_signal_5601), .B1_t (new_AGEMA_signal_5602), .B1_f (new_AGEMA_signal_5603), .Z0_t (LED_128_Instance_state0[26]), .Z0_f (new_AGEMA_signal_6084), .Z1_t (new_AGEMA_signal_6085), .Z1_f (new_AGEMA_signal_6086) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_27_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[27]), .A0_f (new_AGEMA_signal_5598), .A1_t (new_AGEMA_signal_5599), .A1_f (new_AGEMA_signal_5600), .B0_t (LED_128_Instance_addconst_out[27]), .B0_f (new_AGEMA_signal_3717), .B1_t (new_AGEMA_signal_3718), .B1_f (new_AGEMA_signal_3719), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_27_U1_X), .Z0_f (new_AGEMA_signal_5712), .Z1_t (new_AGEMA_signal_5713), .Z1_f (new_AGEMA_signal_5714) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_27_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n22), .A1_f (new_AGEMA_signal_2479), .B0_t (LED_128_Instance_MUX_state0_mux_inst_27_U1_X), .B0_f (new_AGEMA_signal_5712), .B1_t (new_AGEMA_signal_5713), .B1_f (new_AGEMA_signal_5714), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_27_U1_Y), .Z0_f (new_AGEMA_signal_5892), .Z1_t (new_AGEMA_signal_5893), .Z1_f (new_AGEMA_signal_5894) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_27_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_27_U1_Y), .A0_f (new_AGEMA_signal_5892), .A1_t (new_AGEMA_signal_5893), .A1_f (new_AGEMA_signal_5894), .B0_t (LED_128_Instance_mixcolumns_out[27]), .B0_f (new_AGEMA_signal_5598), .B1_t (new_AGEMA_signal_5599), .B1_f (new_AGEMA_signal_5600), .Z0_t (LED_128_Instance_state0[27]), .Z0_f (new_AGEMA_signal_6087), .Z1_t (new_AGEMA_signal_6088), .Z1_f (new_AGEMA_signal_6089) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_28_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[28]), .A0_f (new_AGEMA_signal_5448), .A1_t (new_AGEMA_signal_5449), .A1_f (new_AGEMA_signal_5450), .B0_t (LED_128_Instance_addconst_out[28]), .B0_f (new_AGEMA_signal_3720), .B1_t (new_AGEMA_signal_3721), .B1_f (new_AGEMA_signal_3722), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_28_U1_X), .Z0_f (new_AGEMA_signal_5514), .Z1_t (new_AGEMA_signal_5515), .Z1_f (new_AGEMA_signal_5516) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_28_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n22), .A1_f (new_AGEMA_signal_2479), .B0_t (LED_128_Instance_MUX_state0_mux_inst_28_U1_X), .B0_f (new_AGEMA_signal_5514), .B1_t (new_AGEMA_signal_5515), .B1_f (new_AGEMA_signal_5516), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_28_U1_Y), .Z0_f (new_AGEMA_signal_5715), .Z1_t (new_AGEMA_signal_5716), .Z1_f (new_AGEMA_signal_5717) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_28_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_28_U1_Y), .A0_f (new_AGEMA_signal_5715), .A1_t (new_AGEMA_signal_5716), .A1_f (new_AGEMA_signal_5717), .B0_t (LED_128_Instance_mixcolumns_out[28]), .B0_f (new_AGEMA_signal_5448), .B1_t (new_AGEMA_signal_5449), .B1_f (new_AGEMA_signal_5450), .Z0_t (LED_128_Instance_state0[28]), .Z0_f (new_AGEMA_signal_5895), .Z1_t (new_AGEMA_signal_5896), .Z1_f (new_AGEMA_signal_5897) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_29_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[29]), .A0_f (new_AGEMA_signal_5445), .A1_t (new_AGEMA_signal_5446), .A1_f (new_AGEMA_signal_5447), .B0_t (LED_128_Instance_addconst_out[29]), .B0_f (new_AGEMA_signal_3723), .B1_t (new_AGEMA_signal_3724), .B1_f (new_AGEMA_signal_3725), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_29_U1_X), .Z0_f (new_AGEMA_signal_5517), .Z1_t (new_AGEMA_signal_5518), .Z1_f (new_AGEMA_signal_5519) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_29_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n22), .A1_f (new_AGEMA_signal_2479), .B0_t (LED_128_Instance_MUX_state0_mux_inst_29_U1_X), .B0_f (new_AGEMA_signal_5517), .B1_t (new_AGEMA_signal_5518), .B1_f (new_AGEMA_signal_5519), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_29_U1_Y), .Z0_f (new_AGEMA_signal_5718), .Z1_t (new_AGEMA_signal_5719), .Z1_f (new_AGEMA_signal_5720) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_29_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_29_U1_Y), .A0_f (new_AGEMA_signal_5718), .A1_t (new_AGEMA_signal_5719), .A1_f (new_AGEMA_signal_5720), .B0_t (LED_128_Instance_mixcolumns_out[29]), .B0_f (new_AGEMA_signal_5445), .B1_t (new_AGEMA_signal_5446), .B1_f (new_AGEMA_signal_5447), .Z0_t (LED_128_Instance_state0[29]), .Z0_f (new_AGEMA_signal_5898), .Z1_t (new_AGEMA_signal_5899), .Z1_f (new_AGEMA_signal_5900) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_30_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[30]), .A0_f (new_AGEMA_signal_5838), .A1_t (new_AGEMA_signal_5839), .A1_f (new_AGEMA_signal_5840), .B0_t (LED_128_Instance_addconst_out[30]), .B0_f (new_AGEMA_signal_3726), .B1_t (new_AGEMA_signal_3727), .B1_f (new_AGEMA_signal_3728), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_30_U1_X), .Z0_f (new_AGEMA_signal_5901), .Z1_t (new_AGEMA_signal_5902), .Z1_f (new_AGEMA_signal_5903) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_30_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n22), .A1_f (new_AGEMA_signal_2479), .B0_t (LED_128_Instance_MUX_state0_mux_inst_30_U1_X), .B0_f (new_AGEMA_signal_5901), .B1_t (new_AGEMA_signal_5902), .B1_f (new_AGEMA_signal_5903), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_30_U1_Y), .Z0_f (new_AGEMA_signal_6090), .Z1_t (new_AGEMA_signal_6091), .Z1_f (new_AGEMA_signal_6092) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_30_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_30_U1_Y), .A0_f (new_AGEMA_signal_6090), .A1_t (new_AGEMA_signal_6091), .A1_f (new_AGEMA_signal_6092), .B0_t (LED_128_Instance_mixcolumns_out[30]), .B0_f (new_AGEMA_signal_5838), .B1_t (new_AGEMA_signal_5839), .B1_f (new_AGEMA_signal_5840), .Z0_t (LED_128_Instance_state0[30]), .Z0_f (new_AGEMA_signal_6309), .Z1_t (new_AGEMA_signal_6310), .Z1_f (new_AGEMA_signal_6311) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_31_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[31]), .A0_f (new_AGEMA_signal_5835), .A1_t (new_AGEMA_signal_5836), .A1_f (new_AGEMA_signal_5837), .B0_t (LED_128_Instance_addconst_out[31]), .B0_f (new_AGEMA_signal_3729), .B1_t (new_AGEMA_signal_3730), .B1_f (new_AGEMA_signal_3731), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_31_U1_X), .Z0_f (new_AGEMA_signal_5904), .Z1_t (new_AGEMA_signal_5905), .Z1_f (new_AGEMA_signal_5906) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_31_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n22), .A1_f (new_AGEMA_signal_2479), .B0_t (LED_128_Instance_MUX_state0_mux_inst_31_U1_X), .B0_f (new_AGEMA_signal_5904), .B1_t (new_AGEMA_signal_5905), .B1_f (new_AGEMA_signal_5906), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_31_U1_Y), .Z0_f (new_AGEMA_signal_6093), .Z1_t (new_AGEMA_signal_6094), .Z1_f (new_AGEMA_signal_6095) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_31_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_31_U1_Y), .A0_f (new_AGEMA_signal_6093), .A1_t (new_AGEMA_signal_6094), .A1_f (new_AGEMA_signal_6095), .B0_t (LED_128_Instance_mixcolumns_out[31]), .B0_f (new_AGEMA_signal_5835), .B1_t (new_AGEMA_signal_5836), .B1_f (new_AGEMA_signal_5837), .Z0_t (LED_128_Instance_state0[31]), .Z0_f (new_AGEMA_signal_6312), .Z1_t (new_AGEMA_signal_6313), .Z1_f (new_AGEMA_signal_6314) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_32_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[32]), .A0_f (new_AGEMA_signal_5820), .A1_t (new_AGEMA_signal_5821), .A1_f (new_AGEMA_signal_5822), .B0_t (LED_128_Instance_addconst_out[32]), .B0_f (new_AGEMA_signal_3732), .B1_t (new_AGEMA_signal_3733), .B1_f (new_AGEMA_signal_3734), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_32_U1_X), .Z0_f (new_AGEMA_signal_5907), .Z1_t (new_AGEMA_signal_5908), .Z1_f (new_AGEMA_signal_5909) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_32_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n22), .A1_f (new_AGEMA_signal_2479), .B0_t (LED_128_Instance_MUX_state0_mux_inst_32_U1_X), .B0_f (new_AGEMA_signal_5907), .B1_t (new_AGEMA_signal_5908), .B1_f (new_AGEMA_signal_5909), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_32_U1_Y), .Z0_f (new_AGEMA_signal_6096), .Z1_t (new_AGEMA_signal_6097), .Z1_f (new_AGEMA_signal_6098) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_32_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_32_U1_Y), .A0_f (new_AGEMA_signal_6096), .A1_t (new_AGEMA_signal_6097), .A1_f (new_AGEMA_signal_6098), .B0_t (LED_128_Instance_mixcolumns_out[32]), .B0_f (new_AGEMA_signal_5820), .B1_t (new_AGEMA_signal_5821), .B1_f (new_AGEMA_signal_5822), .Z0_t (LED_128_Instance_state0[32]), .Z0_f (new_AGEMA_signal_6315), .Z1_t (new_AGEMA_signal_6316), .Z1_f (new_AGEMA_signal_6317) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_33_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[33]), .A0_f (new_AGEMA_signal_5562), .A1_t (new_AGEMA_signal_5563), .A1_f (new_AGEMA_signal_5564), .B0_t (LED_128_Instance_addroundkey_out[33]), .B0_f (new_AGEMA_signal_3735), .B1_t (new_AGEMA_signal_3736), .B1_f (new_AGEMA_signal_3737), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_33_U1_X), .Z0_f (new_AGEMA_signal_5721), .Z1_t (new_AGEMA_signal_5722), .Z1_f (new_AGEMA_signal_5723) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_33_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n22), .A1_f (new_AGEMA_signal_2479), .B0_t (LED_128_Instance_MUX_state0_mux_inst_33_U1_X), .B0_f (new_AGEMA_signal_5721), .B1_t (new_AGEMA_signal_5722), .B1_f (new_AGEMA_signal_5723), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_33_U1_Y), .Z0_f (new_AGEMA_signal_5910), .Z1_t (new_AGEMA_signal_5911), .Z1_f (new_AGEMA_signal_5912) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_33_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_33_U1_Y), .A0_f (new_AGEMA_signal_5910), .A1_t (new_AGEMA_signal_5911), .A1_f (new_AGEMA_signal_5912), .B0_t (LED_128_Instance_mixcolumns_out[33]), .B0_f (new_AGEMA_signal_5562), .B1_t (new_AGEMA_signal_5563), .B1_f (new_AGEMA_signal_5564), .Z0_t (LED_128_Instance_state0[33]), .Z0_f (new_AGEMA_signal_6099), .Z1_t (new_AGEMA_signal_6100), .Z1_f (new_AGEMA_signal_6101) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_34_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[34]), .A0_f (new_AGEMA_signal_5328), .A1_t (new_AGEMA_signal_5329), .A1_f (new_AGEMA_signal_5330), .B0_t (LED_128_Instance_addconst_out[34]), .B0_f (new_AGEMA_signal_3738), .B1_t (new_AGEMA_signal_3739), .B1_f (new_AGEMA_signal_3740), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_34_U1_X), .Z0_f (new_AGEMA_signal_5520), .Z1_t (new_AGEMA_signal_5521), .Z1_f (new_AGEMA_signal_5522) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_34_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n22), .A1_f (new_AGEMA_signal_2479), .B0_t (LED_128_Instance_MUX_state0_mux_inst_34_U1_X), .B0_f (new_AGEMA_signal_5520), .B1_t (new_AGEMA_signal_5521), .B1_f (new_AGEMA_signal_5522), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_34_U1_Y), .Z0_f (new_AGEMA_signal_5724), .Z1_t (new_AGEMA_signal_5725), .Z1_f (new_AGEMA_signal_5726) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_34_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_34_U1_Y), .A0_f (new_AGEMA_signal_5724), .A1_t (new_AGEMA_signal_5725), .A1_f (new_AGEMA_signal_5726), .B0_t (LED_128_Instance_mixcolumns_out[34]), .B0_f (new_AGEMA_signal_5328), .B1_t (new_AGEMA_signal_5329), .B1_f (new_AGEMA_signal_5330), .Z0_t (LED_128_Instance_state0[34]), .Z0_f (new_AGEMA_signal_5913), .Z1_t (new_AGEMA_signal_5914), .Z1_f (new_AGEMA_signal_5915) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_35_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[35]), .A0_f (new_AGEMA_signal_5325), .A1_t (new_AGEMA_signal_5326), .A1_f (new_AGEMA_signal_5327), .B0_t (LED_128_Instance_addconst_out[35]), .B0_f (new_AGEMA_signal_3741), .B1_t (new_AGEMA_signal_3742), .B1_f (new_AGEMA_signal_3743), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_35_U1_X), .Z0_f (new_AGEMA_signal_5523), .Z1_t (new_AGEMA_signal_5524), .Z1_f (new_AGEMA_signal_5525) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_35_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n22), .A1_f (new_AGEMA_signal_2479), .B0_t (LED_128_Instance_MUX_state0_mux_inst_35_U1_X), .B0_f (new_AGEMA_signal_5523), .B1_t (new_AGEMA_signal_5524), .B1_f (new_AGEMA_signal_5525), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_35_U1_Y), .Z0_f (new_AGEMA_signal_5727), .Z1_t (new_AGEMA_signal_5728), .Z1_f (new_AGEMA_signal_5729) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_35_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_35_U1_Y), .A0_f (new_AGEMA_signal_5727), .A1_t (new_AGEMA_signal_5728), .A1_f (new_AGEMA_signal_5729), .B0_t (LED_128_Instance_mixcolumns_out[35]), .B0_f (new_AGEMA_signal_5325), .B1_t (new_AGEMA_signal_5326), .B1_f (new_AGEMA_signal_5327), .Z0_t (LED_128_Instance_state0[35]), .Z0_f (new_AGEMA_signal_5916), .Z1_t (new_AGEMA_signal_5917), .Z1_f (new_AGEMA_signal_5918) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_36_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[36]), .A0_f (new_AGEMA_signal_5823), .A1_t (new_AGEMA_signal_5824), .A1_f (new_AGEMA_signal_5825), .B0_t (LED_128_Instance_addroundkey_out[36]), .B0_f (new_AGEMA_signal_3744), .B1_t (new_AGEMA_signal_3745), .B1_f (new_AGEMA_signal_3746), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_36_U1_X), .Z0_f (new_AGEMA_signal_5919), .Z1_t (new_AGEMA_signal_5920), .Z1_f (new_AGEMA_signal_5921) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_36_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n22), .A1_f (new_AGEMA_signal_2479), .B0_t (LED_128_Instance_MUX_state0_mux_inst_36_U1_X), .B0_f (new_AGEMA_signal_5919), .B1_t (new_AGEMA_signal_5920), .B1_f (new_AGEMA_signal_5921), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_36_U1_Y), .Z0_f (new_AGEMA_signal_6102), .Z1_t (new_AGEMA_signal_6103), .Z1_f (new_AGEMA_signal_6104) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_36_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_36_U1_Y), .A0_f (new_AGEMA_signal_6102), .A1_t (new_AGEMA_signal_6103), .A1_f (new_AGEMA_signal_6104), .B0_t (LED_128_Instance_mixcolumns_out[36]), .B0_f (new_AGEMA_signal_5823), .B1_t (new_AGEMA_signal_5824), .B1_f (new_AGEMA_signal_5825), .Z0_t (LED_128_Instance_state0[36]), .Z0_f (new_AGEMA_signal_6318), .Z1_t (new_AGEMA_signal_6319), .Z1_f (new_AGEMA_signal_6320) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_37_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[37]), .A0_f (new_AGEMA_signal_5586), .A1_t (new_AGEMA_signal_5587), .A1_f (new_AGEMA_signal_5588), .B0_t (LED_128_Instance_addroundkey_out[37]), .B0_f (new_AGEMA_signal_3747), .B1_t (new_AGEMA_signal_3748), .B1_f (new_AGEMA_signal_3749), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_37_U1_X), .Z0_f (new_AGEMA_signal_5730), .Z1_t (new_AGEMA_signal_5731), .Z1_f (new_AGEMA_signal_5732) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_37_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n22), .A1_f (new_AGEMA_signal_2479), .B0_t (LED_128_Instance_MUX_state0_mux_inst_37_U1_X), .B0_f (new_AGEMA_signal_5730), .B1_t (new_AGEMA_signal_5731), .B1_f (new_AGEMA_signal_5732), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_37_U1_Y), .Z0_f (new_AGEMA_signal_5922), .Z1_t (new_AGEMA_signal_5923), .Z1_f (new_AGEMA_signal_5924) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_37_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_37_U1_Y), .A0_f (new_AGEMA_signal_5922), .A1_t (new_AGEMA_signal_5923), .A1_f (new_AGEMA_signal_5924), .B0_t (LED_128_Instance_mixcolumns_out[37]), .B0_f (new_AGEMA_signal_5586), .B1_t (new_AGEMA_signal_5587), .B1_f (new_AGEMA_signal_5588), .Z0_t (LED_128_Instance_state0[37]), .Z0_f (new_AGEMA_signal_6105), .Z1_t (new_AGEMA_signal_6106), .Z1_f (new_AGEMA_signal_6107) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_38_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[38]), .A0_f (new_AGEMA_signal_5367), .A1_t (new_AGEMA_signal_5368), .A1_f (new_AGEMA_signal_5369), .B0_t (LED_128_Instance_addroundkey_out[38]), .B0_f (new_AGEMA_signal_3750), .B1_t (new_AGEMA_signal_3751), .B1_f (new_AGEMA_signal_3752), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_38_U1_X), .Z0_f (new_AGEMA_signal_5526), .Z1_t (new_AGEMA_signal_5527), .Z1_f (new_AGEMA_signal_5528) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_38_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n22), .A1_f (new_AGEMA_signal_2479), .B0_t (LED_128_Instance_MUX_state0_mux_inst_38_U1_X), .B0_f (new_AGEMA_signal_5526), .B1_t (new_AGEMA_signal_5527), .B1_f (new_AGEMA_signal_5528), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_38_U1_Y), .Z0_f (new_AGEMA_signal_5733), .Z1_t (new_AGEMA_signal_5734), .Z1_f (new_AGEMA_signal_5735) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_38_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_38_U1_Y), .A0_f (new_AGEMA_signal_5733), .A1_t (new_AGEMA_signal_5734), .A1_f (new_AGEMA_signal_5735), .B0_t (LED_128_Instance_mixcolumns_out[38]), .B0_f (new_AGEMA_signal_5367), .B1_t (new_AGEMA_signal_5368), .B1_f (new_AGEMA_signal_5369), .Z0_t (LED_128_Instance_state0[38]), .Z0_f (new_AGEMA_signal_5925), .Z1_t (new_AGEMA_signal_5926), .Z1_f (new_AGEMA_signal_5927) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_39_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[39]), .A0_f (new_AGEMA_signal_5583), .A1_t (new_AGEMA_signal_5584), .A1_f (new_AGEMA_signal_5585), .B0_t (LED_128_Instance_addconst_out[39]), .B0_f (new_AGEMA_signal_3753), .B1_t (new_AGEMA_signal_3754), .B1_f (new_AGEMA_signal_3755), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_39_U1_X), .Z0_f (new_AGEMA_signal_5736), .Z1_t (new_AGEMA_signal_5737), .Z1_f (new_AGEMA_signal_5738) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_39_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n22), .A1_f (new_AGEMA_signal_2479), .B0_t (LED_128_Instance_MUX_state0_mux_inst_39_U1_X), .B0_f (new_AGEMA_signal_5736), .B1_t (new_AGEMA_signal_5737), .B1_f (new_AGEMA_signal_5738), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_39_U1_Y), .Z0_f (new_AGEMA_signal_5928), .Z1_t (new_AGEMA_signal_5929), .Z1_f (new_AGEMA_signal_5930) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_39_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_39_U1_Y), .A0_f (new_AGEMA_signal_5928), .A1_t (new_AGEMA_signal_5929), .A1_f (new_AGEMA_signal_5930), .B0_t (LED_128_Instance_mixcolumns_out[39]), .B0_f (new_AGEMA_signal_5583), .B1_t (new_AGEMA_signal_5584), .B1_f (new_AGEMA_signal_5585), .Z0_t (LED_128_Instance_state0[39]), .Z0_f (new_AGEMA_signal_6108), .Z1_t (new_AGEMA_signal_6109), .Z1_f (new_AGEMA_signal_6110) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_40_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[40]), .A0_f (new_AGEMA_signal_5826), .A1_t (new_AGEMA_signal_5827), .A1_f (new_AGEMA_signal_5828), .B0_t (LED_128_Instance_addconst_out[40]), .B0_f (new_AGEMA_signal_3756), .B1_t (new_AGEMA_signal_3757), .B1_f (new_AGEMA_signal_3758), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_40_U1_X), .Z0_f (new_AGEMA_signal_5931), .Z1_t (new_AGEMA_signal_5932), .Z1_f (new_AGEMA_signal_5933) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_40_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n22), .A1_f (new_AGEMA_signal_2479), .B0_t (LED_128_Instance_MUX_state0_mux_inst_40_U1_X), .B0_f (new_AGEMA_signal_5931), .B1_t (new_AGEMA_signal_5932), .B1_f (new_AGEMA_signal_5933), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_40_U1_Y), .Z0_f (new_AGEMA_signal_6111), .Z1_t (new_AGEMA_signal_6112), .Z1_f (new_AGEMA_signal_6113) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_40_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_40_U1_Y), .A0_f (new_AGEMA_signal_6111), .A1_t (new_AGEMA_signal_6112), .A1_f (new_AGEMA_signal_6113), .B0_t (LED_128_Instance_mixcolumns_out[40]), .B0_f (new_AGEMA_signal_5826), .B1_t (new_AGEMA_signal_5827), .B1_f (new_AGEMA_signal_5828), .Z0_t (LED_128_Instance_state0[40]), .Z0_f (new_AGEMA_signal_6321), .Z1_t (new_AGEMA_signal_6322), .Z1_f (new_AGEMA_signal_6323) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_41_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[41]), .A0_f (new_AGEMA_signal_5604), .A1_t (new_AGEMA_signal_5605), .A1_f (new_AGEMA_signal_5606), .B0_t (LED_128_Instance_addconst_out[41]), .B0_f (new_AGEMA_signal_3759), .B1_t (new_AGEMA_signal_3760), .B1_f (new_AGEMA_signal_3761), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_41_U1_X), .Z0_f (new_AGEMA_signal_5739), .Z1_t (new_AGEMA_signal_5740), .Z1_f (new_AGEMA_signal_5741) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_41_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n22), .A1_f (new_AGEMA_signal_2479), .B0_t (LED_128_Instance_MUX_state0_mux_inst_41_U1_X), .B0_f (new_AGEMA_signal_5739), .B1_t (new_AGEMA_signal_5740), .B1_f (new_AGEMA_signal_5741), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_41_U1_Y), .Z0_f (new_AGEMA_signal_5934), .Z1_t (new_AGEMA_signal_5935), .Z1_f (new_AGEMA_signal_5936) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_41_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_41_U1_Y), .A0_f (new_AGEMA_signal_5934), .A1_t (new_AGEMA_signal_5935), .A1_f (new_AGEMA_signal_5936), .B0_t (LED_128_Instance_mixcolumns_out[41]), .B0_f (new_AGEMA_signal_5604), .B1_t (new_AGEMA_signal_5605), .B1_f (new_AGEMA_signal_5606), .Z0_t (LED_128_Instance_state0[41]), .Z0_f (new_AGEMA_signal_6114), .Z1_t (new_AGEMA_signal_6115), .Z1_f (new_AGEMA_signal_6116) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_42_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[42]), .A0_f (new_AGEMA_signal_5397), .A1_t (new_AGEMA_signal_5398), .A1_f (new_AGEMA_signal_5399), .B0_t (LED_128_Instance_addconst_out[42]), .B0_f (new_AGEMA_signal_3762), .B1_t (new_AGEMA_signal_3763), .B1_f (new_AGEMA_signal_3764), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_42_U1_X), .Z0_f (new_AGEMA_signal_5529), .Z1_t (new_AGEMA_signal_5530), .Z1_f (new_AGEMA_signal_5531) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_42_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n22), .A1_f (new_AGEMA_signal_2479), .B0_t (LED_128_Instance_MUX_state0_mux_inst_42_U1_X), .B0_f (new_AGEMA_signal_5529), .B1_t (new_AGEMA_signal_5530), .B1_f (new_AGEMA_signal_5531), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_42_U1_Y), .Z0_f (new_AGEMA_signal_5742), .Z1_t (new_AGEMA_signal_5743), .Z1_f (new_AGEMA_signal_5744) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_42_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_42_U1_Y), .A0_f (new_AGEMA_signal_5742), .A1_t (new_AGEMA_signal_5743), .A1_f (new_AGEMA_signal_5744), .B0_t (LED_128_Instance_mixcolumns_out[42]), .B0_f (new_AGEMA_signal_5397), .B1_t (new_AGEMA_signal_5398), .B1_f (new_AGEMA_signal_5399), .Z0_t (LED_128_Instance_state0[42]), .Z0_f (new_AGEMA_signal_5937), .Z1_t (new_AGEMA_signal_5938), .Z1_f (new_AGEMA_signal_5939) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_43_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[43]), .A0_f (new_AGEMA_signal_5394), .A1_t (new_AGEMA_signal_5395), .A1_f (new_AGEMA_signal_5396), .B0_t (LED_128_Instance_addconst_out[43]), .B0_f (new_AGEMA_signal_3765), .B1_t (new_AGEMA_signal_3766), .B1_f (new_AGEMA_signal_3767), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_43_U1_X), .Z0_f (new_AGEMA_signal_5532), .Z1_t (new_AGEMA_signal_5533), .Z1_f (new_AGEMA_signal_5534) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_43_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n22), .A1_f (new_AGEMA_signal_2479), .B0_t (LED_128_Instance_MUX_state0_mux_inst_43_U1_X), .B0_f (new_AGEMA_signal_5532), .B1_t (new_AGEMA_signal_5533), .B1_f (new_AGEMA_signal_5534), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_43_U1_Y), .Z0_f (new_AGEMA_signal_5745), .Z1_t (new_AGEMA_signal_5746), .Z1_f (new_AGEMA_signal_5747) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_43_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_43_U1_Y), .A0_f (new_AGEMA_signal_5745), .A1_t (new_AGEMA_signal_5746), .A1_f (new_AGEMA_signal_5747), .B0_t (LED_128_Instance_mixcolumns_out[43]), .B0_f (new_AGEMA_signal_5394), .B1_t (new_AGEMA_signal_5395), .B1_f (new_AGEMA_signal_5396), .Z0_t (LED_128_Instance_state0[43]), .Z0_f (new_AGEMA_signal_5940), .Z1_t (new_AGEMA_signal_5941), .Z1_f (new_AGEMA_signal_5942) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_44_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[44]), .A0_f (new_AGEMA_signal_6063), .A1_t (new_AGEMA_signal_6064), .A1_f (new_AGEMA_signal_6065), .B0_t (LED_128_Instance_addconst_out[44]), .B0_f (new_AGEMA_signal_3768), .B1_t (new_AGEMA_signal_3769), .B1_f (new_AGEMA_signal_3770), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_44_U1_X), .Z0_f (new_AGEMA_signal_6117), .Z1_t (new_AGEMA_signal_6118), .Z1_f (new_AGEMA_signal_6119) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_44_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n22), .A1_f (new_AGEMA_signal_2479), .B0_t (LED_128_Instance_MUX_state0_mux_inst_44_U1_X), .B0_f (new_AGEMA_signal_6117), .B1_t (new_AGEMA_signal_6118), .B1_f (new_AGEMA_signal_6119), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_44_U1_Y), .Z0_f (new_AGEMA_signal_6324), .Z1_t (new_AGEMA_signal_6325), .Z1_f (new_AGEMA_signal_6326) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_44_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_44_U1_Y), .A0_f (new_AGEMA_signal_6324), .A1_t (new_AGEMA_signal_6325), .A1_f (new_AGEMA_signal_6326), .B0_t (LED_128_Instance_mixcolumns_out[44]), .B0_f (new_AGEMA_signal_6063), .B1_t (new_AGEMA_signal_6064), .B1_f (new_AGEMA_signal_6065), .Z0_t (LED_128_Instance_state0[44]), .Z0_f (new_AGEMA_signal_6525), .Z1_t (new_AGEMA_signal_6526), .Z1_f (new_AGEMA_signal_6527) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_45_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[45]), .A0_f (new_AGEMA_signal_5841), .A1_t (new_AGEMA_signal_5842), .A1_f (new_AGEMA_signal_5843), .B0_t (LED_128_Instance_addconst_out[45]), .B0_f (new_AGEMA_signal_3771), .B1_t (new_AGEMA_signal_3772), .B1_f (new_AGEMA_signal_3773), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_45_U1_X), .Z0_f (new_AGEMA_signal_5943), .Z1_t (new_AGEMA_signal_5944), .Z1_f (new_AGEMA_signal_5945) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_45_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n22), .A1_f (new_AGEMA_signal_2479), .B0_t (LED_128_Instance_MUX_state0_mux_inst_45_U1_X), .B0_f (new_AGEMA_signal_5943), .B1_t (new_AGEMA_signal_5944), .B1_f (new_AGEMA_signal_5945), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_45_U1_Y), .Z0_f (new_AGEMA_signal_6120), .Z1_t (new_AGEMA_signal_6121), .Z1_f (new_AGEMA_signal_6122) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_45_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_45_U1_Y), .A0_f (new_AGEMA_signal_6120), .A1_t (new_AGEMA_signal_6121), .A1_f (new_AGEMA_signal_6122), .B0_t (LED_128_Instance_mixcolumns_out[45]), .B0_f (new_AGEMA_signal_5841), .B1_t (new_AGEMA_signal_5842), .B1_f (new_AGEMA_signal_5843), .Z0_t (LED_128_Instance_state0[45]), .Z0_f (new_AGEMA_signal_6327), .Z1_t (new_AGEMA_signal_6328), .Z1_f (new_AGEMA_signal_6329) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_46_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[46]), .A0_f (new_AGEMA_signal_5628), .A1_t (new_AGEMA_signal_5629), .A1_f (new_AGEMA_signal_5630), .B0_t (LED_128_Instance_addconst_out[46]), .B0_f (new_AGEMA_signal_3774), .B1_t (new_AGEMA_signal_3775), .B1_f (new_AGEMA_signal_3776), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_46_U1_X), .Z0_f (new_AGEMA_signal_5748), .Z1_t (new_AGEMA_signal_5749), .Z1_f (new_AGEMA_signal_5750) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_46_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n22), .A1_f (new_AGEMA_signal_2479), .B0_t (LED_128_Instance_MUX_state0_mux_inst_46_U1_X), .B0_f (new_AGEMA_signal_5748), .B1_t (new_AGEMA_signal_5749), .B1_f (new_AGEMA_signal_5750), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_46_U1_Y), .Z0_f (new_AGEMA_signal_5946), .Z1_t (new_AGEMA_signal_5947), .Z1_f (new_AGEMA_signal_5948) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_46_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_46_U1_Y), .A0_f (new_AGEMA_signal_5946), .A1_t (new_AGEMA_signal_5947), .A1_f (new_AGEMA_signal_5948), .B0_t (LED_128_Instance_mixcolumns_out[46]), .B0_f (new_AGEMA_signal_5628), .B1_t (new_AGEMA_signal_5629), .B1_f (new_AGEMA_signal_5630), .Z0_t (LED_128_Instance_state0[46]), .Z0_f (new_AGEMA_signal_6123), .Z1_t (new_AGEMA_signal_6124), .Z1_f (new_AGEMA_signal_6125) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_47_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[47]), .A0_f (new_AGEMA_signal_5625), .A1_t (new_AGEMA_signal_5626), .A1_f (new_AGEMA_signal_5627), .B0_t (LED_128_Instance_addconst_out[47]), .B0_f (new_AGEMA_signal_3777), .B1_t (new_AGEMA_signal_3778), .B1_f (new_AGEMA_signal_3779), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_47_U1_X), .Z0_f (new_AGEMA_signal_5751), .Z1_t (new_AGEMA_signal_5752), .Z1_f (new_AGEMA_signal_5753) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_47_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n22), .A1_f (new_AGEMA_signal_2479), .B0_t (LED_128_Instance_MUX_state0_mux_inst_47_U1_X), .B0_f (new_AGEMA_signal_5751), .B1_t (new_AGEMA_signal_5752), .B1_f (new_AGEMA_signal_5753), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_47_U1_Y), .Z0_f (new_AGEMA_signal_5949), .Z1_t (new_AGEMA_signal_5950), .Z1_f (new_AGEMA_signal_5951) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_47_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_47_U1_Y), .A0_f (new_AGEMA_signal_5949), .A1_t (new_AGEMA_signal_5950), .A1_f (new_AGEMA_signal_5951), .B0_t (LED_128_Instance_mixcolumns_out[47]), .B0_f (new_AGEMA_signal_5625), .B1_t (new_AGEMA_signal_5626), .B1_f (new_AGEMA_signal_5627), .Z0_t (LED_128_Instance_state0[47]), .Z0_f (new_AGEMA_signal_6126), .Z1_t (new_AGEMA_signal_6127), .Z1_f (new_AGEMA_signal_6128) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_48_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[48]), .A0_f (new_AGEMA_signal_5571), .A1_t (new_AGEMA_signal_5572), .A1_f (new_AGEMA_signal_5573), .B0_t (LED_128_Instance_addroundkey_out[48]), .B0_f (new_AGEMA_signal_3780), .B1_t (new_AGEMA_signal_3781), .B1_f (new_AGEMA_signal_3782), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_48_U1_X), .Z0_f (new_AGEMA_signal_5754), .Z1_t (new_AGEMA_signal_5755), .Z1_f (new_AGEMA_signal_5756) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_48_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n22), .A1_f (new_AGEMA_signal_2479), .B0_t (LED_128_Instance_MUX_state0_mux_inst_48_U1_X), .B0_f (new_AGEMA_signal_5754), .B1_t (new_AGEMA_signal_5755), .B1_f (new_AGEMA_signal_5756), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_48_U1_Y), .Z0_f (new_AGEMA_signal_5952), .Z1_t (new_AGEMA_signal_5953), .Z1_f (new_AGEMA_signal_5954) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_48_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_48_U1_Y), .A0_f (new_AGEMA_signal_5952), .A1_t (new_AGEMA_signal_5953), .A1_f (new_AGEMA_signal_5954), .B0_t (LED_128_Instance_mixcolumns_out[48]), .B0_f (new_AGEMA_signal_5571), .B1_t (new_AGEMA_signal_5572), .B1_f (new_AGEMA_signal_5573), .Z0_t (LED_128_Instance_state0[48]), .Z0_f (new_AGEMA_signal_6129), .Z1_t (new_AGEMA_signal_6130), .Z1_f (new_AGEMA_signal_6131) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_49_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[49]), .A0_f (new_AGEMA_signal_5568), .A1_t (new_AGEMA_signal_5569), .A1_f (new_AGEMA_signal_5570), .B0_t (LED_128_Instance_addroundkey_out[49]), .B0_f (new_AGEMA_signal_3783), .B1_t (new_AGEMA_signal_3784), .B1_f (new_AGEMA_signal_3785), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_49_U1_X), .Z0_f (new_AGEMA_signal_5757), .Z1_t (new_AGEMA_signal_5758), .Z1_f (new_AGEMA_signal_5759) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_49_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n22), .A1_f (new_AGEMA_signal_2479), .B0_t (LED_128_Instance_MUX_state0_mux_inst_49_U1_X), .B0_f (new_AGEMA_signal_5757), .B1_t (new_AGEMA_signal_5758), .B1_f (new_AGEMA_signal_5759), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_49_U1_Y), .Z0_f (new_AGEMA_signal_5955), .Z1_t (new_AGEMA_signal_5956), .Z1_f (new_AGEMA_signal_5957) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_49_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_49_U1_Y), .A0_f (new_AGEMA_signal_5955), .A1_t (new_AGEMA_signal_5956), .A1_f (new_AGEMA_signal_5957), .B0_t (LED_128_Instance_mixcolumns_out[49]), .B0_f (new_AGEMA_signal_5568), .B1_t (new_AGEMA_signal_5569), .B1_f (new_AGEMA_signal_5570), .Z0_t (LED_128_Instance_state0[49]), .Z0_f (new_AGEMA_signal_6132), .Z1_t (new_AGEMA_signal_6133), .Z1_f (new_AGEMA_signal_6134) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_50_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[50]), .A0_f (new_AGEMA_signal_5355), .A1_t (new_AGEMA_signal_5356), .A1_f (new_AGEMA_signal_5357), .B0_t (LED_128_Instance_addconst_out[50]), .B0_f (new_AGEMA_signal_3786), .B1_t (new_AGEMA_signal_3787), .B1_f (new_AGEMA_signal_3788), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_50_U1_X), .Z0_f (new_AGEMA_signal_5535), .Z1_t (new_AGEMA_signal_5536), .Z1_f (new_AGEMA_signal_5537) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_50_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n22), .A1_f (new_AGEMA_signal_2479), .B0_t (LED_128_Instance_MUX_state0_mux_inst_50_U1_X), .B0_f (new_AGEMA_signal_5535), .B1_t (new_AGEMA_signal_5536), .B1_f (new_AGEMA_signal_5537), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_50_U1_Y), .Z0_f (new_AGEMA_signal_5760), .Z1_t (new_AGEMA_signal_5761), .Z1_f (new_AGEMA_signal_5762) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_50_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_50_U1_Y), .A0_f (new_AGEMA_signal_5760), .A1_t (new_AGEMA_signal_5761), .A1_f (new_AGEMA_signal_5762), .B0_t (LED_128_Instance_mixcolumns_out[50]), .B0_f (new_AGEMA_signal_5355), .B1_t (new_AGEMA_signal_5356), .B1_f (new_AGEMA_signal_5357), .Z0_t (LED_128_Instance_state0[50]), .Z0_f (new_AGEMA_signal_5958), .Z1_t (new_AGEMA_signal_5959), .Z1_f (new_AGEMA_signal_5960) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_51_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[51]), .A0_f (new_AGEMA_signal_5337), .A1_t (new_AGEMA_signal_5338), .A1_f (new_AGEMA_signal_5339), .B0_t (LED_128_Instance_addconst_out[51]), .B0_f (new_AGEMA_signal_3789), .B1_t (new_AGEMA_signal_3790), .B1_f (new_AGEMA_signal_3791), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_51_U1_X), .Z0_f (new_AGEMA_signal_5538), .Z1_t (new_AGEMA_signal_5539), .Z1_f (new_AGEMA_signal_5540) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_51_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n22), .A1_f (new_AGEMA_signal_2479), .B0_t (LED_128_Instance_MUX_state0_mux_inst_51_U1_X), .B0_f (new_AGEMA_signal_5538), .B1_t (new_AGEMA_signal_5539), .B1_f (new_AGEMA_signal_5540), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_51_U1_Y), .Z0_f (new_AGEMA_signal_5763), .Z1_t (new_AGEMA_signal_5764), .Z1_f (new_AGEMA_signal_5765) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_51_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_51_U1_Y), .A0_f (new_AGEMA_signal_5763), .A1_t (new_AGEMA_signal_5764), .A1_f (new_AGEMA_signal_5765), .B0_t (LED_128_Instance_mixcolumns_out[51]), .B0_f (new_AGEMA_signal_5337), .B1_t (new_AGEMA_signal_5338), .B1_f (new_AGEMA_signal_5339), .Z0_t (LED_128_Instance_state0[51]), .Z0_f (new_AGEMA_signal_5961), .Z1_t (new_AGEMA_signal_5962), .Z1_f (new_AGEMA_signal_5963) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_52_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[52]), .A0_f (new_AGEMA_signal_5595), .A1_t (new_AGEMA_signal_5596), .A1_f (new_AGEMA_signal_5597), .B0_t (LED_128_Instance_addroundkey_out[52]), .B0_f (new_AGEMA_signal_3792), .B1_t (new_AGEMA_signal_3793), .B1_f (new_AGEMA_signal_3794), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_52_U1_X), .Z0_f (new_AGEMA_signal_5766), .Z1_t (new_AGEMA_signal_5767), .Z1_f (new_AGEMA_signal_5768) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_52_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n22), .A1_f (new_AGEMA_signal_2479), .B0_t (LED_128_Instance_MUX_state0_mux_inst_52_U1_X), .B0_f (new_AGEMA_signal_5766), .B1_t (new_AGEMA_signal_5767), .B1_f (new_AGEMA_signal_5768), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_52_U1_Y), .Z0_f (new_AGEMA_signal_5964), .Z1_t (new_AGEMA_signal_5965), .Z1_f (new_AGEMA_signal_5966) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_52_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_52_U1_Y), .A0_f (new_AGEMA_signal_5964), .A1_t (new_AGEMA_signal_5965), .A1_f (new_AGEMA_signal_5966), .B0_t (LED_128_Instance_mixcolumns_out[52]), .B0_f (new_AGEMA_signal_5595), .B1_t (new_AGEMA_signal_5596), .B1_f (new_AGEMA_signal_5597), .Z0_t (LED_128_Instance_state0[52]), .Z0_f (new_AGEMA_signal_6135), .Z1_t (new_AGEMA_signal_6136), .Z1_f (new_AGEMA_signal_6137) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_53_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[53]), .A0_f (new_AGEMA_signal_5592), .A1_t (new_AGEMA_signal_5593), .A1_f (new_AGEMA_signal_5594), .B0_t (LED_128_Instance_addroundkey_out[53]), .B0_f (new_AGEMA_signal_3795), .B1_t (new_AGEMA_signal_3796), .B1_f (new_AGEMA_signal_3797), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_53_U1_X), .Z0_f (new_AGEMA_signal_5769), .Z1_t (new_AGEMA_signal_5770), .Z1_f (new_AGEMA_signal_5771) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_53_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n22), .A1_f (new_AGEMA_signal_2479), .B0_t (LED_128_Instance_MUX_state0_mux_inst_53_U1_X), .B0_f (new_AGEMA_signal_5769), .B1_t (new_AGEMA_signal_5770), .B1_f (new_AGEMA_signal_5771), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_53_U1_Y), .Z0_f (new_AGEMA_signal_5967), .Z1_t (new_AGEMA_signal_5968), .Z1_f (new_AGEMA_signal_5969) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_53_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_53_U1_Y), .A0_f (new_AGEMA_signal_5967), .A1_t (new_AGEMA_signal_5968), .A1_f (new_AGEMA_signal_5969), .B0_t (LED_128_Instance_mixcolumns_out[53]), .B0_f (new_AGEMA_signal_5592), .B1_t (new_AGEMA_signal_5593), .B1_f (new_AGEMA_signal_5594), .Z0_t (LED_128_Instance_state0[53]), .Z0_f (new_AGEMA_signal_6138), .Z1_t (new_AGEMA_signal_6139), .Z1_f (new_AGEMA_signal_6140) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_54_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[54]), .A0_f (new_AGEMA_signal_5385), .A1_t (new_AGEMA_signal_5386), .A1_f (new_AGEMA_signal_5387), .B0_t (LED_128_Instance_addroundkey_out[54]), .B0_f (new_AGEMA_signal_3798), .B1_t (new_AGEMA_signal_3799), .B1_f (new_AGEMA_signal_3800), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_54_U1_X), .Z0_f (new_AGEMA_signal_5541), .Z1_t (new_AGEMA_signal_5542), .Z1_f (new_AGEMA_signal_5543) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_54_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n22), .A1_f (new_AGEMA_signal_2479), .B0_t (LED_128_Instance_MUX_state0_mux_inst_54_U1_X), .B0_f (new_AGEMA_signal_5541), .B1_t (new_AGEMA_signal_5542), .B1_f (new_AGEMA_signal_5543), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_54_U1_Y), .Z0_f (new_AGEMA_signal_5772), .Z1_t (new_AGEMA_signal_5773), .Z1_f (new_AGEMA_signal_5774) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_54_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_54_U1_Y), .A0_f (new_AGEMA_signal_5772), .A1_t (new_AGEMA_signal_5773), .A1_f (new_AGEMA_signal_5774), .B0_t (LED_128_Instance_mixcolumns_out[54]), .B0_f (new_AGEMA_signal_5385), .B1_t (new_AGEMA_signal_5386), .B1_f (new_AGEMA_signal_5387), .Z0_t (LED_128_Instance_state0[54]), .Z0_f (new_AGEMA_signal_5970), .Z1_t (new_AGEMA_signal_5971), .Z1_f (new_AGEMA_signal_5972) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_55_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[55]), .A0_f (new_AGEMA_signal_5187), .A1_t (new_AGEMA_signal_5188), .A1_f (new_AGEMA_signal_5189), .B0_t (LED_128_Instance_addconst_out[55]), .B0_f (new_AGEMA_signal_3801), .B1_t (new_AGEMA_signal_3802), .B1_f (new_AGEMA_signal_3803), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_55_U1_X), .Z0_f (new_AGEMA_signal_5316), .Z1_t (new_AGEMA_signal_5317), .Z1_f (new_AGEMA_signal_5318) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_55_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n22), .A1_f (new_AGEMA_signal_2479), .B0_t (LED_128_Instance_MUX_state0_mux_inst_55_U1_X), .B0_f (new_AGEMA_signal_5316), .B1_t (new_AGEMA_signal_5317), .B1_f (new_AGEMA_signal_5318), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_55_U1_Y), .Z0_f (new_AGEMA_signal_5544), .Z1_t (new_AGEMA_signal_5545), .Z1_f (new_AGEMA_signal_5546) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_55_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_55_U1_Y), .A0_f (new_AGEMA_signal_5544), .A1_t (new_AGEMA_signal_5545), .A1_f (new_AGEMA_signal_5546), .B0_t (LED_128_Instance_mixcolumns_out[55]), .B0_f (new_AGEMA_signal_5187), .B1_t (new_AGEMA_signal_5188), .B1_f (new_AGEMA_signal_5189), .Z0_t (LED_128_Instance_state0[55]), .Z0_f (new_AGEMA_signal_5775), .Z1_t (new_AGEMA_signal_5776), .Z1_f (new_AGEMA_signal_5777) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_56_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[56]), .A0_f (new_AGEMA_signal_5832), .A1_t (new_AGEMA_signal_5833), .A1_f (new_AGEMA_signal_5834), .B0_t (LED_128_Instance_addconst_out[56]), .B0_f (new_AGEMA_signal_3804), .B1_t (new_AGEMA_signal_3805), .B1_f (new_AGEMA_signal_3806), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_56_U1_X), .Z0_f (new_AGEMA_signal_5973), .Z1_t (new_AGEMA_signal_5974), .Z1_f (new_AGEMA_signal_5975) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_56_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n22), .A1_f (new_AGEMA_signal_2479), .B0_t (LED_128_Instance_MUX_state0_mux_inst_56_U1_X), .B0_f (new_AGEMA_signal_5973), .B1_t (new_AGEMA_signal_5974), .B1_f (new_AGEMA_signal_5975), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_56_U1_Y), .Z0_f (new_AGEMA_signal_6141), .Z1_t (new_AGEMA_signal_6142), .Z1_f (new_AGEMA_signal_6143) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_56_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_56_U1_Y), .A0_f (new_AGEMA_signal_6141), .A1_t (new_AGEMA_signal_6142), .A1_f (new_AGEMA_signal_6143), .B0_t (LED_128_Instance_mixcolumns_out[56]), .B0_f (new_AGEMA_signal_5832), .B1_t (new_AGEMA_signal_5833), .B1_f (new_AGEMA_signal_5834), .Z0_t (LED_128_Instance_state0[56]), .Z0_f (new_AGEMA_signal_6330), .Z1_t (new_AGEMA_signal_6331), .Z1_f (new_AGEMA_signal_6332) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_57_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[57]), .A0_f (new_AGEMA_signal_5829), .A1_t (new_AGEMA_signal_5830), .A1_f (new_AGEMA_signal_5831), .B0_t (LED_128_Instance_addconst_out[57]), .B0_f (new_AGEMA_signal_3807), .B1_t (new_AGEMA_signal_3808), .B1_f (new_AGEMA_signal_3809), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_57_U1_X), .Z0_f (new_AGEMA_signal_5976), .Z1_t (new_AGEMA_signal_5977), .Z1_f (new_AGEMA_signal_5978) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_57_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n22), .A1_f (new_AGEMA_signal_2479), .B0_t (LED_128_Instance_MUX_state0_mux_inst_57_U1_X), .B0_f (new_AGEMA_signal_5976), .B1_t (new_AGEMA_signal_5977), .B1_f (new_AGEMA_signal_5978), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_57_U1_Y), .Z0_f (new_AGEMA_signal_6144), .Z1_t (new_AGEMA_signal_6145), .Z1_f (new_AGEMA_signal_6146) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_57_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_57_U1_Y), .A0_f (new_AGEMA_signal_6144), .A1_t (new_AGEMA_signal_6145), .A1_f (new_AGEMA_signal_6146), .B0_t (LED_128_Instance_mixcolumns_out[57]), .B0_f (new_AGEMA_signal_5829), .B1_t (new_AGEMA_signal_5830), .B1_f (new_AGEMA_signal_5831), .Z0_t (LED_128_Instance_state0[57]), .Z0_f (new_AGEMA_signal_6333), .Z1_t (new_AGEMA_signal_6334), .Z1_f (new_AGEMA_signal_6335) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_58_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[58]), .A0_f (new_AGEMA_signal_5616), .A1_t (new_AGEMA_signal_5617), .A1_f (new_AGEMA_signal_5618), .B0_t (LED_128_Instance_addconst_out[58]), .B0_f (new_AGEMA_signal_3810), .B1_t (new_AGEMA_signal_3811), .B1_f (new_AGEMA_signal_3812), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_58_U1_X), .Z0_f (new_AGEMA_signal_5778), .Z1_t (new_AGEMA_signal_5779), .Z1_f (new_AGEMA_signal_5780) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_58_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n22), .A1_f (new_AGEMA_signal_2479), .B0_t (LED_128_Instance_MUX_state0_mux_inst_58_U1_X), .B0_f (new_AGEMA_signal_5778), .B1_t (new_AGEMA_signal_5779), .B1_f (new_AGEMA_signal_5780), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_58_U1_Y), .Z0_f (new_AGEMA_signal_5979), .Z1_t (new_AGEMA_signal_5980), .Z1_f (new_AGEMA_signal_5981) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_58_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_58_U1_Y), .A0_f (new_AGEMA_signal_5979), .A1_t (new_AGEMA_signal_5980), .A1_f (new_AGEMA_signal_5981), .B0_t (LED_128_Instance_mixcolumns_out[58]), .B0_f (new_AGEMA_signal_5616), .B1_t (new_AGEMA_signal_5617), .B1_f (new_AGEMA_signal_5618), .Z0_t (LED_128_Instance_state0[58]), .Z0_f (new_AGEMA_signal_6147), .Z1_t (new_AGEMA_signal_6148), .Z1_f (new_AGEMA_signal_6149) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_59_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[59]), .A0_f (new_AGEMA_signal_5406), .A1_t (new_AGEMA_signal_5407), .A1_f (new_AGEMA_signal_5408), .B0_t (LED_128_Instance_addconst_out[59]), .B0_f (new_AGEMA_signal_3813), .B1_t (new_AGEMA_signal_3814), .B1_f (new_AGEMA_signal_3815), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_59_U1_X), .Z0_f (new_AGEMA_signal_5547), .Z1_t (new_AGEMA_signal_5548), .Z1_f (new_AGEMA_signal_5549) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_59_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n22), .A1_f (new_AGEMA_signal_2479), .B0_t (LED_128_Instance_MUX_state0_mux_inst_59_U1_X), .B0_f (new_AGEMA_signal_5547), .B1_t (new_AGEMA_signal_5548), .B1_f (new_AGEMA_signal_5549), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_59_U1_Y), .Z0_f (new_AGEMA_signal_5781), .Z1_t (new_AGEMA_signal_5782), .Z1_f (new_AGEMA_signal_5783) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_59_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_59_U1_Y), .A0_f (new_AGEMA_signal_5781), .A1_t (new_AGEMA_signal_5782), .A1_f (new_AGEMA_signal_5783), .B0_t (LED_128_Instance_mixcolumns_out[59]), .B0_f (new_AGEMA_signal_5406), .B1_t (new_AGEMA_signal_5407), .B1_f (new_AGEMA_signal_5408), .Z0_t (LED_128_Instance_state0[59]), .Z0_f (new_AGEMA_signal_5982), .Z1_t (new_AGEMA_signal_5983), .Z1_f (new_AGEMA_signal_5984) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_60_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[60]), .A0_f (new_AGEMA_signal_5640), .A1_t (new_AGEMA_signal_5641), .A1_f (new_AGEMA_signal_5642), .B0_t (LED_128_Instance_addconst_out[60]), .B0_f (new_AGEMA_signal_3816), .B1_t (new_AGEMA_signal_3817), .B1_f (new_AGEMA_signal_3818), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_60_U1_X), .Z0_f (new_AGEMA_signal_5784), .Z1_t (new_AGEMA_signal_5785), .Z1_f (new_AGEMA_signal_5786) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_60_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n22), .A1_f (new_AGEMA_signal_2479), .B0_t (LED_128_Instance_MUX_state0_mux_inst_60_U1_X), .B0_f (new_AGEMA_signal_5784), .B1_t (new_AGEMA_signal_5785), .B1_f (new_AGEMA_signal_5786), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_60_U1_Y), .Z0_f (new_AGEMA_signal_5985), .Z1_t (new_AGEMA_signal_5986), .Z1_f (new_AGEMA_signal_5987) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_60_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_60_U1_Y), .A0_f (new_AGEMA_signal_5985), .A1_t (new_AGEMA_signal_5986), .A1_f (new_AGEMA_signal_5987), .B0_t (LED_128_Instance_mixcolumns_out[60]), .B0_f (new_AGEMA_signal_5640), .B1_t (new_AGEMA_signal_5641), .B1_f (new_AGEMA_signal_5642), .Z0_t (LED_128_Instance_state0[60]), .Z0_f (new_AGEMA_signal_6150), .Z1_t (new_AGEMA_signal_6151), .Z1_f (new_AGEMA_signal_6152) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_61_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[61]), .A0_f (new_AGEMA_signal_5637), .A1_t (new_AGEMA_signal_5638), .A1_f (new_AGEMA_signal_5639), .B0_t (LED_128_Instance_addconst_out[61]), .B0_f (new_AGEMA_signal_3819), .B1_t (new_AGEMA_signal_3820), .B1_f (new_AGEMA_signal_3821), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_61_U1_X), .Z0_f (new_AGEMA_signal_5787), .Z1_t (new_AGEMA_signal_5788), .Z1_f (new_AGEMA_signal_5789) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_61_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n22), .A1_f (new_AGEMA_signal_2479), .B0_t (LED_128_Instance_MUX_state0_mux_inst_61_U1_X), .B0_f (new_AGEMA_signal_5787), .B1_t (new_AGEMA_signal_5788), .B1_f (new_AGEMA_signal_5789), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_61_U1_Y), .Z0_f (new_AGEMA_signal_5988), .Z1_t (new_AGEMA_signal_5989), .Z1_f (new_AGEMA_signal_5990) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_61_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_61_U1_Y), .A0_f (new_AGEMA_signal_5988), .A1_t (new_AGEMA_signal_5989), .A1_f (new_AGEMA_signal_5990), .B0_t (LED_128_Instance_mixcolumns_out[61]), .B0_f (new_AGEMA_signal_5637), .B1_t (new_AGEMA_signal_5638), .B1_f (new_AGEMA_signal_5639), .Z0_t (LED_128_Instance_state0[61]), .Z0_f (new_AGEMA_signal_6153), .Z1_t (new_AGEMA_signal_6154), .Z1_f (new_AGEMA_signal_6155) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_62_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[62]), .A0_f (new_AGEMA_signal_5451), .A1_t (new_AGEMA_signal_5452), .A1_f (new_AGEMA_signal_5453), .B0_t (LED_128_Instance_addconst_out[62]), .B0_f (new_AGEMA_signal_3822), .B1_t (new_AGEMA_signal_3823), .B1_f (new_AGEMA_signal_3824), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_62_U1_X), .Z0_f (new_AGEMA_signal_5550), .Z1_t (new_AGEMA_signal_5551), .Z1_f (new_AGEMA_signal_5552) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_62_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n22), .A1_f (new_AGEMA_signal_2479), .B0_t (LED_128_Instance_MUX_state0_mux_inst_62_U1_X), .B0_f (new_AGEMA_signal_5550), .B1_t (new_AGEMA_signal_5551), .B1_f (new_AGEMA_signal_5552), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_62_U1_Y), .Z0_f (new_AGEMA_signal_5790), .Z1_t (new_AGEMA_signal_5791), .Z1_f (new_AGEMA_signal_5792) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_62_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_62_U1_Y), .A0_f (new_AGEMA_signal_5790), .A1_t (new_AGEMA_signal_5791), .A1_f (new_AGEMA_signal_5792), .B0_t (LED_128_Instance_mixcolumns_out[62]), .B0_f (new_AGEMA_signal_5451), .B1_t (new_AGEMA_signal_5452), .B1_f (new_AGEMA_signal_5453), .Z0_t (LED_128_Instance_state0[62]), .Z0_f (new_AGEMA_signal_5991), .Z1_t (new_AGEMA_signal_5992), .Z1_f (new_AGEMA_signal_5993) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_63_U1_XOR1_U1 ( .A0_t (LED_128_Instance_mixcolumns_out[63]), .A0_f (new_AGEMA_signal_5436), .A1_t (new_AGEMA_signal_5437), .A1_f (new_AGEMA_signal_5438), .B0_t (LED_128_Instance_addconst_out[63]), .B0_f (new_AGEMA_signal_3825), .B1_t (new_AGEMA_signal_3826), .B1_f (new_AGEMA_signal_3827), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_63_U1_X), .Z0_f (new_AGEMA_signal_5553), .Z1_t (new_AGEMA_signal_5554), .Z1_f (new_AGEMA_signal_5555) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_63_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n22), .A1_f (new_AGEMA_signal_2479), .B0_t (LED_128_Instance_MUX_state0_mux_inst_63_U1_X), .B0_f (new_AGEMA_signal_5553), .B1_t (new_AGEMA_signal_5554), .B1_f (new_AGEMA_signal_5555), .Z0_t (LED_128_Instance_MUX_state0_mux_inst_63_U1_Y), .Z0_f (new_AGEMA_signal_5793), .Z1_t (new_AGEMA_signal_5794), .Z1_f (new_AGEMA_signal_5795) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state0_mux_inst_63_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state0_mux_inst_63_U1_Y), .A0_f (new_AGEMA_signal_5793), .A1_t (new_AGEMA_signal_5794), .A1_f (new_AGEMA_signal_5795), .B0_t (LED_128_Instance_mixcolumns_out[63]), .B0_f (new_AGEMA_signal_5436), .B1_t (new_AGEMA_signal_5437), .B1_f (new_AGEMA_signal_5438), .Z0_t (LED_128_Instance_state0[63]), .Z0_f (new_AGEMA_signal_5994), .Z1_t (new_AGEMA_signal_5995), .Z1_f (new_AGEMA_signal_5996) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_0_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[0]), .A0_f (new_AGEMA_signal_5454), .A1_t (new_AGEMA_signal_5455), .A1_f (new_AGEMA_signal_5456), .B0_t (IN_plaintext_s0_t[0]), .B0_f (IN_plaintext_s0_f[0]), .B1_t (IN_plaintext_s1_t[0]), .B1_f (IN_plaintext_s1_f[0]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_0_U1_X), .Z0_f (new_AGEMA_signal_5799), .Z1_t (new_AGEMA_signal_5800), .Z1_f (new_AGEMA_signal_5801) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_0_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (IN_reset_t), .A1_f (IN_reset_f), .B0_t (LED_128_Instance_MUX_state1_mux_inst_0_U1_X), .B0_f (new_AGEMA_signal_5799), .B1_t (new_AGEMA_signal_5800), .B1_f (new_AGEMA_signal_5801), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_0_U1_Y), .Z0_f (new_AGEMA_signal_5997), .Z1_t (new_AGEMA_signal_5998), .Z1_f (new_AGEMA_signal_5999) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_0_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_0_U1_Y), .A0_f (new_AGEMA_signal_5997), .A1_t (new_AGEMA_signal_5998), .A1_f (new_AGEMA_signal_5999), .B0_t (LED_128_Instance_state0[0]), .B0_f (new_AGEMA_signal_5454), .B1_t (new_AGEMA_signal_5455), .B1_f (new_AGEMA_signal_5456), .Z0_t (OUT_ciphertext_s0_t[0]), .Z0_f (OUT_ciphertext_s0_f[0]), .Z1_t (OUT_ciphertext_s1_t[0]), .Z1_f (OUT_ciphertext_s1_f[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_1_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[1]), .A0_f (new_AGEMA_signal_5847), .A1_t (new_AGEMA_signal_5848), .A1_f (new_AGEMA_signal_5849), .B0_t (IN_plaintext_s0_t[1]), .B0_f (IN_plaintext_s0_f[1]), .B1_t (IN_plaintext_s1_t[1]), .B1_f (IN_plaintext_s1_f[1]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_1_U1_X), .Z0_f (new_AGEMA_signal_6159), .Z1_t (new_AGEMA_signal_6160), .Z1_f (new_AGEMA_signal_6161) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_1_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (IN_reset_t), .A1_f (IN_reset_f), .B0_t (LED_128_Instance_MUX_state1_mux_inst_1_U1_X), .B0_f (new_AGEMA_signal_6159), .B1_t (new_AGEMA_signal_6160), .B1_f (new_AGEMA_signal_6161), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_1_U1_Y), .Z0_f (new_AGEMA_signal_6336), .Z1_t (new_AGEMA_signal_6337), .Z1_f (new_AGEMA_signal_6338) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_1_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_1_U1_Y), .A0_f (new_AGEMA_signal_6336), .A1_t (new_AGEMA_signal_6337), .A1_f (new_AGEMA_signal_6338), .B0_t (LED_128_Instance_state0[1]), .B0_f (new_AGEMA_signal_5847), .B1_t (new_AGEMA_signal_5848), .B1_f (new_AGEMA_signal_5849), .Z0_t (OUT_ciphertext_s0_t[1]), .Z0_f (OUT_ciphertext_s0_f[1]), .Z1_t (OUT_ciphertext_s1_t[1]), .Z1_f (OUT_ciphertext_s1_f[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_2_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[2]), .A0_f (new_AGEMA_signal_5460), .A1_t (new_AGEMA_signal_5461), .A1_f (new_AGEMA_signal_5462), .B0_t (IN_plaintext_s0_t[2]), .B0_f (IN_plaintext_s0_f[2]), .B1_t (IN_plaintext_s1_t[2]), .B1_f (IN_plaintext_s1_f[2]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_2_U1_X), .Z0_f (new_AGEMA_signal_5805), .Z1_t (new_AGEMA_signal_5806), .Z1_f (new_AGEMA_signal_5807) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_2_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (IN_reset_t), .A1_f (IN_reset_f), .B0_t (LED_128_Instance_MUX_state1_mux_inst_2_U1_X), .B0_f (new_AGEMA_signal_5805), .B1_t (new_AGEMA_signal_5806), .B1_f (new_AGEMA_signal_5807), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_2_U1_Y), .Z0_f (new_AGEMA_signal_6000), .Z1_t (new_AGEMA_signal_6001), .Z1_f (new_AGEMA_signal_6002) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_2_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_2_U1_Y), .A0_f (new_AGEMA_signal_6000), .A1_t (new_AGEMA_signal_6001), .A1_f (new_AGEMA_signal_6002), .B0_t (LED_128_Instance_state0[2]), .B0_f (new_AGEMA_signal_5460), .B1_t (new_AGEMA_signal_5461), .B1_f (new_AGEMA_signal_5462), .Z0_t (OUT_ciphertext_s0_t[2]), .Z0_f (OUT_ciphertext_s0_f[2]), .Z1_t (OUT_ciphertext_s1_t[2]), .Z1_f (OUT_ciphertext_s1_f[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_3_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[3]), .A0_f (new_AGEMA_signal_5850), .A1_t (new_AGEMA_signal_5851), .A1_f (new_AGEMA_signal_5852), .B0_t (IN_plaintext_s0_t[3]), .B0_f (IN_plaintext_s0_f[3]), .B1_t (IN_plaintext_s1_t[3]), .B1_f (IN_plaintext_s1_f[3]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_3_U1_X), .Z0_f (new_AGEMA_signal_6165), .Z1_t (new_AGEMA_signal_6166), .Z1_f (new_AGEMA_signal_6167) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_3_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (IN_reset_t), .A1_f (IN_reset_f), .B0_t (LED_128_Instance_MUX_state1_mux_inst_3_U1_X), .B0_f (new_AGEMA_signal_6165), .B1_t (new_AGEMA_signal_6166), .B1_f (new_AGEMA_signal_6167), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_3_U1_Y), .Z0_f (new_AGEMA_signal_6339), .Z1_t (new_AGEMA_signal_6340), .Z1_f (new_AGEMA_signal_6341) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_3_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_3_U1_Y), .A0_f (new_AGEMA_signal_6339), .A1_t (new_AGEMA_signal_6340), .A1_f (new_AGEMA_signal_6341), .B0_t (LED_128_Instance_state0[3]), .B0_f (new_AGEMA_signal_5850), .B1_t (new_AGEMA_signal_5851), .B1_f (new_AGEMA_signal_5852), .Z0_t (OUT_ciphertext_s0_t[3]), .Z0_f (OUT_ciphertext_s0_f[3]), .Z1_t (OUT_ciphertext_s1_t[3]), .Z1_f (OUT_ciphertext_s1_f[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_4_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[4]), .A0_f (new_AGEMA_signal_5649), .A1_t (new_AGEMA_signal_5650), .A1_f (new_AGEMA_signal_5651), .B0_t (IN_plaintext_s0_t[4]), .B0_f (IN_plaintext_s0_f[4]), .B1_t (IN_plaintext_s1_t[4]), .B1_f (IN_plaintext_s1_f[4]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_4_U1_X), .Z0_f (new_AGEMA_signal_6006), .Z1_t (new_AGEMA_signal_6007), .Z1_f (new_AGEMA_signal_6008) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_4_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (IN_reset_t), .A1_f (IN_reset_f), .B0_t (LED_128_Instance_MUX_state1_mux_inst_4_U1_X), .B0_f (new_AGEMA_signal_6006), .B1_t (new_AGEMA_signal_6007), .B1_f (new_AGEMA_signal_6008), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_4_U1_Y), .Z0_f (new_AGEMA_signal_6168), .Z1_t (new_AGEMA_signal_6169), .Z1_f (new_AGEMA_signal_6170) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_4_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_4_U1_Y), .A0_f (new_AGEMA_signal_6168), .A1_t (new_AGEMA_signal_6169), .A1_f (new_AGEMA_signal_6170), .B0_t (LED_128_Instance_state0[4]), .B0_f (new_AGEMA_signal_5649), .B1_t (new_AGEMA_signal_5650), .B1_f (new_AGEMA_signal_5651), .Z0_t (OUT_ciphertext_s0_t[4]), .Z0_f (OUT_ciphertext_s0_f[4]), .Z1_t (OUT_ciphertext_s1_t[4]), .Z1_f (OUT_ciphertext_s1_f[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_5_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[5]), .A0_f (new_AGEMA_signal_5853), .A1_t (new_AGEMA_signal_5854), .A1_f (new_AGEMA_signal_5855), .B0_t (IN_plaintext_s0_t[5]), .B0_f (IN_plaintext_s0_f[5]), .B1_t (IN_plaintext_s1_t[5]), .B1_f (IN_plaintext_s1_f[5]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_5_U1_X), .Z0_f (new_AGEMA_signal_6174), .Z1_t (new_AGEMA_signal_6175), .Z1_f (new_AGEMA_signal_6176) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_5_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (IN_reset_t), .A1_f (IN_reset_f), .B0_t (LED_128_Instance_MUX_state1_mux_inst_5_U1_X), .B0_f (new_AGEMA_signal_6174), .B1_t (new_AGEMA_signal_6175), .B1_f (new_AGEMA_signal_6176), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_5_U1_Y), .Z0_f (new_AGEMA_signal_6342), .Z1_t (new_AGEMA_signal_6343), .Z1_f (new_AGEMA_signal_6344) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_5_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_5_U1_Y), .A0_f (new_AGEMA_signal_6342), .A1_t (new_AGEMA_signal_6343), .A1_f (new_AGEMA_signal_6344), .B0_t (LED_128_Instance_state0[5]), .B0_f (new_AGEMA_signal_5853), .B1_t (new_AGEMA_signal_5854), .B1_f (new_AGEMA_signal_5855), .Z0_t (OUT_ciphertext_s0_t[5]), .Z0_f (OUT_ciphertext_s0_f[5]), .Z1_t (OUT_ciphertext_s1_t[5]), .Z1_f (OUT_ciphertext_s1_f[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_6_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[6]), .A0_f (new_AGEMA_signal_5655), .A1_t (new_AGEMA_signal_5656), .A1_f (new_AGEMA_signal_5657), .B0_t (IN_plaintext_s0_t[6]), .B0_f (IN_plaintext_s0_f[6]), .B1_t (IN_plaintext_s1_t[6]), .B1_f (IN_plaintext_s1_f[6]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_6_U1_X), .Z0_f (new_AGEMA_signal_6012), .Z1_t (new_AGEMA_signal_6013), .Z1_f (new_AGEMA_signal_6014) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_6_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (IN_reset_t), .A1_f (IN_reset_f), .B0_t (LED_128_Instance_MUX_state1_mux_inst_6_U1_X), .B0_f (new_AGEMA_signal_6012), .B1_t (new_AGEMA_signal_6013), .B1_f (new_AGEMA_signal_6014), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_6_U1_Y), .Z0_f (new_AGEMA_signal_6177), .Z1_t (new_AGEMA_signal_6178), .Z1_f (new_AGEMA_signal_6179) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_6_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_6_U1_Y), .A0_f (new_AGEMA_signal_6177), .A1_t (new_AGEMA_signal_6178), .A1_f (new_AGEMA_signal_6179), .B0_t (LED_128_Instance_state0[6]), .B0_f (new_AGEMA_signal_5655), .B1_t (new_AGEMA_signal_5656), .B1_f (new_AGEMA_signal_5657), .Z0_t (OUT_ciphertext_s0_t[6]), .Z0_f (OUT_ciphertext_s0_f[6]), .Z1_t (OUT_ciphertext_s1_t[6]), .Z1_f (OUT_ciphertext_s1_f[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_7_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[7]), .A0_f (new_AGEMA_signal_5658), .A1_t (new_AGEMA_signal_5659), .A1_f (new_AGEMA_signal_5660), .B0_t (IN_plaintext_s0_t[7]), .B0_f (IN_plaintext_s0_f[7]), .B1_t (IN_plaintext_s1_t[7]), .B1_f (IN_plaintext_s1_f[7]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_7_U1_X), .Z0_f (new_AGEMA_signal_6018), .Z1_t (new_AGEMA_signal_6019), .Z1_f (new_AGEMA_signal_6020) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_7_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (IN_reset_t), .A1_f (IN_reset_f), .B0_t (LED_128_Instance_MUX_state1_mux_inst_7_U1_X), .B0_f (new_AGEMA_signal_6018), .B1_t (new_AGEMA_signal_6019), .B1_f (new_AGEMA_signal_6020), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_7_U1_Y), .Z0_f (new_AGEMA_signal_6180), .Z1_t (new_AGEMA_signal_6181), .Z1_f (new_AGEMA_signal_6182) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_7_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_7_U1_Y), .A0_f (new_AGEMA_signal_6180), .A1_t (new_AGEMA_signal_6181), .A1_f (new_AGEMA_signal_6182), .B0_t (LED_128_Instance_state0[7]), .B0_f (new_AGEMA_signal_5658), .B1_t (new_AGEMA_signal_5659), .B1_f (new_AGEMA_signal_5660), .Z0_t (OUT_ciphertext_s0_t[7]), .Z0_f (OUT_ciphertext_s0_f[7]), .Z1_t (OUT_ciphertext_s1_t[7]), .Z1_f (OUT_ciphertext_s1_f[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_8_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[8]), .A0_f (new_AGEMA_signal_5478), .A1_t (new_AGEMA_signal_5479), .A1_f (new_AGEMA_signal_5480), .B0_t (IN_plaintext_s0_t[8]), .B0_f (IN_plaintext_s0_f[8]), .B1_t (IN_plaintext_s1_t[8]), .B1_f (IN_plaintext_s1_f[8]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_8_U1_X), .Z0_f (new_AGEMA_signal_5811), .Z1_t (new_AGEMA_signal_5812), .Z1_f (new_AGEMA_signal_5813) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_8_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (IN_reset_t), .A1_f (IN_reset_f), .B0_t (LED_128_Instance_MUX_state1_mux_inst_8_U1_X), .B0_f (new_AGEMA_signal_5811), .B1_t (new_AGEMA_signal_5812), .B1_f (new_AGEMA_signal_5813), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_8_U1_Y), .Z0_f (new_AGEMA_signal_6021), .Z1_t (new_AGEMA_signal_6022), .Z1_f (new_AGEMA_signal_6023) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_8_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_8_U1_Y), .A0_f (new_AGEMA_signal_6021), .A1_t (new_AGEMA_signal_6022), .A1_f (new_AGEMA_signal_6023), .B0_t (LED_128_Instance_state0[8]), .B0_f (new_AGEMA_signal_5478), .B1_t (new_AGEMA_signal_5479), .B1_f (new_AGEMA_signal_5480), .Z0_t (OUT_ciphertext_s0_t[8]), .Z0_f (OUT_ciphertext_s0_f[8]), .Z1_t (OUT_ciphertext_s1_t[8]), .Z1_f (OUT_ciphertext_s1_f[8]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_9_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[9]), .A0_f (new_AGEMA_signal_5856), .A1_t (new_AGEMA_signal_5857), .A1_f (new_AGEMA_signal_5858), .B0_t (IN_plaintext_s0_t[9]), .B0_f (IN_plaintext_s0_f[9]), .B1_t (IN_plaintext_s1_t[9]), .B1_f (IN_plaintext_s1_f[9]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_9_U1_X), .Z0_f (new_AGEMA_signal_6186), .Z1_t (new_AGEMA_signal_6187), .Z1_f (new_AGEMA_signal_6188) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_9_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (IN_reset_t), .A1_f (IN_reset_f), .B0_t (LED_128_Instance_MUX_state1_mux_inst_9_U1_X), .B0_f (new_AGEMA_signal_6186), .B1_t (new_AGEMA_signal_6187), .B1_f (new_AGEMA_signal_6188), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_9_U1_Y), .Z0_f (new_AGEMA_signal_6345), .Z1_t (new_AGEMA_signal_6346), .Z1_f (new_AGEMA_signal_6347) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_9_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_9_U1_Y), .A0_f (new_AGEMA_signal_6345), .A1_t (new_AGEMA_signal_6346), .A1_f (new_AGEMA_signal_6347), .B0_t (LED_128_Instance_state0[9]), .B0_f (new_AGEMA_signal_5856), .B1_t (new_AGEMA_signal_5857), .B1_f (new_AGEMA_signal_5858), .Z0_t (OUT_ciphertext_s0_t[9]), .Z0_f (OUT_ciphertext_s0_f[9]), .Z1_t (OUT_ciphertext_s1_t[9]), .Z1_f (OUT_ciphertext_s1_f[9]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_10_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[10]), .A0_f (new_AGEMA_signal_5664), .A1_t (new_AGEMA_signal_5665), .A1_f (new_AGEMA_signal_5666), .B0_t (IN_plaintext_s0_t[10]), .B0_f (IN_plaintext_s0_f[10]), .B1_t (IN_plaintext_s1_t[10]), .B1_f (IN_plaintext_s1_f[10]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_10_U1_X), .Z0_f (new_AGEMA_signal_6027), .Z1_t (new_AGEMA_signal_6028), .Z1_f (new_AGEMA_signal_6029) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_10_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (IN_reset_t), .A1_f (IN_reset_f), .B0_t (LED_128_Instance_MUX_state1_mux_inst_10_U1_X), .B0_f (new_AGEMA_signal_6027), .B1_t (new_AGEMA_signal_6028), .B1_f (new_AGEMA_signal_6029), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_10_U1_Y), .Z0_f (new_AGEMA_signal_6189), .Z1_t (new_AGEMA_signal_6190), .Z1_f (new_AGEMA_signal_6191) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_10_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_10_U1_Y), .A0_f (new_AGEMA_signal_6189), .A1_t (new_AGEMA_signal_6190), .A1_f (new_AGEMA_signal_6191), .B0_t (LED_128_Instance_state0[10]), .B0_f (new_AGEMA_signal_5664), .B1_t (new_AGEMA_signal_5665), .B1_f (new_AGEMA_signal_5666), .Z0_t (OUT_ciphertext_s0_t[10]), .Z0_f (OUT_ciphertext_s0_f[10]), .Z1_t (OUT_ciphertext_s1_t[10]), .Z1_f (OUT_ciphertext_s1_f[10]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_11_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[11]), .A0_f (new_AGEMA_signal_5667), .A1_t (new_AGEMA_signal_5668), .A1_f (new_AGEMA_signal_5669), .B0_t (IN_plaintext_s0_t[11]), .B0_f (IN_plaintext_s0_f[11]), .B1_t (IN_plaintext_s1_t[11]), .B1_f (IN_plaintext_s1_f[11]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_11_U1_X), .Z0_f (new_AGEMA_signal_6033), .Z1_t (new_AGEMA_signal_6034), .Z1_f (new_AGEMA_signal_6035) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_11_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (IN_reset_t), .A1_f (IN_reset_f), .B0_t (LED_128_Instance_MUX_state1_mux_inst_11_U1_X), .B0_f (new_AGEMA_signal_6033), .B1_t (new_AGEMA_signal_6034), .B1_f (new_AGEMA_signal_6035), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_11_U1_Y), .Z0_f (new_AGEMA_signal_6192), .Z1_t (new_AGEMA_signal_6193), .Z1_f (new_AGEMA_signal_6194) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_11_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_11_U1_Y), .A0_f (new_AGEMA_signal_6192), .A1_t (new_AGEMA_signal_6193), .A1_f (new_AGEMA_signal_6194), .B0_t (LED_128_Instance_state0[11]), .B0_f (new_AGEMA_signal_5667), .B1_t (new_AGEMA_signal_5668), .B1_f (new_AGEMA_signal_5669), .Z0_t (OUT_ciphertext_s0_t[11]), .Z0_f (OUT_ciphertext_s0_f[11]), .Z1_t (OUT_ciphertext_s1_t[11]), .Z1_f (OUT_ciphertext_s1_f[11]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_12_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[12]), .A0_f (new_AGEMA_signal_5670), .A1_t (new_AGEMA_signal_5671), .A1_f (new_AGEMA_signal_5672), .B0_t (IN_plaintext_s0_t[12]), .B0_f (IN_plaintext_s0_f[12]), .B1_t (IN_plaintext_s1_t[12]), .B1_f (IN_plaintext_s1_f[12]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_12_U1_X), .Z0_f (new_AGEMA_signal_6039), .Z1_t (new_AGEMA_signal_6040), .Z1_f (new_AGEMA_signal_6041) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_12_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (IN_reset_t), .A1_f (IN_reset_f), .B0_t (LED_128_Instance_MUX_state1_mux_inst_12_U1_X), .B0_f (new_AGEMA_signal_6039), .B1_t (new_AGEMA_signal_6040), .B1_f (new_AGEMA_signal_6041), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_12_U1_Y), .Z0_f (new_AGEMA_signal_6195), .Z1_t (new_AGEMA_signal_6196), .Z1_f (new_AGEMA_signal_6197) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_12_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_12_U1_Y), .A0_f (new_AGEMA_signal_6195), .A1_t (new_AGEMA_signal_6196), .A1_f (new_AGEMA_signal_6197), .B0_t (LED_128_Instance_state0[12]), .B0_f (new_AGEMA_signal_5670), .B1_t (new_AGEMA_signal_5671), .B1_f (new_AGEMA_signal_5672), .Z0_t (OUT_ciphertext_s0_t[12]), .Z0_f (OUT_ciphertext_s0_f[12]), .Z1_t (OUT_ciphertext_s1_t[12]), .Z1_f (OUT_ciphertext_s1_f[12]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_13_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[13]), .A0_f (new_AGEMA_signal_6066), .A1_t (new_AGEMA_signal_6067), .A1_f (new_AGEMA_signal_6068), .B0_t (IN_plaintext_s0_t[13]), .B0_f (IN_plaintext_s0_f[13]), .B1_t (IN_plaintext_s1_t[13]), .B1_f (IN_plaintext_s1_f[13]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_13_U1_X), .Z0_f (new_AGEMA_signal_6351), .Z1_t (new_AGEMA_signal_6352), .Z1_f (new_AGEMA_signal_6353) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_13_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (IN_reset_t), .A1_f (IN_reset_f), .B0_t (LED_128_Instance_MUX_state1_mux_inst_13_U1_X), .B0_f (new_AGEMA_signal_6351), .B1_t (new_AGEMA_signal_6352), .B1_f (new_AGEMA_signal_6353), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_13_U1_Y), .Z0_f (new_AGEMA_signal_6528), .Z1_t (new_AGEMA_signal_6529), .Z1_f (new_AGEMA_signal_6530) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_13_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_13_U1_Y), .A0_f (new_AGEMA_signal_6528), .A1_t (new_AGEMA_signal_6529), .A1_f (new_AGEMA_signal_6530), .B0_t (LED_128_Instance_state0[13]), .B0_f (new_AGEMA_signal_6066), .B1_t (new_AGEMA_signal_6067), .B1_f (new_AGEMA_signal_6068), .Z0_t (OUT_ciphertext_s0_t[13]), .Z0_f (OUT_ciphertext_s0_f[13]), .Z1_t (OUT_ciphertext_s1_t[13]), .Z1_f (OUT_ciphertext_s1_f[13]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_14_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[14]), .A0_f (new_AGEMA_signal_5493), .A1_t (new_AGEMA_signal_5494), .A1_f (new_AGEMA_signal_5495), .B0_t (IN_plaintext_s0_t[14]), .B0_f (IN_plaintext_s0_f[14]), .B1_t (IN_plaintext_s1_t[14]), .B1_f (IN_plaintext_s1_f[14]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_14_U1_X), .Z0_f (new_AGEMA_signal_5817), .Z1_t (new_AGEMA_signal_5818), .Z1_f (new_AGEMA_signal_5819) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_14_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (IN_reset_t), .A1_f (IN_reset_f), .B0_t (LED_128_Instance_MUX_state1_mux_inst_14_U1_X), .B0_f (new_AGEMA_signal_5817), .B1_t (new_AGEMA_signal_5818), .B1_f (new_AGEMA_signal_5819), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_14_U1_Y), .Z0_f (new_AGEMA_signal_6042), .Z1_t (new_AGEMA_signal_6043), .Z1_f (new_AGEMA_signal_6044) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_14_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_14_U1_Y), .A0_f (new_AGEMA_signal_6042), .A1_t (new_AGEMA_signal_6043), .A1_f (new_AGEMA_signal_6044), .B0_t (LED_128_Instance_state0[14]), .B0_f (new_AGEMA_signal_5493), .B1_t (new_AGEMA_signal_5494), .B1_f (new_AGEMA_signal_5495), .Z0_t (OUT_ciphertext_s0_t[14]), .Z0_f (OUT_ciphertext_s0_f[14]), .Z1_t (OUT_ciphertext_s1_t[14]), .Z1_f (OUT_ciphertext_s1_f[14]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_15_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[15]), .A0_f (new_AGEMA_signal_5676), .A1_t (new_AGEMA_signal_5677), .A1_f (new_AGEMA_signal_5678), .B0_t (IN_plaintext_s0_t[15]), .B0_f (IN_plaintext_s0_f[15]), .B1_t (IN_plaintext_s1_t[15]), .B1_f (IN_plaintext_s1_f[15]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_15_U1_X), .Z0_f (new_AGEMA_signal_6048), .Z1_t (new_AGEMA_signal_6049), .Z1_f (new_AGEMA_signal_6050) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_15_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (IN_reset_t), .A1_f (IN_reset_f), .B0_t (LED_128_Instance_MUX_state1_mux_inst_15_U1_X), .B0_f (new_AGEMA_signal_6048), .B1_t (new_AGEMA_signal_6049), .B1_f (new_AGEMA_signal_6050), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_15_U1_Y), .Z0_f (new_AGEMA_signal_6198), .Z1_t (new_AGEMA_signal_6199), .Z1_f (new_AGEMA_signal_6200) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_15_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_15_U1_Y), .A0_f (new_AGEMA_signal_6198), .A1_t (new_AGEMA_signal_6199), .A1_f (new_AGEMA_signal_6200), .B0_t (LED_128_Instance_state0[15]), .B0_f (new_AGEMA_signal_5676), .B1_t (new_AGEMA_signal_5677), .B1_f (new_AGEMA_signal_5678), .Z0_t (OUT_ciphertext_s0_t[15]), .Z0_f (OUT_ciphertext_s0_f[15]), .Z1_t (OUT_ciphertext_s1_t[15]), .Z1_f (OUT_ciphertext_s1_f[15]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_16_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[16]), .A0_f (new_AGEMA_signal_6069), .A1_t (new_AGEMA_signal_6070), .A1_f (new_AGEMA_signal_6071), .B0_t (IN_plaintext_s0_t[16]), .B0_f (IN_plaintext_s0_f[16]), .B1_t (IN_plaintext_s1_t[16]), .B1_f (IN_plaintext_s1_f[16]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_16_U1_X), .Z0_f (new_AGEMA_signal_6357), .Z1_t (new_AGEMA_signal_6358), .Z1_f (new_AGEMA_signal_6359) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_16_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (IN_reset_t), .A1_f (IN_reset_f), .B0_t (LED_128_Instance_MUX_state1_mux_inst_16_U1_X), .B0_f (new_AGEMA_signal_6357), .B1_t (new_AGEMA_signal_6358), .B1_f (new_AGEMA_signal_6359), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_16_U1_Y), .Z0_f (new_AGEMA_signal_6531), .Z1_t (new_AGEMA_signal_6532), .Z1_f (new_AGEMA_signal_6533) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_16_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_16_U1_Y), .A0_f (new_AGEMA_signal_6531), .A1_t (new_AGEMA_signal_6532), .A1_f (new_AGEMA_signal_6533), .B0_t (LED_128_Instance_state0[16]), .B0_f (new_AGEMA_signal_6069), .B1_t (new_AGEMA_signal_6070), .B1_f (new_AGEMA_signal_6071), .Z0_t (OUT_ciphertext_s0_t[16]), .Z0_f (OUT_ciphertext_s0_f[16]), .Z1_t (OUT_ciphertext_s1_t[16]), .Z1_f (OUT_ciphertext_s1_f[16]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_17_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[17]), .A0_f (new_AGEMA_signal_5865), .A1_t (new_AGEMA_signal_5866), .A1_f (new_AGEMA_signal_5867), .B0_t (IN_plaintext_s0_t[17]), .B0_f (IN_plaintext_s0_f[17]), .B1_t (IN_plaintext_s1_t[17]), .B1_f (IN_plaintext_s1_f[17]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_17_U1_X), .Z0_f (new_AGEMA_signal_6204), .Z1_t (new_AGEMA_signal_6205), .Z1_f (new_AGEMA_signal_6206) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_17_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (IN_reset_t), .A1_f (IN_reset_f), .B0_t (LED_128_Instance_MUX_state1_mux_inst_17_U1_X), .B0_f (new_AGEMA_signal_6204), .B1_t (new_AGEMA_signal_6205), .B1_f (new_AGEMA_signal_6206), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_17_U1_Y), .Z0_f (new_AGEMA_signal_6360), .Z1_t (new_AGEMA_signal_6361), .Z1_f (new_AGEMA_signal_6362) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_17_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_17_U1_Y), .A0_f (new_AGEMA_signal_6360), .A1_t (new_AGEMA_signal_6361), .A1_f (new_AGEMA_signal_6362), .B0_t (LED_128_Instance_state0[17]), .B0_f (new_AGEMA_signal_5865), .B1_t (new_AGEMA_signal_5866), .B1_f (new_AGEMA_signal_5867), .Z0_t (OUT_ciphertext_s0_t[17]), .Z0_f (OUT_ciphertext_s0_f[17]), .Z1_t (OUT_ciphertext_s1_t[17]), .Z1_f (OUT_ciphertext_s1_f[17]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_18_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[18]), .A0_f (new_AGEMA_signal_6072), .A1_t (new_AGEMA_signal_6073), .A1_f (new_AGEMA_signal_6074), .B0_t (IN_plaintext_s0_t[18]), .B0_f (IN_plaintext_s0_f[18]), .B1_t (IN_plaintext_s1_t[18]), .B1_f (IN_plaintext_s1_f[18]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_18_U1_X), .Z0_f (new_AGEMA_signal_6366), .Z1_t (new_AGEMA_signal_6367), .Z1_f (new_AGEMA_signal_6368) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_18_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (IN_reset_t), .A1_f (IN_reset_f), .B0_t (LED_128_Instance_MUX_state1_mux_inst_18_U1_X), .B0_f (new_AGEMA_signal_6366), .B1_t (new_AGEMA_signal_6367), .B1_f (new_AGEMA_signal_6368), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_18_U1_Y), .Z0_f (new_AGEMA_signal_6534), .Z1_t (new_AGEMA_signal_6535), .Z1_f (new_AGEMA_signal_6536) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_18_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_18_U1_Y), .A0_f (new_AGEMA_signal_6534), .A1_t (new_AGEMA_signal_6535), .A1_f (new_AGEMA_signal_6536), .B0_t (LED_128_Instance_state0[18]), .B0_f (new_AGEMA_signal_6072), .B1_t (new_AGEMA_signal_6073), .B1_f (new_AGEMA_signal_6074), .Z0_t (OUT_ciphertext_s0_t[18]), .Z0_f (OUT_ciphertext_s0_f[18]), .Z1_t (OUT_ciphertext_s1_t[18]), .Z1_f (OUT_ciphertext_s1_f[18]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_19_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[19]), .A0_f (new_AGEMA_signal_6075), .A1_t (new_AGEMA_signal_6076), .A1_f (new_AGEMA_signal_6077), .B0_t (IN_plaintext_s0_t[19]), .B0_f (IN_plaintext_s0_f[19]), .B1_t (IN_plaintext_s1_t[19]), .B1_f (IN_plaintext_s1_f[19]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_19_U1_X), .Z0_f (new_AGEMA_signal_6372), .Z1_t (new_AGEMA_signal_6373), .Z1_f (new_AGEMA_signal_6374) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_19_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (IN_reset_t), .A1_f (IN_reset_f), .B0_t (LED_128_Instance_MUX_state1_mux_inst_19_U1_X), .B0_f (new_AGEMA_signal_6372), .B1_t (new_AGEMA_signal_6373), .B1_f (new_AGEMA_signal_6374), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_19_U1_Y), .Z0_f (new_AGEMA_signal_6537), .Z1_t (new_AGEMA_signal_6538), .Z1_f (new_AGEMA_signal_6539) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_19_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_19_U1_Y), .A0_f (new_AGEMA_signal_6537), .A1_t (new_AGEMA_signal_6538), .A1_f (new_AGEMA_signal_6539), .B0_t (LED_128_Instance_state0[19]), .B0_f (new_AGEMA_signal_6075), .B1_t (new_AGEMA_signal_6076), .B1_f (new_AGEMA_signal_6077), .Z0_t (OUT_ciphertext_s0_t[19]), .Z0_f (OUT_ciphertext_s0_f[19]), .Z1_t (OUT_ciphertext_s1_t[19]), .Z1_f (OUT_ciphertext_s1_f[19]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_20_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[20]), .A0_f (new_AGEMA_signal_5874), .A1_t (new_AGEMA_signal_5875), .A1_f (new_AGEMA_signal_5876), .B0_t (IN_plaintext_s0_t[20]), .B0_f (IN_plaintext_s0_f[20]), .B1_t (IN_plaintext_s1_t[20]), .B1_f (IN_plaintext_s1_f[20]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_20_U1_X), .Z0_f (new_AGEMA_signal_6210), .Z1_t (new_AGEMA_signal_6211), .Z1_f (new_AGEMA_signal_6212) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_20_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (IN_reset_t), .A1_f (IN_reset_f), .B0_t (LED_128_Instance_MUX_state1_mux_inst_20_U1_X), .B0_f (new_AGEMA_signal_6210), .B1_t (new_AGEMA_signal_6211), .B1_f (new_AGEMA_signal_6212), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_20_U1_Y), .Z0_f (new_AGEMA_signal_6375), .Z1_t (new_AGEMA_signal_6376), .Z1_f (new_AGEMA_signal_6377) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_20_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_20_U1_Y), .A0_f (new_AGEMA_signal_6375), .A1_t (new_AGEMA_signal_6376), .A1_f (new_AGEMA_signal_6377), .B0_t (LED_128_Instance_state0[20]), .B0_f (new_AGEMA_signal_5874), .B1_t (new_AGEMA_signal_5875), .B1_f (new_AGEMA_signal_5876), .Z0_t (OUT_ciphertext_s0_t[20]), .Z0_f (OUT_ciphertext_s0_f[20]), .Z1_t (OUT_ciphertext_s1_t[20]), .Z1_f (OUT_ciphertext_s1_f[20]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_21_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[21]), .A0_f (new_AGEMA_signal_5694), .A1_t (new_AGEMA_signal_5695), .A1_f (new_AGEMA_signal_5696), .B0_t (IN_plaintext_s0_t[21]), .B0_f (IN_plaintext_s0_f[21]), .B1_t (IN_plaintext_s1_t[21]), .B1_f (IN_plaintext_s1_f[21]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_21_U1_X), .Z0_f (new_AGEMA_signal_6054), .Z1_t (new_AGEMA_signal_6055), .Z1_f (new_AGEMA_signal_6056) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_21_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (IN_reset_t), .A1_f (IN_reset_f), .B0_t (LED_128_Instance_MUX_state1_mux_inst_21_U1_X), .B0_f (new_AGEMA_signal_6054), .B1_t (new_AGEMA_signal_6055), .B1_f (new_AGEMA_signal_6056), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_21_U1_Y), .Z0_f (new_AGEMA_signal_6213), .Z1_t (new_AGEMA_signal_6214), .Z1_f (new_AGEMA_signal_6215) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_21_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_21_U1_Y), .A0_f (new_AGEMA_signal_6213), .A1_t (new_AGEMA_signal_6214), .A1_f (new_AGEMA_signal_6215), .B0_t (LED_128_Instance_state0[21]), .B0_f (new_AGEMA_signal_5694), .B1_t (new_AGEMA_signal_5695), .B1_f (new_AGEMA_signal_5696), .Z0_t (OUT_ciphertext_s0_t[21]), .Z0_f (OUT_ciphertext_s0_f[21]), .Z1_t (OUT_ciphertext_s1_t[21]), .Z1_f (OUT_ciphertext_s1_f[21]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_22_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[22]), .A0_f (new_AGEMA_signal_6078), .A1_t (new_AGEMA_signal_6079), .A1_f (new_AGEMA_signal_6080), .B0_t (IN_plaintext_s0_t[22]), .B0_f (IN_plaintext_s0_f[22]), .B1_t (IN_plaintext_s1_t[22]), .B1_f (IN_plaintext_s1_f[22]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_22_U1_X), .Z0_f (new_AGEMA_signal_6381), .Z1_t (new_AGEMA_signal_6382), .Z1_f (new_AGEMA_signal_6383) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_22_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (IN_reset_t), .A1_f (IN_reset_f), .B0_t (LED_128_Instance_MUX_state1_mux_inst_22_U1_X), .B0_f (new_AGEMA_signal_6381), .B1_t (new_AGEMA_signal_6382), .B1_f (new_AGEMA_signal_6383), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_22_U1_Y), .Z0_f (new_AGEMA_signal_6540), .Z1_t (new_AGEMA_signal_6541), .Z1_f (new_AGEMA_signal_6542) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_22_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_22_U1_Y), .A0_f (new_AGEMA_signal_6540), .A1_t (new_AGEMA_signal_6541), .A1_f (new_AGEMA_signal_6542), .B0_t (LED_128_Instance_state0[22]), .B0_f (new_AGEMA_signal_6078), .B1_t (new_AGEMA_signal_6079), .B1_f (new_AGEMA_signal_6080), .Z0_t (OUT_ciphertext_s0_t[22]), .Z0_f (OUT_ciphertext_s0_f[22]), .Z1_t (OUT_ciphertext_s1_t[22]), .Z1_f (OUT_ciphertext_s1_f[22]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_23_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[23]), .A0_f (new_AGEMA_signal_6081), .A1_t (new_AGEMA_signal_6082), .A1_f (new_AGEMA_signal_6083), .B0_t (IN_plaintext_s0_t[23]), .B0_f (IN_plaintext_s0_f[23]), .B1_t (IN_plaintext_s1_t[23]), .B1_f (IN_plaintext_s1_f[23]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_23_U1_X), .Z0_f (new_AGEMA_signal_6387), .Z1_t (new_AGEMA_signal_6388), .Z1_f (new_AGEMA_signal_6389) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_23_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (IN_reset_t), .A1_f (IN_reset_f), .B0_t (LED_128_Instance_MUX_state1_mux_inst_23_U1_X), .B0_f (new_AGEMA_signal_6387), .B1_t (new_AGEMA_signal_6388), .B1_f (new_AGEMA_signal_6389), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_23_U1_Y), .Z0_f (new_AGEMA_signal_6543), .Z1_t (new_AGEMA_signal_6544), .Z1_f (new_AGEMA_signal_6545) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_23_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_23_U1_Y), .A0_f (new_AGEMA_signal_6543), .A1_t (new_AGEMA_signal_6544), .A1_f (new_AGEMA_signal_6545), .B0_t (LED_128_Instance_state0[23]), .B0_f (new_AGEMA_signal_6081), .B1_t (new_AGEMA_signal_6082), .B1_f (new_AGEMA_signal_6083), .Z0_t (OUT_ciphertext_s0_t[23]), .Z0_f (OUT_ciphertext_s0_f[23]), .Z1_t (OUT_ciphertext_s1_t[23]), .Z1_f (OUT_ciphertext_s1_f[23]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_24_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[24]), .A0_f (new_AGEMA_signal_5883), .A1_t (new_AGEMA_signal_5884), .A1_f (new_AGEMA_signal_5885), .B0_t (IN_plaintext_s0_t[24]), .B0_f (IN_plaintext_s0_f[24]), .B1_t (IN_plaintext_s1_t[24]), .B1_f (IN_plaintext_s1_f[24]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_24_U1_X), .Z0_f (new_AGEMA_signal_6219), .Z1_t (new_AGEMA_signal_6220), .Z1_f (new_AGEMA_signal_6221) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_24_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (IN_reset_t), .A1_f (IN_reset_f), .B0_t (LED_128_Instance_MUX_state1_mux_inst_24_U1_X), .B0_f (new_AGEMA_signal_6219), .B1_t (new_AGEMA_signal_6220), .B1_f (new_AGEMA_signal_6221), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_24_U1_Y), .Z0_f (new_AGEMA_signal_6390), .Z1_t (new_AGEMA_signal_6391), .Z1_f (new_AGEMA_signal_6392) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_24_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_24_U1_Y), .A0_f (new_AGEMA_signal_6390), .A1_t (new_AGEMA_signal_6391), .A1_f (new_AGEMA_signal_6392), .B0_t (LED_128_Instance_state0[24]), .B0_f (new_AGEMA_signal_5883), .B1_t (new_AGEMA_signal_5884), .B1_f (new_AGEMA_signal_5885), .Z0_t (OUT_ciphertext_s0_t[24]), .Z0_f (OUT_ciphertext_s0_f[24]), .Z1_t (OUT_ciphertext_s1_t[24]), .Z1_f (OUT_ciphertext_s1_f[24]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_25_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[25]), .A0_f (new_AGEMA_signal_5886), .A1_t (new_AGEMA_signal_5887), .A1_f (new_AGEMA_signal_5888), .B0_t (IN_plaintext_s0_t[25]), .B0_f (IN_plaintext_s0_f[25]), .B1_t (IN_plaintext_s1_t[25]), .B1_f (IN_plaintext_s1_f[25]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_25_U1_X), .Z0_f (new_AGEMA_signal_6225), .Z1_t (new_AGEMA_signal_6226), .Z1_f (new_AGEMA_signal_6227) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_25_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (IN_reset_t), .A1_f (IN_reset_f), .B0_t (LED_128_Instance_MUX_state1_mux_inst_25_U1_X), .B0_f (new_AGEMA_signal_6225), .B1_t (new_AGEMA_signal_6226), .B1_f (new_AGEMA_signal_6227), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_25_U1_Y), .Z0_f (new_AGEMA_signal_6393), .Z1_t (new_AGEMA_signal_6394), .Z1_f (new_AGEMA_signal_6395) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_25_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_25_U1_Y), .A0_f (new_AGEMA_signal_6393), .A1_t (new_AGEMA_signal_6394), .A1_f (new_AGEMA_signal_6395), .B0_t (LED_128_Instance_state0[25]), .B0_f (new_AGEMA_signal_5886), .B1_t (new_AGEMA_signal_5887), .B1_f (new_AGEMA_signal_5888), .Z0_t (OUT_ciphertext_s0_t[25]), .Z0_f (OUT_ciphertext_s0_f[25]), .Z1_t (OUT_ciphertext_s1_t[25]), .Z1_f (OUT_ciphertext_s1_f[25]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_26_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[26]), .A0_f (new_AGEMA_signal_6084), .A1_t (new_AGEMA_signal_6085), .A1_f (new_AGEMA_signal_6086), .B0_t (IN_plaintext_s0_t[26]), .B0_f (IN_plaintext_s0_f[26]), .B1_t (IN_plaintext_s1_t[26]), .B1_f (IN_plaintext_s1_f[26]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_26_U1_X), .Z0_f (new_AGEMA_signal_6399), .Z1_t (new_AGEMA_signal_6400), .Z1_f (new_AGEMA_signal_6401) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_26_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (IN_reset_t), .A1_f (IN_reset_f), .B0_t (LED_128_Instance_MUX_state1_mux_inst_26_U1_X), .B0_f (new_AGEMA_signal_6399), .B1_t (new_AGEMA_signal_6400), .B1_f (new_AGEMA_signal_6401), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_26_U1_Y), .Z0_f (new_AGEMA_signal_6546), .Z1_t (new_AGEMA_signal_6547), .Z1_f (new_AGEMA_signal_6548) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_26_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_26_U1_Y), .A0_f (new_AGEMA_signal_6546), .A1_t (new_AGEMA_signal_6547), .A1_f (new_AGEMA_signal_6548), .B0_t (LED_128_Instance_state0[26]), .B0_f (new_AGEMA_signal_6084), .B1_t (new_AGEMA_signal_6085), .B1_f (new_AGEMA_signal_6086), .Z0_t (OUT_ciphertext_s0_t[26]), .Z0_f (OUT_ciphertext_s0_f[26]), .Z1_t (OUT_ciphertext_s1_t[26]), .Z1_f (OUT_ciphertext_s1_f[26]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_27_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[27]), .A0_f (new_AGEMA_signal_6087), .A1_t (new_AGEMA_signal_6088), .A1_f (new_AGEMA_signal_6089), .B0_t (IN_plaintext_s0_t[27]), .B0_f (IN_plaintext_s0_f[27]), .B1_t (IN_plaintext_s1_t[27]), .B1_f (IN_plaintext_s1_f[27]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_27_U1_X), .Z0_f (new_AGEMA_signal_6405), .Z1_t (new_AGEMA_signal_6406), .Z1_f (new_AGEMA_signal_6407) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_27_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (IN_reset_t), .A1_f (IN_reset_f), .B0_t (LED_128_Instance_MUX_state1_mux_inst_27_U1_X), .B0_f (new_AGEMA_signal_6405), .B1_t (new_AGEMA_signal_6406), .B1_f (new_AGEMA_signal_6407), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_27_U1_Y), .Z0_f (new_AGEMA_signal_6549), .Z1_t (new_AGEMA_signal_6550), .Z1_f (new_AGEMA_signal_6551) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_27_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_27_U1_Y), .A0_f (new_AGEMA_signal_6549), .A1_t (new_AGEMA_signal_6550), .A1_f (new_AGEMA_signal_6551), .B0_t (LED_128_Instance_state0[27]), .B0_f (new_AGEMA_signal_6087), .B1_t (new_AGEMA_signal_6088), .B1_f (new_AGEMA_signal_6089), .Z0_t (OUT_ciphertext_s0_t[27]), .Z0_f (OUT_ciphertext_s0_f[27]), .Z1_t (OUT_ciphertext_s1_t[27]), .Z1_f (OUT_ciphertext_s1_f[27]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_28_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[28]), .A0_f (new_AGEMA_signal_5895), .A1_t (new_AGEMA_signal_5896), .A1_f (new_AGEMA_signal_5897), .B0_t (IN_plaintext_s0_t[28]), .B0_f (IN_plaintext_s0_f[28]), .B1_t (IN_plaintext_s1_t[28]), .B1_f (IN_plaintext_s1_f[28]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_28_U1_X), .Z0_f (new_AGEMA_signal_6231), .Z1_t (new_AGEMA_signal_6232), .Z1_f (new_AGEMA_signal_6233) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_28_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (IN_reset_t), .A1_f (IN_reset_f), .B0_t (LED_128_Instance_MUX_state1_mux_inst_28_U1_X), .B0_f (new_AGEMA_signal_6231), .B1_t (new_AGEMA_signal_6232), .B1_f (new_AGEMA_signal_6233), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_28_U1_Y), .Z0_f (new_AGEMA_signal_6408), .Z1_t (new_AGEMA_signal_6409), .Z1_f (new_AGEMA_signal_6410) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_28_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_28_U1_Y), .A0_f (new_AGEMA_signal_6408), .A1_t (new_AGEMA_signal_6409), .A1_f (new_AGEMA_signal_6410), .B0_t (LED_128_Instance_state0[28]), .B0_f (new_AGEMA_signal_5895), .B1_t (new_AGEMA_signal_5896), .B1_f (new_AGEMA_signal_5897), .Z0_t (OUT_ciphertext_s0_t[28]), .Z0_f (OUT_ciphertext_s0_f[28]), .Z1_t (OUT_ciphertext_s1_t[28]), .Z1_f (OUT_ciphertext_s1_f[28]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_29_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[29]), .A0_f (new_AGEMA_signal_5898), .A1_t (new_AGEMA_signal_5899), .A1_f (new_AGEMA_signal_5900), .B0_t (IN_plaintext_s0_t[29]), .B0_f (IN_plaintext_s0_f[29]), .B1_t (IN_plaintext_s1_t[29]), .B1_f (IN_plaintext_s1_f[29]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_29_U1_X), .Z0_f (new_AGEMA_signal_6237), .Z1_t (new_AGEMA_signal_6238), .Z1_f (new_AGEMA_signal_6239) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_29_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (IN_reset_t), .A1_f (IN_reset_f), .B0_t (LED_128_Instance_MUX_state1_mux_inst_29_U1_X), .B0_f (new_AGEMA_signal_6237), .B1_t (new_AGEMA_signal_6238), .B1_f (new_AGEMA_signal_6239), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_29_U1_Y), .Z0_f (new_AGEMA_signal_6411), .Z1_t (new_AGEMA_signal_6412), .Z1_f (new_AGEMA_signal_6413) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_29_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_29_U1_Y), .A0_f (new_AGEMA_signal_6411), .A1_t (new_AGEMA_signal_6412), .A1_f (new_AGEMA_signal_6413), .B0_t (LED_128_Instance_state0[29]), .B0_f (new_AGEMA_signal_5898), .B1_t (new_AGEMA_signal_5899), .B1_f (new_AGEMA_signal_5900), .Z0_t (OUT_ciphertext_s0_t[29]), .Z0_f (OUT_ciphertext_s0_f[29]), .Z1_t (OUT_ciphertext_s1_t[29]), .Z1_f (OUT_ciphertext_s1_f[29]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_30_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[30]), .A0_f (new_AGEMA_signal_6309), .A1_t (new_AGEMA_signal_6310), .A1_f (new_AGEMA_signal_6311), .B0_t (IN_plaintext_s0_t[30]), .B0_f (IN_plaintext_s0_f[30]), .B1_t (IN_plaintext_s1_t[30]), .B1_f (IN_plaintext_s1_f[30]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_30_U1_X), .Z0_f (new_AGEMA_signal_6555), .Z1_t (new_AGEMA_signal_6556), .Z1_f (new_AGEMA_signal_6557) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_30_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (IN_reset_t), .A1_f (IN_reset_f), .B0_t (LED_128_Instance_MUX_state1_mux_inst_30_U1_X), .B0_f (new_AGEMA_signal_6555), .B1_t (new_AGEMA_signal_6556), .B1_f (new_AGEMA_signal_6557), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_30_U1_Y), .Z0_f (new_AGEMA_signal_6639), .Z1_t (new_AGEMA_signal_6640), .Z1_f (new_AGEMA_signal_6641) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_30_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_30_U1_Y), .A0_f (new_AGEMA_signal_6639), .A1_t (new_AGEMA_signal_6640), .A1_f (new_AGEMA_signal_6641), .B0_t (LED_128_Instance_state0[30]), .B0_f (new_AGEMA_signal_6309), .B1_t (new_AGEMA_signal_6310), .B1_f (new_AGEMA_signal_6311), .Z0_t (OUT_ciphertext_s0_t[30]), .Z0_f (OUT_ciphertext_s0_f[30]), .Z1_t (OUT_ciphertext_s1_t[30]), .Z1_f (OUT_ciphertext_s1_f[30]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_31_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[31]), .A0_f (new_AGEMA_signal_6312), .A1_t (new_AGEMA_signal_6313), .A1_f (new_AGEMA_signal_6314), .B0_t (IN_plaintext_s0_t[31]), .B0_f (IN_plaintext_s0_f[31]), .B1_t (IN_plaintext_s1_t[31]), .B1_f (IN_plaintext_s1_f[31]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_31_U1_X), .Z0_f (new_AGEMA_signal_6561), .Z1_t (new_AGEMA_signal_6562), .Z1_f (new_AGEMA_signal_6563) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_31_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (IN_reset_t), .A1_f (IN_reset_f), .B0_t (LED_128_Instance_MUX_state1_mux_inst_31_U1_X), .B0_f (new_AGEMA_signal_6561), .B1_t (new_AGEMA_signal_6562), .B1_f (new_AGEMA_signal_6563), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_31_U1_Y), .Z0_f (new_AGEMA_signal_6642), .Z1_t (new_AGEMA_signal_6643), .Z1_f (new_AGEMA_signal_6644) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_31_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_31_U1_Y), .A0_f (new_AGEMA_signal_6642), .A1_t (new_AGEMA_signal_6643), .A1_f (new_AGEMA_signal_6644), .B0_t (LED_128_Instance_state0[31]), .B0_f (new_AGEMA_signal_6312), .B1_t (new_AGEMA_signal_6313), .B1_f (new_AGEMA_signal_6314), .Z0_t (OUT_ciphertext_s0_t[31]), .Z0_f (OUT_ciphertext_s0_f[31]), .Z1_t (OUT_ciphertext_s1_t[31]), .Z1_f (OUT_ciphertext_s1_f[31]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_32_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[32]), .A0_f (new_AGEMA_signal_6315), .A1_t (new_AGEMA_signal_6316), .A1_f (new_AGEMA_signal_6317), .B0_t (IN_plaintext_s0_t[32]), .B0_f (IN_plaintext_s0_f[32]), .B1_t (IN_plaintext_s1_t[32]), .B1_f (IN_plaintext_s1_f[32]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_32_U1_X), .Z0_f (new_AGEMA_signal_6567), .Z1_t (new_AGEMA_signal_6568), .Z1_f (new_AGEMA_signal_6569) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_32_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (IN_reset_t), .A1_f (IN_reset_f), .B0_t (LED_128_Instance_MUX_state1_mux_inst_32_U1_X), .B0_f (new_AGEMA_signal_6567), .B1_t (new_AGEMA_signal_6568), .B1_f (new_AGEMA_signal_6569), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_32_U1_Y), .Z0_f (new_AGEMA_signal_6645), .Z1_t (new_AGEMA_signal_6646), .Z1_f (new_AGEMA_signal_6647) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_32_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_32_U1_Y), .A0_f (new_AGEMA_signal_6645), .A1_t (new_AGEMA_signal_6646), .A1_f (new_AGEMA_signal_6647), .B0_t (LED_128_Instance_state0[32]), .B0_f (new_AGEMA_signal_6315), .B1_t (new_AGEMA_signal_6316), .B1_f (new_AGEMA_signal_6317), .Z0_t (OUT_ciphertext_s0_t[32]), .Z0_f (OUT_ciphertext_s0_f[32]), .Z1_t (OUT_ciphertext_s1_t[32]), .Z1_f (OUT_ciphertext_s1_f[32]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_33_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[33]), .A0_f (new_AGEMA_signal_6099), .A1_t (new_AGEMA_signal_6100), .A1_f (new_AGEMA_signal_6101), .B0_t (IN_plaintext_s0_t[33]), .B0_f (IN_plaintext_s0_f[33]), .B1_t (IN_plaintext_s1_t[33]), .B1_f (IN_plaintext_s1_f[33]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_33_U1_X), .Z0_f (new_AGEMA_signal_6417), .Z1_t (new_AGEMA_signal_6418), .Z1_f (new_AGEMA_signal_6419) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_33_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (IN_reset_t), .A1_f (IN_reset_f), .B0_t (LED_128_Instance_MUX_state1_mux_inst_33_U1_X), .B0_f (new_AGEMA_signal_6417), .B1_t (new_AGEMA_signal_6418), .B1_f (new_AGEMA_signal_6419), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_33_U1_Y), .Z0_f (new_AGEMA_signal_6570), .Z1_t (new_AGEMA_signal_6571), .Z1_f (new_AGEMA_signal_6572) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_33_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_33_U1_Y), .A0_f (new_AGEMA_signal_6570), .A1_t (new_AGEMA_signal_6571), .A1_f (new_AGEMA_signal_6572), .B0_t (LED_128_Instance_state0[33]), .B0_f (new_AGEMA_signal_6099), .B1_t (new_AGEMA_signal_6100), .B1_f (new_AGEMA_signal_6101), .Z0_t (OUT_ciphertext_s0_t[33]), .Z0_f (OUT_ciphertext_s0_f[33]), .Z1_t (OUT_ciphertext_s1_t[33]), .Z1_f (OUT_ciphertext_s1_f[33]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_34_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[34]), .A0_f (new_AGEMA_signal_5913), .A1_t (new_AGEMA_signal_5914), .A1_f (new_AGEMA_signal_5915), .B0_t (IN_plaintext_s0_t[34]), .B0_f (IN_plaintext_s0_f[34]), .B1_t (IN_plaintext_s1_t[34]), .B1_f (IN_plaintext_s1_f[34]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_34_U1_X), .Z0_f (new_AGEMA_signal_6243), .Z1_t (new_AGEMA_signal_6244), .Z1_f (new_AGEMA_signal_6245) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_34_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (IN_reset_t), .A1_f (IN_reset_f), .B0_t (LED_128_Instance_MUX_state1_mux_inst_34_U1_X), .B0_f (new_AGEMA_signal_6243), .B1_t (new_AGEMA_signal_6244), .B1_f (new_AGEMA_signal_6245), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_34_U1_Y), .Z0_f (new_AGEMA_signal_6420), .Z1_t (new_AGEMA_signal_6421), .Z1_f (new_AGEMA_signal_6422) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_34_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_34_U1_Y), .A0_f (new_AGEMA_signal_6420), .A1_t (new_AGEMA_signal_6421), .A1_f (new_AGEMA_signal_6422), .B0_t (LED_128_Instance_state0[34]), .B0_f (new_AGEMA_signal_5913), .B1_t (new_AGEMA_signal_5914), .B1_f (new_AGEMA_signal_5915), .Z0_t (OUT_ciphertext_s0_t[34]), .Z0_f (OUT_ciphertext_s0_f[34]), .Z1_t (OUT_ciphertext_s1_t[34]), .Z1_f (OUT_ciphertext_s1_f[34]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_35_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[35]), .A0_f (new_AGEMA_signal_5916), .A1_t (new_AGEMA_signal_5917), .A1_f (new_AGEMA_signal_5918), .B0_t (IN_plaintext_s0_t[35]), .B0_f (IN_plaintext_s0_f[35]), .B1_t (IN_plaintext_s1_t[35]), .B1_f (IN_plaintext_s1_f[35]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_35_U1_X), .Z0_f (new_AGEMA_signal_6249), .Z1_t (new_AGEMA_signal_6250), .Z1_f (new_AGEMA_signal_6251) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_35_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (IN_reset_t), .A1_f (IN_reset_f), .B0_t (LED_128_Instance_MUX_state1_mux_inst_35_U1_X), .B0_f (new_AGEMA_signal_6249), .B1_t (new_AGEMA_signal_6250), .B1_f (new_AGEMA_signal_6251), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_35_U1_Y), .Z0_f (new_AGEMA_signal_6423), .Z1_t (new_AGEMA_signal_6424), .Z1_f (new_AGEMA_signal_6425) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_35_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_35_U1_Y), .A0_f (new_AGEMA_signal_6423), .A1_t (new_AGEMA_signal_6424), .A1_f (new_AGEMA_signal_6425), .B0_t (LED_128_Instance_state0[35]), .B0_f (new_AGEMA_signal_5916), .B1_t (new_AGEMA_signal_5917), .B1_f (new_AGEMA_signal_5918), .Z0_t (OUT_ciphertext_s0_t[35]), .Z0_f (OUT_ciphertext_s0_f[35]), .Z1_t (OUT_ciphertext_s1_t[35]), .Z1_f (OUT_ciphertext_s1_f[35]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_36_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[36]), .A0_f (new_AGEMA_signal_6318), .A1_t (new_AGEMA_signal_6319), .A1_f (new_AGEMA_signal_6320), .B0_t (IN_plaintext_s0_t[36]), .B0_f (IN_plaintext_s0_f[36]), .B1_t (IN_plaintext_s1_t[36]), .B1_f (IN_plaintext_s1_f[36]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_36_U1_X), .Z0_f (new_AGEMA_signal_6576), .Z1_t (new_AGEMA_signal_6577), .Z1_f (new_AGEMA_signal_6578) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_36_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (IN_reset_t), .A1_f (IN_reset_f), .B0_t (LED_128_Instance_MUX_state1_mux_inst_36_U1_X), .B0_f (new_AGEMA_signal_6576), .B1_t (new_AGEMA_signal_6577), .B1_f (new_AGEMA_signal_6578), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_36_U1_Y), .Z0_f (new_AGEMA_signal_6648), .Z1_t (new_AGEMA_signal_6649), .Z1_f (new_AGEMA_signal_6650) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_36_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_36_U1_Y), .A0_f (new_AGEMA_signal_6648), .A1_t (new_AGEMA_signal_6649), .A1_f (new_AGEMA_signal_6650), .B0_t (LED_128_Instance_state0[36]), .B0_f (new_AGEMA_signal_6318), .B1_t (new_AGEMA_signal_6319), .B1_f (new_AGEMA_signal_6320), .Z0_t (OUT_ciphertext_s0_t[36]), .Z0_f (OUT_ciphertext_s0_f[36]), .Z1_t (OUT_ciphertext_s1_t[36]), .Z1_f (OUT_ciphertext_s1_f[36]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_37_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[37]), .A0_f (new_AGEMA_signal_6105), .A1_t (new_AGEMA_signal_6106), .A1_f (new_AGEMA_signal_6107), .B0_t (IN_plaintext_s0_t[37]), .B0_f (IN_plaintext_s0_f[37]), .B1_t (IN_plaintext_s1_t[37]), .B1_f (IN_plaintext_s1_f[37]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_37_U1_X), .Z0_f (new_AGEMA_signal_6429), .Z1_t (new_AGEMA_signal_6430), .Z1_f (new_AGEMA_signal_6431) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_37_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (IN_reset_t), .A1_f (IN_reset_f), .B0_t (LED_128_Instance_MUX_state1_mux_inst_37_U1_X), .B0_f (new_AGEMA_signal_6429), .B1_t (new_AGEMA_signal_6430), .B1_f (new_AGEMA_signal_6431), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_37_U1_Y), .Z0_f (new_AGEMA_signal_6579), .Z1_t (new_AGEMA_signal_6580), .Z1_f (new_AGEMA_signal_6581) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_37_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_37_U1_Y), .A0_f (new_AGEMA_signal_6579), .A1_t (new_AGEMA_signal_6580), .A1_f (new_AGEMA_signal_6581), .B0_t (LED_128_Instance_state0[37]), .B0_f (new_AGEMA_signal_6105), .B1_t (new_AGEMA_signal_6106), .B1_f (new_AGEMA_signal_6107), .Z0_t (OUT_ciphertext_s0_t[37]), .Z0_f (OUT_ciphertext_s0_f[37]), .Z1_t (OUT_ciphertext_s1_t[37]), .Z1_f (OUT_ciphertext_s1_f[37]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_38_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[38]), .A0_f (new_AGEMA_signal_5925), .A1_t (new_AGEMA_signal_5926), .A1_f (new_AGEMA_signal_5927), .B0_t (IN_plaintext_s0_t[38]), .B0_f (IN_plaintext_s0_f[38]), .B1_t (IN_plaintext_s1_t[38]), .B1_f (IN_plaintext_s1_f[38]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_38_U1_X), .Z0_f (new_AGEMA_signal_6255), .Z1_t (new_AGEMA_signal_6256), .Z1_f (new_AGEMA_signal_6257) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_38_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (IN_reset_t), .A1_f (IN_reset_f), .B0_t (LED_128_Instance_MUX_state1_mux_inst_38_U1_X), .B0_f (new_AGEMA_signal_6255), .B1_t (new_AGEMA_signal_6256), .B1_f (new_AGEMA_signal_6257), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_38_U1_Y), .Z0_f (new_AGEMA_signal_6432), .Z1_t (new_AGEMA_signal_6433), .Z1_f (new_AGEMA_signal_6434) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_38_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_38_U1_Y), .A0_f (new_AGEMA_signal_6432), .A1_t (new_AGEMA_signal_6433), .A1_f (new_AGEMA_signal_6434), .B0_t (LED_128_Instance_state0[38]), .B0_f (new_AGEMA_signal_5925), .B1_t (new_AGEMA_signal_5926), .B1_f (new_AGEMA_signal_5927), .Z0_t (OUT_ciphertext_s0_t[38]), .Z0_f (OUT_ciphertext_s0_f[38]), .Z1_t (OUT_ciphertext_s1_t[38]), .Z1_f (OUT_ciphertext_s1_f[38]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_39_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[39]), .A0_f (new_AGEMA_signal_6108), .A1_t (new_AGEMA_signal_6109), .A1_f (new_AGEMA_signal_6110), .B0_t (IN_plaintext_s0_t[39]), .B0_f (IN_plaintext_s0_f[39]), .B1_t (IN_plaintext_s1_t[39]), .B1_f (IN_plaintext_s1_f[39]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_39_U1_X), .Z0_f (new_AGEMA_signal_6438), .Z1_t (new_AGEMA_signal_6439), .Z1_f (new_AGEMA_signal_6440) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_39_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (IN_reset_t), .A1_f (IN_reset_f), .B0_t (LED_128_Instance_MUX_state1_mux_inst_39_U1_X), .B0_f (new_AGEMA_signal_6438), .B1_t (new_AGEMA_signal_6439), .B1_f (new_AGEMA_signal_6440), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_39_U1_Y), .Z0_f (new_AGEMA_signal_6582), .Z1_t (new_AGEMA_signal_6583), .Z1_f (new_AGEMA_signal_6584) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_39_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_39_U1_Y), .A0_f (new_AGEMA_signal_6582), .A1_t (new_AGEMA_signal_6583), .A1_f (new_AGEMA_signal_6584), .B0_t (LED_128_Instance_state0[39]), .B0_f (new_AGEMA_signal_6108), .B1_t (new_AGEMA_signal_6109), .B1_f (new_AGEMA_signal_6110), .Z0_t (OUT_ciphertext_s0_t[39]), .Z0_f (OUT_ciphertext_s0_f[39]), .Z1_t (OUT_ciphertext_s1_t[39]), .Z1_f (OUT_ciphertext_s1_f[39]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_40_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[40]), .A0_f (new_AGEMA_signal_6321), .A1_t (new_AGEMA_signal_6322), .A1_f (new_AGEMA_signal_6323), .B0_t (IN_plaintext_s0_t[40]), .B0_f (IN_plaintext_s0_f[40]), .B1_t (IN_plaintext_s1_t[40]), .B1_f (IN_plaintext_s1_f[40]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_40_U1_X), .Z0_f (new_AGEMA_signal_6588), .Z1_t (new_AGEMA_signal_6589), .Z1_f (new_AGEMA_signal_6590) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_40_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (IN_reset_t), .A1_f (IN_reset_f), .B0_t (LED_128_Instance_MUX_state1_mux_inst_40_U1_X), .B0_f (new_AGEMA_signal_6588), .B1_t (new_AGEMA_signal_6589), .B1_f (new_AGEMA_signal_6590), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_40_U1_Y), .Z0_f (new_AGEMA_signal_6651), .Z1_t (new_AGEMA_signal_6652), .Z1_f (new_AGEMA_signal_6653) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_40_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_40_U1_Y), .A0_f (new_AGEMA_signal_6651), .A1_t (new_AGEMA_signal_6652), .A1_f (new_AGEMA_signal_6653), .B0_t (LED_128_Instance_state0[40]), .B0_f (new_AGEMA_signal_6321), .B1_t (new_AGEMA_signal_6322), .B1_f (new_AGEMA_signal_6323), .Z0_t (OUT_ciphertext_s0_t[40]), .Z0_f (OUT_ciphertext_s0_f[40]), .Z1_t (OUT_ciphertext_s1_t[40]), .Z1_f (OUT_ciphertext_s1_f[40]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_41_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[41]), .A0_f (new_AGEMA_signal_6114), .A1_t (new_AGEMA_signal_6115), .A1_f (new_AGEMA_signal_6116), .B0_t (IN_plaintext_s0_t[41]), .B0_f (IN_plaintext_s0_f[41]), .B1_t (IN_plaintext_s1_t[41]), .B1_f (IN_plaintext_s1_f[41]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_41_U1_X), .Z0_f (new_AGEMA_signal_6444), .Z1_t (new_AGEMA_signal_6445), .Z1_f (new_AGEMA_signal_6446) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_41_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (IN_reset_t), .A1_f (IN_reset_f), .B0_t (LED_128_Instance_MUX_state1_mux_inst_41_U1_X), .B0_f (new_AGEMA_signal_6444), .B1_t (new_AGEMA_signal_6445), .B1_f (new_AGEMA_signal_6446), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_41_U1_Y), .Z0_f (new_AGEMA_signal_6591), .Z1_t (new_AGEMA_signal_6592), .Z1_f (new_AGEMA_signal_6593) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_41_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_41_U1_Y), .A0_f (new_AGEMA_signal_6591), .A1_t (new_AGEMA_signal_6592), .A1_f (new_AGEMA_signal_6593), .B0_t (LED_128_Instance_state0[41]), .B0_f (new_AGEMA_signal_6114), .B1_t (new_AGEMA_signal_6115), .B1_f (new_AGEMA_signal_6116), .Z0_t (OUT_ciphertext_s0_t[41]), .Z0_f (OUT_ciphertext_s0_f[41]), .Z1_t (OUT_ciphertext_s1_t[41]), .Z1_f (OUT_ciphertext_s1_f[41]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_42_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[42]), .A0_f (new_AGEMA_signal_5937), .A1_t (new_AGEMA_signal_5938), .A1_f (new_AGEMA_signal_5939), .B0_t (IN_plaintext_s0_t[42]), .B0_f (IN_plaintext_s0_f[42]), .B1_t (IN_plaintext_s1_t[42]), .B1_f (IN_plaintext_s1_f[42]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_42_U1_X), .Z0_f (new_AGEMA_signal_6261), .Z1_t (new_AGEMA_signal_6262), .Z1_f (new_AGEMA_signal_6263) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_42_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (IN_reset_t), .A1_f (IN_reset_f), .B0_t (LED_128_Instance_MUX_state1_mux_inst_42_U1_X), .B0_f (new_AGEMA_signal_6261), .B1_t (new_AGEMA_signal_6262), .B1_f (new_AGEMA_signal_6263), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_42_U1_Y), .Z0_f (new_AGEMA_signal_6447), .Z1_t (new_AGEMA_signal_6448), .Z1_f (new_AGEMA_signal_6449) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_42_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_42_U1_Y), .A0_f (new_AGEMA_signal_6447), .A1_t (new_AGEMA_signal_6448), .A1_f (new_AGEMA_signal_6449), .B0_t (LED_128_Instance_state0[42]), .B0_f (new_AGEMA_signal_5937), .B1_t (new_AGEMA_signal_5938), .B1_f (new_AGEMA_signal_5939), .Z0_t (OUT_ciphertext_s0_t[42]), .Z0_f (OUT_ciphertext_s0_f[42]), .Z1_t (OUT_ciphertext_s1_t[42]), .Z1_f (OUT_ciphertext_s1_f[42]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_43_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[43]), .A0_f (new_AGEMA_signal_5940), .A1_t (new_AGEMA_signal_5941), .A1_f (new_AGEMA_signal_5942), .B0_t (IN_plaintext_s0_t[43]), .B0_f (IN_plaintext_s0_f[43]), .B1_t (IN_plaintext_s1_t[43]), .B1_f (IN_plaintext_s1_f[43]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_43_U1_X), .Z0_f (new_AGEMA_signal_6267), .Z1_t (new_AGEMA_signal_6268), .Z1_f (new_AGEMA_signal_6269) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_43_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (IN_reset_t), .A1_f (IN_reset_f), .B0_t (LED_128_Instance_MUX_state1_mux_inst_43_U1_X), .B0_f (new_AGEMA_signal_6267), .B1_t (new_AGEMA_signal_6268), .B1_f (new_AGEMA_signal_6269), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_43_U1_Y), .Z0_f (new_AGEMA_signal_6450), .Z1_t (new_AGEMA_signal_6451), .Z1_f (new_AGEMA_signal_6452) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_43_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_43_U1_Y), .A0_f (new_AGEMA_signal_6450), .A1_t (new_AGEMA_signal_6451), .A1_f (new_AGEMA_signal_6452), .B0_t (LED_128_Instance_state0[43]), .B0_f (new_AGEMA_signal_5940), .B1_t (new_AGEMA_signal_5941), .B1_f (new_AGEMA_signal_5942), .Z0_t (OUT_ciphertext_s0_t[43]), .Z0_f (OUT_ciphertext_s0_f[43]), .Z1_t (OUT_ciphertext_s1_t[43]), .Z1_f (OUT_ciphertext_s1_f[43]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_44_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[44]), .A0_f (new_AGEMA_signal_6525), .A1_t (new_AGEMA_signal_6526), .A1_f (new_AGEMA_signal_6527), .B0_t (IN_plaintext_s0_t[44]), .B0_f (IN_plaintext_s0_f[44]), .B1_t (IN_plaintext_s1_t[44]), .B1_f (IN_plaintext_s1_f[44]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_44_U1_X), .Z0_f (new_AGEMA_signal_6657), .Z1_t (new_AGEMA_signal_6658), .Z1_f (new_AGEMA_signal_6659) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_44_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (IN_reset_t), .A1_f (IN_reset_f), .B0_t (LED_128_Instance_MUX_state1_mux_inst_44_U1_X), .B0_f (new_AGEMA_signal_6657), .B1_t (new_AGEMA_signal_6658), .B1_f (new_AGEMA_signal_6659), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_44_U1_Y), .Z0_f (new_AGEMA_signal_6669), .Z1_t (new_AGEMA_signal_6670), .Z1_f (new_AGEMA_signal_6671) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_44_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_44_U1_Y), .A0_f (new_AGEMA_signal_6669), .A1_t (new_AGEMA_signal_6670), .A1_f (new_AGEMA_signal_6671), .B0_t (LED_128_Instance_state0[44]), .B0_f (new_AGEMA_signal_6525), .B1_t (new_AGEMA_signal_6526), .B1_f (new_AGEMA_signal_6527), .Z0_t (OUT_ciphertext_s0_t[44]), .Z0_f (OUT_ciphertext_s0_f[44]), .Z1_t (OUT_ciphertext_s1_t[44]), .Z1_f (OUT_ciphertext_s1_f[44]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_45_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[45]), .A0_f (new_AGEMA_signal_6327), .A1_t (new_AGEMA_signal_6328), .A1_f (new_AGEMA_signal_6329), .B0_t (IN_plaintext_s0_t[45]), .B0_f (IN_plaintext_s0_f[45]), .B1_t (IN_plaintext_s1_t[45]), .B1_f (IN_plaintext_s1_f[45]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_45_U1_X), .Z0_f (new_AGEMA_signal_6597), .Z1_t (new_AGEMA_signal_6598), .Z1_f (new_AGEMA_signal_6599) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_45_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (IN_reset_t), .A1_f (IN_reset_f), .B0_t (LED_128_Instance_MUX_state1_mux_inst_45_U1_X), .B0_f (new_AGEMA_signal_6597), .B1_t (new_AGEMA_signal_6598), .B1_f (new_AGEMA_signal_6599), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_45_U1_Y), .Z0_f (new_AGEMA_signal_6660), .Z1_t (new_AGEMA_signal_6661), .Z1_f (new_AGEMA_signal_6662) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_45_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_45_U1_Y), .A0_f (new_AGEMA_signal_6660), .A1_t (new_AGEMA_signal_6661), .A1_f (new_AGEMA_signal_6662), .B0_t (LED_128_Instance_state0[45]), .B0_f (new_AGEMA_signal_6327), .B1_t (new_AGEMA_signal_6328), .B1_f (new_AGEMA_signal_6329), .Z0_t (OUT_ciphertext_s0_t[45]), .Z0_f (OUT_ciphertext_s0_f[45]), .Z1_t (OUT_ciphertext_s1_t[45]), .Z1_f (OUT_ciphertext_s1_f[45]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_46_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[46]), .A0_f (new_AGEMA_signal_6123), .A1_t (new_AGEMA_signal_6124), .A1_f (new_AGEMA_signal_6125), .B0_t (IN_plaintext_s0_t[46]), .B0_f (IN_plaintext_s0_f[46]), .B1_t (IN_plaintext_s1_t[46]), .B1_f (IN_plaintext_s1_f[46]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_46_U1_X), .Z0_f (new_AGEMA_signal_6456), .Z1_t (new_AGEMA_signal_6457), .Z1_f (new_AGEMA_signal_6458) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_46_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (IN_reset_t), .A1_f (IN_reset_f), .B0_t (LED_128_Instance_MUX_state1_mux_inst_46_U1_X), .B0_f (new_AGEMA_signal_6456), .B1_t (new_AGEMA_signal_6457), .B1_f (new_AGEMA_signal_6458), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_46_U1_Y), .Z0_f (new_AGEMA_signal_6600), .Z1_t (new_AGEMA_signal_6601), .Z1_f (new_AGEMA_signal_6602) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_46_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_46_U1_Y), .A0_f (new_AGEMA_signal_6600), .A1_t (new_AGEMA_signal_6601), .A1_f (new_AGEMA_signal_6602), .B0_t (LED_128_Instance_state0[46]), .B0_f (new_AGEMA_signal_6123), .B1_t (new_AGEMA_signal_6124), .B1_f (new_AGEMA_signal_6125), .Z0_t (OUT_ciphertext_s0_t[46]), .Z0_f (OUT_ciphertext_s0_f[46]), .Z1_t (OUT_ciphertext_s1_t[46]), .Z1_f (OUT_ciphertext_s1_f[46]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_47_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[47]), .A0_f (new_AGEMA_signal_6126), .A1_t (new_AGEMA_signal_6127), .A1_f (new_AGEMA_signal_6128), .B0_t (IN_plaintext_s0_t[47]), .B0_f (IN_plaintext_s0_f[47]), .B1_t (IN_plaintext_s1_t[47]), .B1_f (IN_plaintext_s1_f[47]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_47_U1_X), .Z0_f (new_AGEMA_signal_6462), .Z1_t (new_AGEMA_signal_6463), .Z1_f (new_AGEMA_signal_6464) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_47_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (IN_reset_t), .A1_f (IN_reset_f), .B0_t (LED_128_Instance_MUX_state1_mux_inst_47_U1_X), .B0_f (new_AGEMA_signal_6462), .B1_t (new_AGEMA_signal_6463), .B1_f (new_AGEMA_signal_6464), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_47_U1_Y), .Z0_f (new_AGEMA_signal_6603), .Z1_t (new_AGEMA_signal_6604), .Z1_f (new_AGEMA_signal_6605) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_47_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_47_U1_Y), .A0_f (new_AGEMA_signal_6603), .A1_t (new_AGEMA_signal_6604), .A1_f (new_AGEMA_signal_6605), .B0_t (LED_128_Instance_state0[47]), .B0_f (new_AGEMA_signal_6126), .B1_t (new_AGEMA_signal_6127), .B1_f (new_AGEMA_signal_6128), .Z0_t (OUT_ciphertext_s0_t[47]), .Z0_f (OUT_ciphertext_s0_f[47]), .Z1_t (OUT_ciphertext_s1_t[47]), .Z1_f (OUT_ciphertext_s1_f[47]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_48_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[48]), .A0_f (new_AGEMA_signal_6129), .A1_t (new_AGEMA_signal_6130), .A1_f (new_AGEMA_signal_6131), .B0_t (IN_plaintext_s0_t[48]), .B0_f (IN_plaintext_s0_f[48]), .B1_t (IN_plaintext_s1_t[48]), .B1_f (IN_plaintext_s1_f[48]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_48_U1_X), .Z0_f (new_AGEMA_signal_6468), .Z1_t (new_AGEMA_signal_6469), .Z1_f (new_AGEMA_signal_6470) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_48_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (IN_reset_t), .A1_f (IN_reset_f), .B0_t (LED_128_Instance_MUX_state1_mux_inst_48_U1_X), .B0_f (new_AGEMA_signal_6468), .B1_t (new_AGEMA_signal_6469), .B1_f (new_AGEMA_signal_6470), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_48_U1_Y), .Z0_f (new_AGEMA_signal_6606), .Z1_t (new_AGEMA_signal_6607), .Z1_f (new_AGEMA_signal_6608) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_48_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_48_U1_Y), .A0_f (new_AGEMA_signal_6606), .A1_t (new_AGEMA_signal_6607), .A1_f (new_AGEMA_signal_6608), .B0_t (LED_128_Instance_state0[48]), .B0_f (new_AGEMA_signal_6129), .B1_t (new_AGEMA_signal_6130), .B1_f (new_AGEMA_signal_6131), .Z0_t (OUT_ciphertext_s0_t[48]), .Z0_f (OUT_ciphertext_s0_f[48]), .Z1_t (OUT_ciphertext_s1_t[48]), .Z1_f (OUT_ciphertext_s1_f[48]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_49_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[49]), .A0_f (new_AGEMA_signal_6132), .A1_t (new_AGEMA_signal_6133), .A1_f (new_AGEMA_signal_6134), .B0_t (IN_plaintext_s0_t[49]), .B0_f (IN_plaintext_s0_f[49]), .B1_t (IN_plaintext_s1_t[49]), .B1_f (IN_plaintext_s1_f[49]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_49_U1_X), .Z0_f (new_AGEMA_signal_6474), .Z1_t (new_AGEMA_signal_6475), .Z1_f (new_AGEMA_signal_6476) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_49_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (IN_reset_t), .A1_f (IN_reset_f), .B0_t (LED_128_Instance_MUX_state1_mux_inst_49_U1_X), .B0_f (new_AGEMA_signal_6474), .B1_t (new_AGEMA_signal_6475), .B1_f (new_AGEMA_signal_6476), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_49_U1_Y), .Z0_f (new_AGEMA_signal_6609), .Z1_t (new_AGEMA_signal_6610), .Z1_f (new_AGEMA_signal_6611) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_49_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_49_U1_Y), .A0_f (new_AGEMA_signal_6609), .A1_t (new_AGEMA_signal_6610), .A1_f (new_AGEMA_signal_6611), .B0_t (LED_128_Instance_state0[49]), .B0_f (new_AGEMA_signal_6132), .B1_t (new_AGEMA_signal_6133), .B1_f (new_AGEMA_signal_6134), .Z0_t (OUT_ciphertext_s0_t[49]), .Z0_f (OUT_ciphertext_s0_f[49]), .Z1_t (OUT_ciphertext_s1_t[49]), .Z1_f (OUT_ciphertext_s1_f[49]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_50_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[50]), .A0_f (new_AGEMA_signal_5958), .A1_t (new_AGEMA_signal_5959), .A1_f (new_AGEMA_signal_5960), .B0_t (IN_plaintext_s0_t[50]), .B0_f (IN_plaintext_s0_f[50]), .B1_t (IN_plaintext_s1_t[50]), .B1_f (IN_plaintext_s1_f[50]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_50_U1_X), .Z0_f (new_AGEMA_signal_6273), .Z1_t (new_AGEMA_signal_6274), .Z1_f (new_AGEMA_signal_6275) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_50_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (IN_reset_t), .A1_f (IN_reset_f), .B0_t (LED_128_Instance_MUX_state1_mux_inst_50_U1_X), .B0_f (new_AGEMA_signal_6273), .B1_t (new_AGEMA_signal_6274), .B1_f (new_AGEMA_signal_6275), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_50_U1_Y), .Z0_f (new_AGEMA_signal_6477), .Z1_t (new_AGEMA_signal_6478), .Z1_f (new_AGEMA_signal_6479) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_50_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_50_U1_Y), .A0_f (new_AGEMA_signal_6477), .A1_t (new_AGEMA_signal_6478), .A1_f (new_AGEMA_signal_6479), .B0_t (LED_128_Instance_state0[50]), .B0_f (new_AGEMA_signal_5958), .B1_t (new_AGEMA_signal_5959), .B1_f (new_AGEMA_signal_5960), .Z0_t (OUT_ciphertext_s0_t[50]), .Z0_f (OUT_ciphertext_s0_f[50]), .Z1_t (OUT_ciphertext_s1_t[50]), .Z1_f (OUT_ciphertext_s1_f[50]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_51_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[51]), .A0_f (new_AGEMA_signal_5961), .A1_t (new_AGEMA_signal_5962), .A1_f (new_AGEMA_signal_5963), .B0_t (IN_plaintext_s0_t[51]), .B0_f (IN_plaintext_s0_f[51]), .B1_t (IN_plaintext_s1_t[51]), .B1_f (IN_plaintext_s1_f[51]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_51_U1_X), .Z0_f (new_AGEMA_signal_6279), .Z1_t (new_AGEMA_signal_6280), .Z1_f (new_AGEMA_signal_6281) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_51_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (IN_reset_t), .A1_f (IN_reset_f), .B0_t (LED_128_Instance_MUX_state1_mux_inst_51_U1_X), .B0_f (new_AGEMA_signal_6279), .B1_t (new_AGEMA_signal_6280), .B1_f (new_AGEMA_signal_6281), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_51_U1_Y), .Z0_f (new_AGEMA_signal_6480), .Z1_t (new_AGEMA_signal_6481), .Z1_f (new_AGEMA_signal_6482) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_51_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_51_U1_Y), .A0_f (new_AGEMA_signal_6480), .A1_t (new_AGEMA_signal_6481), .A1_f (new_AGEMA_signal_6482), .B0_t (LED_128_Instance_state0[51]), .B0_f (new_AGEMA_signal_5961), .B1_t (new_AGEMA_signal_5962), .B1_f (new_AGEMA_signal_5963), .Z0_t (OUT_ciphertext_s0_t[51]), .Z0_f (OUT_ciphertext_s0_f[51]), .Z1_t (OUT_ciphertext_s1_t[51]), .Z1_f (OUT_ciphertext_s1_f[51]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_52_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[52]), .A0_f (new_AGEMA_signal_6135), .A1_t (new_AGEMA_signal_6136), .A1_f (new_AGEMA_signal_6137), .B0_t (IN_plaintext_s0_t[52]), .B0_f (IN_plaintext_s0_f[52]), .B1_t (IN_plaintext_s1_t[52]), .B1_f (IN_plaintext_s1_f[52]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_52_U1_X), .Z0_f (new_AGEMA_signal_6486), .Z1_t (new_AGEMA_signal_6487), .Z1_f (new_AGEMA_signal_6488) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_52_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (IN_reset_t), .A1_f (IN_reset_f), .B0_t (LED_128_Instance_MUX_state1_mux_inst_52_U1_X), .B0_f (new_AGEMA_signal_6486), .B1_t (new_AGEMA_signal_6487), .B1_f (new_AGEMA_signal_6488), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_52_U1_Y), .Z0_f (new_AGEMA_signal_6612), .Z1_t (new_AGEMA_signal_6613), .Z1_f (new_AGEMA_signal_6614) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_52_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_52_U1_Y), .A0_f (new_AGEMA_signal_6612), .A1_t (new_AGEMA_signal_6613), .A1_f (new_AGEMA_signal_6614), .B0_t (LED_128_Instance_state0[52]), .B0_f (new_AGEMA_signal_6135), .B1_t (new_AGEMA_signal_6136), .B1_f (new_AGEMA_signal_6137), .Z0_t (OUT_ciphertext_s0_t[52]), .Z0_f (OUT_ciphertext_s0_f[52]), .Z1_t (OUT_ciphertext_s1_t[52]), .Z1_f (OUT_ciphertext_s1_f[52]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_53_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[53]), .A0_f (new_AGEMA_signal_6138), .A1_t (new_AGEMA_signal_6139), .A1_f (new_AGEMA_signal_6140), .B0_t (IN_plaintext_s0_t[53]), .B0_f (IN_plaintext_s0_f[53]), .B1_t (IN_plaintext_s1_t[53]), .B1_f (IN_plaintext_s1_f[53]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_53_U1_X), .Z0_f (new_AGEMA_signal_6492), .Z1_t (new_AGEMA_signal_6493), .Z1_f (new_AGEMA_signal_6494) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_53_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (IN_reset_t), .A1_f (IN_reset_f), .B0_t (LED_128_Instance_MUX_state1_mux_inst_53_U1_X), .B0_f (new_AGEMA_signal_6492), .B1_t (new_AGEMA_signal_6493), .B1_f (new_AGEMA_signal_6494), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_53_U1_Y), .Z0_f (new_AGEMA_signal_6615), .Z1_t (new_AGEMA_signal_6616), .Z1_f (new_AGEMA_signal_6617) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_53_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_53_U1_Y), .A0_f (new_AGEMA_signal_6615), .A1_t (new_AGEMA_signal_6616), .A1_f (new_AGEMA_signal_6617), .B0_t (LED_128_Instance_state0[53]), .B0_f (new_AGEMA_signal_6138), .B1_t (new_AGEMA_signal_6139), .B1_f (new_AGEMA_signal_6140), .Z0_t (OUT_ciphertext_s0_t[53]), .Z0_f (OUT_ciphertext_s0_f[53]), .Z1_t (OUT_ciphertext_s1_t[53]), .Z1_f (OUT_ciphertext_s1_f[53]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_54_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[54]), .A0_f (new_AGEMA_signal_5970), .A1_t (new_AGEMA_signal_5971), .A1_f (new_AGEMA_signal_5972), .B0_t (IN_plaintext_s0_t[54]), .B0_f (IN_plaintext_s0_f[54]), .B1_t (IN_plaintext_s1_t[54]), .B1_f (IN_plaintext_s1_f[54]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_54_U1_X), .Z0_f (new_AGEMA_signal_6285), .Z1_t (new_AGEMA_signal_6286), .Z1_f (new_AGEMA_signal_6287) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_54_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (IN_reset_t), .A1_f (IN_reset_f), .B0_t (LED_128_Instance_MUX_state1_mux_inst_54_U1_X), .B0_f (new_AGEMA_signal_6285), .B1_t (new_AGEMA_signal_6286), .B1_f (new_AGEMA_signal_6287), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_54_U1_Y), .Z0_f (new_AGEMA_signal_6495), .Z1_t (new_AGEMA_signal_6496), .Z1_f (new_AGEMA_signal_6497) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_54_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_54_U1_Y), .A0_f (new_AGEMA_signal_6495), .A1_t (new_AGEMA_signal_6496), .A1_f (new_AGEMA_signal_6497), .B0_t (LED_128_Instance_state0[54]), .B0_f (new_AGEMA_signal_5970), .B1_t (new_AGEMA_signal_5971), .B1_f (new_AGEMA_signal_5972), .Z0_t (OUT_ciphertext_s0_t[54]), .Z0_f (OUT_ciphertext_s0_f[54]), .Z1_t (OUT_ciphertext_s1_t[54]), .Z1_f (OUT_ciphertext_s1_f[54]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_55_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[55]), .A0_f (new_AGEMA_signal_5775), .A1_t (new_AGEMA_signal_5776), .A1_f (new_AGEMA_signal_5777), .B0_t (IN_plaintext_s0_t[55]), .B0_f (IN_plaintext_s0_f[55]), .B1_t (IN_plaintext_s1_t[55]), .B1_f (IN_plaintext_s1_f[55]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_55_U1_X), .Z0_f (new_AGEMA_signal_6060), .Z1_t (new_AGEMA_signal_6061), .Z1_f (new_AGEMA_signal_6062) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_55_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (IN_reset_t), .A1_f (IN_reset_f), .B0_t (LED_128_Instance_MUX_state1_mux_inst_55_U1_X), .B0_f (new_AGEMA_signal_6060), .B1_t (new_AGEMA_signal_6061), .B1_f (new_AGEMA_signal_6062), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_55_U1_Y), .Z0_f (new_AGEMA_signal_6288), .Z1_t (new_AGEMA_signal_6289), .Z1_f (new_AGEMA_signal_6290) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_55_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_55_U1_Y), .A0_f (new_AGEMA_signal_6288), .A1_t (new_AGEMA_signal_6289), .A1_f (new_AGEMA_signal_6290), .B0_t (LED_128_Instance_state0[55]), .B0_f (new_AGEMA_signal_5775), .B1_t (new_AGEMA_signal_5776), .B1_f (new_AGEMA_signal_5777), .Z0_t (OUT_ciphertext_s0_t[55]), .Z0_f (OUT_ciphertext_s0_f[55]), .Z1_t (OUT_ciphertext_s1_t[55]), .Z1_f (OUT_ciphertext_s1_f[55]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_56_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[56]), .A0_f (new_AGEMA_signal_6330), .A1_t (new_AGEMA_signal_6331), .A1_f (new_AGEMA_signal_6332), .B0_t (IN_plaintext_s0_t[56]), .B0_f (IN_plaintext_s0_f[56]), .B1_t (IN_plaintext_s1_t[56]), .B1_f (IN_plaintext_s1_f[56]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_56_U1_X), .Z0_f (new_AGEMA_signal_6621), .Z1_t (new_AGEMA_signal_6622), .Z1_f (new_AGEMA_signal_6623) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_56_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (IN_reset_t), .A1_f (IN_reset_f), .B0_t (LED_128_Instance_MUX_state1_mux_inst_56_U1_X), .B0_f (new_AGEMA_signal_6621), .B1_t (new_AGEMA_signal_6622), .B1_f (new_AGEMA_signal_6623), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_56_U1_Y), .Z0_f (new_AGEMA_signal_6663), .Z1_t (new_AGEMA_signal_6664), .Z1_f (new_AGEMA_signal_6665) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_56_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_56_U1_Y), .A0_f (new_AGEMA_signal_6663), .A1_t (new_AGEMA_signal_6664), .A1_f (new_AGEMA_signal_6665), .B0_t (LED_128_Instance_state0[56]), .B0_f (new_AGEMA_signal_6330), .B1_t (new_AGEMA_signal_6331), .B1_f (new_AGEMA_signal_6332), .Z0_t (OUT_ciphertext_s0_t[56]), .Z0_f (OUT_ciphertext_s0_f[56]), .Z1_t (OUT_ciphertext_s1_t[56]), .Z1_f (OUT_ciphertext_s1_f[56]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_57_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[57]), .A0_f (new_AGEMA_signal_6333), .A1_t (new_AGEMA_signal_6334), .A1_f (new_AGEMA_signal_6335), .B0_t (IN_plaintext_s0_t[57]), .B0_f (IN_plaintext_s0_f[57]), .B1_t (IN_plaintext_s1_t[57]), .B1_f (IN_plaintext_s1_f[57]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_57_U1_X), .Z0_f (new_AGEMA_signal_6627), .Z1_t (new_AGEMA_signal_6628), .Z1_f (new_AGEMA_signal_6629) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_57_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (IN_reset_t), .A1_f (IN_reset_f), .B0_t (LED_128_Instance_MUX_state1_mux_inst_57_U1_X), .B0_f (new_AGEMA_signal_6627), .B1_t (new_AGEMA_signal_6628), .B1_f (new_AGEMA_signal_6629), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_57_U1_Y), .Z0_f (new_AGEMA_signal_6666), .Z1_t (new_AGEMA_signal_6667), .Z1_f (new_AGEMA_signal_6668) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_57_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_57_U1_Y), .A0_f (new_AGEMA_signal_6666), .A1_t (new_AGEMA_signal_6667), .A1_f (new_AGEMA_signal_6668), .B0_t (LED_128_Instance_state0[57]), .B0_f (new_AGEMA_signal_6333), .B1_t (new_AGEMA_signal_6334), .B1_f (new_AGEMA_signal_6335), .Z0_t (OUT_ciphertext_s0_t[57]), .Z0_f (OUT_ciphertext_s0_f[57]), .Z1_t (OUT_ciphertext_s1_t[57]), .Z1_f (OUT_ciphertext_s1_f[57]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_58_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[58]), .A0_f (new_AGEMA_signal_6147), .A1_t (new_AGEMA_signal_6148), .A1_f (new_AGEMA_signal_6149), .B0_t (IN_plaintext_s0_t[58]), .B0_f (IN_plaintext_s0_f[58]), .B1_t (IN_plaintext_s1_t[58]), .B1_f (IN_plaintext_s1_f[58]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_58_U1_X), .Z0_f (new_AGEMA_signal_6501), .Z1_t (new_AGEMA_signal_6502), .Z1_f (new_AGEMA_signal_6503) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_58_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (IN_reset_t), .A1_f (IN_reset_f), .B0_t (LED_128_Instance_MUX_state1_mux_inst_58_U1_X), .B0_f (new_AGEMA_signal_6501), .B1_t (new_AGEMA_signal_6502), .B1_f (new_AGEMA_signal_6503), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_58_U1_Y), .Z0_f (new_AGEMA_signal_6630), .Z1_t (new_AGEMA_signal_6631), .Z1_f (new_AGEMA_signal_6632) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_58_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_58_U1_Y), .A0_f (new_AGEMA_signal_6630), .A1_t (new_AGEMA_signal_6631), .A1_f (new_AGEMA_signal_6632), .B0_t (LED_128_Instance_state0[58]), .B0_f (new_AGEMA_signal_6147), .B1_t (new_AGEMA_signal_6148), .B1_f (new_AGEMA_signal_6149), .Z0_t (OUT_ciphertext_s0_t[58]), .Z0_f (OUT_ciphertext_s0_f[58]), .Z1_t (OUT_ciphertext_s1_t[58]), .Z1_f (OUT_ciphertext_s1_f[58]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_59_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[59]), .A0_f (new_AGEMA_signal_5982), .A1_t (new_AGEMA_signal_5983), .A1_f (new_AGEMA_signal_5984), .B0_t (IN_plaintext_s0_t[59]), .B0_f (IN_plaintext_s0_f[59]), .B1_t (IN_plaintext_s1_t[59]), .B1_f (IN_plaintext_s1_f[59]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_59_U1_X), .Z0_f (new_AGEMA_signal_6294), .Z1_t (new_AGEMA_signal_6295), .Z1_f (new_AGEMA_signal_6296) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_59_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (IN_reset_t), .A1_f (IN_reset_f), .B0_t (LED_128_Instance_MUX_state1_mux_inst_59_U1_X), .B0_f (new_AGEMA_signal_6294), .B1_t (new_AGEMA_signal_6295), .B1_f (new_AGEMA_signal_6296), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_59_U1_Y), .Z0_f (new_AGEMA_signal_6504), .Z1_t (new_AGEMA_signal_6505), .Z1_f (new_AGEMA_signal_6506) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_59_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_59_U1_Y), .A0_f (new_AGEMA_signal_6504), .A1_t (new_AGEMA_signal_6505), .A1_f (new_AGEMA_signal_6506), .B0_t (LED_128_Instance_state0[59]), .B0_f (new_AGEMA_signal_5982), .B1_t (new_AGEMA_signal_5983), .B1_f (new_AGEMA_signal_5984), .Z0_t (OUT_ciphertext_s0_t[59]), .Z0_f (OUT_ciphertext_s0_f[59]), .Z1_t (OUT_ciphertext_s1_t[59]), .Z1_f (OUT_ciphertext_s1_f[59]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_60_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[60]), .A0_f (new_AGEMA_signal_6150), .A1_t (new_AGEMA_signal_6151), .A1_f (new_AGEMA_signal_6152), .B0_t (IN_plaintext_s0_t[60]), .B0_f (IN_plaintext_s0_f[60]), .B1_t (IN_plaintext_s1_t[60]), .B1_f (IN_plaintext_s1_f[60]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_60_U1_X), .Z0_f (new_AGEMA_signal_6510), .Z1_t (new_AGEMA_signal_6511), .Z1_f (new_AGEMA_signal_6512) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_60_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (IN_reset_t), .A1_f (IN_reset_f), .B0_t (LED_128_Instance_MUX_state1_mux_inst_60_U1_X), .B0_f (new_AGEMA_signal_6510), .B1_t (new_AGEMA_signal_6511), .B1_f (new_AGEMA_signal_6512), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_60_U1_Y), .Z0_f (new_AGEMA_signal_6633), .Z1_t (new_AGEMA_signal_6634), .Z1_f (new_AGEMA_signal_6635) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_60_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_60_U1_Y), .A0_f (new_AGEMA_signal_6633), .A1_t (new_AGEMA_signal_6634), .A1_f (new_AGEMA_signal_6635), .B0_t (LED_128_Instance_state0[60]), .B0_f (new_AGEMA_signal_6150), .B1_t (new_AGEMA_signal_6151), .B1_f (new_AGEMA_signal_6152), .Z0_t (OUT_ciphertext_s0_t[60]), .Z0_f (OUT_ciphertext_s0_f[60]), .Z1_t (OUT_ciphertext_s1_t[60]), .Z1_f (OUT_ciphertext_s1_f[60]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_61_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[61]), .A0_f (new_AGEMA_signal_6153), .A1_t (new_AGEMA_signal_6154), .A1_f (new_AGEMA_signal_6155), .B0_t (IN_plaintext_s0_t[61]), .B0_f (IN_plaintext_s0_f[61]), .B1_t (IN_plaintext_s1_t[61]), .B1_f (IN_plaintext_s1_f[61]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_61_U1_X), .Z0_f (new_AGEMA_signal_6516), .Z1_t (new_AGEMA_signal_6517), .Z1_f (new_AGEMA_signal_6518) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_61_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (IN_reset_t), .A1_f (IN_reset_f), .B0_t (LED_128_Instance_MUX_state1_mux_inst_61_U1_X), .B0_f (new_AGEMA_signal_6516), .B1_t (new_AGEMA_signal_6517), .B1_f (new_AGEMA_signal_6518), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_61_U1_Y), .Z0_f (new_AGEMA_signal_6636), .Z1_t (new_AGEMA_signal_6637), .Z1_f (new_AGEMA_signal_6638) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_61_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_61_U1_Y), .A0_f (new_AGEMA_signal_6636), .A1_t (new_AGEMA_signal_6637), .A1_f (new_AGEMA_signal_6638), .B0_t (LED_128_Instance_state0[61]), .B0_f (new_AGEMA_signal_6153), .B1_t (new_AGEMA_signal_6154), .B1_f (new_AGEMA_signal_6155), .Z0_t (OUT_ciphertext_s0_t[61]), .Z0_f (OUT_ciphertext_s0_f[61]), .Z1_t (OUT_ciphertext_s1_t[61]), .Z1_f (OUT_ciphertext_s1_f[61]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_62_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[62]), .A0_f (new_AGEMA_signal_5991), .A1_t (new_AGEMA_signal_5992), .A1_f (new_AGEMA_signal_5993), .B0_t (IN_plaintext_s0_t[62]), .B0_f (IN_plaintext_s0_f[62]), .B1_t (IN_plaintext_s1_t[62]), .B1_f (IN_plaintext_s1_f[62]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_62_U1_X), .Z0_f (new_AGEMA_signal_6300), .Z1_t (new_AGEMA_signal_6301), .Z1_f (new_AGEMA_signal_6302) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_62_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (IN_reset_t), .A1_f (IN_reset_f), .B0_t (LED_128_Instance_MUX_state1_mux_inst_62_U1_X), .B0_f (new_AGEMA_signal_6300), .B1_t (new_AGEMA_signal_6301), .B1_f (new_AGEMA_signal_6302), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_62_U1_Y), .Z0_f (new_AGEMA_signal_6519), .Z1_t (new_AGEMA_signal_6520), .Z1_f (new_AGEMA_signal_6521) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_62_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_62_U1_Y), .A0_f (new_AGEMA_signal_6519), .A1_t (new_AGEMA_signal_6520), .A1_f (new_AGEMA_signal_6521), .B0_t (LED_128_Instance_state0[62]), .B0_f (new_AGEMA_signal_5991), .B1_t (new_AGEMA_signal_5992), .B1_f (new_AGEMA_signal_5993), .Z0_t (OUT_ciphertext_s0_t[62]), .Z0_f (OUT_ciphertext_s0_f[62]), .Z1_t (OUT_ciphertext_s1_t[62]), .Z1_f (OUT_ciphertext_s1_f[62]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_63_U1_XOR1_U1 ( .A0_t (LED_128_Instance_state0[63]), .A0_f (new_AGEMA_signal_5994), .A1_t (new_AGEMA_signal_5995), .A1_f (new_AGEMA_signal_5996), .B0_t (IN_plaintext_s0_t[63]), .B0_f (IN_plaintext_s0_f[63]), .B1_t (IN_plaintext_s1_t[63]), .B1_f (IN_plaintext_s1_f[63]), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_63_U1_X), .Z0_f (new_AGEMA_signal_6306), .Z1_t (new_AGEMA_signal_6307), .Z1_f (new_AGEMA_signal_6308) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_state1_mux_inst_63_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (IN_reset_t), .A1_f (IN_reset_f), .B0_t (LED_128_Instance_MUX_state1_mux_inst_63_U1_X), .B0_f (new_AGEMA_signal_6306), .B1_t (new_AGEMA_signal_6307), .B1_f (new_AGEMA_signal_6308), .Z0_t (LED_128_Instance_MUX_state1_mux_inst_63_U1_Y), .Z0_f (new_AGEMA_signal_6522), .Z1_t (new_AGEMA_signal_6523), .Z1_f (new_AGEMA_signal_6524) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) LED_128_Instance_MUX_state1_mux_inst_63_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_state1_mux_inst_63_U1_Y), .A0_f (new_AGEMA_signal_6522), .A1_t (new_AGEMA_signal_6523), .A1_f (new_AGEMA_signal_6524), .B0_t (LED_128_Instance_state0[63]), .B0_f (new_AGEMA_signal_5994), .B1_t (new_AGEMA_signal_5995), .B1_f (new_AGEMA_signal_5996), .Z0_t (OUT_ciphertext_s0_t[63]), .Z0_f (OUT_ciphertext_s0_f[63]), .Z1_t (OUT_ciphertext_s1_t[63]), .Z1_f (OUT_ciphertext_s1_f[63]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_0_U1_XOR1_U1 ( .A0_t (IN_key_s0_t[64]), .A0_f (IN_key_s0_f[64]), .A1_t (IN_key_s1_t[64]), .A1_f (IN_key_s1_f[64]), .B0_t (IN_key_s0_t[0]), .B0_f (IN_key_s0_f[0]), .B1_t (IN_key_s1_t[0]), .B1_f (IN_key_s1_f[0]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_0_U1_X), .Z0_f (new_AGEMA_signal_1900), .Z1_t (new_AGEMA_signal_1901), .Z1_f (new_AGEMA_signal_1902) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_0_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n31), .A1_f (new_AGEMA_signal_2477), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_0_U1_X), .B0_f (new_AGEMA_signal_1900), .B1_t (new_AGEMA_signal_1901), .B1_f (new_AGEMA_signal_1902), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_0_U1_Y), .Z0_f (new_AGEMA_signal_2481), .Z1_t (new_AGEMA_signal_2482), .Z1_f (new_AGEMA_signal_2483) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_0_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_0_U1_Y), .A0_f (new_AGEMA_signal_2481), .A1_t (new_AGEMA_signal_2482), .A1_f (new_AGEMA_signal_2483), .B0_t (IN_key_s0_t[64]), .B0_f (IN_key_s0_f[64]), .B1_t (IN_key_s1_t[64]), .B1_f (IN_key_s1_f[64]), .Z0_t (LED_128_Instance_current_roundkey[0]), .Z0_f (new_AGEMA_signal_2674), .Z1_t (new_AGEMA_signal_2675), .Z1_f (new_AGEMA_signal_2676) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_1_U1_XOR1_U1 ( .A0_t (IN_key_s0_t[65]), .A0_f (IN_key_s0_f[65]), .A1_t (IN_key_s1_t[65]), .A1_f (IN_key_s1_f[65]), .B0_t (IN_key_s0_t[1]), .B0_f (IN_key_s0_f[1]), .B1_t (IN_key_s1_t[1]), .B1_f (IN_key_s1_f[1]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_1_U1_X), .Z0_f (new_AGEMA_signal_1909), .Z1_t (new_AGEMA_signal_1910), .Z1_f (new_AGEMA_signal_1911) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_1_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n31), .A1_f (new_AGEMA_signal_2477), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_1_U1_X), .B0_f (new_AGEMA_signal_1909), .B1_t (new_AGEMA_signal_1910), .B1_f (new_AGEMA_signal_1911), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_1_U1_Y), .Z0_f (new_AGEMA_signal_2484), .Z1_t (new_AGEMA_signal_2485), .Z1_f (new_AGEMA_signal_2486) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_1_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_1_U1_Y), .A0_f (new_AGEMA_signal_2484), .A1_t (new_AGEMA_signal_2485), .A1_f (new_AGEMA_signal_2486), .B0_t (IN_key_s0_t[65]), .B0_f (IN_key_s0_f[65]), .B1_t (IN_key_s1_t[65]), .B1_f (IN_key_s1_f[65]), .Z0_t (LED_128_Instance_current_roundkey[1]), .Z0_f (new_AGEMA_signal_2677), .Z1_t (new_AGEMA_signal_2678), .Z1_f (new_AGEMA_signal_2679) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_2_U1_XOR1_U1 ( .A0_t (IN_key_s0_t[66]), .A0_f (IN_key_s0_f[66]), .A1_t (IN_key_s1_t[66]), .A1_f (IN_key_s1_f[66]), .B0_t (IN_key_s0_t[2]), .B0_f (IN_key_s0_f[2]), .B1_t (IN_key_s1_t[2]), .B1_f (IN_key_s1_f[2]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_2_U1_X), .Z0_f (new_AGEMA_signal_1918), .Z1_t (new_AGEMA_signal_1919), .Z1_f (new_AGEMA_signal_1920) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_2_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n31), .A1_f (new_AGEMA_signal_2477), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_2_U1_X), .B0_f (new_AGEMA_signal_1918), .B1_t (new_AGEMA_signal_1919), .B1_f (new_AGEMA_signal_1920), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_2_U1_Y), .Z0_f (new_AGEMA_signal_2487), .Z1_t (new_AGEMA_signal_2488), .Z1_f (new_AGEMA_signal_2489) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_2_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_2_U1_Y), .A0_f (new_AGEMA_signal_2487), .A1_t (new_AGEMA_signal_2488), .A1_f (new_AGEMA_signal_2489), .B0_t (IN_key_s0_t[66]), .B0_f (IN_key_s0_f[66]), .B1_t (IN_key_s1_t[66]), .B1_f (IN_key_s1_f[66]), .Z0_t (LED_128_Instance_current_roundkey[2]), .Z0_f (new_AGEMA_signal_2680), .Z1_t (new_AGEMA_signal_2681), .Z1_f (new_AGEMA_signal_2682) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_3_U1_XOR1_U1 ( .A0_t (IN_key_s0_t[67]), .A0_f (IN_key_s0_f[67]), .A1_t (IN_key_s1_t[67]), .A1_f (IN_key_s1_f[67]), .B0_t (IN_key_s0_t[3]), .B0_f (IN_key_s0_f[3]), .B1_t (IN_key_s1_t[3]), .B1_f (IN_key_s1_f[3]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_3_U1_X), .Z0_f (new_AGEMA_signal_1927), .Z1_t (new_AGEMA_signal_1928), .Z1_f (new_AGEMA_signal_1929) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_3_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n31), .A1_f (new_AGEMA_signal_2477), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_3_U1_X), .B0_f (new_AGEMA_signal_1927), .B1_t (new_AGEMA_signal_1928), .B1_f (new_AGEMA_signal_1929), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_3_U1_Y), .Z0_f (new_AGEMA_signal_2490), .Z1_t (new_AGEMA_signal_2491), .Z1_f (new_AGEMA_signal_2492) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_3_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_3_U1_Y), .A0_f (new_AGEMA_signal_2490), .A1_t (new_AGEMA_signal_2491), .A1_f (new_AGEMA_signal_2492), .B0_t (IN_key_s0_t[67]), .B0_f (IN_key_s0_f[67]), .B1_t (IN_key_s1_t[67]), .B1_f (IN_key_s1_f[67]), .Z0_t (LED_128_Instance_current_roundkey[3]), .Z0_f (new_AGEMA_signal_2683), .Z1_t (new_AGEMA_signal_2684), .Z1_f (new_AGEMA_signal_2685) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_4_U1_XOR1_U1 ( .A0_t (IN_key_s0_t[68]), .A0_f (IN_key_s0_f[68]), .A1_t (IN_key_s1_t[68]), .A1_f (IN_key_s1_f[68]), .B0_t (IN_key_s0_t[4]), .B0_f (IN_key_s0_f[4]), .B1_t (IN_key_s1_t[4]), .B1_f (IN_key_s1_f[4]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_4_U1_X), .Z0_f (new_AGEMA_signal_1936), .Z1_t (new_AGEMA_signal_1937), .Z1_f (new_AGEMA_signal_1938) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_4_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n31), .A1_f (new_AGEMA_signal_2477), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_4_U1_X), .B0_f (new_AGEMA_signal_1936), .B1_t (new_AGEMA_signal_1937), .B1_f (new_AGEMA_signal_1938), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_4_U1_Y), .Z0_f (new_AGEMA_signal_2493), .Z1_t (new_AGEMA_signal_2494), .Z1_f (new_AGEMA_signal_2495) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_4_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_4_U1_Y), .A0_f (new_AGEMA_signal_2493), .A1_t (new_AGEMA_signal_2494), .A1_f (new_AGEMA_signal_2495), .B0_t (IN_key_s0_t[68]), .B0_f (IN_key_s0_f[68]), .B1_t (IN_key_s1_t[68]), .B1_f (IN_key_s1_f[68]), .Z0_t (LED_128_Instance_current_roundkey[4]), .Z0_f (new_AGEMA_signal_2686), .Z1_t (new_AGEMA_signal_2687), .Z1_f (new_AGEMA_signal_2688) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_5_U1_XOR1_U1 ( .A0_t (IN_key_s0_t[69]), .A0_f (IN_key_s0_f[69]), .A1_t (IN_key_s1_t[69]), .A1_f (IN_key_s1_f[69]), .B0_t (IN_key_s0_t[5]), .B0_f (IN_key_s0_f[5]), .B1_t (IN_key_s1_t[5]), .B1_f (IN_key_s1_f[5]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_5_U1_X), .Z0_f (new_AGEMA_signal_1945), .Z1_t (new_AGEMA_signal_1946), .Z1_f (new_AGEMA_signal_1947) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_5_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n31), .A1_f (new_AGEMA_signal_2477), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_5_U1_X), .B0_f (new_AGEMA_signal_1945), .B1_t (new_AGEMA_signal_1946), .B1_f (new_AGEMA_signal_1947), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_5_U1_Y), .Z0_f (new_AGEMA_signal_2496), .Z1_t (new_AGEMA_signal_2497), .Z1_f (new_AGEMA_signal_2498) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_5_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_5_U1_Y), .A0_f (new_AGEMA_signal_2496), .A1_t (new_AGEMA_signal_2497), .A1_f (new_AGEMA_signal_2498), .B0_t (IN_key_s0_t[69]), .B0_f (IN_key_s0_f[69]), .B1_t (IN_key_s1_t[69]), .B1_f (IN_key_s1_f[69]), .Z0_t (LED_128_Instance_current_roundkey[5]), .Z0_f (new_AGEMA_signal_2689), .Z1_t (new_AGEMA_signal_2690), .Z1_f (new_AGEMA_signal_2691) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_6_U1_XOR1_U1 ( .A0_t (IN_key_s0_t[70]), .A0_f (IN_key_s0_f[70]), .A1_t (IN_key_s1_t[70]), .A1_f (IN_key_s1_f[70]), .B0_t (IN_key_s0_t[6]), .B0_f (IN_key_s0_f[6]), .B1_t (IN_key_s1_t[6]), .B1_f (IN_key_s1_f[6]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_6_U1_X), .Z0_f (new_AGEMA_signal_1954), .Z1_t (new_AGEMA_signal_1955), .Z1_f (new_AGEMA_signal_1956) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_6_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n31), .A1_f (new_AGEMA_signal_2477), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_6_U1_X), .B0_f (new_AGEMA_signal_1954), .B1_t (new_AGEMA_signal_1955), .B1_f (new_AGEMA_signal_1956), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_6_U1_Y), .Z0_f (new_AGEMA_signal_2499), .Z1_t (new_AGEMA_signal_2500), .Z1_f (new_AGEMA_signal_2501) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_6_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_6_U1_Y), .A0_f (new_AGEMA_signal_2499), .A1_t (new_AGEMA_signal_2500), .A1_f (new_AGEMA_signal_2501), .B0_t (IN_key_s0_t[70]), .B0_f (IN_key_s0_f[70]), .B1_t (IN_key_s1_t[70]), .B1_f (IN_key_s1_f[70]), .Z0_t (LED_128_Instance_current_roundkey[6]), .Z0_f (new_AGEMA_signal_2692), .Z1_t (new_AGEMA_signal_2693), .Z1_f (new_AGEMA_signal_2694) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_7_U1_XOR1_U1 ( .A0_t (IN_key_s0_t[71]), .A0_f (IN_key_s0_f[71]), .A1_t (IN_key_s1_t[71]), .A1_f (IN_key_s1_f[71]), .B0_t (IN_key_s0_t[7]), .B0_f (IN_key_s0_f[7]), .B1_t (IN_key_s1_t[7]), .B1_f (IN_key_s1_f[7]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_7_U1_X), .Z0_f (new_AGEMA_signal_1963), .Z1_t (new_AGEMA_signal_1964), .Z1_f (new_AGEMA_signal_1965) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_7_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n31), .A1_f (new_AGEMA_signal_2477), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_7_U1_X), .B0_f (new_AGEMA_signal_1963), .B1_t (new_AGEMA_signal_1964), .B1_f (new_AGEMA_signal_1965), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_7_U1_Y), .Z0_f (new_AGEMA_signal_2502), .Z1_t (new_AGEMA_signal_2503), .Z1_f (new_AGEMA_signal_2504) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_7_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_7_U1_Y), .A0_f (new_AGEMA_signal_2502), .A1_t (new_AGEMA_signal_2503), .A1_f (new_AGEMA_signal_2504), .B0_t (IN_key_s0_t[71]), .B0_f (IN_key_s0_f[71]), .B1_t (IN_key_s1_t[71]), .B1_f (IN_key_s1_f[71]), .Z0_t (LED_128_Instance_current_roundkey[7]), .Z0_f (new_AGEMA_signal_2695), .Z1_t (new_AGEMA_signal_2696), .Z1_f (new_AGEMA_signal_2697) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_8_U1_XOR1_U1 ( .A0_t (IN_key_s0_t[72]), .A0_f (IN_key_s0_f[72]), .A1_t (IN_key_s1_t[72]), .A1_f (IN_key_s1_f[72]), .B0_t (IN_key_s0_t[8]), .B0_f (IN_key_s0_f[8]), .B1_t (IN_key_s1_t[8]), .B1_f (IN_key_s1_f[8]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_8_U1_X), .Z0_f (new_AGEMA_signal_1972), .Z1_t (new_AGEMA_signal_1973), .Z1_f (new_AGEMA_signal_1974) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_8_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n31), .A1_f (new_AGEMA_signal_2477), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_8_U1_X), .B0_f (new_AGEMA_signal_1972), .B1_t (new_AGEMA_signal_1973), .B1_f (new_AGEMA_signal_1974), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_8_U1_Y), .Z0_f (new_AGEMA_signal_2505), .Z1_t (new_AGEMA_signal_2506), .Z1_f (new_AGEMA_signal_2507) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_8_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_8_U1_Y), .A0_f (new_AGEMA_signal_2505), .A1_t (new_AGEMA_signal_2506), .A1_f (new_AGEMA_signal_2507), .B0_t (IN_key_s0_t[72]), .B0_f (IN_key_s0_f[72]), .B1_t (IN_key_s1_t[72]), .B1_f (IN_key_s1_f[72]), .Z0_t (LED_128_Instance_current_roundkey[8]), .Z0_f (new_AGEMA_signal_2698), .Z1_t (new_AGEMA_signal_2699), .Z1_f (new_AGEMA_signal_2700) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_9_U1_XOR1_U1 ( .A0_t (IN_key_s0_t[73]), .A0_f (IN_key_s0_f[73]), .A1_t (IN_key_s1_t[73]), .A1_f (IN_key_s1_f[73]), .B0_t (IN_key_s0_t[9]), .B0_f (IN_key_s0_f[9]), .B1_t (IN_key_s1_t[9]), .B1_f (IN_key_s1_f[9]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_9_U1_X), .Z0_f (new_AGEMA_signal_1981), .Z1_t (new_AGEMA_signal_1982), .Z1_f (new_AGEMA_signal_1983) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_9_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n31), .A1_f (new_AGEMA_signal_2477), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_9_U1_X), .B0_f (new_AGEMA_signal_1981), .B1_t (new_AGEMA_signal_1982), .B1_f (new_AGEMA_signal_1983), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_9_U1_Y), .Z0_f (new_AGEMA_signal_2508), .Z1_t (new_AGEMA_signal_2509), .Z1_f (new_AGEMA_signal_2510) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_9_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_9_U1_Y), .A0_f (new_AGEMA_signal_2508), .A1_t (new_AGEMA_signal_2509), .A1_f (new_AGEMA_signal_2510), .B0_t (IN_key_s0_t[73]), .B0_f (IN_key_s0_f[73]), .B1_t (IN_key_s1_t[73]), .B1_f (IN_key_s1_f[73]), .Z0_t (LED_128_Instance_current_roundkey[9]), .Z0_f (new_AGEMA_signal_2701), .Z1_t (new_AGEMA_signal_2702), .Z1_f (new_AGEMA_signal_2703) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_10_U1_XOR1_U1 ( .A0_t (IN_key_s0_t[74]), .A0_f (IN_key_s0_f[74]), .A1_t (IN_key_s1_t[74]), .A1_f (IN_key_s1_f[74]), .B0_t (IN_key_s0_t[10]), .B0_f (IN_key_s0_f[10]), .B1_t (IN_key_s1_t[10]), .B1_f (IN_key_s1_f[10]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_10_U1_X), .Z0_f (new_AGEMA_signal_1990), .Z1_t (new_AGEMA_signal_1991), .Z1_f (new_AGEMA_signal_1992) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_10_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n31), .A1_f (new_AGEMA_signal_2477), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_10_U1_X), .B0_f (new_AGEMA_signal_1990), .B1_t (new_AGEMA_signal_1991), .B1_f (new_AGEMA_signal_1992), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_10_U1_Y), .Z0_f (new_AGEMA_signal_2511), .Z1_t (new_AGEMA_signal_2512), .Z1_f (new_AGEMA_signal_2513) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_10_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_10_U1_Y), .A0_f (new_AGEMA_signal_2511), .A1_t (new_AGEMA_signal_2512), .A1_f (new_AGEMA_signal_2513), .B0_t (IN_key_s0_t[74]), .B0_f (IN_key_s0_f[74]), .B1_t (IN_key_s1_t[74]), .B1_f (IN_key_s1_f[74]), .Z0_t (LED_128_Instance_current_roundkey[10]), .Z0_f (new_AGEMA_signal_2704), .Z1_t (new_AGEMA_signal_2705), .Z1_f (new_AGEMA_signal_2706) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_11_U1_XOR1_U1 ( .A0_t (IN_key_s0_t[75]), .A0_f (IN_key_s0_f[75]), .A1_t (IN_key_s1_t[75]), .A1_f (IN_key_s1_f[75]), .B0_t (IN_key_s0_t[11]), .B0_f (IN_key_s0_f[11]), .B1_t (IN_key_s1_t[11]), .B1_f (IN_key_s1_f[11]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_11_U1_X), .Z0_f (new_AGEMA_signal_1999), .Z1_t (new_AGEMA_signal_2000), .Z1_f (new_AGEMA_signal_2001) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_11_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n31), .A1_f (new_AGEMA_signal_2477), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_11_U1_X), .B0_f (new_AGEMA_signal_1999), .B1_t (new_AGEMA_signal_2000), .B1_f (new_AGEMA_signal_2001), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_11_U1_Y), .Z0_f (new_AGEMA_signal_2514), .Z1_t (new_AGEMA_signal_2515), .Z1_f (new_AGEMA_signal_2516) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_11_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_11_U1_Y), .A0_f (new_AGEMA_signal_2514), .A1_t (new_AGEMA_signal_2515), .A1_f (new_AGEMA_signal_2516), .B0_t (IN_key_s0_t[75]), .B0_f (IN_key_s0_f[75]), .B1_t (IN_key_s1_t[75]), .B1_f (IN_key_s1_f[75]), .Z0_t (LED_128_Instance_current_roundkey[11]), .Z0_f (new_AGEMA_signal_2707), .Z1_t (new_AGEMA_signal_2708), .Z1_f (new_AGEMA_signal_2709) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_12_U1_XOR1_U1 ( .A0_t (IN_key_s0_t[76]), .A0_f (IN_key_s0_f[76]), .A1_t (IN_key_s1_t[76]), .A1_f (IN_key_s1_f[76]), .B0_t (IN_key_s0_t[12]), .B0_f (IN_key_s0_f[12]), .B1_t (IN_key_s1_t[12]), .B1_f (IN_key_s1_f[12]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_12_U1_X), .Z0_f (new_AGEMA_signal_2008), .Z1_t (new_AGEMA_signal_2009), .Z1_f (new_AGEMA_signal_2010) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_12_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n31), .A1_f (new_AGEMA_signal_2477), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_12_U1_X), .B0_f (new_AGEMA_signal_2008), .B1_t (new_AGEMA_signal_2009), .B1_f (new_AGEMA_signal_2010), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_12_U1_Y), .Z0_f (new_AGEMA_signal_2517), .Z1_t (new_AGEMA_signal_2518), .Z1_f (new_AGEMA_signal_2519) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_12_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_12_U1_Y), .A0_f (new_AGEMA_signal_2517), .A1_t (new_AGEMA_signal_2518), .A1_f (new_AGEMA_signal_2519), .B0_t (IN_key_s0_t[76]), .B0_f (IN_key_s0_f[76]), .B1_t (IN_key_s1_t[76]), .B1_f (IN_key_s1_f[76]), .Z0_t (LED_128_Instance_current_roundkey[12]), .Z0_f (new_AGEMA_signal_2710), .Z1_t (new_AGEMA_signal_2711), .Z1_f (new_AGEMA_signal_2712) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_13_U1_XOR1_U1 ( .A0_t (IN_key_s0_t[77]), .A0_f (IN_key_s0_f[77]), .A1_t (IN_key_s1_t[77]), .A1_f (IN_key_s1_f[77]), .B0_t (IN_key_s0_t[13]), .B0_f (IN_key_s0_f[13]), .B1_t (IN_key_s1_t[13]), .B1_f (IN_key_s1_f[13]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_13_U1_X), .Z0_f (new_AGEMA_signal_2017), .Z1_t (new_AGEMA_signal_2018), .Z1_f (new_AGEMA_signal_2019) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_13_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n31), .A1_f (new_AGEMA_signal_2477), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_13_U1_X), .B0_f (new_AGEMA_signal_2017), .B1_t (new_AGEMA_signal_2018), .B1_f (new_AGEMA_signal_2019), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_13_U1_Y), .Z0_f (new_AGEMA_signal_2520), .Z1_t (new_AGEMA_signal_2521), .Z1_f (new_AGEMA_signal_2522) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_13_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_13_U1_Y), .A0_f (new_AGEMA_signal_2520), .A1_t (new_AGEMA_signal_2521), .A1_f (new_AGEMA_signal_2522), .B0_t (IN_key_s0_t[77]), .B0_f (IN_key_s0_f[77]), .B1_t (IN_key_s1_t[77]), .B1_f (IN_key_s1_f[77]), .Z0_t (LED_128_Instance_current_roundkey[13]), .Z0_f (new_AGEMA_signal_2713), .Z1_t (new_AGEMA_signal_2714), .Z1_f (new_AGEMA_signal_2715) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_14_U1_XOR1_U1 ( .A0_t (IN_key_s0_t[78]), .A0_f (IN_key_s0_f[78]), .A1_t (IN_key_s1_t[78]), .A1_f (IN_key_s1_f[78]), .B0_t (IN_key_s0_t[14]), .B0_f (IN_key_s0_f[14]), .B1_t (IN_key_s1_t[14]), .B1_f (IN_key_s1_f[14]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_14_U1_X), .Z0_f (new_AGEMA_signal_2026), .Z1_t (new_AGEMA_signal_2027), .Z1_f (new_AGEMA_signal_2028) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_14_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n31), .A1_f (new_AGEMA_signal_2477), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_14_U1_X), .B0_f (new_AGEMA_signal_2026), .B1_t (new_AGEMA_signal_2027), .B1_f (new_AGEMA_signal_2028), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_14_U1_Y), .Z0_f (new_AGEMA_signal_2523), .Z1_t (new_AGEMA_signal_2524), .Z1_f (new_AGEMA_signal_2525) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_14_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_14_U1_Y), .A0_f (new_AGEMA_signal_2523), .A1_t (new_AGEMA_signal_2524), .A1_f (new_AGEMA_signal_2525), .B0_t (IN_key_s0_t[78]), .B0_f (IN_key_s0_f[78]), .B1_t (IN_key_s1_t[78]), .B1_f (IN_key_s1_f[78]), .Z0_t (LED_128_Instance_current_roundkey[14]), .Z0_f (new_AGEMA_signal_2716), .Z1_t (new_AGEMA_signal_2717), .Z1_f (new_AGEMA_signal_2718) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_15_U1_XOR1_U1 ( .A0_t (IN_key_s0_t[79]), .A0_f (IN_key_s0_f[79]), .A1_t (IN_key_s1_t[79]), .A1_f (IN_key_s1_f[79]), .B0_t (IN_key_s0_t[15]), .B0_f (IN_key_s0_f[15]), .B1_t (IN_key_s1_t[15]), .B1_f (IN_key_s1_f[15]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_15_U1_X), .Z0_f (new_AGEMA_signal_2035), .Z1_t (new_AGEMA_signal_2036), .Z1_f (new_AGEMA_signal_2037) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_15_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n31), .A1_f (new_AGEMA_signal_2477), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_15_U1_X), .B0_f (new_AGEMA_signal_2035), .B1_t (new_AGEMA_signal_2036), .B1_f (new_AGEMA_signal_2037), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_15_U1_Y), .Z0_f (new_AGEMA_signal_2526), .Z1_t (new_AGEMA_signal_2527), .Z1_f (new_AGEMA_signal_2528) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_15_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_15_U1_Y), .A0_f (new_AGEMA_signal_2526), .A1_t (new_AGEMA_signal_2527), .A1_f (new_AGEMA_signal_2528), .B0_t (IN_key_s0_t[79]), .B0_f (IN_key_s0_f[79]), .B1_t (IN_key_s1_t[79]), .B1_f (IN_key_s1_f[79]), .Z0_t (LED_128_Instance_current_roundkey[15]), .Z0_f (new_AGEMA_signal_2719), .Z1_t (new_AGEMA_signal_2720), .Z1_f (new_AGEMA_signal_2721) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_16_U1_XOR1_U1 ( .A0_t (IN_key_s0_t[80]), .A0_f (IN_key_s0_f[80]), .A1_t (IN_key_s1_t[80]), .A1_f (IN_key_s1_f[80]), .B0_t (IN_key_s0_t[16]), .B0_f (IN_key_s0_f[16]), .B1_t (IN_key_s1_t[16]), .B1_f (IN_key_s1_f[16]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_16_U1_X), .Z0_f (new_AGEMA_signal_2044), .Z1_t (new_AGEMA_signal_2045), .Z1_f (new_AGEMA_signal_2046) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_16_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n31), .A1_f (new_AGEMA_signal_2477), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_16_U1_X), .B0_f (new_AGEMA_signal_2044), .B1_t (new_AGEMA_signal_2045), .B1_f (new_AGEMA_signal_2046), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_16_U1_Y), .Z0_f (new_AGEMA_signal_2529), .Z1_t (new_AGEMA_signal_2530), .Z1_f (new_AGEMA_signal_2531) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_16_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_16_U1_Y), .A0_f (new_AGEMA_signal_2529), .A1_t (new_AGEMA_signal_2530), .A1_f (new_AGEMA_signal_2531), .B0_t (IN_key_s0_t[80]), .B0_f (IN_key_s0_f[80]), .B1_t (IN_key_s1_t[80]), .B1_f (IN_key_s1_f[80]), .Z0_t (LED_128_Instance_current_roundkey[16]), .Z0_f (new_AGEMA_signal_2722), .Z1_t (new_AGEMA_signal_2723), .Z1_f (new_AGEMA_signal_2724) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_17_U1_XOR1_U1 ( .A0_t (IN_key_s0_t[81]), .A0_f (IN_key_s0_f[81]), .A1_t (IN_key_s1_t[81]), .A1_f (IN_key_s1_f[81]), .B0_t (IN_key_s0_t[17]), .B0_f (IN_key_s0_f[17]), .B1_t (IN_key_s1_t[17]), .B1_f (IN_key_s1_f[17]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_17_U1_X), .Z0_f (new_AGEMA_signal_2053), .Z1_t (new_AGEMA_signal_2054), .Z1_f (new_AGEMA_signal_2055) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_17_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n31), .A1_f (new_AGEMA_signal_2477), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_17_U1_X), .B0_f (new_AGEMA_signal_2053), .B1_t (new_AGEMA_signal_2054), .B1_f (new_AGEMA_signal_2055), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_17_U1_Y), .Z0_f (new_AGEMA_signal_2532), .Z1_t (new_AGEMA_signal_2533), .Z1_f (new_AGEMA_signal_2534) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_17_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_17_U1_Y), .A0_f (new_AGEMA_signal_2532), .A1_t (new_AGEMA_signal_2533), .A1_f (new_AGEMA_signal_2534), .B0_t (IN_key_s0_t[81]), .B0_f (IN_key_s0_f[81]), .B1_t (IN_key_s1_t[81]), .B1_f (IN_key_s1_f[81]), .Z0_t (LED_128_Instance_current_roundkey[17]), .Z0_f (new_AGEMA_signal_2725), .Z1_t (new_AGEMA_signal_2726), .Z1_f (new_AGEMA_signal_2727) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_18_U1_XOR1_U1 ( .A0_t (IN_key_s0_t[82]), .A0_f (IN_key_s0_f[82]), .A1_t (IN_key_s1_t[82]), .A1_f (IN_key_s1_f[82]), .B0_t (IN_key_s0_t[18]), .B0_f (IN_key_s0_f[18]), .B1_t (IN_key_s1_t[18]), .B1_f (IN_key_s1_f[18]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_18_U1_X), .Z0_f (new_AGEMA_signal_2062), .Z1_t (new_AGEMA_signal_2063), .Z1_f (new_AGEMA_signal_2064) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_18_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n31), .A1_f (new_AGEMA_signal_2477), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_18_U1_X), .B0_f (new_AGEMA_signal_2062), .B1_t (new_AGEMA_signal_2063), .B1_f (new_AGEMA_signal_2064), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_18_U1_Y), .Z0_f (new_AGEMA_signal_2535), .Z1_t (new_AGEMA_signal_2536), .Z1_f (new_AGEMA_signal_2537) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_18_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_18_U1_Y), .A0_f (new_AGEMA_signal_2535), .A1_t (new_AGEMA_signal_2536), .A1_f (new_AGEMA_signal_2537), .B0_t (IN_key_s0_t[82]), .B0_f (IN_key_s0_f[82]), .B1_t (IN_key_s1_t[82]), .B1_f (IN_key_s1_f[82]), .Z0_t (LED_128_Instance_current_roundkey[18]), .Z0_f (new_AGEMA_signal_2728), .Z1_t (new_AGEMA_signal_2729), .Z1_f (new_AGEMA_signal_2730) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_19_U1_XOR1_U1 ( .A0_t (IN_key_s0_t[83]), .A0_f (IN_key_s0_f[83]), .A1_t (IN_key_s1_t[83]), .A1_f (IN_key_s1_f[83]), .B0_t (IN_key_s0_t[19]), .B0_f (IN_key_s0_f[19]), .B1_t (IN_key_s1_t[19]), .B1_f (IN_key_s1_f[19]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_19_U1_X), .Z0_f (new_AGEMA_signal_2071), .Z1_t (new_AGEMA_signal_2072), .Z1_f (new_AGEMA_signal_2073) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_19_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n31), .A1_f (new_AGEMA_signal_2477), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_19_U1_X), .B0_f (new_AGEMA_signal_2071), .B1_t (new_AGEMA_signal_2072), .B1_f (new_AGEMA_signal_2073), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_19_U1_Y), .Z0_f (new_AGEMA_signal_2538), .Z1_t (new_AGEMA_signal_2539), .Z1_f (new_AGEMA_signal_2540) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_19_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_19_U1_Y), .A0_f (new_AGEMA_signal_2538), .A1_t (new_AGEMA_signal_2539), .A1_f (new_AGEMA_signal_2540), .B0_t (IN_key_s0_t[83]), .B0_f (IN_key_s0_f[83]), .B1_t (IN_key_s1_t[83]), .B1_f (IN_key_s1_f[83]), .Z0_t (LED_128_Instance_current_roundkey[19]), .Z0_f (new_AGEMA_signal_2731), .Z1_t (new_AGEMA_signal_2732), .Z1_f (new_AGEMA_signal_2733) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_20_U1_XOR1_U1 ( .A0_t (IN_key_s0_t[84]), .A0_f (IN_key_s0_f[84]), .A1_t (IN_key_s1_t[84]), .A1_f (IN_key_s1_f[84]), .B0_t (IN_key_s0_t[20]), .B0_f (IN_key_s0_f[20]), .B1_t (IN_key_s1_t[20]), .B1_f (IN_key_s1_f[20]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_20_U1_X), .Z0_f (new_AGEMA_signal_2080), .Z1_t (new_AGEMA_signal_2081), .Z1_f (new_AGEMA_signal_2082) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_20_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n31), .A1_f (new_AGEMA_signal_2477), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_20_U1_X), .B0_f (new_AGEMA_signal_2080), .B1_t (new_AGEMA_signal_2081), .B1_f (new_AGEMA_signal_2082), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_20_U1_Y), .Z0_f (new_AGEMA_signal_2541), .Z1_t (new_AGEMA_signal_2542), .Z1_f (new_AGEMA_signal_2543) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_20_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_20_U1_Y), .A0_f (new_AGEMA_signal_2541), .A1_t (new_AGEMA_signal_2542), .A1_f (new_AGEMA_signal_2543), .B0_t (IN_key_s0_t[84]), .B0_f (IN_key_s0_f[84]), .B1_t (IN_key_s1_t[84]), .B1_f (IN_key_s1_f[84]), .Z0_t (LED_128_Instance_current_roundkey[20]), .Z0_f (new_AGEMA_signal_2734), .Z1_t (new_AGEMA_signal_2735), .Z1_f (new_AGEMA_signal_2736) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_21_U1_XOR1_U1 ( .A0_t (IN_key_s0_t[85]), .A0_f (IN_key_s0_f[85]), .A1_t (IN_key_s1_t[85]), .A1_f (IN_key_s1_f[85]), .B0_t (IN_key_s0_t[21]), .B0_f (IN_key_s0_f[21]), .B1_t (IN_key_s1_t[21]), .B1_f (IN_key_s1_f[21]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_21_U1_X), .Z0_f (new_AGEMA_signal_2089), .Z1_t (new_AGEMA_signal_2090), .Z1_f (new_AGEMA_signal_2091) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_21_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n31), .A1_f (new_AGEMA_signal_2477), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_21_U1_X), .B0_f (new_AGEMA_signal_2089), .B1_t (new_AGEMA_signal_2090), .B1_f (new_AGEMA_signal_2091), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_21_U1_Y), .Z0_f (new_AGEMA_signal_2544), .Z1_t (new_AGEMA_signal_2545), .Z1_f (new_AGEMA_signal_2546) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_21_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_21_U1_Y), .A0_f (new_AGEMA_signal_2544), .A1_t (new_AGEMA_signal_2545), .A1_f (new_AGEMA_signal_2546), .B0_t (IN_key_s0_t[85]), .B0_f (IN_key_s0_f[85]), .B1_t (IN_key_s1_t[85]), .B1_f (IN_key_s1_f[85]), .Z0_t (LED_128_Instance_current_roundkey[21]), .Z0_f (new_AGEMA_signal_2737), .Z1_t (new_AGEMA_signal_2738), .Z1_f (new_AGEMA_signal_2739) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_22_U1_XOR1_U1 ( .A0_t (IN_key_s0_t[86]), .A0_f (IN_key_s0_f[86]), .A1_t (IN_key_s1_t[86]), .A1_f (IN_key_s1_f[86]), .B0_t (IN_key_s0_t[22]), .B0_f (IN_key_s0_f[22]), .B1_t (IN_key_s1_t[22]), .B1_f (IN_key_s1_f[22]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_22_U1_X), .Z0_f (new_AGEMA_signal_2098), .Z1_t (new_AGEMA_signal_2099), .Z1_f (new_AGEMA_signal_2100) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_22_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n31), .A1_f (new_AGEMA_signal_2477), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_22_U1_X), .B0_f (new_AGEMA_signal_2098), .B1_t (new_AGEMA_signal_2099), .B1_f (new_AGEMA_signal_2100), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_22_U1_Y), .Z0_f (new_AGEMA_signal_2547), .Z1_t (new_AGEMA_signal_2548), .Z1_f (new_AGEMA_signal_2549) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_22_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_22_U1_Y), .A0_f (new_AGEMA_signal_2547), .A1_t (new_AGEMA_signal_2548), .A1_f (new_AGEMA_signal_2549), .B0_t (IN_key_s0_t[86]), .B0_f (IN_key_s0_f[86]), .B1_t (IN_key_s1_t[86]), .B1_f (IN_key_s1_f[86]), .Z0_t (LED_128_Instance_current_roundkey[22]), .Z0_f (new_AGEMA_signal_2740), .Z1_t (new_AGEMA_signal_2741), .Z1_f (new_AGEMA_signal_2742) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_23_U1_XOR1_U1 ( .A0_t (IN_key_s0_t[87]), .A0_f (IN_key_s0_f[87]), .A1_t (IN_key_s1_t[87]), .A1_f (IN_key_s1_f[87]), .B0_t (IN_key_s0_t[23]), .B0_f (IN_key_s0_f[23]), .B1_t (IN_key_s1_t[23]), .B1_f (IN_key_s1_f[23]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_23_U1_X), .Z0_f (new_AGEMA_signal_2107), .Z1_t (new_AGEMA_signal_2108), .Z1_f (new_AGEMA_signal_2109) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_23_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n31), .A1_f (new_AGEMA_signal_2477), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_23_U1_X), .B0_f (new_AGEMA_signal_2107), .B1_t (new_AGEMA_signal_2108), .B1_f (new_AGEMA_signal_2109), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_23_U1_Y), .Z0_f (new_AGEMA_signal_2550), .Z1_t (new_AGEMA_signal_2551), .Z1_f (new_AGEMA_signal_2552) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_23_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_23_U1_Y), .A0_f (new_AGEMA_signal_2550), .A1_t (new_AGEMA_signal_2551), .A1_f (new_AGEMA_signal_2552), .B0_t (IN_key_s0_t[87]), .B0_f (IN_key_s0_f[87]), .B1_t (IN_key_s1_t[87]), .B1_f (IN_key_s1_f[87]), .Z0_t (LED_128_Instance_current_roundkey[23]), .Z0_f (new_AGEMA_signal_2743), .Z1_t (new_AGEMA_signal_2744), .Z1_f (new_AGEMA_signal_2745) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_24_U1_XOR1_U1 ( .A0_t (IN_key_s0_t[88]), .A0_f (IN_key_s0_f[88]), .A1_t (IN_key_s1_t[88]), .A1_f (IN_key_s1_f[88]), .B0_t (IN_key_s0_t[24]), .B0_f (IN_key_s0_f[24]), .B1_t (IN_key_s1_t[24]), .B1_f (IN_key_s1_f[24]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_24_U1_X), .Z0_f (new_AGEMA_signal_2116), .Z1_t (new_AGEMA_signal_2117), .Z1_f (new_AGEMA_signal_2118) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_24_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n31), .A1_f (new_AGEMA_signal_2477), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_24_U1_X), .B0_f (new_AGEMA_signal_2116), .B1_t (new_AGEMA_signal_2117), .B1_f (new_AGEMA_signal_2118), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_24_U1_Y), .Z0_f (new_AGEMA_signal_2553), .Z1_t (new_AGEMA_signal_2554), .Z1_f (new_AGEMA_signal_2555) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_24_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_24_U1_Y), .A0_f (new_AGEMA_signal_2553), .A1_t (new_AGEMA_signal_2554), .A1_f (new_AGEMA_signal_2555), .B0_t (IN_key_s0_t[88]), .B0_f (IN_key_s0_f[88]), .B1_t (IN_key_s1_t[88]), .B1_f (IN_key_s1_f[88]), .Z0_t (LED_128_Instance_current_roundkey[24]), .Z0_f (new_AGEMA_signal_2746), .Z1_t (new_AGEMA_signal_2747), .Z1_f (new_AGEMA_signal_2748) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_25_U1_XOR1_U1 ( .A0_t (IN_key_s0_t[89]), .A0_f (IN_key_s0_f[89]), .A1_t (IN_key_s1_t[89]), .A1_f (IN_key_s1_f[89]), .B0_t (IN_key_s0_t[25]), .B0_f (IN_key_s0_f[25]), .B1_t (IN_key_s1_t[25]), .B1_f (IN_key_s1_f[25]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_25_U1_X), .Z0_f (new_AGEMA_signal_2125), .Z1_t (new_AGEMA_signal_2126), .Z1_f (new_AGEMA_signal_2127) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_25_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n31), .A1_f (new_AGEMA_signal_2477), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_25_U1_X), .B0_f (new_AGEMA_signal_2125), .B1_t (new_AGEMA_signal_2126), .B1_f (new_AGEMA_signal_2127), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_25_U1_Y), .Z0_f (new_AGEMA_signal_2556), .Z1_t (new_AGEMA_signal_2557), .Z1_f (new_AGEMA_signal_2558) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_25_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_25_U1_Y), .A0_f (new_AGEMA_signal_2556), .A1_t (new_AGEMA_signal_2557), .A1_f (new_AGEMA_signal_2558), .B0_t (IN_key_s0_t[89]), .B0_f (IN_key_s0_f[89]), .B1_t (IN_key_s1_t[89]), .B1_f (IN_key_s1_f[89]), .Z0_t (LED_128_Instance_current_roundkey[25]), .Z0_f (new_AGEMA_signal_2749), .Z1_t (new_AGEMA_signal_2750), .Z1_f (new_AGEMA_signal_2751) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_26_U1_XOR1_U1 ( .A0_t (IN_key_s0_t[90]), .A0_f (IN_key_s0_f[90]), .A1_t (IN_key_s1_t[90]), .A1_f (IN_key_s1_f[90]), .B0_t (IN_key_s0_t[26]), .B0_f (IN_key_s0_f[26]), .B1_t (IN_key_s1_t[26]), .B1_f (IN_key_s1_f[26]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_26_U1_X), .Z0_f (new_AGEMA_signal_2134), .Z1_t (new_AGEMA_signal_2135), .Z1_f (new_AGEMA_signal_2136) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_26_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n31), .A1_f (new_AGEMA_signal_2477), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_26_U1_X), .B0_f (new_AGEMA_signal_2134), .B1_t (new_AGEMA_signal_2135), .B1_f (new_AGEMA_signal_2136), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_26_U1_Y), .Z0_f (new_AGEMA_signal_2559), .Z1_t (new_AGEMA_signal_2560), .Z1_f (new_AGEMA_signal_2561) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_26_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_26_U1_Y), .A0_f (new_AGEMA_signal_2559), .A1_t (new_AGEMA_signal_2560), .A1_f (new_AGEMA_signal_2561), .B0_t (IN_key_s0_t[90]), .B0_f (IN_key_s0_f[90]), .B1_t (IN_key_s1_t[90]), .B1_f (IN_key_s1_f[90]), .Z0_t (LED_128_Instance_current_roundkey[26]), .Z0_f (new_AGEMA_signal_2752), .Z1_t (new_AGEMA_signal_2753), .Z1_f (new_AGEMA_signal_2754) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_27_U1_XOR1_U1 ( .A0_t (IN_key_s0_t[91]), .A0_f (IN_key_s0_f[91]), .A1_t (IN_key_s1_t[91]), .A1_f (IN_key_s1_f[91]), .B0_t (IN_key_s0_t[27]), .B0_f (IN_key_s0_f[27]), .B1_t (IN_key_s1_t[27]), .B1_f (IN_key_s1_f[27]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_27_U1_X), .Z0_f (new_AGEMA_signal_2143), .Z1_t (new_AGEMA_signal_2144), .Z1_f (new_AGEMA_signal_2145) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_27_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n31), .A1_f (new_AGEMA_signal_2477), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_27_U1_X), .B0_f (new_AGEMA_signal_2143), .B1_t (new_AGEMA_signal_2144), .B1_f (new_AGEMA_signal_2145), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_27_U1_Y), .Z0_f (new_AGEMA_signal_2562), .Z1_t (new_AGEMA_signal_2563), .Z1_f (new_AGEMA_signal_2564) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_27_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_27_U1_Y), .A0_f (new_AGEMA_signal_2562), .A1_t (new_AGEMA_signal_2563), .A1_f (new_AGEMA_signal_2564), .B0_t (IN_key_s0_t[91]), .B0_f (IN_key_s0_f[91]), .B1_t (IN_key_s1_t[91]), .B1_f (IN_key_s1_f[91]), .Z0_t (LED_128_Instance_current_roundkey[27]), .Z0_f (new_AGEMA_signal_2755), .Z1_t (new_AGEMA_signal_2756), .Z1_f (new_AGEMA_signal_2757) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_28_U1_XOR1_U1 ( .A0_t (IN_key_s0_t[92]), .A0_f (IN_key_s0_f[92]), .A1_t (IN_key_s1_t[92]), .A1_f (IN_key_s1_f[92]), .B0_t (IN_key_s0_t[28]), .B0_f (IN_key_s0_f[28]), .B1_t (IN_key_s1_t[28]), .B1_f (IN_key_s1_f[28]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_28_U1_X), .Z0_f (new_AGEMA_signal_2152), .Z1_t (new_AGEMA_signal_2153), .Z1_f (new_AGEMA_signal_2154) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_28_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n31), .A1_f (new_AGEMA_signal_2477), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_28_U1_X), .B0_f (new_AGEMA_signal_2152), .B1_t (new_AGEMA_signal_2153), .B1_f (new_AGEMA_signal_2154), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_28_U1_Y), .Z0_f (new_AGEMA_signal_2565), .Z1_t (new_AGEMA_signal_2566), .Z1_f (new_AGEMA_signal_2567) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_28_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_28_U1_Y), .A0_f (new_AGEMA_signal_2565), .A1_t (new_AGEMA_signal_2566), .A1_f (new_AGEMA_signal_2567), .B0_t (IN_key_s0_t[92]), .B0_f (IN_key_s0_f[92]), .B1_t (IN_key_s1_t[92]), .B1_f (IN_key_s1_f[92]), .Z0_t (LED_128_Instance_current_roundkey[28]), .Z0_f (new_AGEMA_signal_2758), .Z1_t (new_AGEMA_signal_2759), .Z1_f (new_AGEMA_signal_2760) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_29_U1_XOR1_U1 ( .A0_t (IN_key_s0_t[93]), .A0_f (IN_key_s0_f[93]), .A1_t (IN_key_s1_t[93]), .A1_f (IN_key_s1_f[93]), .B0_t (IN_key_s0_t[29]), .B0_f (IN_key_s0_f[29]), .B1_t (IN_key_s1_t[29]), .B1_f (IN_key_s1_f[29]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_29_U1_X), .Z0_f (new_AGEMA_signal_2161), .Z1_t (new_AGEMA_signal_2162), .Z1_f (new_AGEMA_signal_2163) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_29_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n31), .A1_f (new_AGEMA_signal_2477), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_29_U1_X), .B0_f (new_AGEMA_signal_2161), .B1_t (new_AGEMA_signal_2162), .B1_f (new_AGEMA_signal_2163), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_29_U1_Y), .Z0_f (new_AGEMA_signal_2568), .Z1_t (new_AGEMA_signal_2569), .Z1_f (new_AGEMA_signal_2570) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_29_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_29_U1_Y), .A0_f (new_AGEMA_signal_2568), .A1_t (new_AGEMA_signal_2569), .A1_f (new_AGEMA_signal_2570), .B0_t (IN_key_s0_t[93]), .B0_f (IN_key_s0_f[93]), .B1_t (IN_key_s1_t[93]), .B1_f (IN_key_s1_f[93]), .Z0_t (LED_128_Instance_current_roundkey[29]), .Z0_f (new_AGEMA_signal_2761), .Z1_t (new_AGEMA_signal_2762), .Z1_f (new_AGEMA_signal_2763) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_30_U1_XOR1_U1 ( .A0_t (IN_key_s0_t[94]), .A0_f (IN_key_s0_f[94]), .A1_t (IN_key_s1_t[94]), .A1_f (IN_key_s1_f[94]), .B0_t (IN_key_s0_t[30]), .B0_f (IN_key_s0_f[30]), .B1_t (IN_key_s1_t[30]), .B1_f (IN_key_s1_f[30]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_30_U1_X), .Z0_f (new_AGEMA_signal_2170), .Z1_t (new_AGEMA_signal_2171), .Z1_f (new_AGEMA_signal_2172) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_30_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n31), .A1_f (new_AGEMA_signal_2477), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_30_U1_X), .B0_f (new_AGEMA_signal_2170), .B1_t (new_AGEMA_signal_2171), .B1_f (new_AGEMA_signal_2172), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_30_U1_Y), .Z0_f (new_AGEMA_signal_2571), .Z1_t (new_AGEMA_signal_2572), .Z1_f (new_AGEMA_signal_2573) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_30_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_30_U1_Y), .A0_f (new_AGEMA_signal_2571), .A1_t (new_AGEMA_signal_2572), .A1_f (new_AGEMA_signal_2573), .B0_t (IN_key_s0_t[94]), .B0_f (IN_key_s0_f[94]), .B1_t (IN_key_s1_t[94]), .B1_f (IN_key_s1_f[94]), .Z0_t (LED_128_Instance_current_roundkey[30]), .Z0_f (new_AGEMA_signal_2764), .Z1_t (new_AGEMA_signal_2765), .Z1_f (new_AGEMA_signal_2766) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_31_U1_XOR1_U1 ( .A0_t (IN_key_s0_t[95]), .A0_f (IN_key_s0_f[95]), .A1_t (IN_key_s1_t[95]), .A1_f (IN_key_s1_f[95]), .B0_t (IN_key_s0_t[31]), .B0_f (IN_key_s0_f[31]), .B1_t (IN_key_s1_t[31]), .B1_f (IN_key_s1_f[31]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_31_U1_X), .Z0_f (new_AGEMA_signal_2179), .Z1_t (new_AGEMA_signal_2180), .Z1_f (new_AGEMA_signal_2181) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_31_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n31), .A1_f (new_AGEMA_signal_2477), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_31_U1_X), .B0_f (new_AGEMA_signal_2179), .B1_t (new_AGEMA_signal_2180), .B1_f (new_AGEMA_signal_2181), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_31_U1_Y), .Z0_f (new_AGEMA_signal_2574), .Z1_t (new_AGEMA_signal_2575), .Z1_f (new_AGEMA_signal_2576) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_31_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_31_U1_Y), .A0_f (new_AGEMA_signal_2574), .A1_t (new_AGEMA_signal_2575), .A1_f (new_AGEMA_signal_2576), .B0_t (IN_key_s0_t[95]), .B0_f (IN_key_s0_f[95]), .B1_t (IN_key_s1_t[95]), .B1_f (IN_key_s1_f[95]), .Z0_t (LED_128_Instance_current_roundkey[31]), .Z0_f (new_AGEMA_signal_2767), .Z1_t (new_AGEMA_signal_2768), .Z1_f (new_AGEMA_signal_2769) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_32_U1_XOR1_U1 ( .A0_t (IN_key_s0_t[96]), .A0_f (IN_key_s0_f[96]), .A1_t (IN_key_s1_t[96]), .A1_f (IN_key_s1_f[96]), .B0_t (IN_key_s0_t[32]), .B0_f (IN_key_s0_f[32]), .B1_t (IN_key_s1_t[32]), .B1_f (IN_key_s1_f[32]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_32_U1_X), .Z0_f (new_AGEMA_signal_2188), .Z1_t (new_AGEMA_signal_2189), .Z1_f (new_AGEMA_signal_2190) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_32_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n31), .A1_f (new_AGEMA_signal_2477), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_32_U1_X), .B0_f (new_AGEMA_signal_2188), .B1_t (new_AGEMA_signal_2189), .B1_f (new_AGEMA_signal_2190), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_32_U1_Y), .Z0_f (new_AGEMA_signal_2577), .Z1_t (new_AGEMA_signal_2578), .Z1_f (new_AGEMA_signal_2579) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_32_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_32_U1_Y), .A0_f (new_AGEMA_signal_2577), .A1_t (new_AGEMA_signal_2578), .A1_f (new_AGEMA_signal_2579), .B0_t (IN_key_s0_t[96]), .B0_f (IN_key_s0_f[96]), .B1_t (IN_key_s1_t[96]), .B1_f (IN_key_s1_f[96]), .Z0_t (LED_128_Instance_current_roundkey[32]), .Z0_f (new_AGEMA_signal_2770), .Z1_t (new_AGEMA_signal_2771), .Z1_f (new_AGEMA_signal_2772) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_33_U1_XOR1_U1 ( .A0_t (IN_key_s0_t[97]), .A0_f (IN_key_s0_f[97]), .A1_t (IN_key_s1_t[97]), .A1_f (IN_key_s1_f[97]), .B0_t (IN_key_s0_t[33]), .B0_f (IN_key_s0_f[33]), .B1_t (IN_key_s1_t[33]), .B1_f (IN_key_s1_f[33]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_33_U1_X), .Z0_f (new_AGEMA_signal_2197), .Z1_t (new_AGEMA_signal_2198), .Z1_f (new_AGEMA_signal_2199) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_33_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n31), .A1_f (new_AGEMA_signal_2477), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_33_U1_X), .B0_f (new_AGEMA_signal_2197), .B1_t (new_AGEMA_signal_2198), .B1_f (new_AGEMA_signal_2199), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_33_U1_Y), .Z0_f (new_AGEMA_signal_2580), .Z1_t (new_AGEMA_signal_2581), .Z1_f (new_AGEMA_signal_2582) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_33_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_33_U1_Y), .A0_f (new_AGEMA_signal_2580), .A1_t (new_AGEMA_signal_2581), .A1_f (new_AGEMA_signal_2582), .B0_t (IN_key_s0_t[97]), .B0_f (IN_key_s0_f[97]), .B1_t (IN_key_s1_t[97]), .B1_f (IN_key_s1_f[97]), .Z0_t (LED_128_Instance_current_roundkey[33]), .Z0_f (new_AGEMA_signal_2773), .Z1_t (new_AGEMA_signal_2774), .Z1_f (new_AGEMA_signal_2775) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_34_U1_XOR1_U1 ( .A0_t (IN_key_s0_t[98]), .A0_f (IN_key_s0_f[98]), .A1_t (IN_key_s1_t[98]), .A1_f (IN_key_s1_f[98]), .B0_t (IN_key_s0_t[34]), .B0_f (IN_key_s0_f[34]), .B1_t (IN_key_s1_t[34]), .B1_f (IN_key_s1_f[34]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_34_U1_X), .Z0_f (new_AGEMA_signal_2206), .Z1_t (new_AGEMA_signal_2207), .Z1_f (new_AGEMA_signal_2208) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_34_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n31), .A1_f (new_AGEMA_signal_2477), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_34_U1_X), .B0_f (new_AGEMA_signal_2206), .B1_t (new_AGEMA_signal_2207), .B1_f (new_AGEMA_signal_2208), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_34_U1_Y), .Z0_f (new_AGEMA_signal_2583), .Z1_t (new_AGEMA_signal_2584), .Z1_f (new_AGEMA_signal_2585) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_34_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_34_U1_Y), .A0_f (new_AGEMA_signal_2583), .A1_t (new_AGEMA_signal_2584), .A1_f (new_AGEMA_signal_2585), .B0_t (IN_key_s0_t[98]), .B0_f (IN_key_s0_f[98]), .B1_t (IN_key_s1_t[98]), .B1_f (IN_key_s1_f[98]), .Z0_t (LED_128_Instance_current_roundkey[34]), .Z0_f (new_AGEMA_signal_2776), .Z1_t (new_AGEMA_signal_2777), .Z1_f (new_AGEMA_signal_2778) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_35_U1_XOR1_U1 ( .A0_t (IN_key_s0_t[99]), .A0_f (IN_key_s0_f[99]), .A1_t (IN_key_s1_t[99]), .A1_f (IN_key_s1_f[99]), .B0_t (IN_key_s0_t[35]), .B0_f (IN_key_s0_f[35]), .B1_t (IN_key_s1_t[35]), .B1_f (IN_key_s1_f[35]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_35_U1_X), .Z0_f (new_AGEMA_signal_2215), .Z1_t (new_AGEMA_signal_2216), .Z1_f (new_AGEMA_signal_2217) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_35_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n31), .A1_f (new_AGEMA_signal_2477), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_35_U1_X), .B0_f (new_AGEMA_signal_2215), .B1_t (new_AGEMA_signal_2216), .B1_f (new_AGEMA_signal_2217), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_35_U1_Y), .Z0_f (new_AGEMA_signal_2586), .Z1_t (new_AGEMA_signal_2587), .Z1_f (new_AGEMA_signal_2588) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_35_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_35_U1_Y), .A0_f (new_AGEMA_signal_2586), .A1_t (new_AGEMA_signal_2587), .A1_f (new_AGEMA_signal_2588), .B0_t (IN_key_s0_t[99]), .B0_f (IN_key_s0_f[99]), .B1_t (IN_key_s1_t[99]), .B1_f (IN_key_s1_f[99]), .Z0_t (LED_128_Instance_current_roundkey[35]), .Z0_f (new_AGEMA_signal_2779), .Z1_t (new_AGEMA_signal_2780), .Z1_f (new_AGEMA_signal_2781) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_36_U1_XOR1_U1 ( .A0_t (IN_key_s0_t[100]), .A0_f (IN_key_s0_f[100]), .A1_t (IN_key_s1_t[100]), .A1_f (IN_key_s1_f[100]), .B0_t (IN_key_s0_t[36]), .B0_f (IN_key_s0_f[36]), .B1_t (IN_key_s1_t[36]), .B1_f (IN_key_s1_f[36]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_36_U1_X), .Z0_f (new_AGEMA_signal_2224), .Z1_t (new_AGEMA_signal_2225), .Z1_f (new_AGEMA_signal_2226) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_36_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n31), .A1_f (new_AGEMA_signal_2477), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_36_U1_X), .B0_f (new_AGEMA_signal_2224), .B1_t (new_AGEMA_signal_2225), .B1_f (new_AGEMA_signal_2226), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_36_U1_Y), .Z0_f (new_AGEMA_signal_2589), .Z1_t (new_AGEMA_signal_2590), .Z1_f (new_AGEMA_signal_2591) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_36_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_36_U1_Y), .A0_f (new_AGEMA_signal_2589), .A1_t (new_AGEMA_signal_2590), .A1_f (new_AGEMA_signal_2591), .B0_t (IN_key_s0_t[100]), .B0_f (IN_key_s0_f[100]), .B1_t (IN_key_s1_t[100]), .B1_f (IN_key_s1_f[100]), .Z0_t (LED_128_Instance_current_roundkey[36]), .Z0_f (new_AGEMA_signal_2782), .Z1_t (new_AGEMA_signal_2783), .Z1_f (new_AGEMA_signal_2784) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_37_U1_XOR1_U1 ( .A0_t (IN_key_s0_t[101]), .A0_f (IN_key_s0_f[101]), .A1_t (IN_key_s1_t[101]), .A1_f (IN_key_s1_f[101]), .B0_t (IN_key_s0_t[37]), .B0_f (IN_key_s0_f[37]), .B1_t (IN_key_s1_t[37]), .B1_f (IN_key_s1_f[37]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_37_U1_X), .Z0_f (new_AGEMA_signal_2233), .Z1_t (new_AGEMA_signal_2234), .Z1_f (new_AGEMA_signal_2235) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_37_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n31), .A1_f (new_AGEMA_signal_2477), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_37_U1_X), .B0_f (new_AGEMA_signal_2233), .B1_t (new_AGEMA_signal_2234), .B1_f (new_AGEMA_signal_2235), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_37_U1_Y), .Z0_f (new_AGEMA_signal_2592), .Z1_t (new_AGEMA_signal_2593), .Z1_f (new_AGEMA_signal_2594) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_37_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_37_U1_Y), .A0_f (new_AGEMA_signal_2592), .A1_t (new_AGEMA_signal_2593), .A1_f (new_AGEMA_signal_2594), .B0_t (IN_key_s0_t[101]), .B0_f (IN_key_s0_f[101]), .B1_t (IN_key_s1_t[101]), .B1_f (IN_key_s1_f[101]), .Z0_t (LED_128_Instance_current_roundkey[37]), .Z0_f (new_AGEMA_signal_2785), .Z1_t (new_AGEMA_signal_2786), .Z1_f (new_AGEMA_signal_2787) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_38_U1_XOR1_U1 ( .A0_t (IN_key_s0_t[102]), .A0_f (IN_key_s0_f[102]), .A1_t (IN_key_s1_t[102]), .A1_f (IN_key_s1_f[102]), .B0_t (IN_key_s0_t[38]), .B0_f (IN_key_s0_f[38]), .B1_t (IN_key_s1_t[38]), .B1_f (IN_key_s1_f[38]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_38_U1_X), .Z0_f (new_AGEMA_signal_2242), .Z1_t (new_AGEMA_signal_2243), .Z1_f (new_AGEMA_signal_2244) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_38_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n31), .A1_f (new_AGEMA_signal_2477), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_38_U1_X), .B0_f (new_AGEMA_signal_2242), .B1_t (new_AGEMA_signal_2243), .B1_f (new_AGEMA_signal_2244), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_38_U1_Y), .Z0_f (new_AGEMA_signal_2595), .Z1_t (new_AGEMA_signal_2596), .Z1_f (new_AGEMA_signal_2597) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_38_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_38_U1_Y), .A0_f (new_AGEMA_signal_2595), .A1_t (new_AGEMA_signal_2596), .A1_f (new_AGEMA_signal_2597), .B0_t (IN_key_s0_t[102]), .B0_f (IN_key_s0_f[102]), .B1_t (IN_key_s1_t[102]), .B1_f (IN_key_s1_f[102]), .Z0_t (LED_128_Instance_current_roundkey[38]), .Z0_f (new_AGEMA_signal_2788), .Z1_t (new_AGEMA_signal_2789), .Z1_f (new_AGEMA_signal_2790) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_39_U1_XOR1_U1 ( .A0_t (IN_key_s0_t[103]), .A0_f (IN_key_s0_f[103]), .A1_t (IN_key_s1_t[103]), .A1_f (IN_key_s1_f[103]), .B0_t (IN_key_s0_t[39]), .B0_f (IN_key_s0_f[39]), .B1_t (IN_key_s1_t[39]), .B1_f (IN_key_s1_f[39]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_39_U1_X), .Z0_f (new_AGEMA_signal_2251), .Z1_t (new_AGEMA_signal_2252), .Z1_f (new_AGEMA_signal_2253) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_39_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n31), .A1_f (new_AGEMA_signal_2477), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_39_U1_X), .B0_f (new_AGEMA_signal_2251), .B1_t (new_AGEMA_signal_2252), .B1_f (new_AGEMA_signal_2253), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_39_U1_Y), .Z0_f (new_AGEMA_signal_2598), .Z1_t (new_AGEMA_signal_2599), .Z1_f (new_AGEMA_signal_2600) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_39_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_39_U1_Y), .A0_f (new_AGEMA_signal_2598), .A1_t (new_AGEMA_signal_2599), .A1_f (new_AGEMA_signal_2600), .B0_t (IN_key_s0_t[103]), .B0_f (IN_key_s0_f[103]), .B1_t (IN_key_s1_t[103]), .B1_f (IN_key_s1_f[103]), .Z0_t (LED_128_Instance_current_roundkey[39]), .Z0_f (new_AGEMA_signal_2791), .Z1_t (new_AGEMA_signal_2792), .Z1_f (new_AGEMA_signal_2793) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_40_U1_XOR1_U1 ( .A0_t (IN_key_s0_t[104]), .A0_f (IN_key_s0_f[104]), .A1_t (IN_key_s1_t[104]), .A1_f (IN_key_s1_f[104]), .B0_t (IN_key_s0_t[40]), .B0_f (IN_key_s0_f[40]), .B1_t (IN_key_s1_t[40]), .B1_f (IN_key_s1_f[40]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_40_U1_X), .Z0_f (new_AGEMA_signal_2260), .Z1_t (new_AGEMA_signal_2261), .Z1_f (new_AGEMA_signal_2262) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_40_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n31), .A1_f (new_AGEMA_signal_2477), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_40_U1_X), .B0_f (new_AGEMA_signal_2260), .B1_t (new_AGEMA_signal_2261), .B1_f (new_AGEMA_signal_2262), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_40_U1_Y), .Z0_f (new_AGEMA_signal_2601), .Z1_t (new_AGEMA_signal_2602), .Z1_f (new_AGEMA_signal_2603) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_40_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_40_U1_Y), .A0_f (new_AGEMA_signal_2601), .A1_t (new_AGEMA_signal_2602), .A1_f (new_AGEMA_signal_2603), .B0_t (IN_key_s0_t[104]), .B0_f (IN_key_s0_f[104]), .B1_t (IN_key_s1_t[104]), .B1_f (IN_key_s1_f[104]), .Z0_t (LED_128_Instance_current_roundkey[40]), .Z0_f (new_AGEMA_signal_2794), .Z1_t (new_AGEMA_signal_2795), .Z1_f (new_AGEMA_signal_2796) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_41_U1_XOR1_U1 ( .A0_t (IN_key_s0_t[105]), .A0_f (IN_key_s0_f[105]), .A1_t (IN_key_s1_t[105]), .A1_f (IN_key_s1_f[105]), .B0_t (IN_key_s0_t[41]), .B0_f (IN_key_s0_f[41]), .B1_t (IN_key_s1_t[41]), .B1_f (IN_key_s1_f[41]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_41_U1_X), .Z0_f (new_AGEMA_signal_2269), .Z1_t (new_AGEMA_signal_2270), .Z1_f (new_AGEMA_signal_2271) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_41_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n31), .A1_f (new_AGEMA_signal_2477), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_41_U1_X), .B0_f (new_AGEMA_signal_2269), .B1_t (new_AGEMA_signal_2270), .B1_f (new_AGEMA_signal_2271), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_41_U1_Y), .Z0_f (new_AGEMA_signal_2604), .Z1_t (new_AGEMA_signal_2605), .Z1_f (new_AGEMA_signal_2606) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_41_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_41_U1_Y), .A0_f (new_AGEMA_signal_2604), .A1_t (new_AGEMA_signal_2605), .A1_f (new_AGEMA_signal_2606), .B0_t (IN_key_s0_t[105]), .B0_f (IN_key_s0_f[105]), .B1_t (IN_key_s1_t[105]), .B1_f (IN_key_s1_f[105]), .Z0_t (LED_128_Instance_current_roundkey[41]), .Z0_f (new_AGEMA_signal_2797), .Z1_t (new_AGEMA_signal_2798), .Z1_f (new_AGEMA_signal_2799) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_42_U1_XOR1_U1 ( .A0_t (IN_key_s0_t[106]), .A0_f (IN_key_s0_f[106]), .A1_t (IN_key_s1_t[106]), .A1_f (IN_key_s1_f[106]), .B0_t (IN_key_s0_t[42]), .B0_f (IN_key_s0_f[42]), .B1_t (IN_key_s1_t[42]), .B1_f (IN_key_s1_f[42]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_42_U1_X), .Z0_f (new_AGEMA_signal_2278), .Z1_t (new_AGEMA_signal_2279), .Z1_f (new_AGEMA_signal_2280) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_42_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n31), .A1_f (new_AGEMA_signal_2477), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_42_U1_X), .B0_f (new_AGEMA_signal_2278), .B1_t (new_AGEMA_signal_2279), .B1_f (new_AGEMA_signal_2280), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_42_U1_Y), .Z0_f (new_AGEMA_signal_2607), .Z1_t (new_AGEMA_signal_2608), .Z1_f (new_AGEMA_signal_2609) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_42_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_42_U1_Y), .A0_f (new_AGEMA_signal_2607), .A1_t (new_AGEMA_signal_2608), .A1_f (new_AGEMA_signal_2609), .B0_t (IN_key_s0_t[106]), .B0_f (IN_key_s0_f[106]), .B1_t (IN_key_s1_t[106]), .B1_f (IN_key_s1_f[106]), .Z0_t (LED_128_Instance_current_roundkey[42]), .Z0_f (new_AGEMA_signal_2800), .Z1_t (new_AGEMA_signal_2801), .Z1_f (new_AGEMA_signal_2802) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_43_U1_XOR1_U1 ( .A0_t (IN_key_s0_t[107]), .A0_f (IN_key_s0_f[107]), .A1_t (IN_key_s1_t[107]), .A1_f (IN_key_s1_f[107]), .B0_t (IN_key_s0_t[43]), .B0_f (IN_key_s0_f[43]), .B1_t (IN_key_s1_t[43]), .B1_f (IN_key_s1_f[43]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_43_U1_X), .Z0_f (new_AGEMA_signal_2287), .Z1_t (new_AGEMA_signal_2288), .Z1_f (new_AGEMA_signal_2289) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_43_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n31), .A1_f (new_AGEMA_signal_2477), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_43_U1_X), .B0_f (new_AGEMA_signal_2287), .B1_t (new_AGEMA_signal_2288), .B1_f (new_AGEMA_signal_2289), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_43_U1_Y), .Z0_f (new_AGEMA_signal_2610), .Z1_t (new_AGEMA_signal_2611), .Z1_f (new_AGEMA_signal_2612) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_43_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_43_U1_Y), .A0_f (new_AGEMA_signal_2610), .A1_t (new_AGEMA_signal_2611), .A1_f (new_AGEMA_signal_2612), .B0_t (IN_key_s0_t[107]), .B0_f (IN_key_s0_f[107]), .B1_t (IN_key_s1_t[107]), .B1_f (IN_key_s1_f[107]), .Z0_t (LED_128_Instance_current_roundkey[43]), .Z0_f (new_AGEMA_signal_2803), .Z1_t (new_AGEMA_signal_2804), .Z1_f (new_AGEMA_signal_2805) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_44_U1_XOR1_U1 ( .A0_t (IN_key_s0_t[108]), .A0_f (IN_key_s0_f[108]), .A1_t (IN_key_s1_t[108]), .A1_f (IN_key_s1_f[108]), .B0_t (IN_key_s0_t[44]), .B0_f (IN_key_s0_f[44]), .B1_t (IN_key_s1_t[44]), .B1_f (IN_key_s1_f[44]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_44_U1_X), .Z0_f (new_AGEMA_signal_2296), .Z1_t (new_AGEMA_signal_2297), .Z1_f (new_AGEMA_signal_2298) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_44_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n31), .A1_f (new_AGEMA_signal_2477), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_44_U1_X), .B0_f (new_AGEMA_signal_2296), .B1_t (new_AGEMA_signal_2297), .B1_f (new_AGEMA_signal_2298), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_44_U1_Y), .Z0_f (new_AGEMA_signal_2613), .Z1_t (new_AGEMA_signal_2614), .Z1_f (new_AGEMA_signal_2615) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_44_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_44_U1_Y), .A0_f (new_AGEMA_signal_2613), .A1_t (new_AGEMA_signal_2614), .A1_f (new_AGEMA_signal_2615), .B0_t (IN_key_s0_t[108]), .B0_f (IN_key_s0_f[108]), .B1_t (IN_key_s1_t[108]), .B1_f (IN_key_s1_f[108]), .Z0_t (LED_128_Instance_current_roundkey[44]), .Z0_f (new_AGEMA_signal_2806), .Z1_t (new_AGEMA_signal_2807), .Z1_f (new_AGEMA_signal_2808) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_45_U1_XOR1_U1 ( .A0_t (IN_key_s0_t[109]), .A0_f (IN_key_s0_f[109]), .A1_t (IN_key_s1_t[109]), .A1_f (IN_key_s1_f[109]), .B0_t (IN_key_s0_t[45]), .B0_f (IN_key_s0_f[45]), .B1_t (IN_key_s1_t[45]), .B1_f (IN_key_s1_f[45]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_45_U1_X), .Z0_f (new_AGEMA_signal_2305), .Z1_t (new_AGEMA_signal_2306), .Z1_f (new_AGEMA_signal_2307) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_45_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n31), .A1_f (new_AGEMA_signal_2477), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_45_U1_X), .B0_f (new_AGEMA_signal_2305), .B1_t (new_AGEMA_signal_2306), .B1_f (new_AGEMA_signal_2307), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_45_U1_Y), .Z0_f (new_AGEMA_signal_2616), .Z1_t (new_AGEMA_signal_2617), .Z1_f (new_AGEMA_signal_2618) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_45_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_45_U1_Y), .A0_f (new_AGEMA_signal_2616), .A1_t (new_AGEMA_signal_2617), .A1_f (new_AGEMA_signal_2618), .B0_t (IN_key_s0_t[109]), .B0_f (IN_key_s0_f[109]), .B1_t (IN_key_s1_t[109]), .B1_f (IN_key_s1_f[109]), .Z0_t (LED_128_Instance_current_roundkey[45]), .Z0_f (new_AGEMA_signal_2809), .Z1_t (new_AGEMA_signal_2810), .Z1_f (new_AGEMA_signal_2811) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_46_U1_XOR1_U1 ( .A0_t (IN_key_s0_t[110]), .A0_f (IN_key_s0_f[110]), .A1_t (IN_key_s1_t[110]), .A1_f (IN_key_s1_f[110]), .B0_t (IN_key_s0_t[46]), .B0_f (IN_key_s0_f[46]), .B1_t (IN_key_s1_t[46]), .B1_f (IN_key_s1_f[46]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_46_U1_X), .Z0_f (new_AGEMA_signal_2314), .Z1_t (new_AGEMA_signal_2315), .Z1_f (new_AGEMA_signal_2316) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_46_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n31), .A1_f (new_AGEMA_signal_2477), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_46_U1_X), .B0_f (new_AGEMA_signal_2314), .B1_t (new_AGEMA_signal_2315), .B1_f (new_AGEMA_signal_2316), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_46_U1_Y), .Z0_f (new_AGEMA_signal_2619), .Z1_t (new_AGEMA_signal_2620), .Z1_f (new_AGEMA_signal_2621) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_46_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_46_U1_Y), .A0_f (new_AGEMA_signal_2619), .A1_t (new_AGEMA_signal_2620), .A1_f (new_AGEMA_signal_2621), .B0_t (IN_key_s0_t[110]), .B0_f (IN_key_s0_f[110]), .B1_t (IN_key_s1_t[110]), .B1_f (IN_key_s1_f[110]), .Z0_t (LED_128_Instance_current_roundkey[46]), .Z0_f (new_AGEMA_signal_2812), .Z1_t (new_AGEMA_signal_2813), .Z1_f (new_AGEMA_signal_2814) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_47_U1_XOR1_U1 ( .A0_t (IN_key_s0_t[111]), .A0_f (IN_key_s0_f[111]), .A1_t (IN_key_s1_t[111]), .A1_f (IN_key_s1_f[111]), .B0_t (IN_key_s0_t[47]), .B0_f (IN_key_s0_f[47]), .B1_t (IN_key_s1_t[47]), .B1_f (IN_key_s1_f[47]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_47_U1_X), .Z0_f (new_AGEMA_signal_2323), .Z1_t (new_AGEMA_signal_2324), .Z1_f (new_AGEMA_signal_2325) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_47_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n31), .A1_f (new_AGEMA_signal_2477), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_47_U1_X), .B0_f (new_AGEMA_signal_2323), .B1_t (new_AGEMA_signal_2324), .B1_f (new_AGEMA_signal_2325), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_47_U1_Y), .Z0_f (new_AGEMA_signal_2622), .Z1_t (new_AGEMA_signal_2623), .Z1_f (new_AGEMA_signal_2624) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_47_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_47_U1_Y), .A0_f (new_AGEMA_signal_2622), .A1_t (new_AGEMA_signal_2623), .A1_f (new_AGEMA_signal_2624), .B0_t (IN_key_s0_t[111]), .B0_f (IN_key_s0_f[111]), .B1_t (IN_key_s1_t[111]), .B1_f (IN_key_s1_f[111]), .Z0_t (LED_128_Instance_current_roundkey[47]), .Z0_f (new_AGEMA_signal_2815), .Z1_t (new_AGEMA_signal_2816), .Z1_f (new_AGEMA_signal_2817) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_48_U1_XOR1_U1 ( .A0_t (IN_key_s0_t[112]), .A0_f (IN_key_s0_f[112]), .A1_t (IN_key_s1_t[112]), .A1_f (IN_key_s1_f[112]), .B0_t (IN_key_s0_t[48]), .B0_f (IN_key_s0_f[48]), .B1_t (IN_key_s1_t[48]), .B1_f (IN_key_s1_f[48]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_48_U1_X), .Z0_f (new_AGEMA_signal_2332), .Z1_t (new_AGEMA_signal_2333), .Z1_f (new_AGEMA_signal_2334) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_48_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n31), .A1_f (new_AGEMA_signal_2477), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_48_U1_X), .B0_f (new_AGEMA_signal_2332), .B1_t (new_AGEMA_signal_2333), .B1_f (new_AGEMA_signal_2334), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_48_U1_Y), .Z0_f (new_AGEMA_signal_2625), .Z1_t (new_AGEMA_signal_2626), .Z1_f (new_AGEMA_signal_2627) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_48_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_48_U1_Y), .A0_f (new_AGEMA_signal_2625), .A1_t (new_AGEMA_signal_2626), .A1_f (new_AGEMA_signal_2627), .B0_t (IN_key_s0_t[112]), .B0_f (IN_key_s0_f[112]), .B1_t (IN_key_s1_t[112]), .B1_f (IN_key_s1_f[112]), .Z0_t (LED_128_Instance_current_roundkey[48]), .Z0_f (new_AGEMA_signal_2818), .Z1_t (new_AGEMA_signal_2819), .Z1_f (new_AGEMA_signal_2820) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_49_U1_XOR1_U1 ( .A0_t (IN_key_s0_t[113]), .A0_f (IN_key_s0_f[113]), .A1_t (IN_key_s1_t[113]), .A1_f (IN_key_s1_f[113]), .B0_t (IN_key_s0_t[49]), .B0_f (IN_key_s0_f[49]), .B1_t (IN_key_s1_t[49]), .B1_f (IN_key_s1_f[49]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_49_U1_X), .Z0_f (new_AGEMA_signal_2341), .Z1_t (new_AGEMA_signal_2342), .Z1_f (new_AGEMA_signal_2343) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_49_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n31), .A1_f (new_AGEMA_signal_2477), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_49_U1_X), .B0_f (new_AGEMA_signal_2341), .B1_t (new_AGEMA_signal_2342), .B1_f (new_AGEMA_signal_2343), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_49_U1_Y), .Z0_f (new_AGEMA_signal_2628), .Z1_t (new_AGEMA_signal_2629), .Z1_f (new_AGEMA_signal_2630) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_49_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_49_U1_Y), .A0_f (new_AGEMA_signal_2628), .A1_t (new_AGEMA_signal_2629), .A1_f (new_AGEMA_signal_2630), .B0_t (IN_key_s0_t[113]), .B0_f (IN_key_s0_f[113]), .B1_t (IN_key_s1_t[113]), .B1_f (IN_key_s1_f[113]), .Z0_t (LED_128_Instance_current_roundkey[49]), .Z0_f (new_AGEMA_signal_2821), .Z1_t (new_AGEMA_signal_2822), .Z1_f (new_AGEMA_signal_2823) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_50_U1_XOR1_U1 ( .A0_t (IN_key_s0_t[114]), .A0_f (IN_key_s0_f[114]), .A1_t (IN_key_s1_t[114]), .A1_f (IN_key_s1_f[114]), .B0_t (IN_key_s0_t[50]), .B0_f (IN_key_s0_f[50]), .B1_t (IN_key_s1_t[50]), .B1_f (IN_key_s1_f[50]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_50_U1_X), .Z0_f (new_AGEMA_signal_2350), .Z1_t (new_AGEMA_signal_2351), .Z1_f (new_AGEMA_signal_2352) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_50_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n31), .A1_f (new_AGEMA_signal_2477), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_50_U1_X), .B0_f (new_AGEMA_signal_2350), .B1_t (new_AGEMA_signal_2351), .B1_f (new_AGEMA_signal_2352), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_50_U1_Y), .Z0_f (new_AGEMA_signal_2631), .Z1_t (new_AGEMA_signal_2632), .Z1_f (new_AGEMA_signal_2633) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_50_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_50_U1_Y), .A0_f (new_AGEMA_signal_2631), .A1_t (new_AGEMA_signal_2632), .A1_f (new_AGEMA_signal_2633), .B0_t (IN_key_s0_t[114]), .B0_f (IN_key_s0_f[114]), .B1_t (IN_key_s1_t[114]), .B1_f (IN_key_s1_f[114]), .Z0_t (LED_128_Instance_current_roundkey[50]), .Z0_f (new_AGEMA_signal_2824), .Z1_t (new_AGEMA_signal_2825), .Z1_f (new_AGEMA_signal_2826) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_51_U1_XOR1_U1 ( .A0_t (IN_key_s0_t[115]), .A0_f (IN_key_s0_f[115]), .A1_t (IN_key_s1_t[115]), .A1_f (IN_key_s1_f[115]), .B0_t (IN_key_s0_t[51]), .B0_f (IN_key_s0_f[51]), .B1_t (IN_key_s1_t[51]), .B1_f (IN_key_s1_f[51]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_51_U1_X), .Z0_f (new_AGEMA_signal_2359), .Z1_t (new_AGEMA_signal_2360), .Z1_f (new_AGEMA_signal_2361) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_51_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n31), .A1_f (new_AGEMA_signal_2477), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_51_U1_X), .B0_f (new_AGEMA_signal_2359), .B1_t (new_AGEMA_signal_2360), .B1_f (new_AGEMA_signal_2361), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_51_U1_Y), .Z0_f (new_AGEMA_signal_2634), .Z1_t (new_AGEMA_signal_2635), .Z1_f (new_AGEMA_signal_2636) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_51_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_51_U1_Y), .A0_f (new_AGEMA_signal_2634), .A1_t (new_AGEMA_signal_2635), .A1_f (new_AGEMA_signal_2636), .B0_t (IN_key_s0_t[115]), .B0_f (IN_key_s0_f[115]), .B1_t (IN_key_s1_t[115]), .B1_f (IN_key_s1_f[115]), .Z0_t (LED_128_Instance_current_roundkey[51]), .Z0_f (new_AGEMA_signal_2827), .Z1_t (new_AGEMA_signal_2828), .Z1_f (new_AGEMA_signal_2829) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_52_U1_XOR1_U1 ( .A0_t (IN_key_s0_t[116]), .A0_f (IN_key_s0_f[116]), .A1_t (IN_key_s1_t[116]), .A1_f (IN_key_s1_f[116]), .B0_t (IN_key_s0_t[52]), .B0_f (IN_key_s0_f[52]), .B1_t (IN_key_s1_t[52]), .B1_f (IN_key_s1_f[52]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_52_U1_X), .Z0_f (new_AGEMA_signal_2368), .Z1_t (new_AGEMA_signal_2369), .Z1_f (new_AGEMA_signal_2370) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_52_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n31), .A1_f (new_AGEMA_signal_2477), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_52_U1_X), .B0_f (new_AGEMA_signal_2368), .B1_t (new_AGEMA_signal_2369), .B1_f (new_AGEMA_signal_2370), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_52_U1_Y), .Z0_f (new_AGEMA_signal_2637), .Z1_t (new_AGEMA_signal_2638), .Z1_f (new_AGEMA_signal_2639) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_52_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_52_U1_Y), .A0_f (new_AGEMA_signal_2637), .A1_t (new_AGEMA_signal_2638), .A1_f (new_AGEMA_signal_2639), .B0_t (IN_key_s0_t[116]), .B0_f (IN_key_s0_f[116]), .B1_t (IN_key_s1_t[116]), .B1_f (IN_key_s1_f[116]), .Z0_t (LED_128_Instance_current_roundkey[52]), .Z0_f (new_AGEMA_signal_2830), .Z1_t (new_AGEMA_signal_2831), .Z1_f (new_AGEMA_signal_2832) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_53_U1_XOR1_U1 ( .A0_t (IN_key_s0_t[117]), .A0_f (IN_key_s0_f[117]), .A1_t (IN_key_s1_t[117]), .A1_f (IN_key_s1_f[117]), .B0_t (IN_key_s0_t[53]), .B0_f (IN_key_s0_f[53]), .B1_t (IN_key_s1_t[53]), .B1_f (IN_key_s1_f[53]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_53_U1_X), .Z0_f (new_AGEMA_signal_2377), .Z1_t (new_AGEMA_signal_2378), .Z1_f (new_AGEMA_signal_2379) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_53_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n31), .A1_f (new_AGEMA_signal_2477), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_53_U1_X), .B0_f (new_AGEMA_signal_2377), .B1_t (new_AGEMA_signal_2378), .B1_f (new_AGEMA_signal_2379), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_53_U1_Y), .Z0_f (new_AGEMA_signal_2640), .Z1_t (new_AGEMA_signal_2641), .Z1_f (new_AGEMA_signal_2642) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_53_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_53_U1_Y), .A0_f (new_AGEMA_signal_2640), .A1_t (new_AGEMA_signal_2641), .A1_f (new_AGEMA_signal_2642), .B0_t (IN_key_s0_t[117]), .B0_f (IN_key_s0_f[117]), .B1_t (IN_key_s1_t[117]), .B1_f (IN_key_s1_f[117]), .Z0_t (LED_128_Instance_current_roundkey[53]), .Z0_f (new_AGEMA_signal_2833), .Z1_t (new_AGEMA_signal_2834), .Z1_f (new_AGEMA_signal_2835) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_54_U1_XOR1_U1 ( .A0_t (IN_key_s0_t[118]), .A0_f (IN_key_s0_f[118]), .A1_t (IN_key_s1_t[118]), .A1_f (IN_key_s1_f[118]), .B0_t (IN_key_s0_t[54]), .B0_f (IN_key_s0_f[54]), .B1_t (IN_key_s1_t[54]), .B1_f (IN_key_s1_f[54]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_54_U1_X), .Z0_f (new_AGEMA_signal_2386), .Z1_t (new_AGEMA_signal_2387), .Z1_f (new_AGEMA_signal_2388) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_54_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n31), .A1_f (new_AGEMA_signal_2477), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_54_U1_X), .B0_f (new_AGEMA_signal_2386), .B1_t (new_AGEMA_signal_2387), .B1_f (new_AGEMA_signal_2388), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_54_U1_Y), .Z0_f (new_AGEMA_signal_2643), .Z1_t (new_AGEMA_signal_2644), .Z1_f (new_AGEMA_signal_2645) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_54_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_54_U1_Y), .A0_f (new_AGEMA_signal_2643), .A1_t (new_AGEMA_signal_2644), .A1_f (new_AGEMA_signal_2645), .B0_t (IN_key_s0_t[118]), .B0_f (IN_key_s0_f[118]), .B1_t (IN_key_s1_t[118]), .B1_f (IN_key_s1_f[118]), .Z0_t (LED_128_Instance_current_roundkey[54]), .Z0_f (new_AGEMA_signal_2836), .Z1_t (new_AGEMA_signal_2837), .Z1_f (new_AGEMA_signal_2838) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_55_U1_XOR1_U1 ( .A0_t (IN_key_s0_t[119]), .A0_f (IN_key_s0_f[119]), .A1_t (IN_key_s1_t[119]), .A1_f (IN_key_s1_f[119]), .B0_t (IN_key_s0_t[55]), .B0_f (IN_key_s0_f[55]), .B1_t (IN_key_s1_t[55]), .B1_f (IN_key_s1_f[55]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_55_U1_X), .Z0_f (new_AGEMA_signal_2395), .Z1_t (new_AGEMA_signal_2396), .Z1_f (new_AGEMA_signal_2397) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_55_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n31), .A1_f (new_AGEMA_signal_2477), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_55_U1_X), .B0_f (new_AGEMA_signal_2395), .B1_t (new_AGEMA_signal_2396), .B1_f (new_AGEMA_signal_2397), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_55_U1_Y), .Z0_f (new_AGEMA_signal_2646), .Z1_t (new_AGEMA_signal_2647), .Z1_f (new_AGEMA_signal_2648) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_55_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_55_U1_Y), .A0_f (new_AGEMA_signal_2646), .A1_t (new_AGEMA_signal_2647), .A1_f (new_AGEMA_signal_2648), .B0_t (IN_key_s0_t[119]), .B0_f (IN_key_s0_f[119]), .B1_t (IN_key_s1_t[119]), .B1_f (IN_key_s1_f[119]), .Z0_t (LED_128_Instance_current_roundkey[55]), .Z0_f (new_AGEMA_signal_2839), .Z1_t (new_AGEMA_signal_2840), .Z1_f (new_AGEMA_signal_2841) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_56_U1_XOR1_U1 ( .A0_t (IN_key_s0_t[120]), .A0_f (IN_key_s0_f[120]), .A1_t (IN_key_s1_t[120]), .A1_f (IN_key_s1_f[120]), .B0_t (IN_key_s0_t[56]), .B0_f (IN_key_s0_f[56]), .B1_t (IN_key_s1_t[56]), .B1_f (IN_key_s1_f[56]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_56_U1_X), .Z0_f (new_AGEMA_signal_2404), .Z1_t (new_AGEMA_signal_2405), .Z1_f (new_AGEMA_signal_2406) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_56_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n31), .A1_f (new_AGEMA_signal_2477), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_56_U1_X), .B0_f (new_AGEMA_signal_2404), .B1_t (new_AGEMA_signal_2405), .B1_f (new_AGEMA_signal_2406), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_56_U1_Y), .Z0_f (new_AGEMA_signal_2649), .Z1_t (new_AGEMA_signal_2650), .Z1_f (new_AGEMA_signal_2651) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_56_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_56_U1_Y), .A0_f (new_AGEMA_signal_2649), .A1_t (new_AGEMA_signal_2650), .A1_f (new_AGEMA_signal_2651), .B0_t (IN_key_s0_t[120]), .B0_f (IN_key_s0_f[120]), .B1_t (IN_key_s1_t[120]), .B1_f (IN_key_s1_f[120]), .Z0_t (LED_128_Instance_current_roundkey[56]), .Z0_f (new_AGEMA_signal_2842), .Z1_t (new_AGEMA_signal_2843), .Z1_f (new_AGEMA_signal_2844) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_57_U1_XOR1_U1 ( .A0_t (IN_key_s0_t[121]), .A0_f (IN_key_s0_f[121]), .A1_t (IN_key_s1_t[121]), .A1_f (IN_key_s1_f[121]), .B0_t (IN_key_s0_t[57]), .B0_f (IN_key_s0_f[57]), .B1_t (IN_key_s1_t[57]), .B1_f (IN_key_s1_f[57]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_57_U1_X), .Z0_f (new_AGEMA_signal_2413), .Z1_t (new_AGEMA_signal_2414), .Z1_f (new_AGEMA_signal_2415) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_57_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n31), .A1_f (new_AGEMA_signal_2477), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_57_U1_X), .B0_f (new_AGEMA_signal_2413), .B1_t (new_AGEMA_signal_2414), .B1_f (new_AGEMA_signal_2415), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_57_U1_Y), .Z0_f (new_AGEMA_signal_2652), .Z1_t (new_AGEMA_signal_2653), .Z1_f (new_AGEMA_signal_2654) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_57_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_57_U1_Y), .A0_f (new_AGEMA_signal_2652), .A1_t (new_AGEMA_signal_2653), .A1_f (new_AGEMA_signal_2654), .B0_t (IN_key_s0_t[121]), .B0_f (IN_key_s0_f[121]), .B1_t (IN_key_s1_t[121]), .B1_f (IN_key_s1_f[121]), .Z0_t (LED_128_Instance_current_roundkey[57]), .Z0_f (new_AGEMA_signal_2845), .Z1_t (new_AGEMA_signal_2846), .Z1_f (new_AGEMA_signal_2847) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_58_U1_XOR1_U1 ( .A0_t (IN_key_s0_t[122]), .A0_f (IN_key_s0_f[122]), .A1_t (IN_key_s1_t[122]), .A1_f (IN_key_s1_f[122]), .B0_t (IN_key_s0_t[58]), .B0_f (IN_key_s0_f[58]), .B1_t (IN_key_s1_t[58]), .B1_f (IN_key_s1_f[58]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_58_U1_X), .Z0_f (new_AGEMA_signal_2422), .Z1_t (new_AGEMA_signal_2423), .Z1_f (new_AGEMA_signal_2424) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_58_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n31), .A1_f (new_AGEMA_signal_2477), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_58_U1_X), .B0_f (new_AGEMA_signal_2422), .B1_t (new_AGEMA_signal_2423), .B1_f (new_AGEMA_signal_2424), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_58_U1_Y), .Z0_f (new_AGEMA_signal_2655), .Z1_t (new_AGEMA_signal_2656), .Z1_f (new_AGEMA_signal_2657) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_58_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_58_U1_Y), .A0_f (new_AGEMA_signal_2655), .A1_t (new_AGEMA_signal_2656), .A1_f (new_AGEMA_signal_2657), .B0_t (IN_key_s0_t[122]), .B0_f (IN_key_s0_f[122]), .B1_t (IN_key_s1_t[122]), .B1_f (IN_key_s1_f[122]), .Z0_t (LED_128_Instance_current_roundkey[58]), .Z0_f (new_AGEMA_signal_2848), .Z1_t (new_AGEMA_signal_2849), .Z1_f (new_AGEMA_signal_2850) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_59_U1_XOR1_U1 ( .A0_t (IN_key_s0_t[123]), .A0_f (IN_key_s0_f[123]), .A1_t (IN_key_s1_t[123]), .A1_f (IN_key_s1_f[123]), .B0_t (IN_key_s0_t[59]), .B0_f (IN_key_s0_f[59]), .B1_t (IN_key_s1_t[59]), .B1_f (IN_key_s1_f[59]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_59_U1_X), .Z0_f (new_AGEMA_signal_2431), .Z1_t (new_AGEMA_signal_2432), .Z1_f (new_AGEMA_signal_2433) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_59_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n31), .A1_f (new_AGEMA_signal_2477), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_59_U1_X), .B0_f (new_AGEMA_signal_2431), .B1_t (new_AGEMA_signal_2432), .B1_f (new_AGEMA_signal_2433), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_59_U1_Y), .Z0_f (new_AGEMA_signal_2658), .Z1_t (new_AGEMA_signal_2659), .Z1_f (new_AGEMA_signal_2660) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_59_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_59_U1_Y), .A0_f (new_AGEMA_signal_2658), .A1_t (new_AGEMA_signal_2659), .A1_f (new_AGEMA_signal_2660), .B0_t (IN_key_s0_t[123]), .B0_f (IN_key_s0_f[123]), .B1_t (IN_key_s1_t[123]), .B1_f (IN_key_s1_f[123]), .Z0_t (LED_128_Instance_current_roundkey[59]), .Z0_f (new_AGEMA_signal_2851), .Z1_t (new_AGEMA_signal_2852), .Z1_f (new_AGEMA_signal_2853) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_60_U1_XOR1_U1 ( .A0_t (IN_key_s0_t[124]), .A0_f (IN_key_s0_f[124]), .A1_t (IN_key_s1_t[124]), .A1_f (IN_key_s1_f[124]), .B0_t (IN_key_s0_t[60]), .B0_f (IN_key_s0_f[60]), .B1_t (IN_key_s1_t[60]), .B1_f (IN_key_s1_f[60]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_60_U1_X), .Z0_f (new_AGEMA_signal_2440), .Z1_t (new_AGEMA_signal_2441), .Z1_f (new_AGEMA_signal_2442) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_60_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n31), .A1_f (new_AGEMA_signal_2477), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_60_U1_X), .B0_f (new_AGEMA_signal_2440), .B1_t (new_AGEMA_signal_2441), .B1_f (new_AGEMA_signal_2442), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_60_U1_Y), .Z0_f (new_AGEMA_signal_2661), .Z1_t (new_AGEMA_signal_2662), .Z1_f (new_AGEMA_signal_2663) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_60_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_60_U1_Y), .A0_f (new_AGEMA_signal_2661), .A1_t (new_AGEMA_signal_2662), .A1_f (new_AGEMA_signal_2663), .B0_t (IN_key_s0_t[124]), .B0_f (IN_key_s0_f[124]), .B1_t (IN_key_s1_t[124]), .B1_f (IN_key_s1_f[124]), .Z0_t (LED_128_Instance_current_roundkey[60]), .Z0_f (new_AGEMA_signal_2854), .Z1_t (new_AGEMA_signal_2855), .Z1_f (new_AGEMA_signal_2856) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_61_U1_XOR1_U1 ( .A0_t (IN_key_s0_t[125]), .A0_f (IN_key_s0_f[125]), .A1_t (IN_key_s1_t[125]), .A1_f (IN_key_s1_f[125]), .B0_t (IN_key_s0_t[61]), .B0_f (IN_key_s0_f[61]), .B1_t (IN_key_s1_t[61]), .B1_f (IN_key_s1_f[61]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_61_U1_X), .Z0_f (new_AGEMA_signal_2449), .Z1_t (new_AGEMA_signal_2450), .Z1_f (new_AGEMA_signal_2451) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_61_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n31), .A1_f (new_AGEMA_signal_2477), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_61_U1_X), .B0_f (new_AGEMA_signal_2449), .B1_t (new_AGEMA_signal_2450), .B1_f (new_AGEMA_signal_2451), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_61_U1_Y), .Z0_f (new_AGEMA_signal_2664), .Z1_t (new_AGEMA_signal_2665), .Z1_f (new_AGEMA_signal_2666) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_61_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_61_U1_Y), .A0_f (new_AGEMA_signal_2664), .A1_t (new_AGEMA_signal_2665), .A1_f (new_AGEMA_signal_2666), .B0_t (IN_key_s0_t[125]), .B0_f (IN_key_s0_f[125]), .B1_t (IN_key_s1_t[125]), .B1_f (IN_key_s1_f[125]), .Z0_t (LED_128_Instance_current_roundkey[61]), .Z0_f (new_AGEMA_signal_2857), .Z1_t (new_AGEMA_signal_2858), .Z1_f (new_AGEMA_signal_2859) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_62_U1_XOR1_U1 ( .A0_t (IN_key_s0_t[126]), .A0_f (IN_key_s0_f[126]), .A1_t (IN_key_s1_t[126]), .A1_f (IN_key_s1_f[126]), .B0_t (IN_key_s0_t[62]), .B0_f (IN_key_s0_f[62]), .B1_t (IN_key_s1_t[62]), .B1_f (IN_key_s1_f[62]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_62_U1_X), .Z0_f (new_AGEMA_signal_2458), .Z1_t (new_AGEMA_signal_2459), .Z1_f (new_AGEMA_signal_2460) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_62_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n31), .A1_f (new_AGEMA_signal_2477), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_62_U1_X), .B0_f (new_AGEMA_signal_2458), .B1_t (new_AGEMA_signal_2459), .B1_f (new_AGEMA_signal_2460), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_62_U1_Y), .Z0_f (new_AGEMA_signal_2667), .Z1_t (new_AGEMA_signal_2668), .Z1_f (new_AGEMA_signal_2669) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_62_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_62_U1_Y), .A0_f (new_AGEMA_signal_2667), .A1_t (new_AGEMA_signal_2668), .A1_f (new_AGEMA_signal_2669), .B0_t (IN_key_s0_t[126]), .B0_f (IN_key_s0_f[126]), .B1_t (IN_key_s1_t[126]), .B1_f (IN_key_s1_f[126]), .Z0_t (LED_128_Instance_current_roundkey[62]), .Z0_f (new_AGEMA_signal_2860), .Z1_t (new_AGEMA_signal_2861), .Z1_f (new_AGEMA_signal_2862) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_63_U1_XOR1_U1 ( .A0_t (IN_key_s0_t[127]), .A0_f (IN_key_s0_f[127]), .A1_t (IN_key_s1_t[127]), .A1_f (IN_key_s1_f[127]), .B0_t (IN_key_s0_t[63]), .B0_f (IN_key_s0_f[63]), .B1_t (IN_key_s1_t[63]), .B1_f (IN_key_s1_f[63]), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_63_U1_X), .Z0_f (new_AGEMA_signal_2467), .Z1_t (new_AGEMA_signal_2468), .Z1_f (new_AGEMA_signal_2469) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_63_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n31), .A1_f (new_AGEMA_signal_2477), .B0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_63_U1_X), .B0_f (new_AGEMA_signal_2467), .B1_t (new_AGEMA_signal_2468), .B1_f (new_AGEMA_signal_2469), .Z0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_63_U1_Y), .Z0_f (new_AGEMA_signal_2670), .Z1_t (new_AGEMA_signal_2671), .Z1_f (new_AGEMA_signal_2672) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_current_roundkey_mux_inst_63_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_current_roundkey_mux_inst_63_U1_Y), .A0_f (new_AGEMA_signal_2670), .A1_t (new_AGEMA_signal_2671), .A1_f (new_AGEMA_signal_2672), .B0_t (IN_key_s0_t[127]), .B0_f (IN_key_s0_f[127]), .B1_t (IN_key_s1_t[127]), .B1_f (IN_key_s1_f[127]), .Z0_t (LED_128_Instance_current_roundkey[63]), .Z0_f (new_AGEMA_signal_2863), .Z1_t (new_AGEMA_signal_2864), .Z1_f (new_AGEMA_signal_2865) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U64 ( .A0_t (OUT_ciphertext_s0_t[28]), .A0_f (OUT_ciphertext_s0_f[28]), .A1_t (OUT_ciphertext_s1_t[28]), .A1_f (OUT_ciphertext_s1_f[28]), .B0_t (LED_128_Instance_current_roundkey[28]), .B0_f (new_AGEMA_signal_2758), .B1_t (new_AGEMA_signal_2759), .B1_f (new_AGEMA_signal_2760), .Z0_t (LED_128_Instance_addroundkey_tmp[28]), .Z0_f (new_AGEMA_signal_2871), .Z1_t (new_AGEMA_signal_2872), .Z1_f (new_AGEMA_signal_2873) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U63 ( .A0_t (OUT_ciphertext_s0_t[24]), .A0_f (OUT_ciphertext_s0_f[24]), .A1_t (OUT_ciphertext_s1_t[24]), .A1_f (OUT_ciphertext_s1_f[24]), .B0_t (LED_128_Instance_current_roundkey[24]), .B0_f (new_AGEMA_signal_2746), .B1_t (new_AGEMA_signal_2747), .B1_f (new_AGEMA_signal_2748), .Z0_t (LED_128_Instance_addroundkey_tmp[24]), .Z0_f (new_AGEMA_signal_2877), .Z1_t (new_AGEMA_signal_2878), .Z1_f (new_AGEMA_signal_2879) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U62 ( .A0_t (OUT_ciphertext_s0_t[12]), .A0_f (OUT_ciphertext_s0_f[12]), .A1_t (OUT_ciphertext_s1_t[12]), .A1_f (OUT_ciphertext_s1_f[12]), .B0_t (LED_128_Instance_current_roundkey[12]), .B0_f (new_AGEMA_signal_2710), .B1_t (new_AGEMA_signal_2711), .B1_f (new_AGEMA_signal_2712), .Z0_t (LED_128_Instance_addroundkey_tmp[12]), .Z0_f (new_AGEMA_signal_2883), .Z1_t (new_AGEMA_signal_2884), .Z1_f (new_AGEMA_signal_2885) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U61 ( .A0_t (OUT_ciphertext_s0_t[8]), .A0_f (OUT_ciphertext_s0_f[8]), .A1_t (OUT_ciphertext_s1_t[8]), .A1_f (OUT_ciphertext_s1_f[8]), .B0_t (LED_128_Instance_current_roundkey[8]), .B0_f (new_AGEMA_signal_2698), .B1_t (new_AGEMA_signal_2699), .B1_f (new_AGEMA_signal_2700), .Z0_t (LED_128_Instance_addroundkey_tmp[8]), .Z0_f (new_AGEMA_signal_2889), .Z1_t (new_AGEMA_signal_2890), .Z1_f (new_AGEMA_signal_2891) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U60 ( .A0_t (OUT_ciphertext_s0_t[0]), .A0_f (OUT_ciphertext_s0_f[0]), .A1_t (OUT_ciphertext_s1_t[0]), .A1_f (OUT_ciphertext_s1_f[0]), .B0_t (LED_128_Instance_current_roundkey[0]), .B0_f (new_AGEMA_signal_2674), .B1_t (new_AGEMA_signal_2675), .B1_f (new_AGEMA_signal_2676), .Z0_t (LED_128_Instance_addroundkey_tmp[0]), .Z0_f (new_AGEMA_signal_2895), .Z1_t (new_AGEMA_signal_2896), .Z1_f (new_AGEMA_signal_2897) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U59 ( .A0_t (OUT_ciphertext_s0_t[48]), .A0_f (OUT_ciphertext_s0_f[48]), .A1_t (OUT_ciphertext_s1_t[48]), .A1_f (OUT_ciphertext_s1_f[48]), .B0_t (LED_128_Instance_current_roundkey[48]), .B0_f (new_AGEMA_signal_2818), .B1_t (new_AGEMA_signal_2819), .B1_f (new_AGEMA_signal_2820), .Z0_t (LED_128_Instance_addroundkey_tmp[48]), .Z0_f (new_AGEMA_signal_2901), .Z1_t (new_AGEMA_signal_2902), .Z1_f (new_AGEMA_signal_2903) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U58 ( .A0_t (OUT_ciphertext_s0_t[16]), .A0_f (OUT_ciphertext_s0_f[16]), .A1_t (OUT_ciphertext_s1_t[16]), .A1_f (OUT_ciphertext_s1_f[16]), .B0_t (LED_128_Instance_current_roundkey[16]), .B0_f (new_AGEMA_signal_2722), .B1_t (new_AGEMA_signal_2723), .B1_f (new_AGEMA_signal_2724), .Z0_t (LED_128_Instance_addroundkey_tmp[16]), .Z0_f (new_AGEMA_signal_2907), .Z1_t (new_AGEMA_signal_2908), .Z1_f (new_AGEMA_signal_2909) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U57 ( .A0_t (OUT_ciphertext_s0_t[56]), .A0_f (OUT_ciphertext_s0_f[56]), .A1_t (OUT_ciphertext_s1_t[56]), .A1_f (OUT_ciphertext_s1_f[56]), .B0_t (LED_128_Instance_current_roundkey[56]), .B0_f (new_AGEMA_signal_2842), .B1_t (new_AGEMA_signal_2843), .B1_f (new_AGEMA_signal_2844), .Z0_t (LED_128_Instance_addroundkey_tmp[56]), .Z0_f (new_AGEMA_signal_2913), .Z1_t (new_AGEMA_signal_2914), .Z1_f (new_AGEMA_signal_2915) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U56 ( .A0_t (OUT_ciphertext_s0_t[60]), .A0_f (OUT_ciphertext_s0_f[60]), .A1_t (OUT_ciphertext_s1_t[60]), .A1_f (OUT_ciphertext_s1_f[60]), .B0_t (LED_128_Instance_current_roundkey[60]), .B0_f (new_AGEMA_signal_2854), .B1_t (new_AGEMA_signal_2855), .B1_f (new_AGEMA_signal_2856), .Z0_t (LED_128_Instance_addroundkey_tmp[60]), .Z0_f (new_AGEMA_signal_2919), .Z1_t (new_AGEMA_signal_2920), .Z1_f (new_AGEMA_signal_2921) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U55 ( .A0_t (OUT_ciphertext_s0_t[31]), .A0_f (OUT_ciphertext_s0_f[31]), .A1_t (OUT_ciphertext_s1_t[31]), .A1_f (OUT_ciphertext_s1_f[31]), .B0_t (LED_128_Instance_current_roundkey[31]), .B0_f (new_AGEMA_signal_2767), .B1_t (new_AGEMA_signal_2768), .B1_f (new_AGEMA_signal_2769), .Z0_t (LED_128_Instance_addroundkey_tmp[31]), .Z0_f (new_AGEMA_signal_2925), .Z1_t (new_AGEMA_signal_2926), .Z1_f (new_AGEMA_signal_2927) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U54 ( .A0_t (OUT_ciphertext_s0_t[27]), .A0_f (OUT_ciphertext_s0_f[27]), .A1_t (OUT_ciphertext_s1_t[27]), .A1_f (OUT_ciphertext_s1_f[27]), .B0_t (LED_128_Instance_current_roundkey[27]), .B0_f (new_AGEMA_signal_2755), .B1_t (new_AGEMA_signal_2756), .B1_f (new_AGEMA_signal_2757), .Z0_t (LED_128_Instance_addroundkey_tmp[27]), .Z0_f (new_AGEMA_signal_2931), .Z1_t (new_AGEMA_signal_2932), .Z1_f (new_AGEMA_signal_2933) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U53 ( .A0_t (OUT_ciphertext_s0_t[23]), .A0_f (OUT_ciphertext_s0_f[23]), .A1_t (OUT_ciphertext_s1_t[23]), .A1_f (OUT_ciphertext_s1_f[23]), .B0_t (LED_128_Instance_current_roundkey[23]), .B0_f (new_AGEMA_signal_2743), .B1_t (new_AGEMA_signal_2744), .B1_f (new_AGEMA_signal_2745), .Z0_t (LED_128_Instance_addroundkey_tmp[23]), .Z0_f (new_AGEMA_signal_2937), .Z1_t (new_AGEMA_signal_2938), .Z1_f (new_AGEMA_signal_2939) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U52 ( .A0_t (OUT_ciphertext_s0_t[32]), .A0_f (OUT_ciphertext_s0_f[32]), .A1_t (OUT_ciphertext_s1_t[32]), .A1_f (OUT_ciphertext_s1_f[32]), .B0_t (LED_128_Instance_current_roundkey[32]), .B0_f (new_AGEMA_signal_2770), .B1_t (new_AGEMA_signal_2771), .B1_f (new_AGEMA_signal_2772), .Z0_t (LED_128_Instance_addroundkey_tmp[32]), .Z0_f (new_AGEMA_signal_2943), .Z1_t (new_AGEMA_signal_2944), .Z1_f (new_AGEMA_signal_2945) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U51 ( .A0_t (OUT_ciphertext_s0_t[44]), .A0_f (OUT_ciphertext_s0_f[44]), .A1_t (OUT_ciphertext_s1_t[44]), .A1_f (OUT_ciphertext_s1_f[44]), .B0_t (LED_128_Instance_current_roundkey[44]), .B0_f (new_AGEMA_signal_2806), .B1_t (new_AGEMA_signal_2807), .B1_f (new_AGEMA_signal_2808), .Z0_t (LED_128_Instance_addroundkey_tmp[44]), .Z0_f (new_AGEMA_signal_2949), .Z1_t (new_AGEMA_signal_2950), .Z1_f (new_AGEMA_signal_2951) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U50 ( .A0_t (OUT_ciphertext_s0_t[40]), .A0_f (OUT_ciphertext_s0_f[40]), .A1_t (OUT_ciphertext_s1_t[40]), .A1_f (OUT_ciphertext_s1_f[40]), .B0_t (LED_128_Instance_current_roundkey[40]), .B0_f (new_AGEMA_signal_2794), .B1_t (new_AGEMA_signal_2795), .B1_f (new_AGEMA_signal_2796), .Z0_t (LED_128_Instance_addroundkey_tmp[40]), .Z0_f (new_AGEMA_signal_2955), .Z1_t (new_AGEMA_signal_2956), .Z1_f (new_AGEMA_signal_2957) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U49 ( .A0_t (OUT_ciphertext_s0_t[33]), .A0_f (OUT_ciphertext_s0_f[33]), .A1_t (OUT_ciphertext_s1_t[33]), .A1_f (OUT_ciphertext_s1_f[33]), .B0_t (LED_128_Instance_current_roundkey[33]), .B0_f (new_AGEMA_signal_2773), .B1_t (new_AGEMA_signal_2774), .B1_f (new_AGEMA_signal_2775), .Z0_t (LED_128_Instance_addroundkey_tmp[33]), .Z0_f (new_AGEMA_signal_2961), .Z1_t (new_AGEMA_signal_2962), .Z1_f (new_AGEMA_signal_2963) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U48 ( .A0_t (OUT_ciphertext_s0_t[49]), .A0_f (OUT_ciphertext_s0_f[49]), .A1_t (OUT_ciphertext_s1_t[49]), .A1_f (OUT_ciphertext_s1_f[49]), .B0_t (LED_128_Instance_current_roundkey[49]), .B0_f (new_AGEMA_signal_2821), .B1_t (new_AGEMA_signal_2822), .B1_f (new_AGEMA_signal_2823), .Z0_t (LED_128_Instance_addroundkey_tmp[49]), .Z0_f (new_AGEMA_signal_2967), .Z1_t (new_AGEMA_signal_2968), .Z1_f (new_AGEMA_signal_2969) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U47 ( .A0_t (OUT_ciphertext_s0_t[19]), .A0_f (OUT_ciphertext_s0_f[19]), .A1_t (OUT_ciphertext_s1_t[19]), .A1_f (OUT_ciphertext_s1_f[19]), .B0_t (LED_128_Instance_current_roundkey[19]), .B0_f (new_AGEMA_signal_2731), .B1_t (new_AGEMA_signal_2732), .B1_f (new_AGEMA_signal_2733), .Z0_t (LED_128_Instance_addroundkey_tmp[19]), .Z0_f (new_AGEMA_signal_2973), .Z1_t (new_AGEMA_signal_2974), .Z1_f (new_AGEMA_signal_2975) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U46 ( .A0_t (OUT_ciphertext_s0_t[3]), .A0_f (OUT_ciphertext_s0_f[3]), .A1_t (OUT_ciphertext_s1_t[3]), .A1_f (OUT_ciphertext_s1_f[3]), .B0_t (LED_128_Instance_current_roundkey[3]), .B0_f (new_AGEMA_signal_2683), .B1_t (new_AGEMA_signal_2684), .B1_f (new_AGEMA_signal_2685), .Z0_t (LED_128_Instance_addroundkey_tmp[3]), .Z0_f (new_AGEMA_signal_2979), .Z1_t (new_AGEMA_signal_2980), .Z1_f (new_AGEMA_signal_2981) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U45 ( .A0_t (OUT_ciphertext_s0_t[54]), .A0_f (OUT_ciphertext_s0_f[54]), .A1_t (OUT_ciphertext_s1_t[54]), .A1_f (OUT_ciphertext_s1_f[54]), .B0_t (LED_128_Instance_current_roundkey[54]), .B0_f (new_AGEMA_signal_2836), .B1_t (new_AGEMA_signal_2837), .B1_f (new_AGEMA_signal_2838), .Z0_t (LED_128_Instance_addroundkey_tmp[54]), .Z0_f (new_AGEMA_signal_2985), .Z1_t (new_AGEMA_signal_2986), .Z1_f (new_AGEMA_signal_2987) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U44 ( .A0_t (OUT_ciphertext_s0_t[38]), .A0_f (OUT_ciphertext_s0_f[38]), .A1_t (OUT_ciphertext_s1_t[38]), .A1_f (OUT_ciphertext_s1_f[38]), .B0_t (LED_128_Instance_current_roundkey[38]), .B0_f (new_AGEMA_signal_2788), .B1_t (new_AGEMA_signal_2789), .B1_f (new_AGEMA_signal_2790), .Z0_t (LED_128_Instance_addroundkey_tmp[38]), .Z0_f (new_AGEMA_signal_2991), .Z1_t (new_AGEMA_signal_2992), .Z1_f (new_AGEMA_signal_2993) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U43 ( .A0_t (OUT_ciphertext_s0_t[36]), .A0_f (OUT_ciphertext_s0_f[36]), .A1_t (OUT_ciphertext_s1_t[36]), .A1_f (OUT_ciphertext_s1_f[36]), .B0_t (LED_128_Instance_current_roundkey[36]), .B0_f (new_AGEMA_signal_2782), .B1_t (new_AGEMA_signal_2783), .B1_f (new_AGEMA_signal_2784), .Z0_t (LED_128_Instance_addroundkey_tmp[36]), .Z0_f (new_AGEMA_signal_2997), .Z1_t (new_AGEMA_signal_2998), .Z1_f (new_AGEMA_signal_2999) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U42 ( .A0_t (OUT_ciphertext_s0_t[52]), .A0_f (OUT_ciphertext_s0_f[52]), .A1_t (OUT_ciphertext_s1_t[52]), .A1_f (OUT_ciphertext_s1_f[52]), .B0_t (LED_128_Instance_current_roundkey[52]), .B0_f (new_AGEMA_signal_2830), .B1_t (new_AGEMA_signal_2831), .B1_f (new_AGEMA_signal_2832), .Z0_t (LED_128_Instance_addroundkey_tmp[52]), .Z0_f (new_AGEMA_signal_3003), .Z1_t (new_AGEMA_signal_3004), .Z1_f (new_AGEMA_signal_3005) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U41 ( .A0_t (OUT_ciphertext_s0_t[37]), .A0_f (OUT_ciphertext_s0_f[37]), .A1_t (OUT_ciphertext_s1_t[37]), .A1_f (OUT_ciphertext_s1_f[37]), .B0_t (LED_128_Instance_current_roundkey[37]), .B0_f (new_AGEMA_signal_2785), .B1_t (new_AGEMA_signal_2786), .B1_f (new_AGEMA_signal_2787), .Z0_t (LED_128_Instance_addroundkey_tmp[37]), .Z0_f (new_AGEMA_signal_3009), .Z1_t (new_AGEMA_signal_3010), .Z1_f (new_AGEMA_signal_3011) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U40 ( .A0_t (OUT_ciphertext_s0_t[53]), .A0_f (OUT_ciphertext_s0_f[53]), .A1_t (OUT_ciphertext_s1_t[53]), .A1_f (OUT_ciphertext_s1_f[53]), .B0_t (LED_128_Instance_current_roundkey[53]), .B0_f (new_AGEMA_signal_2833), .B1_t (new_AGEMA_signal_2834), .B1_f (new_AGEMA_signal_2835), .Z0_t (LED_128_Instance_addroundkey_tmp[53]), .Z0_f (new_AGEMA_signal_3015), .Z1_t (new_AGEMA_signal_3016), .Z1_f (new_AGEMA_signal_3017) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U39 ( .A0_t (OUT_ciphertext_s0_t[4]), .A0_f (OUT_ciphertext_s0_f[4]), .A1_t (OUT_ciphertext_s1_t[4]), .A1_f (OUT_ciphertext_s1_f[4]), .B0_t (LED_128_Instance_current_roundkey[4]), .B0_f (new_AGEMA_signal_2686), .B1_t (new_AGEMA_signal_2687), .B1_f (new_AGEMA_signal_2688), .Z0_t (LED_128_Instance_addroundkey_tmp[4]), .Z0_f (new_AGEMA_signal_3021), .Z1_t (new_AGEMA_signal_3022), .Z1_f (new_AGEMA_signal_3023) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U38 ( .A0_t (OUT_ciphertext_s0_t[6]), .A0_f (OUT_ciphertext_s0_f[6]), .A1_t (OUT_ciphertext_s1_t[6]), .A1_f (OUT_ciphertext_s1_f[6]), .B0_t (LED_128_Instance_current_roundkey[6]), .B0_f (new_AGEMA_signal_2692), .B1_t (new_AGEMA_signal_2693), .B1_f (new_AGEMA_signal_2694), .Z0_t (LED_128_Instance_addroundkey_tmp[6]), .Z0_f (new_AGEMA_signal_3027), .Z1_t (new_AGEMA_signal_3028), .Z1_f (new_AGEMA_signal_3029) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U37 ( .A0_t (OUT_ciphertext_s0_t[20]), .A0_f (OUT_ciphertext_s0_f[20]), .A1_t (OUT_ciphertext_s1_t[20]), .A1_f (OUT_ciphertext_s1_f[20]), .B0_t (LED_128_Instance_current_roundkey[20]), .B0_f (new_AGEMA_signal_2734), .B1_t (new_AGEMA_signal_2735), .B1_f (new_AGEMA_signal_2736), .Z0_t (LED_128_Instance_addroundkey_tmp[20]), .Z0_f (new_AGEMA_signal_3033), .Z1_t (new_AGEMA_signal_3034), .Z1_f (new_AGEMA_signal_3035) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U36 ( .A0_t (OUT_ciphertext_s0_t[22]), .A0_f (OUT_ciphertext_s0_f[22]), .A1_t (OUT_ciphertext_s1_t[22]), .A1_f (OUT_ciphertext_s1_f[22]), .B0_t (LED_128_Instance_current_roundkey[22]), .B0_f (new_AGEMA_signal_2740), .B1_t (new_AGEMA_signal_2741), .B1_f (new_AGEMA_signal_2742), .Z0_t (LED_128_Instance_addroundkey_tmp[22]), .Z0_f (new_AGEMA_signal_3039), .Z1_t (new_AGEMA_signal_3040), .Z1_f (new_AGEMA_signal_3041) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U35 ( .A0_t (OUT_ciphertext_s0_t[5]), .A0_f (OUT_ciphertext_s0_f[5]), .A1_t (OUT_ciphertext_s1_t[5]), .A1_f (OUT_ciphertext_s1_f[5]), .B0_t (LED_128_Instance_current_roundkey[5]), .B0_f (new_AGEMA_signal_2689), .B1_t (new_AGEMA_signal_2690), .B1_f (new_AGEMA_signal_2691), .Z0_t (LED_128_Instance_addroundkey_tmp[5]), .Z0_f (new_AGEMA_signal_3045), .Z1_t (new_AGEMA_signal_3046), .Z1_f (new_AGEMA_signal_3047) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U34 ( .A0_t (OUT_ciphertext_s0_t[21]), .A0_f (OUT_ciphertext_s0_f[21]), .A1_t (OUT_ciphertext_s1_t[21]), .A1_f (OUT_ciphertext_s1_f[21]), .B0_t (LED_128_Instance_current_roundkey[21]), .B0_f (new_AGEMA_signal_2737), .B1_t (new_AGEMA_signal_2738), .B1_f (new_AGEMA_signal_2739), .Z0_t (LED_128_Instance_addroundkey_tmp[21]), .Z0_f (new_AGEMA_signal_3051), .Z1_t (new_AGEMA_signal_3052), .Z1_f (new_AGEMA_signal_3053) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U33 ( .A0_t (OUT_ciphertext_s0_t[58]), .A0_f (OUT_ciphertext_s0_f[58]), .A1_t (OUT_ciphertext_s1_t[58]), .A1_f (OUT_ciphertext_s1_f[58]), .B0_t (LED_128_Instance_current_roundkey[58]), .B0_f (new_AGEMA_signal_2848), .B1_t (new_AGEMA_signal_2849), .B1_f (new_AGEMA_signal_2850), .Z0_t (LED_128_Instance_addroundkey_tmp[58]), .Z0_f (new_AGEMA_signal_3057), .Z1_t (new_AGEMA_signal_3058), .Z1_f (new_AGEMA_signal_3059) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U32 ( .A0_t (OUT_ciphertext_s0_t[50]), .A0_f (OUT_ciphertext_s0_f[50]), .A1_t (OUT_ciphertext_s1_t[50]), .A1_f (OUT_ciphertext_s1_f[50]), .B0_t (LED_128_Instance_current_roundkey[50]), .B0_f (new_AGEMA_signal_2824), .B1_t (new_AGEMA_signal_2825), .B1_f (new_AGEMA_signal_2826), .Z0_t (LED_128_Instance_addroundkey_tmp[50]), .Z0_f (new_AGEMA_signal_3063), .Z1_t (new_AGEMA_signal_3064), .Z1_f (new_AGEMA_signal_3065) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U31 ( .A0_t (OUT_ciphertext_s0_t[62]), .A0_f (OUT_ciphertext_s0_f[62]), .A1_t (OUT_ciphertext_s1_t[62]), .A1_f (OUT_ciphertext_s1_f[62]), .B0_t (LED_128_Instance_current_roundkey[62]), .B0_f (new_AGEMA_signal_2860), .B1_t (new_AGEMA_signal_2861), .B1_f (new_AGEMA_signal_2862), .Z0_t (LED_128_Instance_addroundkey_tmp[62]), .Z0_f (new_AGEMA_signal_3069), .Z1_t (new_AGEMA_signal_3070), .Z1_f (new_AGEMA_signal_3071) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U30 ( .A0_t (OUT_ciphertext_s0_t[34]), .A0_f (OUT_ciphertext_s0_f[34]), .A1_t (OUT_ciphertext_s1_t[34]), .A1_f (OUT_ciphertext_s1_f[34]), .B0_t (LED_128_Instance_current_roundkey[34]), .B0_f (new_AGEMA_signal_2776), .B1_t (new_AGEMA_signal_2777), .B1_f (new_AGEMA_signal_2778), .Z0_t (LED_128_Instance_addroundkey_tmp[34]), .Z0_f (new_AGEMA_signal_3075), .Z1_t (new_AGEMA_signal_3076), .Z1_f (new_AGEMA_signal_3077) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U29 ( .A0_t (OUT_ciphertext_s0_t[46]), .A0_f (OUT_ciphertext_s0_f[46]), .A1_t (OUT_ciphertext_s1_t[46]), .A1_f (OUT_ciphertext_s1_f[46]), .B0_t (LED_128_Instance_current_roundkey[46]), .B0_f (new_AGEMA_signal_2812), .B1_t (new_AGEMA_signal_2813), .B1_f (new_AGEMA_signal_2814), .Z0_t (LED_128_Instance_addroundkey_tmp[46]), .Z0_f (new_AGEMA_signal_3081), .Z1_t (new_AGEMA_signal_3082), .Z1_f (new_AGEMA_signal_3083) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U28 ( .A0_t (OUT_ciphertext_s0_t[42]), .A0_f (OUT_ciphertext_s0_f[42]), .A1_t (OUT_ciphertext_s1_t[42]), .A1_f (OUT_ciphertext_s1_f[42]), .B0_t (LED_128_Instance_current_roundkey[42]), .B0_f (new_AGEMA_signal_2800), .B1_t (new_AGEMA_signal_2801), .B1_f (new_AGEMA_signal_2802), .Z0_t (LED_128_Instance_addroundkey_tmp[42]), .Z0_f (new_AGEMA_signal_3087), .Z1_t (new_AGEMA_signal_3088), .Z1_f (new_AGEMA_signal_3089) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U27 ( .A0_t (OUT_ciphertext_s0_t[14]), .A0_f (OUT_ciphertext_s0_f[14]), .A1_t (OUT_ciphertext_s1_t[14]), .A1_f (OUT_ciphertext_s1_f[14]), .B0_t (LED_128_Instance_current_roundkey[14]), .B0_f (new_AGEMA_signal_2716), .B1_t (new_AGEMA_signal_2717), .B1_f (new_AGEMA_signal_2718), .Z0_t (LED_128_Instance_addroundkey_tmp[14]), .Z0_f (new_AGEMA_signal_3093), .Z1_t (new_AGEMA_signal_3094), .Z1_f (new_AGEMA_signal_3095) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U26 ( .A0_t (OUT_ciphertext_s0_t[18]), .A0_f (OUT_ciphertext_s0_f[18]), .A1_t (OUT_ciphertext_s1_t[18]), .A1_f (OUT_ciphertext_s1_f[18]), .B0_t (LED_128_Instance_current_roundkey[18]), .B0_f (new_AGEMA_signal_2728), .B1_t (new_AGEMA_signal_2729), .B1_f (new_AGEMA_signal_2730), .Z0_t (LED_128_Instance_addroundkey_tmp[18]), .Z0_f (new_AGEMA_signal_3099), .Z1_t (new_AGEMA_signal_3100), .Z1_f (new_AGEMA_signal_3101) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U25 ( .A0_t (OUT_ciphertext_s0_t[10]), .A0_f (OUT_ciphertext_s0_f[10]), .A1_t (OUT_ciphertext_s1_t[10]), .A1_f (OUT_ciphertext_s1_f[10]), .B0_t (LED_128_Instance_current_roundkey[10]), .B0_f (new_AGEMA_signal_2704), .B1_t (new_AGEMA_signal_2705), .B1_f (new_AGEMA_signal_2706), .Z0_t (LED_128_Instance_addroundkey_tmp[10]), .Z0_f (new_AGEMA_signal_3105), .Z1_t (new_AGEMA_signal_3106), .Z1_f (new_AGEMA_signal_3107) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U24 ( .A0_t (OUT_ciphertext_s0_t[30]), .A0_f (OUT_ciphertext_s0_f[30]), .A1_t (OUT_ciphertext_s1_t[30]), .A1_f (OUT_ciphertext_s1_f[30]), .B0_t (LED_128_Instance_current_roundkey[30]), .B0_f (new_AGEMA_signal_2764), .B1_t (new_AGEMA_signal_2765), .B1_f (new_AGEMA_signal_2766), .Z0_t (LED_128_Instance_addroundkey_tmp[30]), .Z0_f (new_AGEMA_signal_3111), .Z1_t (new_AGEMA_signal_3112), .Z1_f (new_AGEMA_signal_3113) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U23 ( .A0_t (OUT_ciphertext_s0_t[26]), .A0_f (OUT_ciphertext_s0_f[26]), .A1_t (OUT_ciphertext_s1_t[26]), .A1_f (OUT_ciphertext_s1_f[26]), .B0_t (LED_128_Instance_current_roundkey[26]), .B0_f (new_AGEMA_signal_2752), .B1_t (new_AGEMA_signal_2753), .B1_f (new_AGEMA_signal_2754), .Z0_t (LED_128_Instance_addroundkey_tmp[26]), .Z0_f (new_AGEMA_signal_3117), .Z1_t (new_AGEMA_signal_3118), .Z1_f (new_AGEMA_signal_3119) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U22 ( .A0_t (OUT_ciphertext_s0_t[2]), .A0_f (OUT_ciphertext_s0_f[2]), .A1_t (OUT_ciphertext_s1_t[2]), .A1_f (OUT_ciphertext_s1_f[2]), .B0_t (LED_128_Instance_current_roundkey[2]), .B0_f (new_AGEMA_signal_2680), .B1_t (new_AGEMA_signal_2681), .B1_f (new_AGEMA_signal_2682), .Z0_t (LED_128_Instance_addroundkey_tmp[2]), .Z0_f (new_AGEMA_signal_3123), .Z1_t (new_AGEMA_signal_3124), .Z1_f (new_AGEMA_signal_3125) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U21 ( .A0_t (OUT_ciphertext_s0_t[45]), .A0_f (OUT_ciphertext_s0_f[45]), .A1_t (OUT_ciphertext_s1_t[45]), .A1_f (OUT_ciphertext_s1_f[45]), .B0_t (LED_128_Instance_current_roundkey[45]), .B0_f (new_AGEMA_signal_2809), .B1_t (new_AGEMA_signal_2810), .B1_f (new_AGEMA_signal_2811), .Z0_t (LED_128_Instance_addroundkey_tmp[45]), .Z0_f (new_AGEMA_signal_3129), .Z1_t (new_AGEMA_signal_3130), .Z1_f (new_AGEMA_signal_3131) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U20 ( .A0_t (OUT_ciphertext_s0_t[41]), .A0_f (OUT_ciphertext_s0_f[41]), .A1_t (OUT_ciphertext_s1_t[41]), .A1_f (OUT_ciphertext_s1_f[41]), .B0_t (LED_128_Instance_current_roundkey[41]), .B0_f (new_AGEMA_signal_2797), .B1_t (new_AGEMA_signal_2798), .B1_f (new_AGEMA_signal_2799), .Z0_t (LED_128_Instance_addroundkey_tmp[41]), .Z0_f (new_AGEMA_signal_3135), .Z1_t (new_AGEMA_signal_3136), .Z1_f (new_AGEMA_signal_3137) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U19 ( .A0_t (OUT_ciphertext_s0_t[57]), .A0_f (OUT_ciphertext_s0_f[57]), .A1_t (OUT_ciphertext_s1_t[57]), .A1_f (OUT_ciphertext_s1_f[57]), .B0_t (LED_128_Instance_current_roundkey[57]), .B0_f (new_AGEMA_signal_2845), .B1_t (new_AGEMA_signal_2846), .B1_f (new_AGEMA_signal_2847), .Z0_t (LED_128_Instance_addroundkey_tmp[57]), .Z0_f (new_AGEMA_signal_3141), .Z1_t (new_AGEMA_signal_3142), .Z1_f (new_AGEMA_signal_3143) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U18 ( .A0_t (OUT_ciphertext_s0_t[61]), .A0_f (OUT_ciphertext_s0_f[61]), .A1_t (OUT_ciphertext_s1_t[61]), .A1_f (OUT_ciphertext_s1_f[61]), .B0_t (LED_128_Instance_current_roundkey[61]), .B0_f (new_AGEMA_signal_2857), .B1_t (new_AGEMA_signal_2858), .B1_f (new_AGEMA_signal_2859), .Z0_t (LED_128_Instance_addroundkey_tmp[61]), .Z0_f (new_AGEMA_signal_3147), .Z1_t (new_AGEMA_signal_3148), .Z1_f (new_AGEMA_signal_3149) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U17 ( .A0_t (OUT_ciphertext_s0_t[13]), .A0_f (OUT_ciphertext_s0_f[13]), .A1_t (OUT_ciphertext_s1_t[13]), .A1_f (OUT_ciphertext_s1_f[13]), .B0_t (LED_128_Instance_current_roundkey[13]), .B0_f (new_AGEMA_signal_2713), .B1_t (new_AGEMA_signal_2714), .B1_f (new_AGEMA_signal_2715), .Z0_t (LED_128_Instance_addroundkey_tmp[13]), .Z0_f (new_AGEMA_signal_3153), .Z1_t (new_AGEMA_signal_3154), .Z1_f (new_AGEMA_signal_3155) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U16 ( .A0_t (OUT_ciphertext_s0_t[17]), .A0_f (OUT_ciphertext_s0_f[17]), .A1_t (OUT_ciphertext_s1_t[17]), .A1_f (OUT_ciphertext_s1_f[17]), .B0_t (LED_128_Instance_current_roundkey[17]), .B0_f (new_AGEMA_signal_2725), .B1_t (new_AGEMA_signal_2726), .B1_f (new_AGEMA_signal_2727), .Z0_t (LED_128_Instance_addroundkey_tmp[17]), .Z0_f (new_AGEMA_signal_3159), .Z1_t (new_AGEMA_signal_3160), .Z1_f (new_AGEMA_signal_3161) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U15 ( .A0_t (OUT_ciphertext_s0_t[9]), .A0_f (OUT_ciphertext_s0_f[9]), .A1_t (OUT_ciphertext_s1_t[9]), .A1_f (OUT_ciphertext_s1_f[9]), .B0_t (LED_128_Instance_current_roundkey[9]), .B0_f (new_AGEMA_signal_2701), .B1_t (new_AGEMA_signal_2702), .B1_f (new_AGEMA_signal_2703), .Z0_t (LED_128_Instance_addroundkey_tmp[9]), .Z0_f (new_AGEMA_signal_3165), .Z1_t (new_AGEMA_signal_3166), .Z1_f (new_AGEMA_signal_3167) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U14 ( .A0_t (OUT_ciphertext_s0_t[29]), .A0_f (OUT_ciphertext_s0_f[29]), .A1_t (OUT_ciphertext_s1_t[29]), .A1_f (OUT_ciphertext_s1_f[29]), .B0_t (LED_128_Instance_current_roundkey[29]), .B0_f (new_AGEMA_signal_2761), .B1_t (new_AGEMA_signal_2762), .B1_f (new_AGEMA_signal_2763), .Z0_t (LED_128_Instance_addroundkey_tmp[29]), .Z0_f (new_AGEMA_signal_3171), .Z1_t (new_AGEMA_signal_3172), .Z1_f (new_AGEMA_signal_3173) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U13 ( .A0_t (OUT_ciphertext_s0_t[25]), .A0_f (OUT_ciphertext_s0_f[25]), .A1_t (OUT_ciphertext_s1_t[25]), .A1_f (OUT_ciphertext_s1_f[25]), .B0_t (LED_128_Instance_current_roundkey[25]), .B0_f (new_AGEMA_signal_2749), .B1_t (new_AGEMA_signal_2750), .B1_f (new_AGEMA_signal_2751), .Z0_t (LED_128_Instance_addroundkey_tmp[25]), .Z0_f (new_AGEMA_signal_3177), .Z1_t (new_AGEMA_signal_3178), .Z1_f (new_AGEMA_signal_3179) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U12 ( .A0_t (OUT_ciphertext_s0_t[1]), .A0_f (OUT_ciphertext_s0_f[1]), .A1_t (OUT_ciphertext_s1_t[1]), .A1_f (OUT_ciphertext_s1_f[1]), .B0_t (LED_128_Instance_current_roundkey[1]), .B0_f (new_AGEMA_signal_2677), .B1_t (new_AGEMA_signal_2678), .B1_f (new_AGEMA_signal_2679), .Z0_t (LED_128_Instance_addroundkey_tmp[1]), .Z0_f (new_AGEMA_signal_3183), .Z1_t (new_AGEMA_signal_3184), .Z1_f (new_AGEMA_signal_3185) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U11 ( .A0_t (OUT_ciphertext_s0_t[39]), .A0_f (OUT_ciphertext_s0_f[39]), .A1_t (OUT_ciphertext_s1_t[39]), .A1_f (OUT_ciphertext_s1_f[39]), .B0_t (LED_128_Instance_current_roundkey[39]), .B0_f (new_AGEMA_signal_2791), .B1_t (new_AGEMA_signal_2792), .B1_f (new_AGEMA_signal_2793), .Z0_t (LED_128_Instance_addroundkey_tmp[39]), .Z0_f (new_AGEMA_signal_3189), .Z1_t (new_AGEMA_signal_3190), .Z1_f (new_AGEMA_signal_3191) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U10 ( .A0_t (OUT_ciphertext_s0_t[35]), .A0_f (OUT_ciphertext_s0_f[35]), .A1_t (OUT_ciphertext_s1_t[35]), .A1_f (OUT_ciphertext_s1_f[35]), .B0_t (LED_128_Instance_current_roundkey[35]), .B0_f (new_AGEMA_signal_2779), .B1_t (new_AGEMA_signal_2780), .B1_f (new_AGEMA_signal_2781), .Z0_t (LED_128_Instance_addroundkey_tmp[35]), .Z0_f (new_AGEMA_signal_3195), .Z1_t (new_AGEMA_signal_3196), .Z1_f (new_AGEMA_signal_3197) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U9 ( .A0_t (OUT_ciphertext_s0_t[47]), .A0_f (OUT_ciphertext_s0_f[47]), .A1_t (OUT_ciphertext_s1_t[47]), .A1_f (OUT_ciphertext_s1_f[47]), .B0_t (LED_128_Instance_current_roundkey[47]), .B0_f (new_AGEMA_signal_2815), .B1_t (new_AGEMA_signal_2816), .B1_f (new_AGEMA_signal_2817), .Z0_t (LED_128_Instance_addroundkey_tmp[47]), .Z0_f (new_AGEMA_signal_3201), .Z1_t (new_AGEMA_signal_3202), .Z1_f (new_AGEMA_signal_3203) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U8 ( .A0_t (OUT_ciphertext_s0_t[43]), .A0_f (OUT_ciphertext_s0_f[43]), .A1_t (OUT_ciphertext_s1_t[43]), .A1_f (OUT_ciphertext_s1_f[43]), .B0_t (LED_128_Instance_current_roundkey[43]), .B0_f (new_AGEMA_signal_2803), .B1_t (new_AGEMA_signal_2804), .B1_f (new_AGEMA_signal_2805), .Z0_t (LED_128_Instance_addroundkey_tmp[43]), .Z0_f (new_AGEMA_signal_3207), .Z1_t (new_AGEMA_signal_3208), .Z1_f (new_AGEMA_signal_3209) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U7 ( .A0_t (OUT_ciphertext_s0_t[59]), .A0_f (OUT_ciphertext_s0_f[59]), .A1_t (OUT_ciphertext_s1_t[59]), .A1_f (OUT_ciphertext_s1_f[59]), .B0_t (LED_128_Instance_current_roundkey[59]), .B0_f (new_AGEMA_signal_2851), .B1_t (new_AGEMA_signal_2852), .B1_f (new_AGEMA_signal_2853), .Z0_t (LED_128_Instance_addroundkey_tmp[59]), .Z0_f (new_AGEMA_signal_3213), .Z1_t (new_AGEMA_signal_3214), .Z1_f (new_AGEMA_signal_3215) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U6 ( .A0_t (OUT_ciphertext_s0_t[55]), .A0_f (OUT_ciphertext_s0_f[55]), .A1_t (OUT_ciphertext_s1_t[55]), .A1_f (OUT_ciphertext_s1_f[55]), .B0_t (LED_128_Instance_current_roundkey[55]), .B0_f (new_AGEMA_signal_2839), .B1_t (new_AGEMA_signal_2840), .B1_f (new_AGEMA_signal_2841), .Z0_t (LED_128_Instance_addroundkey_tmp[55]), .Z0_f (new_AGEMA_signal_3219), .Z1_t (new_AGEMA_signal_3220), .Z1_f (new_AGEMA_signal_3221) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U5 ( .A0_t (OUT_ciphertext_s0_t[51]), .A0_f (OUT_ciphertext_s0_f[51]), .A1_t (OUT_ciphertext_s1_t[51]), .A1_f (OUT_ciphertext_s1_f[51]), .B0_t (LED_128_Instance_current_roundkey[51]), .B0_f (new_AGEMA_signal_2827), .B1_t (new_AGEMA_signal_2828), .B1_f (new_AGEMA_signal_2829), .Z0_t (LED_128_Instance_addroundkey_tmp[51]), .Z0_f (new_AGEMA_signal_3225), .Z1_t (new_AGEMA_signal_3226), .Z1_f (new_AGEMA_signal_3227) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U4 ( .A0_t (OUT_ciphertext_s0_t[63]), .A0_f (OUT_ciphertext_s0_f[63]), .A1_t (OUT_ciphertext_s1_t[63]), .A1_f (OUT_ciphertext_s1_f[63]), .B0_t (LED_128_Instance_current_roundkey[63]), .B0_f (new_AGEMA_signal_2863), .B1_t (new_AGEMA_signal_2864), .B1_f (new_AGEMA_signal_2865), .Z0_t (LED_128_Instance_addroundkey_tmp[63]), .Z0_f (new_AGEMA_signal_3231), .Z1_t (new_AGEMA_signal_3232), .Z1_f (new_AGEMA_signal_3233) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U3 ( .A0_t (OUT_ciphertext_s0_t[15]), .A0_f (OUT_ciphertext_s0_f[15]), .A1_t (OUT_ciphertext_s1_t[15]), .A1_f (OUT_ciphertext_s1_f[15]), .B0_t (LED_128_Instance_current_roundkey[15]), .B0_f (new_AGEMA_signal_2719), .B1_t (new_AGEMA_signal_2720), .B1_f (new_AGEMA_signal_2721), .Z0_t (LED_128_Instance_addroundkey_tmp[15]), .Z0_f (new_AGEMA_signal_3237), .Z1_t (new_AGEMA_signal_3238), .Z1_f (new_AGEMA_signal_3239) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U2 ( .A0_t (OUT_ciphertext_s0_t[11]), .A0_f (OUT_ciphertext_s0_f[11]), .A1_t (OUT_ciphertext_s1_t[11]), .A1_f (OUT_ciphertext_s1_f[11]), .B0_t (LED_128_Instance_current_roundkey[11]), .B0_f (new_AGEMA_signal_2707), .B1_t (new_AGEMA_signal_2708), .B1_f (new_AGEMA_signal_2709), .Z0_t (LED_128_Instance_addroundkey_tmp[11]), .Z0_f (new_AGEMA_signal_3243), .Z1_t (new_AGEMA_signal_3244), .Z1_f (new_AGEMA_signal_3245) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_addRoundKey_instance_U1 ( .A0_t (OUT_ciphertext_s0_t[7]), .A0_f (OUT_ciphertext_s0_f[7]), .A1_t (OUT_ciphertext_s1_t[7]), .A1_f (OUT_ciphertext_s1_f[7]), .B0_t (LED_128_Instance_current_roundkey[7]), .B0_f (new_AGEMA_signal_2695), .B1_t (new_AGEMA_signal_2696), .B1_f (new_AGEMA_signal_2697), .Z0_t (LED_128_Instance_addroundkey_tmp[7]), .Z0_f (new_AGEMA_signal_3249), .Z1_t (new_AGEMA_signal_3250), .Z1_f (new_AGEMA_signal_3251) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_0_U1_XOR1_U1 ( .A0_t (OUT_ciphertext_s0_t[0]), .A0_f (OUT_ciphertext_s0_f[0]), .A1_t (OUT_ciphertext_s1_t[0]), .A1_f (OUT_ciphertext_s1_f[0]), .B0_t (LED_128_Instance_addroundkey_tmp[0]), .B0_f (new_AGEMA_signal_2895), .B1_t (new_AGEMA_signal_2896), .B1_f (new_AGEMA_signal_2897), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_0_U1_X), .Z0_f (new_AGEMA_signal_3252), .Z1_t (new_AGEMA_signal_3253), .Z1_f (new_AGEMA_signal_3254) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_0_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n23), .A1_f (new_AGEMA_signal_2480), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_0_U1_X), .B0_f (new_AGEMA_signal_3252), .B1_t (new_AGEMA_signal_3253), .B1_f (new_AGEMA_signal_3254), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_0_U1_Y), .Z0_f (new_AGEMA_signal_3444), .Z1_t (new_AGEMA_signal_3445), .Z1_f (new_AGEMA_signal_3446) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_0_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_0_U1_Y), .A0_f (new_AGEMA_signal_3444), .A1_t (new_AGEMA_signal_3445), .A1_f (new_AGEMA_signal_3446), .B0_t (OUT_ciphertext_s0_t[0]), .B0_f (OUT_ciphertext_s0_f[0]), .B1_t (OUT_ciphertext_s1_t[0]), .B1_f (OUT_ciphertext_s1_f[0]), .Z0_t (LED_128_Instance_addconst_out[0]), .Z0_f (new_AGEMA_signal_3636), .Z1_t (new_AGEMA_signal_3637), .Z1_f (new_AGEMA_signal_3638) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_1_U1_XOR1_U1 ( .A0_t (OUT_ciphertext_s0_t[1]), .A0_f (OUT_ciphertext_s0_f[1]), .A1_t (OUT_ciphertext_s1_t[1]), .A1_f (OUT_ciphertext_s1_f[1]), .B0_t (LED_128_Instance_addroundkey_tmp[1]), .B0_f (new_AGEMA_signal_3183), .B1_t (new_AGEMA_signal_3184), .B1_f (new_AGEMA_signal_3185), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_1_U1_X), .Z0_f (new_AGEMA_signal_3255), .Z1_t (new_AGEMA_signal_3256), .Z1_f (new_AGEMA_signal_3257) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_1_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n23), .A1_f (new_AGEMA_signal_2480), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_1_U1_X), .B0_f (new_AGEMA_signal_3255), .B1_t (new_AGEMA_signal_3256), .B1_f (new_AGEMA_signal_3257), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_1_U1_Y), .Z0_f (new_AGEMA_signal_3447), .Z1_t (new_AGEMA_signal_3448), .Z1_f (new_AGEMA_signal_3449) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_1_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_1_U1_Y), .A0_f (new_AGEMA_signal_3447), .A1_t (new_AGEMA_signal_3448), .A1_f (new_AGEMA_signal_3449), .B0_t (OUT_ciphertext_s0_t[1]), .B0_f (OUT_ciphertext_s0_f[1]), .B1_t (OUT_ciphertext_s1_t[1]), .B1_f (OUT_ciphertext_s1_f[1]), .Z0_t (LED_128_Instance_addconst_out[1]), .Z0_f (new_AGEMA_signal_3639), .Z1_t (new_AGEMA_signal_3640), .Z1_f (new_AGEMA_signal_3641) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_2_U1_XOR1_U1 ( .A0_t (OUT_ciphertext_s0_t[2]), .A0_f (OUT_ciphertext_s0_f[2]), .A1_t (OUT_ciphertext_s1_t[2]), .A1_f (OUT_ciphertext_s1_f[2]), .B0_t (LED_128_Instance_addroundkey_tmp[2]), .B0_f (new_AGEMA_signal_3123), .B1_t (new_AGEMA_signal_3124), .B1_f (new_AGEMA_signal_3125), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_2_U1_X), .Z0_f (new_AGEMA_signal_3258), .Z1_t (new_AGEMA_signal_3259), .Z1_f (new_AGEMA_signal_3260) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_2_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n23), .A1_f (new_AGEMA_signal_2480), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_2_U1_X), .B0_f (new_AGEMA_signal_3258), .B1_t (new_AGEMA_signal_3259), .B1_f (new_AGEMA_signal_3260), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_2_U1_Y), .Z0_f (new_AGEMA_signal_3450), .Z1_t (new_AGEMA_signal_3451), .Z1_f (new_AGEMA_signal_3452) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_2_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_2_U1_Y), .A0_f (new_AGEMA_signal_3450), .A1_t (new_AGEMA_signal_3451), .A1_f (new_AGEMA_signal_3452), .B0_t (OUT_ciphertext_s0_t[2]), .B0_f (OUT_ciphertext_s0_f[2]), .B1_t (OUT_ciphertext_s1_t[2]), .B1_f (OUT_ciphertext_s1_f[2]), .Z0_t (LED_128_Instance_addconst_out[2]), .Z0_f (new_AGEMA_signal_3642), .Z1_t (new_AGEMA_signal_3643), .Z1_f (new_AGEMA_signal_3644) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_3_U1_XOR1_U1 ( .A0_t (OUT_ciphertext_s0_t[3]), .A0_f (OUT_ciphertext_s0_f[3]), .A1_t (OUT_ciphertext_s1_t[3]), .A1_f (OUT_ciphertext_s1_f[3]), .B0_t (LED_128_Instance_addroundkey_tmp[3]), .B0_f (new_AGEMA_signal_2979), .B1_t (new_AGEMA_signal_2980), .B1_f (new_AGEMA_signal_2981), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_3_U1_X), .Z0_f (new_AGEMA_signal_3261), .Z1_t (new_AGEMA_signal_3262), .Z1_f (new_AGEMA_signal_3263) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_3_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n23), .A1_f (new_AGEMA_signal_2480), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_3_U1_X), .B0_f (new_AGEMA_signal_3261), .B1_t (new_AGEMA_signal_3262), .B1_f (new_AGEMA_signal_3263), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_3_U1_Y), .Z0_f (new_AGEMA_signal_3453), .Z1_t (new_AGEMA_signal_3454), .Z1_f (new_AGEMA_signal_3455) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_3_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_3_U1_Y), .A0_f (new_AGEMA_signal_3453), .A1_t (new_AGEMA_signal_3454), .A1_f (new_AGEMA_signal_3455), .B0_t (OUT_ciphertext_s0_t[3]), .B0_f (OUT_ciphertext_s0_f[3]), .B1_t (OUT_ciphertext_s1_t[3]), .B1_f (OUT_ciphertext_s1_f[3]), .Z0_t (LED_128_Instance_addroundkey_out[3]), .Z0_f (new_AGEMA_signal_3645), .Z1_t (new_AGEMA_signal_3646), .Z1_f (new_AGEMA_signal_3647) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_4_U1_XOR1_U1 ( .A0_t (OUT_ciphertext_s0_t[4]), .A0_f (OUT_ciphertext_s0_f[4]), .A1_t (OUT_ciphertext_s1_t[4]), .A1_f (OUT_ciphertext_s1_f[4]), .B0_t (LED_128_Instance_addroundkey_tmp[4]), .B0_f (new_AGEMA_signal_3021), .B1_t (new_AGEMA_signal_3022), .B1_f (new_AGEMA_signal_3023), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_4_U1_X), .Z0_f (new_AGEMA_signal_3264), .Z1_t (new_AGEMA_signal_3265), .Z1_f (new_AGEMA_signal_3266) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_4_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n23), .A1_f (new_AGEMA_signal_2480), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_4_U1_X), .B0_f (new_AGEMA_signal_3264), .B1_t (new_AGEMA_signal_3265), .B1_f (new_AGEMA_signal_3266), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_4_U1_Y), .Z0_f (new_AGEMA_signal_3456), .Z1_t (new_AGEMA_signal_3457), .Z1_f (new_AGEMA_signal_3458) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_4_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_4_U1_Y), .A0_f (new_AGEMA_signal_3456), .A1_t (new_AGEMA_signal_3457), .A1_f (new_AGEMA_signal_3458), .B0_t (OUT_ciphertext_s0_t[4]), .B0_f (OUT_ciphertext_s0_f[4]), .B1_t (OUT_ciphertext_s1_t[4]), .B1_f (OUT_ciphertext_s1_f[4]), .Z0_t (LED_128_Instance_addroundkey_out[4]), .Z0_f (new_AGEMA_signal_3648), .Z1_t (new_AGEMA_signal_3649), .Z1_f (new_AGEMA_signal_3650) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_5_U1_XOR1_U1 ( .A0_t (OUT_ciphertext_s0_t[5]), .A0_f (OUT_ciphertext_s0_f[5]), .A1_t (OUT_ciphertext_s1_t[5]), .A1_f (OUT_ciphertext_s1_f[5]), .B0_t (LED_128_Instance_addroundkey_tmp[5]), .B0_f (new_AGEMA_signal_3045), .B1_t (new_AGEMA_signal_3046), .B1_f (new_AGEMA_signal_3047), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_5_U1_X), .Z0_f (new_AGEMA_signal_3267), .Z1_t (new_AGEMA_signal_3268), .Z1_f (new_AGEMA_signal_3269) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_5_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n23), .A1_f (new_AGEMA_signal_2480), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_5_U1_X), .B0_f (new_AGEMA_signal_3267), .B1_t (new_AGEMA_signal_3268), .B1_f (new_AGEMA_signal_3269), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_5_U1_Y), .Z0_f (new_AGEMA_signal_3459), .Z1_t (new_AGEMA_signal_3460), .Z1_f (new_AGEMA_signal_3461) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_5_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_5_U1_Y), .A0_f (new_AGEMA_signal_3459), .A1_t (new_AGEMA_signal_3460), .A1_f (new_AGEMA_signal_3461), .B0_t (OUT_ciphertext_s0_t[5]), .B0_f (OUT_ciphertext_s0_f[5]), .B1_t (OUT_ciphertext_s1_t[5]), .B1_f (OUT_ciphertext_s1_f[5]), .Z0_t (LED_128_Instance_addroundkey_out[5]), .Z0_f (new_AGEMA_signal_3651), .Z1_t (new_AGEMA_signal_3652), .Z1_f (new_AGEMA_signal_3653) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_6_U1_XOR1_U1 ( .A0_t (OUT_ciphertext_s0_t[6]), .A0_f (OUT_ciphertext_s0_f[6]), .A1_t (OUT_ciphertext_s1_t[6]), .A1_f (OUT_ciphertext_s1_f[6]), .B0_t (LED_128_Instance_addroundkey_tmp[6]), .B0_f (new_AGEMA_signal_3027), .B1_t (new_AGEMA_signal_3028), .B1_f (new_AGEMA_signal_3029), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_6_U1_X), .Z0_f (new_AGEMA_signal_3270), .Z1_t (new_AGEMA_signal_3271), .Z1_f (new_AGEMA_signal_3272) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_6_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n23), .A1_f (new_AGEMA_signal_2480), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_6_U1_X), .B0_f (new_AGEMA_signal_3270), .B1_t (new_AGEMA_signal_3271), .B1_f (new_AGEMA_signal_3272), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_6_U1_Y), .Z0_f (new_AGEMA_signal_3462), .Z1_t (new_AGEMA_signal_3463), .Z1_f (new_AGEMA_signal_3464) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_6_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_6_U1_Y), .A0_f (new_AGEMA_signal_3462), .A1_t (new_AGEMA_signal_3463), .A1_f (new_AGEMA_signal_3464), .B0_t (OUT_ciphertext_s0_t[6]), .B0_f (OUT_ciphertext_s0_f[6]), .B1_t (OUT_ciphertext_s1_t[6]), .B1_f (OUT_ciphertext_s1_f[6]), .Z0_t (LED_128_Instance_addroundkey_out[6]), .Z0_f (new_AGEMA_signal_3654), .Z1_t (new_AGEMA_signal_3655), .Z1_f (new_AGEMA_signal_3656) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_7_U1_XOR1_U1 ( .A0_t (OUT_ciphertext_s0_t[7]), .A0_f (OUT_ciphertext_s0_f[7]), .A1_t (OUT_ciphertext_s1_t[7]), .A1_f (OUT_ciphertext_s1_f[7]), .B0_t (LED_128_Instance_addroundkey_tmp[7]), .B0_f (new_AGEMA_signal_3249), .B1_t (new_AGEMA_signal_3250), .B1_f (new_AGEMA_signal_3251), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_7_U1_X), .Z0_f (new_AGEMA_signal_3273), .Z1_t (new_AGEMA_signal_3274), .Z1_f (new_AGEMA_signal_3275) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_7_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n23), .A1_f (new_AGEMA_signal_2480), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_7_U1_X), .B0_f (new_AGEMA_signal_3273), .B1_t (new_AGEMA_signal_3274), .B1_f (new_AGEMA_signal_3275), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_7_U1_Y), .Z0_f (new_AGEMA_signal_3465), .Z1_t (new_AGEMA_signal_3466), .Z1_f (new_AGEMA_signal_3467) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_7_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_7_U1_Y), .A0_f (new_AGEMA_signal_3465), .A1_t (new_AGEMA_signal_3466), .A1_f (new_AGEMA_signal_3467), .B0_t (OUT_ciphertext_s0_t[7]), .B0_f (OUT_ciphertext_s0_f[7]), .B1_t (OUT_ciphertext_s1_t[7]), .B1_f (OUT_ciphertext_s1_f[7]), .Z0_t (LED_128_Instance_addconst_out[7]), .Z0_f (new_AGEMA_signal_3657), .Z1_t (new_AGEMA_signal_3658), .Z1_f (new_AGEMA_signal_3659) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_8_U1_XOR1_U1 ( .A0_t (OUT_ciphertext_s0_t[8]), .A0_f (OUT_ciphertext_s0_f[8]), .A1_t (OUT_ciphertext_s1_t[8]), .A1_f (OUT_ciphertext_s1_f[8]), .B0_t (LED_128_Instance_addroundkey_tmp[8]), .B0_f (new_AGEMA_signal_2889), .B1_t (new_AGEMA_signal_2890), .B1_f (new_AGEMA_signal_2891), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_8_U1_X), .Z0_f (new_AGEMA_signal_3276), .Z1_t (new_AGEMA_signal_3277), .Z1_f (new_AGEMA_signal_3278) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_8_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n23), .A1_f (new_AGEMA_signal_2480), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_8_U1_X), .B0_f (new_AGEMA_signal_3276), .B1_t (new_AGEMA_signal_3277), .B1_f (new_AGEMA_signal_3278), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_8_U1_Y), .Z0_f (new_AGEMA_signal_3468), .Z1_t (new_AGEMA_signal_3469), .Z1_f (new_AGEMA_signal_3470) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_8_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_8_U1_Y), .A0_f (new_AGEMA_signal_3468), .A1_t (new_AGEMA_signal_3469), .A1_f (new_AGEMA_signal_3470), .B0_t (OUT_ciphertext_s0_t[8]), .B0_f (OUT_ciphertext_s0_f[8]), .B1_t (OUT_ciphertext_s1_t[8]), .B1_f (OUT_ciphertext_s1_f[8]), .Z0_t (LED_128_Instance_addconst_out[8]), .Z0_f (new_AGEMA_signal_3660), .Z1_t (new_AGEMA_signal_3661), .Z1_f (new_AGEMA_signal_3662) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_9_U1_XOR1_U1 ( .A0_t (OUT_ciphertext_s0_t[9]), .A0_f (OUT_ciphertext_s0_f[9]), .A1_t (OUT_ciphertext_s1_t[9]), .A1_f (OUT_ciphertext_s1_f[9]), .B0_t (LED_128_Instance_addroundkey_tmp[9]), .B0_f (new_AGEMA_signal_3165), .B1_t (new_AGEMA_signal_3166), .B1_f (new_AGEMA_signal_3167), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_9_U1_X), .Z0_f (new_AGEMA_signal_3279), .Z1_t (new_AGEMA_signal_3280), .Z1_f (new_AGEMA_signal_3281) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_9_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n23), .A1_f (new_AGEMA_signal_2480), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_9_U1_X), .B0_f (new_AGEMA_signal_3279), .B1_t (new_AGEMA_signal_3280), .B1_f (new_AGEMA_signal_3281), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_9_U1_Y), .Z0_f (new_AGEMA_signal_3471), .Z1_t (new_AGEMA_signal_3472), .Z1_f (new_AGEMA_signal_3473) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_9_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_9_U1_Y), .A0_f (new_AGEMA_signal_3471), .A1_t (new_AGEMA_signal_3472), .A1_f (new_AGEMA_signal_3473), .B0_t (OUT_ciphertext_s0_t[9]), .B0_f (OUT_ciphertext_s0_f[9]), .B1_t (OUT_ciphertext_s1_t[9]), .B1_f (OUT_ciphertext_s1_f[9]), .Z0_t (LED_128_Instance_addconst_out[9]), .Z0_f (new_AGEMA_signal_3663), .Z1_t (new_AGEMA_signal_3664), .Z1_f (new_AGEMA_signal_3665) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_10_U1_XOR1_U1 ( .A0_t (OUT_ciphertext_s0_t[10]), .A0_f (OUT_ciphertext_s0_f[10]), .A1_t (OUT_ciphertext_s1_t[10]), .A1_f (OUT_ciphertext_s1_f[10]), .B0_t (LED_128_Instance_addroundkey_tmp[10]), .B0_f (new_AGEMA_signal_3105), .B1_t (new_AGEMA_signal_3106), .B1_f (new_AGEMA_signal_3107), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_10_U1_X), .Z0_f (new_AGEMA_signal_3282), .Z1_t (new_AGEMA_signal_3283), .Z1_f (new_AGEMA_signal_3284) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_10_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n23), .A1_f (new_AGEMA_signal_2480), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_10_U1_X), .B0_f (new_AGEMA_signal_3282), .B1_t (new_AGEMA_signal_3283), .B1_f (new_AGEMA_signal_3284), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_10_U1_Y), .Z0_f (new_AGEMA_signal_3474), .Z1_t (new_AGEMA_signal_3475), .Z1_f (new_AGEMA_signal_3476) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_10_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_10_U1_Y), .A0_f (new_AGEMA_signal_3474), .A1_t (new_AGEMA_signal_3475), .A1_f (new_AGEMA_signal_3476), .B0_t (OUT_ciphertext_s0_t[10]), .B0_f (OUT_ciphertext_s0_f[10]), .B1_t (OUT_ciphertext_s1_t[10]), .B1_f (OUT_ciphertext_s1_f[10]), .Z0_t (LED_128_Instance_addconst_out[10]), .Z0_f (new_AGEMA_signal_3666), .Z1_t (new_AGEMA_signal_3667), .Z1_f (new_AGEMA_signal_3668) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_11_U1_XOR1_U1 ( .A0_t (OUT_ciphertext_s0_t[11]), .A0_f (OUT_ciphertext_s0_f[11]), .A1_t (OUT_ciphertext_s1_t[11]), .A1_f (OUT_ciphertext_s1_f[11]), .B0_t (LED_128_Instance_addroundkey_tmp[11]), .B0_f (new_AGEMA_signal_3243), .B1_t (new_AGEMA_signal_3244), .B1_f (new_AGEMA_signal_3245), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_11_U1_X), .Z0_f (new_AGEMA_signal_3285), .Z1_t (new_AGEMA_signal_3286), .Z1_f (new_AGEMA_signal_3287) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_11_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n23), .A1_f (new_AGEMA_signal_2480), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_11_U1_X), .B0_f (new_AGEMA_signal_3285), .B1_t (new_AGEMA_signal_3286), .B1_f (new_AGEMA_signal_3287), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_11_U1_Y), .Z0_f (new_AGEMA_signal_3477), .Z1_t (new_AGEMA_signal_3478), .Z1_f (new_AGEMA_signal_3479) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_11_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_11_U1_Y), .A0_f (new_AGEMA_signal_3477), .A1_t (new_AGEMA_signal_3478), .A1_f (new_AGEMA_signal_3479), .B0_t (OUT_ciphertext_s0_t[11]), .B0_f (OUT_ciphertext_s0_f[11]), .B1_t (OUT_ciphertext_s1_t[11]), .B1_f (OUT_ciphertext_s1_f[11]), .Z0_t (LED_128_Instance_addconst_out[11]), .Z0_f (new_AGEMA_signal_3669), .Z1_t (new_AGEMA_signal_3670), .Z1_f (new_AGEMA_signal_3671) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_12_U1_XOR1_U1 ( .A0_t (OUT_ciphertext_s0_t[12]), .A0_f (OUT_ciphertext_s0_f[12]), .A1_t (OUT_ciphertext_s1_t[12]), .A1_f (OUT_ciphertext_s1_f[12]), .B0_t (LED_128_Instance_addroundkey_tmp[12]), .B0_f (new_AGEMA_signal_2883), .B1_t (new_AGEMA_signal_2884), .B1_f (new_AGEMA_signal_2885), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_12_U1_X), .Z0_f (new_AGEMA_signal_3288), .Z1_t (new_AGEMA_signal_3289), .Z1_f (new_AGEMA_signal_3290) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_12_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n23), .A1_f (new_AGEMA_signal_2480), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_12_U1_X), .B0_f (new_AGEMA_signal_3288), .B1_t (new_AGEMA_signal_3289), .B1_f (new_AGEMA_signal_3290), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_12_U1_Y), .Z0_f (new_AGEMA_signal_3480), .Z1_t (new_AGEMA_signal_3481), .Z1_f (new_AGEMA_signal_3482) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_12_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_12_U1_Y), .A0_f (new_AGEMA_signal_3480), .A1_t (new_AGEMA_signal_3481), .A1_f (new_AGEMA_signal_3482), .B0_t (OUT_ciphertext_s0_t[12]), .B0_f (OUT_ciphertext_s0_f[12]), .B1_t (OUT_ciphertext_s1_t[12]), .B1_f (OUT_ciphertext_s1_f[12]), .Z0_t (LED_128_Instance_addconst_out[12]), .Z0_f (new_AGEMA_signal_3672), .Z1_t (new_AGEMA_signal_3673), .Z1_f (new_AGEMA_signal_3674) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_13_U1_XOR1_U1 ( .A0_t (OUT_ciphertext_s0_t[13]), .A0_f (OUT_ciphertext_s0_f[13]), .A1_t (OUT_ciphertext_s1_t[13]), .A1_f (OUT_ciphertext_s1_f[13]), .B0_t (LED_128_Instance_addroundkey_tmp[13]), .B0_f (new_AGEMA_signal_3153), .B1_t (new_AGEMA_signal_3154), .B1_f (new_AGEMA_signal_3155), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_13_U1_X), .Z0_f (new_AGEMA_signal_3291), .Z1_t (new_AGEMA_signal_3292), .Z1_f (new_AGEMA_signal_3293) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_13_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n23), .A1_f (new_AGEMA_signal_2480), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_13_U1_X), .B0_f (new_AGEMA_signal_3291), .B1_t (new_AGEMA_signal_3292), .B1_f (new_AGEMA_signal_3293), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_13_U1_Y), .Z0_f (new_AGEMA_signal_3483), .Z1_t (new_AGEMA_signal_3484), .Z1_f (new_AGEMA_signal_3485) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_13_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_13_U1_Y), .A0_f (new_AGEMA_signal_3483), .A1_t (new_AGEMA_signal_3484), .A1_f (new_AGEMA_signal_3485), .B0_t (OUT_ciphertext_s0_t[13]), .B0_f (OUT_ciphertext_s0_f[13]), .B1_t (OUT_ciphertext_s1_t[13]), .B1_f (OUT_ciphertext_s1_f[13]), .Z0_t (LED_128_Instance_addconst_out[13]), .Z0_f (new_AGEMA_signal_3675), .Z1_t (new_AGEMA_signal_3676), .Z1_f (new_AGEMA_signal_3677) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_14_U1_XOR1_U1 ( .A0_t (OUT_ciphertext_s0_t[14]), .A0_f (OUT_ciphertext_s0_f[14]), .A1_t (OUT_ciphertext_s1_t[14]), .A1_f (OUT_ciphertext_s1_f[14]), .B0_t (LED_128_Instance_addroundkey_tmp[14]), .B0_f (new_AGEMA_signal_3093), .B1_t (new_AGEMA_signal_3094), .B1_f (new_AGEMA_signal_3095), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_14_U1_X), .Z0_f (new_AGEMA_signal_3294), .Z1_t (new_AGEMA_signal_3295), .Z1_f (new_AGEMA_signal_3296) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_14_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n23), .A1_f (new_AGEMA_signal_2480), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_14_U1_X), .B0_f (new_AGEMA_signal_3294), .B1_t (new_AGEMA_signal_3295), .B1_f (new_AGEMA_signal_3296), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_14_U1_Y), .Z0_f (new_AGEMA_signal_3486), .Z1_t (new_AGEMA_signal_3487), .Z1_f (new_AGEMA_signal_3488) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_14_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_14_U1_Y), .A0_f (new_AGEMA_signal_3486), .A1_t (new_AGEMA_signal_3487), .A1_f (new_AGEMA_signal_3488), .B0_t (OUT_ciphertext_s0_t[14]), .B0_f (OUT_ciphertext_s0_f[14]), .B1_t (OUT_ciphertext_s1_t[14]), .B1_f (OUT_ciphertext_s1_f[14]), .Z0_t (LED_128_Instance_addconst_out[14]), .Z0_f (new_AGEMA_signal_3678), .Z1_t (new_AGEMA_signal_3679), .Z1_f (new_AGEMA_signal_3680) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_15_U1_XOR1_U1 ( .A0_t (OUT_ciphertext_s0_t[15]), .A0_f (OUT_ciphertext_s0_f[15]), .A1_t (OUT_ciphertext_s1_t[15]), .A1_f (OUT_ciphertext_s1_f[15]), .B0_t (LED_128_Instance_addroundkey_tmp[15]), .B0_f (new_AGEMA_signal_3237), .B1_t (new_AGEMA_signal_3238), .B1_f (new_AGEMA_signal_3239), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_15_U1_X), .Z0_f (new_AGEMA_signal_3297), .Z1_t (new_AGEMA_signal_3298), .Z1_f (new_AGEMA_signal_3299) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_15_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n23), .A1_f (new_AGEMA_signal_2480), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_15_U1_X), .B0_f (new_AGEMA_signal_3297), .B1_t (new_AGEMA_signal_3298), .B1_f (new_AGEMA_signal_3299), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_15_U1_Y), .Z0_f (new_AGEMA_signal_3489), .Z1_t (new_AGEMA_signal_3490), .Z1_f (new_AGEMA_signal_3491) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_15_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_15_U1_Y), .A0_f (new_AGEMA_signal_3489), .A1_t (new_AGEMA_signal_3490), .A1_f (new_AGEMA_signal_3491), .B0_t (OUT_ciphertext_s0_t[15]), .B0_f (OUT_ciphertext_s0_f[15]), .B1_t (OUT_ciphertext_s1_t[15]), .B1_f (OUT_ciphertext_s1_f[15]), .Z0_t (LED_128_Instance_addconst_out[15]), .Z0_f (new_AGEMA_signal_3681), .Z1_t (new_AGEMA_signal_3682), .Z1_f (new_AGEMA_signal_3683) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_16_U1_XOR1_U1 ( .A0_t (OUT_ciphertext_s0_t[16]), .A0_f (OUT_ciphertext_s0_f[16]), .A1_t (OUT_ciphertext_s1_t[16]), .A1_f (OUT_ciphertext_s1_f[16]), .B0_t (LED_128_Instance_addroundkey_tmp[16]), .B0_f (new_AGEMA_signal_2907), .B1_t (new_AGEMA_signal_2908), .B1_f (new_AGEMA_signal_2909), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_16_U1_X), .Z0_f (new_AGEMA_signal_3300), .Z1_t (new_AGEMA_signal_3301), .Z1_f (new_AGEMA_signal_3302) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_16_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n23), .A1_f (new_AGEMA_signal_2480), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_16_U1_X), .B0_f (new_AGEMA_signal_3300), .B1_t (new_AGEMA_signal_3301), .B1_f (new_AGEMA_signal_3302), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_16_U1_Y), .Z0_f (new_AGEMA_signal_3492), .Z1_t (new_AGEMA_signal_3493), .Z1_f (new_AGEMA_signal_3494) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_16_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_16_U1_Y), .A0_f (new_AGEMA_signal_3492), .A1_t (new_AGEMA_signal_3493), .A1_f (new_AGEMA_signal_3494), .B0_t (OUT_ciphertext_s0_t[16]), .B0_f (OUT_ciphertext_s0_f[16]), .B1_t (OUT_ciphertext_s1_t[16]), .B1_f (OUT_ciphertext_s1_f[16]), .Z0_t (LED_128_Instance_addroundkey_out[16]), .Z0_f (new_AGEMA_signal_3684), .Z1_t (new_AGEMA_signal_3685), .Z1_f (new_AGEMA_signal_3686) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_17_U1_XOR1_U1 ( .A0_t (OUT_ciphertext_s0_t[17]), .A0_f (OUT_ciphertext_s0_f[17]), .A1_t (OUT_ciphertext_s1_t[17]), .A1_f (OUT_ciphertext_s1_f[17]), .B0_t (LED_128_Instance_addroundkey_tmp[17]), .B0_f (new_AGEMA_signal_3159), .B1_t (new_AGEMA_signal_3160), .B1_f (new_AGEMA_signal_3161), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_17_U1_X), .Z0_f (new_AGEMA_signal_3303), .Z1_t (new_AGEMA_signal_3304), .Z1_f (new_AGEMA_signal_3305) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_17_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n23), .A1_f (new_AGEMA_signal_2480), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_17_U1_X), .B0_f (new_AGEMA_signal_3303), .B1_t (new_AGEMA_signal_3304), .B1_f (new_AGEMA_signal_3305), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_17_U1_Y), .Z0_f (new_AGEMA_signal_3495), .Z1_t (new_AGEMA_signal_3496), .Z1_f (new_AGEMA_signal_3497) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_17_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_17_U1_Y), .A0_f (new_AGEMA_signal_3495), .A1_t (new_AGEMA_signal_3496), .A1_f (new_AGEMA_signal_3497), .B0_t (OUT_ciphertext_s0_t[17]), .B0_f (OUT_ciphertext_s0_f[17]), .B1_t (OUT_ciphertext_s1_t[17]), .B1_f (OUT_ciphertext_s1_f[17]), .Z0_t (LED_128_Instance_addconst_out[17]), .Z0_f (new_AGEMA_signal_3687), .Z1_t (new_AGEMA_signal_3688), .Z1_f (new_AGEMA_signal_3689) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_18_U1_XOR1_U1 ( .A0_t (OUT_ciphertext_s0_t[18]), .A0_f (OUT_ciphertext_s0_f[18]), .A1_t (OUT_ciphertext_s1_t[18]), .A1_f (OUT_ciphertext_s1_f[18]), .B0_t (LED_128_Instance_addroundkey_tmp[18]), .B0_f (new_AGEMA_signal_3099), .B1_t (new_AGEMA_signal_3100), .B1_f (new_AGEMA_signal_3101), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_18_U1_X), .Z0_f (new_AGEMA_signal_3306), .Z1_t (new_AGEMA_signal_3307), .Z1_f (new_AGEMA_signal_3308) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_18_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n23), .A1_f (new_AGEMA_signal_2480), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_18_U1_X), .B0_f (new_AGEMA_signal_3306), .B1_t (new_AGEMA_signal_3307), .B1_f (new_AGEMA_signal_3308), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_18_U1_Y), .Z0_f (new_AGEMA_signal_3498), .Z1_t (new_AGEMA_signal_3499), .Z1_f (new_AGEMA_signal_3500) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_18_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_18_U1_Y), .A0_f (new_AGEMA_signal_3498), .A1_t (new_AGEMA_signal_3499), .A1_f (new_AGEMA_signal_3500), .B0_t (OUT_ciphertext_s0_t[18]), .B0_f (OUT_ciphertext_s0_f[18]), .B1_t (OUT_ciphertext_s1_t[18]), .B1_f (OUT_ciphertext_s1_f[18]), .Z0_t (LED_128_Instance_addconst_out[18]), .Z0_f (new_AGEMA_signal_3690), .Z1_t (new_AGEMA_signal_3691), .Z1_f (new_AGEMA_signal_3692) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_19_U1_XOR1_U1 ( .A0_t (OUT_ciphertext_s0_t[19]), .A0_f (OUT_ciphertext_s0_f[19]), .A1_t (OUT_ciphertext_s1_t[19]), .A1_f (OUT_ciphertext_s1_f[19]), .B0_t (LED_128_Instance_addroundkey_tmp[19]), .B0_f (new_AGEMA_signal_2973), .B1_t (new_AGEMA_signal_2974), .B1_f (new_AGEMA_signal_2975), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_19_U1_X), .Z0_f (new_AGEMA_signal_3309), .Z1_t (new_AGEMA_signal_3310), .Z1_f (new_AGEMA_signal_3311) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_19_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n23), .A1_f (new_AGEMA_signal_2480), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_19_U1_X), .B0_f (new_AGEMA_signal_3309), .B1_t (new_AGEMA_signal_3310), .B1_f (new_AGEMA_signal_3311), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_19_U1_Y), .Z0_f (new_AGEMA_signal_3501), .Z1_t (new_AGEMA_signal_3502), .Z1_f (new_AGEMA_signal_3503) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_19_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_19_U1_Y), .A0_f (new_AGEMA_signal_3501), .A1_t (new_AGEMA_signal_3502), .A1_f (new_AGEMA_signal_3503), .B0_t (OUT_ciphertext_s0_t[19]), .B0_f (OUT_ciphertext_s0_f[19]), .B1_t (OUT_ciphertext_s1_t[19]), .B1_f (OUT_ciphertext_s1_f[19]), .Z0_t (LED_128_Instance_addroundkey_out[19]), .Z0_f (new_AGEMA_signal_3693), .Z1_t (new_AGEMA_signal_3694), .Z1_f (new_AGEMA_signal_3695) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_20_U1_XOR1_U1 ( .A0_t (OUT_ciphertext_s0_t[20]), .A0_f (OUT_ciphertext_s0_f[20]), .A1_t (OUT_ciphertext_s1_t[20]), .A1_f (OUT_ciphertext_s1_f[20]), .B0_t (LED_128_Instance_addroundkey_tmp[20]), .B0_f (new_AGEMA_signal_3033), .B1_t (new_AGEMA_signal_3034), .B1_f (new_AGEMA_signal_3035), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_20_U1_X), .Z0_f (new_AGEMA_signal_3312), .Z1_t (new_AGEMA_signal_3313), .Z1_f (new_AGEMA_signal_3314) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_20_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n23), .A1_f (new_AGEMA_signal_2480), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_20_U1_X), .B0_f (new_AGEMA_signal_3312), .B1_t (new_AGEMA_signal_3313), .B1_f (new_AGEMA_signal_3314), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_20_U1_Y), .Z0_f (new_AGEMA_signal_3504), .Z1_t (new_AGEMA_signal_3505), .Z1_f (new_AGEMA_signal_3506) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_20_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_20_U1_Y), .A0_f (new_AGEMA_signal_3504), .A1_t (new_AGEMA_signal_3505), .A1_f (new_AGEMA_signal_3506), .B0_t (OUT_ciphertext_s0_t[20]), .B0_f (OUT_ciphertext_s0_f[20]), .B1_t (OUT_ciphertext_s1_t[20]), .B1_f (OUT_ciphertext_s1_f[20]), .Z0_t (LED_128_Instance_addroundkey_out[20]), .Z0_f (new_AGEMA_signal_3696), .Z1_t (new_AGEMA_signal_3697), .Z1_f (new_AGEMA_signal_3698) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_21_U1_XOR1_U1 ( .A0_t (OUT_ciphertext_s0_t[21]), .A0_f (OUT_ciphertext_s0_f[21]), .A1_t (OUT_ciphertext_s1_t[21]), .A1_f (OUT_ciphertext_s1_f[21]), .B0_t (LED_128_Instance_addroundkey_tmp[21]), .B0_f (new_AGEMA_signal_3051), .B1_t (new_AGEMA_signal_3052), .B1_f (new_AGEMA_signal_3053), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_21_U1_X), .Z0_f (new_AGEMA_signal_3315), .Z1_t (new_AGEMA_signal_3316), .Z1_f (new_AGEMA_signal_3317) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_21_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n23), .A1_f (new_AGEMA_signal_2480), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_21_U1_X), .B0_f (new_AGEMA_signal_3315), .B1_t (new_AGEMA_signal_3316), .B1_f (new_AGEMA_signal_3317), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_21_U1_Y), .Z0_f (new_AGEMA_signal_3507), .Z1_t (new_AGEMA_signal_3508), .Z1_f (new_AGEMA_signal_3509) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_21_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_21_U1_Y), .A0_f (new_AGEMA_signal_3507), .A1_t (new_AGEMA_signal_3508), .A1_f (new_AGEMA_signal_3509), .B0_t (OUT_ciphertext_s0_t[21]), .B0_f (OUT_ciphertext_s0_f[21]), .B1_t (OUT_ciphertext_s1_t[21]), .B1_f (OUT_ciphertext_s1_f[21]), .Z0_t (LED_128_Instance_addroundkey_out[21]), .Z0_f (new_AGEMA_signal_3699), .Z1_t (new_AGEMA_signal_3700), .Z1_f (new_AGEMA_signal_3701) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_22_U1_XOR1_U1 ( .A0_t (OUT_ciphertext_s0_t[22]), .A0_f (OUT_ciphertext_s0_f[22]), .A1_t (OUT_ciphertext_s1_t[22]), .A1_f (OUT_ciphertext_s1_f[22]), .B0_t (LED_128_Instance_addroundkey_tmp[22]), .B0_f (new_AGEMA_signal_3039), .B1_t (new_AGEMA_signal_3040), .B1_f (new_AGEMA_signal_3041), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_22_U1_X), .Z0_f (new_AGEMA_signal_3318), .Z1_t (new_AGEMA_signal_3319), .Z1_f (new_AGEMA_signal_3320) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_22_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n23), .A1_f (new_AGEMA_signal_2480), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_22_U1_X), .B0_f (new_AGEMA_signal_3318), .B1_t (new_AGEMA_signal_3319), .B1_f (new_AGEMA_signal_3320), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_22_U1_Y), .Z0_f (new_AGEMA_signal_3510), .Z1_t (new_AGEMA_signal_3511), .Z1_f (new_AGEMA_signal_3512) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_22_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_22_U1_Y), .A0_f (new_AGEMA_signal_3510), .A1_t (new_AGEMA_signal_3511), .A1_f (new_AGEMA_signal_3512), .B0_t (OUT_ciphertext_s0_t[22]), .B0_f (OUT_ciphertext_s0_f[22]), .B1_t (OUT_ciphertext_s1_t[22]), .B1_f (OUT_ciphertext_s1_f[22]), .Z0_t (LED_128_Instance_addroundkey_out[22]), .Z0_f (new_AGEMA_signal_3702), .Z1_t (new_AGEMA_signal_3703), .Z1_f (new_AGEMA_signal_3704) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_23_U1_XOR1_U1 ( .A0_t (OUT_ciphertext_s0_t[23]), .A0_f (OUT_ciphertext_s0_f[23]), .A1_t (OUT_ciphertext_s1_t[23]), .A1_f (OUT_ciphertext_s1_f[23]), .B0_t (LED_128_Instance_addroundkey_tmp[23]), .B0_f (new_AGEMA_signal_2937), .B1_t (new_AGEMA_signal_2938), .B1_f (new_AGEMA_signal_2939), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_23_U1_X), .Z0_f (new_AGEMA_signal_3321), .Z1_t (new_AGEMA_signal_3322), .Z1_f (new_AGEMA_signal_3323) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_23_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n23), .A1_f (new_AGEMA_signal_2480), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_23_U1_X), .B0_f (new_AGEMA_signal_3321), .B1_t (new_AGEMA_signal_3322), .B1_f (new_AGEMA_signal_3323), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_23_U1_Y), .Z0_f (new_AGEMA_signal_3513), .Z1_t (new_AGEMA_signal_3514), .Z1_f (new_AGEMA_signal_3515) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_23_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_23_U1_Y), .A0_f (new_AGEMA_signal_3513), .A1_t (new_AGEMA_signal_3514), .A1_f (new_AGEMA_signal_3515), .B0_t (OUT_ciphertext_s0_t[23]), .B0_f (OUT_ciphertext_s0_f[23]), .B1_t (OUT_ciphertext_s1_t[23]), .B1_f (OUT_ciphertext_s1_f[23]), .Z0_t (LED_128_Instance_addconst_out[23]), .Z0_f (new_AGEMA_signal_3705), .Z1_t (new_AGEMA_signal_3706), .Z1_f (new_AGEMA_signal_3707) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_24_U1_XOR1_U1 ( .A0_t (OUT_ciphertext_s0_t[24]), .A0_f (OUT_ciphertext_s0_f[24]), .A1_t (OUT_ciphertext_s1_t[24]), .A1_f (OUT_ciphertext_s1_f[24]), .B0_t (LED_128_Instance_addroundkey_tmp[24]), .B0_f (new_AGEMA_signal_2877), .B1_t (new_AGEMA_signal_2878), .B1_f (new_AGEMA_signal_2879), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_24_U1_X), .Z0_f (new_AGEMA_signal_3324), .Z1_t (new_AGEMA_signal_3325), .Z1_f (new_AGEMA_signal_3326) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_24_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n23), .A1_f (new_AGEMA_signal_2480), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_24_U1_X), .B0_f (new_AGEMA_signal_3324), .B1_t (new_AGEMA_signal_3325), .B1_f (new_AGEMA_signal_3326), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_24_U1_Y), .Z0_f (new_AGEMA_signal_3516), .Z1_t (new_AGEMA_signal_3517), .Z1_f (new_AGEMA_signal_3518) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_24_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_24_U1_Y), .A0_f (new_AGEMA_signal_3516), .A1_t (new_AGEMA_signal_3517), .A1_f (new_AGEMA_signal_3518), .B0_t (OUT_ciphertext_s0_t[24]), .B0_f (OUT_ciphertext_s0_f[24]), .B1_t (OUT_ciphertext_s1_t[24]), .B1_f (OUT_ciphertext_s1_f[24]), .Z0_t (LED_128_Instance_addconst_out[24]), .Z0_f (new_AGEMA_signal_3708), .Z1_t (new_AGEMA_signal_3709), .Z1_f (new_AGEMA_signal_3710) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_25_U1_XOR1_U1 ( .A0_t (OUT_ciphertext_s0_t[25]), .A0_f (OUT_ciphertext_s0_f[25]), .A1_t (OUT_ciphertext_s1_t[25]), .A1_f (OUT_ciphertext_s1_f[25]), .B0_t (LED_128_Instance_addroundkey_tmp[25]), .B0_f (new_AGEMA_signal_3177), .B1_t (new_AGEMA_signal_3178), .B1_f (new_AGEMA_signal_3179), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_25_U1_X), .Z0_f (new_AGEMA_signal_3327), .Z1_t (new_AGEMA_signal_3328), .Z1_f (new_AGEMA_signal_3329) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_25_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n23), .A1_f (new_AGEMA_signal_2480), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_25_U1_X), .B0_f (new_AGEMA_signal_3327), .B1_t (new_AGEMA_signal_3328), .B1_f (new_AGEMA_signal_3329), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_25_U1_Y), .Z0_f (new_AGEMA_signal_3519), .Z1_t (new_AGEMA_signal_3520), .Z1_f (new_AGEMA_signal_3521) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_25_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_25_U1_Y), .A0_f (new_AGEMA_signal_3519), .A1_t (new_AGEMA_signal_3520), .A1_f (new_AGEMA_signal_3521), .B0_t (OUT_ciphertext_s0_t[25]), .B0_f (OUT_ciphertext_s0_f[25]), .B1_t (OUT_ciphertext_s1_t[25]), .B1_f (OUT_ciphertext_s1_f[25]), .Z0_t (LED_128_Instance_addconst_out[25]), .Z0_f (new_AGEMA_signal_3711), .Z1_t (new_AGEMA_signal_3712), .Z1_f (new_AGEMA_signal_3713) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_26_U1_XOR1_U1 ( .A0_t (OUT_ciphertext_s0_t[26]), .A0_f (OUT_ciphertext_s0_f[26]), .A1_t (OUT_ciphertext_s1_t[26]), .A1_f (OUT_ciphertext_s1_f[26]), .B0_t (LED_128_Instance_addroundkey_tmp[26]), .B0_f (new_AGEMA_signal_3117), .B1_t (new_AGEMA_signal_3118), .B1_f (new_AGEMA_signal_3119), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_26_U1_X), .Z0_f (new_AGEMA_signal_3330), .Z1_t (new_AGEMA_signal_3331), .Z1_f (new_AGEMA_signal_3332) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_26_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n23), .A1_f (new_AGEMA_signal_2480), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_26_U1_X), .B0_f (new_AGEMA_signal_3330), .B1_t (new_AGEMA_signal_3331), .B1_f (new_AGEMA_signal_3332), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_26_U1_Y), .Z0_f (new_AGEMA_signal_3522), .Z1_t (new_AGEMA_signal_3523), .Z1_f (new_AGEMA_signal_3524) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_26_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_26_U1_Y), .A0_f (new_AGEMA_signal_3522), .A1_t (new_AGEMA_signal_3523), .A1_f (new_AGEMA_signal_3524), .B0_t (OUT_ciphertext_s0_t[26]), .B0_f (OUT_ciphertext_s0_f[26]), .B1_t (OUT_ciphertext_s1_t[26]), .B1_f (OUT_ciphertext_s1_f[26]), .Z0_t (LED_128_Instance_addconst_out[26]), .Z0_f (new_AGEMA_signal_3714), .Z1_t (new_AGEMA_signal_3715), .Z1_f (new_AGEMA_signal_3716) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_27_U1_XOR1_U1 ( .A0_t (OUT_ciphertext_s0_t[27]), .A0_f (OUT_ciphertext_s0_f[27]), .A1_t (OUT_ciphertext_s1_t[27]), .A1_f (OUT_ciphertext_s1_f[27]), .B0_t (LED_128_Instance_addroundkey_tmp[27]), .B0_f (new_AGEMA_signal_2931), .B1_t (new_AGEMA_signal_2932), .B1_f (new_AGEMA_signal_2933), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_27_U1_X), .Z0_f (new_AGEMA_signal_3333), .Z1_t (new_AGEMA_signal_3334), .Z1_f (new_AGEMA_signal_3335) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_27_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n23), .A1_f (new_AGEMA_signal_2480), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_27_U1_X), .B0_f (new_AGEMA_signal_3333), .B1_t (new_AGEMA_signal_3334), .B1_f (new_AGEMA_signal_3335), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_27_U1_Y), .Z0_f (new_AGEMA_signal_3525), .Z1_t (new_AGEMA_signal_3526), .Z1_f (new_AGEMA_signal_3527) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_27_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_27_U1_Y), .A0_f (new_AGEMA_signal_3525), .A1_t (new_AGEMA_signal_3526), .A1_f (new_AGEMA_signal_3527), .B0_t (OUT_ciphertext_s0_t[27]), .B0_f (OUT_ciphertext_s0_f[27]), .B1_t (OUT_ciphertext_s1_t[27]), .B1_f (OUT_ciphertext_s1_f[27]), .Z0_t (LED_128_Instance_addconst_out[27]), .Z0_f (new_AGEMA_signal_3717), .Z1_t (new_AGEMA_signal_3718), .Z1_f (new_AGEMA_signal_3719) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_28_U1_XOR1_U1 ( .A0_t (OUT_ciphertext_s0_t[28]), .A0_f (OUT_ciphertext_s0_f[28]), .A1_t (OUT_ciphertext_s1_t[28]), .A1_f (OUT_ciphertext_s1_f[28]), .B0_t (LED_128_Instance_addroundkey_tmp[28]), .B0_f (new_AGEMA_signal_2871), .B1_t (new_AGEMA_signal_2872), .B1_f (new_AGEMA_signal_2873), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_28_U1_X), .Z0_f (new_AGEMA_signal_3336), .Z1_t (new_AGEMA_signal_3337), .Z1_f (new_AGEMA_signal_3338) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_28_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n23), .A1_f (new_AGEMA_signal_2480), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_28_U1_X), .B0_f (new_AGEMA_signal_3336), .B1_t (new_AGEMA_signal_3337), .B1_f (new_AGEMA_signal_3338), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_28_U1_Y), .Z0_f (new_AGEMA_signal_3528), .Z1_t (new_AGEMA_signal_3529), .Z1_f (new_AGEMA_signal_3530) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_28_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_28_U1_Y), .A0_f (new_AGEMA_signal_3528), .A1_t (new_AGEMA_signal_3529), .A1_f (new_AGEMA_signal_3530), .B0_t (OUT_ciphertext_s0_t[28]), .B0_f (OUT_ciphertext_s0_f[28]), .B1_t (OUT_ciphertext_s1_t[28]), .B1_f (OUT_ciphertext_s1_f[28]), .Z0_t (LED_128_Instance_addconst_out[28]), .Z0_f (new_AGEMA_signal_3720), .Z1_t (new_AGEMA_signal_3721), .Z1_f (new_AGEMA_signal_3722) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_29_U1_XOR1_U1 ( .A0_t (OUT_ciphertext_s0_t[29]), .A0_f (OUT_ciphertext_s0_f[29]), .A1_t (OUT_ciphertext_s1_t[29]), .A1_f (OUT_ciphertext_s1_f[29]), .B0_t (LED_128_Instance_addroundkey_tmp[29]), .B0_f (new_AGEMA_signal_3171), .B1_t (new_AGEMA_signal_3172), .B1_f (new_AGEMA_signal_3173), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_29_U1_X), .Z0_f (new_AGEMA_signal_3339), .Z1_t (new_AGEMA_signal_3340), .Z1_f (new_AGEMA_signal_3341) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_29_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n23), .A1_f (new_AGEMA_signal_2480), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_29_U1_X), .B0_f (new_AGEMA_signal_3339), .B1_t (new_AGEMA_signal_3340), .B1_f (new_AGEMA_signal_3341), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_29_U1_Y), .Z0_f (new_AGEMA_signal_3531), .Z1_t (new_AGEMA_signal_3532), .Z1_f (new_AGEMA_signal_3533) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_29_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_29_U1_Y), .A0_f (new_AGEMA_signal_3531), .A1_t (new_AGEMA_signal_3532), .A1_f (new_AGEMA_signal_3533), .B0_t (OUT_ciphertext_s0_t[29]), .B0_f (OUT_ciphertext_s0_f[29]), .B1_t (OUT_ciphertext_s1_t[29]), .B1_f (OUT_ciphertext_s1_f[29]), .Z0_t (LED_128_Instance_addconst_out[29]), .Z0_f (new_AGEMA_signal_3723), .Z1_t (new_AGEMA_signal_3724), .Z1_f (new_AGEMA_signal_3725) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_30_U1_XOR1_U1 ( .A0_t (OUT_ciphertext_s0_t[30]), .A0_f (OUT_ciphertext_s0_f[30]), .A1_t (OUT_ciphertext_s1_t[30]), .A1_f (OUT_ciphertext_s1_f[30]), .B0_t (LED_128_Instance_addroundkey_tmp[30]), .B0_f (new_AGEMA_signal_3111), .B1_t (new_AGEMA_signal_3112), .B1_f (new_AGEMA_signal_3113), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_30_U1_X), .Z0_f (new_AGEMA_signal_3342), .Z1_t (new_AGEMA_signal_3343), .Z1_f (new_AGEMA_signal_3344) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_30_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n23), .A1_f (new_AGEMA_signal_2480), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_30_U1_X), .B0_f (new_AGEMA_signal_3342), .B1_t (new_AGEMA_signal_3343), .B1_f (new_AGEMA_signal_3344), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_30_U1_Y), .Z0_f (new_AGEMA_signal_3534), .Z1_t (new_AGEMA_signal_3535), .Z1_f (new_AGEMA_signal_3536) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_30_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_30_U1_Y), .A0_f (new_AGEMA_signal_3534), .A1_t (new_AGEMA_signal_3535), .A1_f (new_AGEMA_signal_3536), .B0_t (OUT_ciphertext_s0_t[30]), .B0_f (OUT_ciphertext_s0_f[30]), .B1_t (OUT_ciphertext_s1_t[30]), .B1_f (OUT_ciphertext_s1_f[30]), .Z0_t (LED_128_Instance_addconst_out[30]), .Z0_f (new_AGEMA_signal_3726), .Z1_t (new_AGEMA_signal_3727), .Z1_f (new_AGEMA_signal_3728) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_31_U1_XOR1_U1 ( .A0_t (OUT_ciphertext_s0_t[31]), .A0_f (OUT_ciphertext_s0_f[31]), .A1_t (OUT_ciphertext_s1_t[31]), .A1_f (OUT_ciphertext_s1_f[31]), .B0_t (LED_128_Instance_addroundkey_tmp[31]), .B0_f (new_AGEMA_signal_2925), .B1_t (new_AGEMA_signal_2926), .B1_f (new_AGEMA_signal_2927), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_31_U1_X), .Z0_f (new_AGEMA_signal_3345), .Z1_t (new_AGEMA_signal_3346), .Z1_f (new_AGEMA_signal_3347) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_31_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n23), .A1_f (new_AGEMA_signal_2480), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_31_U1_X), .B0_f (new_AGEMA_signal_3345), .B1_t (new_AGEMA_signal_3346), .B1_f (new_AGEMA_signal_3347), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_31_U1_Y), .Z0_f (new_AGEMA_signal_3537), .Z1_t (new_AGEMA_signal_3538), .Z1_f (new_AGEMA_signal_3539) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_31_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_31_U1_Y), .A0_f (new_AGEMA_signal_3537), .A1_t (new_AGEMA_signal_3538), .A1_f (new_AGEMA_signal_3539), .B0_t (OUT_ciphertext_s0_t[31]), .B0_f (OUT_ciphertext_s0_f[31]), .B1_t (OUT_ciphertext_s1_t[31]), .B1_f (OUT_ciphertext_s1_f[31]), .Z0_t (LED_128_Instance_addconst_out[31]), .Z0_f (new_AGEMA_signal_3729), .Z1_t (new_AGEMA_signal_3730), .Z1_f (new_AGEMA_signal_3731) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_32_U1_XOR1_U1 ( .A0_t (OUT_ciphertext_s0_t[32]), .A0_f (OUT_ciphertext_s0_f[32]), .A1_t (OUT_ciphertext_s1_t[32]), .A1_f (OUT_ciphertext_s1_f[32]), .B0_t (LED_128_Instance_addroundkey_tmp[32]), .B0_f (new_AGEMA_signal_2943), .B1_t (new_AGEMA_signal_2944), .B1_f (new_AGEMA_signal_2945), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_32_U1_X), .Z0_f (new_AGEMA_signal_3348), .Z1_t (new_AGEMA_signal_3349), .Z1_f (new_AGEMA_signal_3350) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_32_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n23), .A1_f (new_AGEMA_signal_2480), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_32_U1_X), .B0_f (new_AGEMA_signal_3348), .B1_t (new_AGEMA_signal_3349), .B1_f (new_AGEMA_signal_3350), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_32_U1_Y), .Z0_f (new_AGEMA_signal_3540), .Z1_t (new_AGEMA_signal_3541), .Z1_f (new_AGEMA_signal_3542) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_32_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_32_U1_Y), .A0_f (new_AGEMA_signal_3540), .A1_t (new_AGEMA_signal_3541), .A1_f (new_AGEMA_signal_3542), .B0_t (OUT_ciphertext_s0_t[32]), .B0_f (OUT_ciphertext_s0_f[32]), .B1_t (OUT_ciphertext_s1_t[32]), .B1_f (OUT_ciphertext_s1_f[32]), .Z0_t (LED_128_Instance_addconst_out[32]), .Z0_f (new_AGEMA_signal_3732), .Z1_t (new_AGEMA_signal_3733), .Z1_f (new_AGEMA_signal_3734) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_33_U1_XOR1_U1 ( .A0_t (OUT_ciphertext_s0_t[33]), .A0_f (OUT_ciphertext_s0_f[33]), .A1_t (OUT_ciphertext_s1_t[33]), .A1_f (OUT_ciphertext_s1_f[33]), .B0_t (LED_128_Instance_addroundkey_tmp[33]), .B0_f (new_AGEMA_signal_2961), .B1_t (new_AGEMA_signal_2962), .B1_f (new_AGEMA_signal_2963), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_33_U1_X), .Z0_f (new_AGEMA_signal_3351), .Z1_t (new_AGEMA_signal_3352), .Z1_f (new_AGEMA_signal_3353) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_33_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n23), .A1_f (new_AGEMA_signal_2480), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_33_U1_X), .B0_f (new_AGEMA_signal_3351), .B1_t (new_AGEMA_signal_3352), .B1_f (new_AGEMA_signal_3353), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_33_U1_Y), .Z0_f (new_AGEMA_signal_3543), .Z1_t (new_AGEMA_signal_3544), .Z1_f (new_AGEMA_signal_3545) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_33_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_33_U1_Y), .A0_f (new_AGEMA_signal_3543), .A1_t (new_AGEMA_signal_3544), .A1_f (new_AGEMA_signal_3545), .B0_t (OUT_ciphertext_s0_t[33]), .B0_f (OUT_ciphertext_s0_f[33]), .B1_t (OUT_ciphertext_s1_t[33]), .B1_f (OUT_ciphertext_s1_f[33]), .Z0_t (LED_128_Instance_addroundkey_out[33]), .Z0_f (new_AGEMA_signal_3735), .Z1_t (new_AGEMA_signal_3736), .Z1_f (new_AGEMA_signal_3737) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_34_U1_XOR1_U1 ( .A0_t (OUT_ciphertext_s0_t[34]), .A0_f (OUT_ciphertext_s0_f[34]), .A1_t (OUT_ciphertext_s1_t[34]), .A1_f (OUT_ciphertext_s1_f[34]), .B0_t (LED_128_Instance_addroundkey_tmp[34]), .B0_f (new_AGEMA_signal_3075), .B1_t (new_AGEMA_signal_3076), .B1_f (new_AGEMA_signal_3077), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_34_U1_X), .Z0_f (new_AGEMA_signal_3354), .Z1_t (new_AGEMA_signal_3355), .Z1_f (new_AGEMA_signal_3356) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_34_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n23), .A1_f (new_AGEMA_signal_2480), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_34_U1_X), .B0_f (new_AGEMA_signal_3354), .B1_t (new_AGEMA_signal_3355), .B1_f (new_AGEMA_signal_3356), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_34_U1_Y), .Z0_f (new_AGEMA_signal_3546), .Z1_t (new_AGEMA_signal_3547), .Z1_f (new_AGEMA_signal_3548) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_34_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_34_U1_Y), .A0_f (new_AGEMA_signal_3546), .A1_t (new_AGEMA_signal_3547), .A1_f (new_AGEMA_signal_3548), .B0_t (OUT_ciphertext_s0_t[34]), .B0_f (OUT_ciphertext_s0_f[34]), .B1_t (OUT_ciphertext_s1_t[34]), .B1_f (OUT_ciphertext_s1_f[34]), .Z0_t (LED_128_Instance_addconst_out[34]), .Z0_f (new_AGEMA_signal_3738), .Z1_t (new_AGEMA_signal_3739), .Z1_f (new_AGEMA_signal_3740) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_35_U1_XOR1_U1 ( .A0_t (OUT_ciphertext_s0_t[35]), .A0_f (OUT_ciphertext_s0_f[35]), .A1_t (OUT_ciphertext_s1_t[35]), .A1_f (OUT_ciphertext_s1_f[35]), .B0_t (LED_128_Instance_addroundkey_tmp[35]), .B0_f (new_AGEMA_signal_3195), .B1_t (new_AGEMA_signal_3196), .B1_f (new_AGEMA_signal_3197), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_35_U1_X), .Z0_f (new_AGEMA_signal_3357), .Z1_t (new_AGEMA_signal_3358), .Z1_f (new_AGEMA_signal_3359) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_35_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n23), .A1_f (new_AGEMA_signal_2480), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_35_U1_X), .B0_f (new_AGEMA_signal_3357), .B1_t (new_AGEMA_signal_3358), .B1_f (new_AGEMA_signal_3359), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_35_U1_Y), .Z0_f (new_AGEMA_signal_3549), .Z1_t (new_AGEMA_signal_3550), .Z1_f (new_AGEMA_signal_3551) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_35_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_35_U1_Y), .A0_f (new_AGEMA_signal_3549), .A1_t (new_AGEMA_signal_3550), .A1_f (new_AGEMA_signal_3551), .B0_t (OUT_ciphertext_s0_t[35]), .B0_f (OUT_ciphertext_s0_f[35]), .B1_t (OUT_ciphertext_s1_t[35]), .B1_f (OUT_ciphertext_s1_f[35]), .Z0_t (LED_128_Instance_addconst_out[35]), .Z0_f (new_AGEMA_signal_3741), .Z1_t (new_AGEMA_signal_3742), .Z1_f (new_AGEMA_signal_3743) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_36_U1_XOR1_U1 ( .A0_t (OUT_ciphertext_s0_t[36]), .A0_f (OUT_ciphertext_s0_f[36]), .A1_t (OUT_ciphertext_s1_t[36]), .A1_f (OUT_ciphertext_s1_f[36]), .B0_t (LED_128_Instance_addroundkey_tmp[36]), .B0_f (new_AGEMA_signal_2997), .B1_t (new_AGEMA_signal_2998), .B1_f (new_AGEMA_signal_2999), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_36_U1_X), .Z0_f (new_AGEMA_signal_3360), .Z1_t (new_AGEMA_signal_3361), .Z1_f (new_AGEMA_signal_3362) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_36_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n23), .A1_f (new_AGEMA_signal_2480), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_36_U1_X), .B0_f (new_AGEMA_signal_3360), .B1_t (new_AGEMA_signal_3361), .B1_f (new_AGEMA_signal_3362), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_36_U1_Y), .Z0_f (new_AGEMA_signal_3552), .Z1_t (new_AGEMA_signal_3553), .Z1_f (new_AGEMA_signal_3554) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_36_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_36_U1_Y), .A0_f (new_AGEMA_signal_3552), .A1_t (new_AGEMA_signal_3553), .A1_f (new_AGEMA_signal_3554), .B0_t (OUT_ciphertext_s0_t[36]), .B0_f (OUT_ciphertext_s0_f[36]), .B1_t (OUT_ciphertext_s1_t[36]), .B1_f (OUT_ciphertext_s1_f[36]), .Z0_t (LED_128_Instance_addroundkey_out[36]), .Z0_f (new_AGEMA_signal_3744), .Z1_t (new_AGEMA_signal_3745), .Z1_f (new_AGEMA_signal_3746) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_37_U1_XOR1_U1 ( .A0_t (OUT_ciphertext_s0_t[37]), .A0_f (OUT_ciphertext_s0_f[37]), .A1_t (OUT_ciphertext_s1_t[37]), .A1_f (OUT_ciphertext_s1_f[37]), .B0_t (LED_128_Instance_addroundkey_tmp[37]), .B0_f (new_AGEMA_signal_3009), .B1_t (new_AGEMA_signal_3010), .B1_f (new_AGEMA_signal_3011), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_37_U1_X), .Z0_f (new_AGEMA_signal_3363), .Z1_t (new_AGEMA_signal_3364), .Z1_f (new_AGEMA_signal_3365) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_37_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n23), .A1_f (new_AGEMA_signal_2480), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_37_U1_X), .B0_f (new_AGEMA_signal_3363), .B1_t (new_AGEMA_signal_3364), .B1_f (new_AGEMA_signal_3365), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_37_U1_Y), .Z0_f (new_AGEMA_signal_3555), .Z1_t (new_AGEMA_signal_3556), .Z1_f (new_AGEMA_signal_3557) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_37_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_37_U1_Y), .A0_f (new_AGEMA_signal_3555), .A1_t (new_AGEMA_signal_3556), .A1_f (new_AGEMA_signal_3557), .B0_t (OUT_ciphertext_s0_t[37]), .B0_f (OUT_ciphertext_s0_f[37]), .B1_t (OUT_ciphertext_s1_t[37]), .B1_f (OUT_ciphertext_s1_f[37]), .Z0_t (LED_128_Instance_addroundkey_out[37]), .Z0_f (new_AGEMA_signal_3747), .Z1_t (new_AGEMA_signal_3748), .Z1_f (new_AGEMA_signal_3749) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_38_U1_XOR1_U1 ( .A0_t (OUT_ciphertext_s0_t[38]), .A0_f (OUT_ciphertext_s0_f[38]), .A1_t (OUT_ciphertext_s1_t[38]), .A1_f (OUT_ciphertext_s1_f[38]), .B0_t (LED_128_Instance_addroundkey_tmp[38]), .B0_f (new_AGEMA_signal_2991), .B1_t (new_AGEMA_signal_2992), .B1_f (new_AGEMA_signal_2993), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_38_U1_X), .Z0_f (new_AGEMA_signal_3366), .Z1_t (new_AGEMA_signal_3367), .Z1_f (new_AGEMA_signal_3368) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_38_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n23), .A1_f (new_AGEMA_signal_2480), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_38_U1_X), .B0_f (new_AGEMA_signal_3366), .B1_t (new_AGEMA_signal_3367), .B1_f (new_AGEMA_signal_3368), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_38_U1_Y), .Z0_f (new_AGEMA_signal_3558), .Z1_t (new_AGEMA_signal_3559), .Z1_f (new_AGEMA_signal_3560) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_38_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_38_U1_Y), .A0_f (new_AGEMA_signal_3558), .A1_t (new_AGEMA_signal_3559), .A1_f (new_AGEMA_signal_3560), .B0_t (OUT_ciphertext_s0_t[38]), .B0_f (OUT_ciphertext_s0_f[38]), .B1_t (OUT_ciphertext_s1_t[38]), .B1_f (OUT_ciphertext_s1_f[38]), .Z0_t (LED_128_Instance_addroundkey_out[38]), .Z0_f (new_AGEMA_signal_3750), .Z1_t (new_AGEMA_signal_3751), .Z1_f (new_AGEMA_signal_3752) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_39_U1_XOR1_U1 ( .A0_t (OUT_ciphertext_s0_t[39]), .A0_f (OUT_ciphertext_s0_f[39]), .A1_t (OUT_ciphertext_s1_t[39]), .A1_f (OUT_ciphertext_s1_f[39]), .B0_t (LED_128_Instance_addroundkey_tmp[39]), .B0_f (new_AGEMA_signal_3189), .B1_t (new_AGEMA_signal_3190), .B1_f (new_AGEMA_signal_3191), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_39_U1_X), .Z0_f (new_AGEMA_signal_3369), .Z1_t (new_AGEMA_signal_3370), .Z1_f (new_AGEMA_signal_3371) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_39_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n23), .A1_f (new_AGEMA_signal_2480), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_39_U1_X), .B0_f (new_AGEMA_signal_3369), .B1_t (new_AGEMA_signal_3370), .B1_f (new_AGEMA_signal_3371), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_39_U1_Y), .Z0_f (new_AGEMA_signal_3561), .Z1_t (new_AGEMA_signal_3562), .Z1_f (new_AGEMA_signal_3563) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_39_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_39_U1_Y), .A0_f (new_AGEMA_signal_3561), .A1_t (new_AGEMA_signal_3562), .A1_f (new_AGEMA_signal_3563), .B0_t (OUT_ciphertext_s0_t[39]), .B0_f (OUT_ciphertext_s0_f[39]), .B1_t (OUT_ciphertext_s1_t[39]), .B1_f (OUT_ciphertext_s1_f[39]), .Z0_t (LED_128_Instance_addconst_out[39]), .Z0_f (new_AGEMA_signal_3753), .Z1_t (new_AGEMA_signal_3754), .Z1_f (new_AGEMA_signal_3755) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_40_U1_XOR1_U1 ( .A0_t (OUT_ciphertext_s0_t[40]), .A0_f (OUT_ciphertext_s0_f[40]), .A1_t (OUT_ciphertext_s1_t[40]), .A1_f (OUT_ciphertext_s1_f[40]), .B0_t (LED_128_Instance_addroundkey_tmp[40]), .B0_f (new_AGEMA_signal_2955), .B1_t (new_AGEMA_signal_2956), .B1_f (new_AGEMA_signal_2957), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_40_U1_X), .Z0_f (new_AGEMA_signal_3372), .Z1_t (new_AGEMA_signal_3373), .Z1_f (new_AGEMA_signal_3374) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_40_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n23), .A1_f (new_AGEMA_signal_2480), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_40_U1_X), .B0_f (new_AGEMA_signal_3372), .B1_t (new_AGEMA_signal_3373), .B1_f (new_AGEMA_signal_3374), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_40_U1_Y), .Z0_f (new_AGEMA_signal_3564), .Z1_t (new_AGEMA_signal_3565), .Z1_f (new_AGEMA_signal_3566) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_40_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_40_U1_Y), .A0_f (new_AGEMA_signal_3564), .A1_t (new_AGEMA_signal_3565), .A1_f (new_AGEMA_signal_3566), .B0_t (OUT_ciphertext_s0_t[40]), .B0_f (OUT_ciphertext_s0_f[40]), .B1_t (OUT_ciphertext_s1_t[40]), .B1_f (OUT_ciphertext_s1_f[40]), .Z0_t (LED_128_Instance_addconst_out[40]), .Z0_f (new_AGEMA_signal_3756), .Z1_t (new_AGEMA_signal_3757), .Z1_f (new_AGEMA_signal_3758) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_41_U1_XOR1_U1 ( .A0_t (OUT_ciphertext_s0_t[41]), .A0_f (OUT_ciphertext_s0_f[41]), .A1_t (OUT_ciphertext_s1_t[41]), .A1_f (OUT_ciphertext_s1_f[41]), .B0_t (LED_128_Instance_addroundkey_tmp[41]), .B0_f (new_AGEMA_signal_3135), .B1_t (new_AGEMA_signal_3136), .B1_f (new_AGEMA_signal_3137), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_41_U1_X), .Z0_f (new_AGEMA_signal_3375), .Z1_t (new_AGEMA_signal_3376), .Z1_f (new_AGEMA_signal_3377) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_41_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n23), .A1_f (new_AGEMA_signal_2480), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_41_U1_X), .B0_f (new_AGEMA_signal_3375), .B1_t (new_AGEMA_signal_3376), .B1_f (new_AGEMA_signal_3377), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_41_U1_Y), .Z0_f (new_AGEMA_signal_3567), .Z1_t (new_AGEMA_signal_3568), .Z1_f (new_AGEMA_signal_3569) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_41_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_41_U1_Y), .A0_f (new_AGEMA_signal_3567), .A1_t (new_AGEMA_signal_3568), .A1_f (new_AGEMA_signal_3569), .B0_t (OUT_ciphertext_s0_t[41]), .B0_f (OUT_ciphertext_s0_f[41]), .B1_t (OUT_ciphertext_s1_t[41]), .B1_f (OUT_ciphertext_s1_f[41]), .Z0_t (LED_128_Instance_addconst_out[41]), .Z0_f (new_AGEMA_signal_3759), .Z1_t (new_AGEMA_signal_3760), .Z1_f (new_AGEMA_signal_3761) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_42_U1_XOR1_U1 ( .A0_t (OUT_ciphertext_s0_t[42]), .A0_f (OUT_ciphertext_s0_f[42]), .A1_t (OUT_ciphertext_s1_t[42]), .A1_f (OUT_ciphertext_s1_f[42]), .B0_t (LED_128_Instance_addroundkey_tmp[42]), .B0_f (new_AGEMA_signal_3087), .B1_t (new_AGEMA_signal_3088), .B1_f (new_AGEMA_signal_3089), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_42_U1_X), .Z0_f (new_AGEMA_signal_3378), .Z1_t (new_AGEMA_signal_3379), .Z1_f (new_AGEMA_signal_3380) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_42_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n23), .A1_f (new_AGEMA_signal_2480), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_42_U1_X), .B0_f (new_AGEMA_signal_3378), .B1_t (new_AGEMA_signal_3379), .B1_f (new_AGEMA_signal_3380), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_42_U1_Y), .Z0_f (new_AGEMA_signal_3570), .Z1_t (new_AGEMA_signal_3571), .Z1_f (new_AGEMA_signal_3572) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_42_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_42_U1_Y), .A0_f (new_AGEMA_signal_3570), .A1_t (new_AGEMA_signal_3571), .A1_f (new_AGEMA_signal_3572), .B0_t (OUT_ciphertext_s0_t[42]), .B0_f (OUT_ciphertext_s0_f[42]), .B1_t (OUT_ciphertext_s1_t[42]), .B1_f (OUT_ciphertext_s1_f[42]), .Z0_t (LED_128_Instance_addconst_out[42]), .Z0_f (new_AGEMA_signal_3762), .Z1_t (new_AGEMA_signal_3763), .Z1_f (new_AGEMA_signal_3764) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_43_U1_XOR1_U1 ( .A0_t (OUT_ciphertext_s0_t[43]), .A0_f (OUT_ciphertext_s0_f[43]), .A1_t (OUT_ciphertext_s1_t[43]), .A1_f (OUT_ciphertext_s1_f[43]), .B0_t (LED_128_Instance_addroundkey_tmp[43]), .B0_f (new_AGEMA_signal_3207), .B1_t (new_AGEMA_signal_3208), .B1_f (new_AGEMA_signal_3209), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_43_U1_X), .Z0_f (new_AGEMA_signal_3381), .Z1_t (new_AGEMA_signal_3382), .Z1_f (new_AGEMA_signal_3383) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_43_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n23), .A1_f (new_AGEMA_signal_2480), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_43_U1_X), .B0_f (new_AGEMA_signal_3381), .B1_t (new_AGEMA_signal_3382), .B1_f (new_AGEMA_signal_3383), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_43_U1_Y), .Z0_f (new_AGEMA_signal_3573), .Z1_t (new_AGEMA_signal_3574), .Z1_f (new_AGEMA_signal_3575) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_43_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_43_U1_Y), .A0_f (new_AGEMA_signal_3573), .A1_t (new_AGEMA_signal_3574), .A1_f (new_AGEMA_signal_3575), .B0_t (OUT_ciphertext_s0_t[43]), .B0_f (OUT_ciphertext_s0_f[43]), .B1_t (OUT_ciphertext_s1_t[43]), .B1_f (OUT_ciphertext_s1_f[43]), .Z0_t (LED_128_Instance_addconst_out[43]), .Z0_f (new_AGEMA_signal_3765), .Z1_t (new_AGEMA_signal_3766), .Z1_f (new_AGEMA_signal_3767) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_44_U1_XOR1_U1 ( .A0_t (OUT_ciphertext_s0_t[44]), .A0_f (OUT_ciphertext_s0_f[44]), .A1_t (OUT_ciphertext_s1_t[44]), .A1_f (OUT_ciphertext_s1_f[44]), .B0_t (LED_128_Instance_addroundkey_tmp[44]), .B0_f (new_AGEMA_signal_2949), .B1_t (new_AGEMA_signal_2950), .B1_f (new_AGEMA_signal_2951), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_44_U1_X), .Z0_f (new_AGEMA_signal_3384), .Z1_t (new_AGEMA_signal_3385), .Z1_f (new_AGEMA_signal_3386) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_44_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n23), .A1_f (new_AGEMA_signal_2480), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_44_U1_X), .B0_f (new_AGEMA_signal_3384), .B1_t (new_AGEMA_signal_3385), .B1_f (new_AGEMA_signal_3386), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_44_U1_Y), .Z0_f (new_AGEMA_signal_3576), .Z1_t (new_AGEMA_signal_3577), .Z1_f (new_AGEMA_signal_3578) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_44_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_44_U1_Y), .A0_f (new_AGEMA_signal_3576), .A1_t (new_AGEMA_signal_3577), .A1_f (new_AGEMA_signal_3578), .B0_t (OUT_ciphertext_s0_t[44]), .B0_f (OUT_ciphertext_s0_f[44]), .B1_t (OUT_ciphertext_s1_t[44]), .B1_f (OUT_ciphertext_s1_f[44]), .Z0_t (LED_128_Instance_addconst_out[44]), .Z0_f (new_AGEMA_signal_3768), .Z1_t (new_AGEMA_signal_3769), .Z1_f (new_AGEMA_signal_3770) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_45_U1_XOR1_U1 ( .A0_t (OUT_ciphertext_s0_t[45]), .A0_f (OUT_ciphertext_s0_f[45]), .A1_t (OUT_ciphertext_s1_t[45]), .A1_f (OUT_ciphertext_s1_f[45]), .B0_t (LED_128_Instance_addroundkey_tmp[45]), .B0_f (new_AGEMA_signal_3129), .B1_t (new_AGEMA_signal_3130), .B1_f (new_AGEMA_signal_3131), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_45_U1_X), .Z0_f (new_AGEMA_signal_3387), .Z1_t (new_AGEMA_signal_3388), .Z1_f (new_AGEMA_signal_3389) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_45_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n23), .A1_f (new_AGEMA_signal_2480), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_45_U1_X), .B0_f (new_AGEMA_signal_3387), .B1_t (new_AGEMA_signal_3388), .B1_f (new_AGEMA_signal_3389), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_45_U1_Y), .Z0_f (new_AGEMA_signal_3579), .Z1_t (new_AGEMA_signal_3580), .Z1_f (new_AGEMA_signal_3581) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_45_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_45_U1_Y), .A0_f (new_AGEMA_signal_3579), .A1_t (new_AGEMA_signal_3580), .A1_f (new_AGEMA_signal_3581), .B0_t (OUT_ciphertext_s0_t[45]), .B0_f (OUT_ciphertext_s0_f[45]), .B1_t (OUT_ciphertext_s1_t[45]), .B1_f (OUT_ciphertext_s1_f[45]), .Z0_t (LED_128_Instance_addconst_out[45]), .Z0_f (new_AGEMA_signal_3771), .Z1_t (new_AGEMA_signal_3772), .Z1_f (new_AGEMA_signal_3773) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_46_U1_XOR1_U1 ( .A0_t (OUT_ciphertext_s0_t[46]), .A0_f (OUT_ciphertext_s0_f[46]), .A1_t (OUT_ciphertext_s1_t[46]), .A1_f (OUT_ciphertext_s1_f[46]), .B0_t (LED_128_Instance_addroundkey_tmp[46]), .B0_f (new_AGEMA_signal_3081), .B1_t (new_AGEMA_signal_3082), .B1_f (new_AGEMA_signal_3083), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_46_U1_X), .Z0_f (new_AGEMA_signal_3390), .Z1_t (new_AGEMA_signal_3391), .Z1_f (new_AGEMA_signal_3392) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_46_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n23), .A1_f (new_AGEMA_signal_2480), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_46_U1_X), .B0_f (new_AGEMA_signal_3390), .B1_t (new_AGEMA_signal_3391), .B1_f (new_AGEMA_signal_3392), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_46_U1_Y), .Z0_f (new_AGEMA_signal_3582), .Z1_t (new_AGEMA_signal_3583), .Z1_f (new_AGEMA_signal_3584) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_46_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_46_U1_Y), .A0_f (new_AGEMA_signal_3582), .A1_t (new_AGEMA_signal_3583), .A1_f (new_AGEMA_signal_3584), .B0_t (OUT_ciphertext_s0_t[46]), .B0_f (OUT_ciphertext_s0_f[46]), .B1_t (OUT_ciphertext_s1_t[46]), .B1_f (OUT_ciphertext_s1_f[46]), .Z0_t (LED_128_Instance_addconst_out[46]), .Z0_f (new_AGEMA_signal_3774), .Z1_t (new_AGEMA_signal_3775), .Z1_f (new_AGEMA_signal_3776) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_47_U1_XOR1_U1 ( .A0_t (OUT_ciphertext_s0_t[47]), .A0_f (OUT_ciphertext_s0_f[47]), .A1_t (OUT_ciphertext_s1_t[47]), .A1_f (OUT_ciphertext_s1_f[47]), .B0_t (LED_128_Instance_addroundkey_tmp[47]), .B0_f (new_AGEMA_signal_3201), .B1_t (new_AGEMA_signal_3202), .B1_f (new_AGEMA_signal_3203), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_47_U1_X), .Z0_f (new_AGEMA_signal_3393), .Z1_t (new_AGEMA_signal_3394), .Z1_f (new_AGEMA_signal_3395) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_47_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n23), .A1_f (new_AGEMA_signal_2480), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_47_U1_X), .B0_f (new_AGEMA_signal_3393), .B1_t (new_AGEMA_signal_3394), .B1_f (new_AGEMA_signal_3395), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_47_U1_Y), .Z0_f (new_AGEMA_signal_3585), .Z1_t (new_AGEMA_signal_3586), .Z1_f (new_AGEMA_signal_3587) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_47_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_47_U1_Y), .A0_f (new_AGEMA_signal_3585), .A1_t (new_AGEMA_signal_3586), .A1_f (new_AGEMA_signal_3587), .B0_t (OUT_ciphertext_s0_t[47]), .B0_f (OUT_ciphertext_s0_f[47]), .B1_t (OUT_ciphertext_s1_t[47]), .B1_f (OUT_ciphertext_s1_f[47]), .Z0_t (LED_128_Instance_addconst_out[47]), .Z0_f (new_AGEMA_signal_3777), .Z1_t (new_AGEMA_signal_3778), .Z1_f (new_AGEMA_signal_3779) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_48_U1_XOR1_U1 ( .A0_t (OUT_ciphertext_s0_t[48]), .A0_f (OUT_ciphertext_s0_f[48]), .A1_t (OUT_ciphertext_s1_t[48]), .A1_f (OUT_ciphertext_s1_f[48]), .B0_t (LED_128_Instance_addroundkey_tmp[48]), .B0_f (new_AGEMA_signal_2901), .B1_t (new_AGEMA_signal_2902), .B1_f (new_AGEMA_signal_2903), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_48_U1_X), .Z0_f (new_AGEMA_signal_3396), .Z1_t (new_AGEMA_signal_3397), .Z1_f (new_AGEMA_signal_3398) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_48_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n23), .A1_f (new_AGEMA_signal_2480), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_48_U1_X), .B0_f (new_AGEMA_signal_3396), .B1_t (new_AGEMA_signal_3397), .B1_f (new_AGEMA_signal_3398), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_48_U1_Y), .Z0_f (new_AGEMA_signal_3588), .Z1_t (new_AGEMA_signal_3589), .Z1_f (new_AGEMA_signal_3590) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_48_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_48_U1_Y), .A0_f (new_AGEMA_signal_3588), .A1_t (new_AGEMA_signal_3589), .A1_f (new_AGEMA_signal_3590), .B0_t (OUT_ciphertext_s0_t[48]), .B0_f (OUT_ciphertext_s0_f[48]), .B1_t (OUT_ciphertext_s1_t[48]), .B1_f (OUT_ciphertext_s1_f[48]), .Z0_t (LED_128_Instance_addroundkey_out[48]), .Z0_f (new_AGEMA_signal_3780), .Z1_t (new_AGEMA_signal_3781), .Z1_f (new_AGEMA_signal_3782) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_49_U1_XOR1_U1 ( .A0_t (OUT_ciphertext_s0_t[49]), .A0_f (OUT_ciphertext_s0_f[49]), .A1_t (OUT_ciphertext_s1_t[49]), .A1_f (OUT_ciphertext_s1_f[49]), .B0_t (LED_128_Instance_addroundkey_tmp[49]), .B0_f (new_AGEMA_signal_2967), .B1_t (new_AGEMA_signal_2968), .B1_f (new_AGEMA_signal_2969), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_49_U1_X), .Z0_f (new_AGEMA_signal_3399), .Z1_t (new_AGEMA_signal_3400), .Z1_f (new_AGEMA_signal_3401) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_49_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n23), .A1_f (new_AGEMA_signal_2480), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_49_U1_X), .B0_f (new_AGEMA_signal_3399), .B1_t (new_AGEMA_signal_3400), .B1_f (new_AGEMA_signal_3401), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_49_U1_Y), .Z0_f (new_AGEMA_signal_3591), .Z1_t (new_AGEMA_signal_3592), .Z1_f (new_AGEMA_signal_3593) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_49_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_49_U1_Y), .A0_f (new_AGEMA_signal_3591), .A1_t (new_AGEMA_signal_3592), .A1_f (new_AGEMA_signal_3593), .B0_t (OUT_ciphertext_s0_t[49]), .B0_f (OUT_ciphertext_s0_f[49]), .B1_t (OUT_ciphertext_s1_t[49]), .B1_f (OUT_ciphertext_s1_f[49]), .Z0_t (LED_128_Instance_addroundkey_out[49]), .Z0_f (new_AGEMA_signal_3783), .Z1_t (new_AGEMA_signal_3784), .Z1_f (new_AGEMA_signal_3785) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_50_U1_XOR1_U1 ( .A0_t (OUT_ciphertext_s0_t[50]), .A0_f (OUT_ciphertext_s0_f[50]), .A1_t (OUT_ciphertext_s1_t[50]), .A1_f (OUT_ciphertext_s1_f[50]), .B0_t (LED_128_Instance_addroundkey_tmp[50]), .B0_f (new_AGEMA_signal_3063), .B1_t (new_AGEMA_signal_3064), .B1_f (new_AGEMA_signal_3065), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_50_U1_X), .Z0_f (new_AGEMA_signal_3402), .Z1_t (new_AGEMA_signal_3403), .Z1_f (new_AGEMA_signal_3404) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_50_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n23), .A1_f (new_AGEMA_signal_2480), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_50_U1_X), .B0_f (new_AGEMA_signal_3402), .B1_t (new_AGEMA_signal_3403), .B1_f (new_AGEMA_signal_3404), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_50_U1_Y), .Z0_f (new_AGEMA_signal_3594), .Z1_t (new_AGEMA_signal_3595), .Z1_f (new_AGEMA_signal_3596) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_50_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_50_U1_Y), .A0_f (new_AGEMA_signal_3594), .A1_t (new_AGEMA_signal_3595), .A1_f (new_AGEMA_signal_3596), .B0_t (OUT_ciphertext_s0_t[50]), .B0_f (OUT_ciphertext_s0_f[50]), .B1_t (OUT_ciphertext_s1_t[50]), .B1_f (OUT_ciphertext_s1_f[50]), .Z0_t (LED_128_Instance_addconst_out[50]), .Z0_f (new_AGEMA_signal_3786), .Z1_t (new_AGEMA_signal_3787), .Z1_f (new_AGEMA_signal_3788) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_51_U1_XOR1_U1 ( .A0_t (OUT_ciphertext_s0_t[51]), .A0_f (OUT_ciphertext_s0_f[51]), .A1_t (OUT_ciphertext_s1_t[51]), .A1_f (OUT_ciphertext_s1_f[51]), .B0_t (LED_128_Instance_addroundkey_tmp[51]), .B0_f (new_AGEMA_signal_3225), .B1_t (new_AGEMA_signal_3226), .B1_f (new_AGEMA_signal_3227), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_51_U1_X), .Z0_f (new_AGEMA_signal_3405), .Z1_t (new_AGEMA_signal_3406), .Z1_f (new_AGEMA_signal_3407) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_51_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n23), .A1_f (new_AGEMA_signal_2480), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_51_U1_X), .B0_f (new_AGEMA_signal_3405), .B1_t (new_AGEMA_signal_3406), .B1_f (new_AGEMA_signal_3407), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_51_U1_Y), .Z0_f (new_AGEMA_signal_3597), .Z1_t (new_AGEMA_signal_3598), .Z1_f (new_AGEMA_signal_3599) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_51_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_51_U1_Y), .A0_f (new_AGEMA_signal_3597), .A1_t (new_AGEMA_signal_3598), .A1_f (new_AGEMA_signal_3599), .B0_t (OUT_ciphertext_s0_t[51]), .B0_f (OUT_ciphertext_s0_f[51]), .B1_t (OUT_ciphertext_s1_t[51]), .B1_f (OUT_ciphertext_s1_f[51]), .Z0_t (LED_128_Instance_addconst_out[51]), .Z0_f (new_AGEMA_signal_3789), .Z1_t (new_AGEMA_signal_3790), .Z1_f (new_AGEMA_signal_3791) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_52_U1_XOR1_U1 ( .A0_t (OUT_ciphertext_s0_t[52]), .A0_f (OUT_ciphertext_s0_f[52]), .A1_t (OUT_ciphertext_s1_t[52]), .A1_f (OUT_ciphertext_s1_f[52]), .B0_t (LED_128_Instance_addroundkey_tmp[52]), .B0_f (new_AGEMA_signal_3003), .B1_t (new_AGEMA_signal_3004), .B1_f (new_AGEMA_signal_3005), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_52_U1_X), .Z0_f (new_AGEMA_signal_3408), .Z1_t (new_AGEMA_signal_3409), .Z1_f (new_AGEMA_signal_3410) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_52_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n23), .A1_f (new_AGEMA_signal_2480), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_52_U1_X), .B0_f (new_AGEMA_signal_3408), .B1_t (new_AGEMA_signal_3409), .B1_f (new_AGEMA_signal_3410), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_52_U1_Y), .Z0_f (new_AGEMA_signal_3600), .Z1_t (new_AGEMA_signal_3601), .Z1_f (new_AGEMA_signal_3602) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_52_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_52_U1_Y), .A0_f (new_AGEMA_signal_3600), .A1_t (new_AGEMA_signal_3601), .A1_f (new_AGEMA_signal_3602), .B0_t (OUT_ciphertext_s0_t[52]), .B0_f (OUT_ciphertext_s0_f[52]), .B1_t (OUT_ciphertext_s1_t[52]), .B1_f (OUT_ciphertext_s1_f[52]), .Z0_t (LED_128_Instance_addroundkey_out[52]), .Z0_f (new_AGEMA_signal_3792), .Z1_t (new_AGEMA_signal_3793), .Z1_f (new_AGEMA_signal_3794) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_53_U1_XOR1_U1 ( .A0_t (OUT_ciphertext_s0_t[53]), .A0_f (OUT_ciphertext_s0_f[53]), .A1_t (OUT_ciphertext_s1_t[53]), .A1_f (OUT_ciphertext_s1_f[53]), .B0_t (LED_128_Instance_addroundkey_tmp[53]), .B0_f (new_AGEMA_signal_3015), .B1_t (new_AGEMA_signal_3016), .B1_f (new_AGEMA_signal_3017), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_53_U1_X), .Z0_f (new_AGEMA_signal_3411), .Z1_t (new_AGEMA_signal_3412), .Z1_f (new_AGEMA_signal_3413) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_53_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n23), .A1_f (new_AGEMA_signal_2480), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_53_U1_X), .B0_f (new_AGEMA_signal_3411), .B1_t (new_AGEMA_signal_3412), .B1_f (new_AGEMA_signal_3413), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_53_U1_Y), .Z0_f (new_AGEMA_signal_3603), .Z1_t (new_AGEMA_signal_3604), .Z1_f (new_AGEMA_signal_3605) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_53_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_53_U1_Y), .A0_f (new_AGEMA_signal_3603), .A1_t (new_AGEMA_signal_3604), .A1_f (new_AGEMA_signal_3605), .B0_t (OUT_ciphertext_s0_t[53]), .B0_f (OUT_ciphertext_s0_f[53]), .B1_t (OUT_ciphertext_s1_t[53]), .B1_f (OUT_ciphertext_s1_f[53]), .Z0_t (LED_128_Instance_addroundkey_out[53]), .Z0_f (new_AGEMA_signal_3795), .Z1_t (new_AGEMA_signal_3796), .Z1_f (new_AGEMA_signal_3797) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_54_U1_XOR1_U1 ( .A0_t (OUT_ciphertext_s0_t[54]), .A0_f (OUT_ciphertext_s0_f[54]), .A1_t (OUT_ciphertext_s1_t[54]), .A1_f (OUT_ciphertext_s1_f[54]), .B0_t (LED_128_Instance_addroundkey_tmp[54]), .B0_f (new_AGEMA_signal_2985), .B1_t (new_AGEMA_signal_2986), .B1_f (new_AGEMA_signal_2987), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_54_U1_X), .Z0_f (new_AGEMA_signal_3414), .Z1_t (new_AGEMA_signal_3415), .Z1_f (new_AGEMA_signal_3416) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_54_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n23), .A1_f (new_AGEMA_signal_2480), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_54_U1_X), .B0_f (new_AGEMA_signal_3414), .B1_t (new_AGEMA_signal_3415), .B1_f (new_AGEMA_signal_3416), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_54_U1_Y), .Z0_f (new_AGEMA_signal_3606), .Z1_t (new_AGEMA_signal_3607), .Z1_f (new_AGEMA_signal_3608) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_54_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_54_U1_Y), .A0_f (new_AGEMA_signal_3606), .A1_t (new_AGEMA_signal_3607), .A1_f (new_AGEMA_signal_3608), .B0_t (OUT_ciphertext_s0_t[54]), .B0_f (OUT_ciphertext_s0_f[54]), .B1_t (OUT_ciphertext_s1_t[54]), .B1_f (OUT_ciphertext_s1_f[54]), .Z0_t (LED_128_Instance_addroundkey_out[54]), .Z0_f (new_AGEMA_signal_3798), .Z1_t (new_AGEMA_signal_3799), .Z1_f (new_AGEMA_signal_3800) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_55_U1_XOR1_U1 ( .A0_t (OUT_ciphertext_s0_t[55]), .A0_f (OUT_ciphertext_s0_f[55]), .A1_t (OUT_ciphertext_s1_t[55]), .A1_f (OUT_ciphertext_s1_f[55]), .B0_t (LED_128_Instance_addroundkey_tmp[55]), .B0_f (new_AGEMA_signal_3219), .B1_t (new_AGEMA_signal_3220), .B1_f (new_AGEMA_signal_3221), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_55_U1_X), .Z0_f (new_AGEMA_signal_3417), .Z1_t (new_AGEMA_signal_3418), .Z1_f (new_AGEMA_signal_3419) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_55_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n23), .A1_f (new_AGEMA_signal_2480), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_55_U1_X), .B0_f (new_AGEMA_signal_3417), .B1_t (new_AGEMA_signal_3418), .B1_f (new_AGEMA_signal_3419), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_55_U1_Y), .Z0_f (new_AGEMA_signal_3609), .Z1_t (new_AGEMA_signal_3610), .Z1_f (new_AGEMA_signal_3611) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_55_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_55_U1_Y), .A0_f (new_AGEMA_signal_3609), .A1_t (new_AGEMA_signal_3610), .A1_f (new_AGEMA_signal_3611), .B0_t (OUT_ciphertext_s0_t[55]), .B0_f (OUT_ciphertext_s0_f[55]), .B1_t (OUT_ciphertext_s1_t[55]), .B1_f (OUT_ciphertext_s1_f[55]), .Z0_t (LED_128_Instance_addconst_out[55]), .Z0_f (new_AGEMA_signal_3801), .Z1_t (new_AGEMA_signal_3802), .Z1_f (new_AGEMA_signal_3803) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_56_U1_XOR1_U1 ( .A0_t (OUT_ciphertext_s0_t[56]), .A0_f (OUT_ciphertext_s0_f[56]), .A1_t (OUT_ciphertext_s1_t[56]), .A1_f (OUT_ciphertext_s1_f[56]), .B0_t (LED_128_Instance_addroundkey_tmp[56]), .B0_f (new_AGEMA_signal_2913), .B1_t (new_AGEMA_signal_2914), .B1_f (new_AGEMA_signal_2915), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_56_U1_X), .Z0_f (new_AGEMA_signal_3420), .Z1_t (new_AGEMA_signal_3421), .Z1_f (new_AGEMA_signal_3422) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_56_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n23), .A1_f (new_AGEMA_signal_2480), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_56_U1_X), .B0_f (new_AGEMA_signal_3420), .B1_t (new_AGEMA_signal_3421), .B1_f (new_AGEMA_signal_3422), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_56_U1_Y), .Z0_f (new_AGEMA_signal_3612), .Z1_t (new_AGEMA_signal_3613), .Z1_f (new_AGEMA_signal_3614) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_56_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_56_U1_Y), .A0_f (new_AGEMA_signal_3612), .A1_t (new_AGEMA_signal_3613), .A1_f (new_AGEMA_signal_3614), .B0_t (OUT_ciphertext_s0_t[56]), .B0_f (OUT_ciphertext_s0_f[56]), .B1_t (OUT_ciphertext_s1_t[56]), .B1_f (OUT_ciphertext_s1_f[56]), .Z0_t (LED_128_Instance_addconst_out[56]), .Z0_f (new_AGEMA_signal_3804), .Z1_t (new_AGEMA_signal_3805), .Z1_f (new_AGEMA_signal_3806) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_57_U1_XOR1_U1 ( .A0_t (OUT_ciphertext_s0_t[57]), .A0_f (OUT_ciphertext_s0_f[57]), .A1_t (OUT_ciphertext_s1_t[57]), .A1_f (OUT_ciphertext_s1_f[57]), .B0_t (LED_128_Instance_addroundkey_tmp[57]), .B0_f (new_AGEMA_signal_3141), .B1_t (new_AGEMA_signal_3142), .B1_f (new_AGEMA_signal_3143), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_57_U1_X), .Z0_f (new_AGEMA_signal_3423), .Z1_t (new_AGEMA_signal_3424), .Z1_f (new_AGEMA_signal_3425) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_57_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n23), .A1_f (new_AGEMA_signal_2480), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_57_U1_X), .B0_f (new_AGEMA_signal_3423), .B1_t (new_AGEMA_signal_3424), .B1_f (new_AGEMA_signal_3425), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_57_U1_Y), .Z0_f (new_AGEMA_signal_3615), .Z1_t (new_AGEMA_signal_3616), .Z1_f (new_AGEMA_signal_3617) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_57_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_57_U1_Y), .A0_f (new_AGEMA_signal_3615), .A1_t (new_AGEMA_signal_3616), .A1_f (new_AGEMA_signal_3617), .B0_t (OUT_ciphertext_s0_t[57]), .B0_f (OUT_ciphertext_s0_f[57]), .B1_t (OUT_ciphertext_s1_t[57]), .B1_f (OUT_ciphertext_s1_f[57]), .Z0_t (LED_128_Instance_addconst_out[57]), .Z0_f (new_AGEMA_signal_3807), .Z1_t (new_AGEMA_signal_3808), .Z1_f (new_AGEMA_signal_3809) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_58_U1_XOR1_U1 ( .A0_t (OUT_ciphertext_s0_t[58]), .A0_f (OUT_ciphertext_s0_f[58]), .A1_t (OUT_ciphertext_s1_t[58]), .A1_f (OUT_ciphertext_s1_f[58]), .B0_t (LED_128_Instance_addroundkey_tmp[58]), .B0_f (new_AGEMA_signal_3057), .B1_t (new_AGEMA_signal_3058), .B1_f (new_AGEMA_signal_3059), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_58_U1_X), .Z0_f (new_AGEMA_signal_3426), .Z1_t (new_AGEMA_signal_3427), .Z1_f (new_AGEMA_signal_3428) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_58_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n23), .A1_f (new_AGEMA_signal_2480), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_58_U1_X), .B0_f (new_AGEMA_signal_3426), .B1_t (new_AGEMA_signal_3427), .B1_f (new_AGEMA_signal_3428), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_58_U1_Y), .Z0_f (new_AGEMA_signal_3618), .Z1_t (new_AGEMA_signal_3619), .Z1_f (new_AGEMA_signal_3620) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_58_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_58_U1_Y), .A0_f (new_AGEMA_signal_3618), .A1_t (new_AGEMA_signal_3619), .A1_f (new_AGEMA_signal_3620), .B0_t (OUT_ciphertext_s0_t[58]), .B0_f (OUT_ciphertext_s0_f[58]), .B1_t (OUT_ciphertext_s1_t[58]), .B1_f (OUT_ciphertext_s1_f[58]), .Z0_t (LED_128_Instance_addconst_out[58]), .Z0_f (new_AGEMA_signal_3810), .Z1_t (new_AGEMA_signal_3811), .Z1_f (new_AGEMA_signal_3812) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_59_U1_XOR1_U1 ( .A0_t (OUT_ciphertext_s0_t[59]), .A0_f (OUT_ciphertext_s0_f[59]), .A1_t (OUT_ciphertext_s1_t[59]), .A1_f (OUT_ciphertext_s1_f[59]), .B0_t (LED_128_Instance_addroundkey_tmp[59]), .B0_f (new_AGEMA_signal_3213), .B1_t (new_AGEMA_signal_3214), .B1_f (new_AGEMA_signal_3215), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_59_U1_X), .Z0_f (new_AGEMA_signal_3429), .Z1_t (new_AGEMA_signal_3430), .Z1_f (new_AGEMA_signal_3431) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_59_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n23), .A1_f (new_AGEMA_signal_2480), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_59_U1_X), .B0_f (new_AGEMA_signal_3429), .B1_t (new_AGEMA_signal_3430), .B1_f (new_AGEMA_signal_3431), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_59_U1_Y), .Z0_f (new_AGEMA_signal_3621), .Z1_t (new_AGEMA_signal_3622), .Z1_f (new_AGEMA_signal_3623) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_59_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_59_U1_Y), .A0_f (new_AGEMA_signal_3621), .A1_t (new_AGEMA_signal_3622), .A1_f (new_AGEMA_signal_3623), .B0_t (OUT_ciphertext_s0_t[59]), .B0_f (OUT_ciphertext_s0_f[59]), .B1_t (OUT_ciphertext_s1_t[59]), .B1_f (OUT_ciphertext_s1_f[59]), .Z0_t (LED_128_Instance_addconst_out[59]), .Z0_f (new_AGEMA_signal_3813), .Z1_t (new_AGEMA_signal_3814), .Z1_f (new_AGEMA_signal_3815) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_60_U1_XOR1_U1 ( .A0_t (OUT_ciphertext_s0_t[60]), .A0_f (OUT_ciphertext_s0_f[60]), .A1_t (OUT_ciphertext_s1_t[60]), .A1_f (OUT_ciphertext_s1_f[60]), .B0_t (LED_128_Instance_addroundkey_tmp[60]), .B0_f (new_AGEMA_signal_2919), .B1_t (new_AGEMA_signal_2920), .B1_f (new_AGEMA_signal_2921), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_60_U1_X), .Z0_f (new_AGEMA_signal_3432), .Z1_t (new_AGEMA_signal_3433), .Z1_f (new_AGEMA_signal_3434) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_60_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n23), .A1_f (new_AGEMA_signal_2480), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_60_U1_X), .B0_f (new_AGEMA_signal_3432), .B1_t (new_AGEMA_signal_3433), .B1_f (new_AGEMA_signal_3434), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_60_U1_Y), .Z0_f (new_AGEMA_signal_3624), .Z1_t (new_AGEMA_signal_3625), .Z1_f (new_AGEMA_signal_3626) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_60_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_60_U1_Y), .A0_f (new_AGEMA_signal_3624), .A1_t (new_AGEMA_signal_3625), .A1_f (new_AGEMA_signal_3626), .B0_t (OUT_ciphertext_s0_t[60]), .B0_f (OUT_ciphertext_s0_f[60]), .B1_t (OUT_ciphertext_s1_t[60]), .B1_f (OUT_ciphertext_s1_f[60]), .Z0_t (LED_128_Instance_addconst_out[60]), .Z0_f (new_AGEMA_signal_3816), .Z1_t (new_AGEMA_signal_3817), .Z1_f (new_AGEMA_signal_3818) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_61_U1_XOR1_U1 ( .A0_t (OUT_ciphertext_s0_t[61]), .A0_f (OUT_ciphertext_s0_f[61]), .A1_t (OUT_ciphertext_s1_t[61]), .A1_f (OUT_ciphertext_s1_f[61]), .B0_t (LED_128_Instance_addroundkey_tmp[61]), .B0_f (new_AGEMA_signal_3147), .B1_t (new_AGEMA_signal_3148), .B1_f (new_AGEMA_signal_3149), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_61_U1_X), .Z0_f (new_AGEMA_signal_3435), .Z1_t (new_AGEMA_signal_3436), .Z1_f (new_AGEMA_signal_3437) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_61_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n23), .A1_f (new_AGEMA_signal_2480), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_61_U1_X), .B0_f (new_AGEMA_signal_3435), .B1_t (new_AGEMA_signal_3436), .B1_f (new_AGEMA_signal_3437), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_61_U1_Y), .Z0_f (new_AGEMA_signal_3627), .Z1_t (new_AGEMA_signal_3628), .Z1_f (new_AGEMA_signal_3629) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_61_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_61_U1_Y), .A0_f (new_AGEMA_signal_3627), .A1_t (new_AGEMA_signal_3628), .A1_f (new_AGEMA_signal_3629), .B0_t (OUT_ciphertext_s0_t[61]), .B0_f (OUT_ciphertext_s0_f[61]), .B1_t (OUT_ciphertext_s1_t[61]), .B1_f (OUT_ciphertext_s1_f[61]), .Z0_t (LED_128_Instance_addconst_out[61]), .Z0_f (new_AGEMA_signal_3819), .Z1_t (new_AGEMA_signal_3820), .Z1_f (new_AGEMA_signal_3821) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_62_U1_XOR1_U1 ( .A0_t (OUT_ciphertext_s0_t[62]), .A0_f (OUT_ciphertext_s0_f[62]), .A1_t (OUT_ciphertext_s1_t[62]), .A1_f (OUT_ciphertext_s1_f[62]), .B0_t (LED_128_Instance_addroundkey_tmp[62]), .B0_f (new_AGEMA_signal_3069), .B1_t (new_AGEMA_signal_3070), .B1_f (new_AGEMA_signal_3071), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_62_U1_X), .Z0_f (new_AGEMA_signal_3438), .Z1_t (new_AGEMA_signal_3439), .Z1_f (new_AGEMA_signal_3440) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_62_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n23), .A1_f (new_AGEMA_signal_2480), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_62_U1_X), .B0_f (new_AGEMA_signal_3438), .B1_t (new_AGEMA_signal_3439), .B1_f (new_AGEMA_signal_3440), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_62_U1_Y), .Z0_f (new_AGEMA_signal_3630), .Z1_t (new_AGEMA_signal_3631), .Z1_f (new_AGEMA_signal_3632) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_62_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_62_U1_Y), .A0_f (new_AGEMA_signal_3630), .A1_t (new_AGEMA_signal_3631), .A1_f (new_AGEMA_signal_3632), .B0_t (OUT_ciphertext_s0_t[62]), .B0_f (OUT_ciphertext_s0_f[62]), .B1_t (OUT_ciphertext_s1_t[62]), .B1_f (OUT_ciphertext_s1_f[62]), .Z0_t (LED_128_Instance_addconst_out[62]), .Z0_f (new_AGEMA_signal_3822), .Z1_t (new_AGEMA_signal_3823), .Z1_f (new_AGEMA_signal_3824) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_63_U1_XOR1_U1 ( .A0_t (OUT_ciphertext_s0_t[63]), .A0_f (OUT_ciphertext_s0_f[63]), .A1_t (OUT_ciphertext_s1_t[63]), .A1_f (OUT_ciphertext_s1_f[63]), .B0_t (LED_128_Instance_addroundkey_tmp[63]), .B0_f (new_AGEMA_signal_3231), .B1_t (new_AGEMA_signal_3232), .B1_f (new_AGEMA_signal_3233), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_63_U1_X), .Z0_f (new_AGEMA_signal_3441), .Z1_t (new_AGEMA_signal_3442), .Z1_f (new_AGEMA_signal_3443) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_63_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (LED_128_Instance_n23), .A1_f (new_AGEMA_signal_2480), .B0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_63_U1_X), .B0_f (new_AGEMA_signal_3441), .B1_t (new_AGEMA_signal_3442), .B1_f (new_AGEMA_signal_3443), .Z0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_63_U1_Y), .Z0_f (new_AGEMA_signal_3633), .Z1_t (new_AGEMA_signal_3634), .Z1_f (new_AGEMA_signal_3635) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MUX_addroundkey_out_mux_inst_63_U1_XOR2_U1 ( .A0_t (LED_128_Instance_MUX_addroundkey_out_mux_inst_63_U1_Y), .A0_f (new_AGEMA_signal_3633), .A1_t (new_AGEMA_signal_3634), .A1_f (new_AGEMA_signal_3635), .B0_t (OUT_ciphertext_s0_t[63]), .B0_f (OUT_ciphertext_s0_f[63]), .B1_t (OUT_ciphertext_s1_t[63]), .B1_f (OUT_ciphertext_s1_f[63]), .Z0_t (LED_128_Instance_addconst_out[63]), .Z0_f (new_AGEMA_signal_3825), .Z1_t (new_AGEMA_signal_3826), .Z1_f (new_AGEMA_signal_3827) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_AddConstants_instance_U14 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (roundconstant[2]), .A1_f (new_AGEMA_signal_1887), .B0_t (LED_128_Instance_addroundkey_out[54]), .B0_f (new_AGEMA_signal_3798), .B1_t (new_AGEMA_signal_3799), .B1_f (new_AGEMA_signal_3800), .Z0_t (LED_128_Instance_addconst_out[54]), .Z0_f (new_AGEMA_signal_3828), .Z1_t (new_AGEMA_signal_3829), .Z1_f (new_AGEMA_signal_3830) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_AddConstants_instance_U13 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (roundconstant[5]), .A1_f (new_AGEMA_signal_1877), .B0_t (LED_128_Instance_addroundkey_out[38]), .B0_f (new_AGEMA_signal_3750), .B1_t (new_AGEMA_signal_3751), .B1_f (new_AGEMA_signal_3752), .Z0_t (LED_128_Instance_addconst_out[38]), .Z0_f (new_AGEMA_signal_3831), .Z1_t (new_AGEMA_signal_3832), .Z1_f (new_AGEMA_signal_3833) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_AddConstants_instance_U12 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (roundconstant[5]), .A1_f (new_AGEMA_signal_1877), .B0_t (LED_128_Instance_addroundkey_out[6]), .B0_f (new_AGEMA_signal_3654), .B1_t (new_AGEMA_signal_3655), .B1_f (new_AGEMA_signal_3656), .Z0_t (LED_128_Instance_addconst_out[6]), .Z0_f (new_AGEMA_signal_3834), .Z1_t (new_AGEMA_signal_3835), .Z1_f (new_AGEMA_signal_3836) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_AddConstants_instance_U11 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (roundconstant[2]), .A1_f (new_AGEMA_signal_1887), .B0_t (LED_128_Instance_addroundkey_out[22]), .B0_f (new_AGEMA_signal_3702), .B1_t (new_AGEMA_signal_3703), .B1_f (new_AGEMA_signal_3704), .Z0_t (LED_128_Instance_addconst_out[22]), .Z0_f (new_AGEMA_signal_3837), .Z1_t (new_AGEMA_signal_3838), .Z1_f (new_AGEMA_signal_3839) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_AddConstants_instance_U10 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (roundconstant[3]), .A1_f (new_AGEMA_signal_1880), .B0_t (LED_128_Instance_addroundkey_out[36]), .B0_f (new_AGEMA_signal_3744), .B1_t (new_AGEMA_signal_3745), .B1_f (new_AGEMA_signal_3746), .Z0_t (LED_128_Instance_addconst_out[36]), .Z0_f (new_AGEMA_signal_3840), .Z1_t (new_AGEMA_signal_3841), .Z1_f (new_AGEMA_signal_3842) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_AddConstants_instance_U9 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (roundconstant[3]), .A1_f (new_AGEMA_signal_1880), .B0_t (LED_128_Instance_addroundkey_out[4]), .B0_f (new_AGEMA_signal_3648), .B1_t (new_AGEMA_signal_3649), .B1_f (new_AGEMA_signal_3650), .Z0_t (LED_128_Instance_addconst_out[4]), .Z0_f (new_AGEMA_signal_3843), .Z1_t (new_AGEMA_signal_3844), .Z1_f (new_AGEMA_signal_3845) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_AddConstants_instance_U8 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (roundconstant[0]), .A1_f (new_AGEMA_signal_1888), .B0_t (LED_128_Instance_addroundkey_out[52]), .B0_f (new_AGEMA_signal_3792), .B1_t (new_AGEMA_signal_3793), .B1_f (new_AGEMA_signal_3794), .Z0_t (LED_128_Instance_addconst_out[52]), .Z0_f (new_AGEMA_signal_3846), .Z1_t (new_AGEMA_signal_3847), .Z1_f (new_AGEMA_signal_3848) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_AddConstants_instance_U7 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (roundconstant[0]), .A1_f (new_AGEMA_signal_1888), .B0_t (LED_128_Instance_addroundkey_out[20]), .B0_f (new_AGEMA_signal_3696), .B1_t (new_AGEMA_signal_3697), .B1_f (new_AGEMA_signal_3698), .Z0_t (LED_128_Instance_addconst_out[20]), .Z0_f (new_AGEMA_signal_3849), .Z1_t (new_AGEMA_signal_3850), .Z1_f (new_AGEMA_signal_3851) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_AddConstants_instance_U6 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (roundconstant[1]), .A1_f (new_AGEMA_signal_1878), .B0_t (LED_128_Instance_addroundkey_out[53]), .B0_f (new_AGEMA_signal_3795), .B1_t (new_AGEMA_signal_3796), .B1_f (new_AGEMA_signal_3797), .Z0_t (LED_128_Instance_addconst_out[53]), .Z0_f (new_AGEMA_signal_3852), .Z1_t (new_AGEMA_signal_3853), .Z1_f (new_AGEMA_signal_3854) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_AddConstants_instance_U5 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (roundconstant[1]), .A1_f (new_AGEMA_signal_1878), .B0_t (LED_128_Instance_addroundkey_out[21]), .B0_f (new_AGEMA_signal_3699), .B1_t (new_AGEMA_signal_3700), .B1_f (new_AGEMA_signal_3701), .Z0_t (LED_128_Instance_addconst_out[21]), .Z0_f (new_AGEMA_signal_3855), .Z1_t (new_AGEMA_signal_3856), .Z1_f (new_AGEMA_signal_3857) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_AddConstants_instance_U4 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (roundconstant[4]), .A1_f (new_AGEMA_signal_1882), .B0_t (LED_128_Instance_addroundkey_out[37]), .B0_f (new_AGEMA_signal_3747), .B1_t (new_AGEMA_signal_3748), .B1_f (new_AGEMA_signal_3749), .Z0_t (LED_128_Instance_addconst_out[37]), .Z0_f (new_AGEMA_signal_3858), .Z1_t (new_AGEMA_signal_3859), .Z1_f (new_AGEMA_signal_3860) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_AddConstants_instance_U3 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (roundconstant[4]), .A1_f (new_AGEMA_signal_1882), .B0_t (LED_128_Instance_addroundkey_out[5]), .B0_f (new_AGEMA_signal_3651), .B1_t (new_AGEMA_signal_3652), .B1_f (new_AGEMA_signal_3653), .Z0_t (LED_128_Instance_addconst_out[5]), .Z0_f (new_AGEMA_signal_3861), .Z1_t (new_AGEMA_signal_3862), .Z1_f (new_AGEMA_signal_3863) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_0_XOR1_U1 ( .A0_t (LED_128_Instance_addconst_out[2]), .A0_f (new_AGEMA_signal_3642), .A1_t (new_AGEMA_signal_3643), .A1_f (new_AGEMA_signal_3644), .B0_t (LED_128_Instance_addconst_out[1]), .B0_f (new_AGEMA_signal_3639), .B1_t (new_AGEMA_signal_3640), .B1_f (new_AGEMA_signal_3641), .Z0_t (LED_128_Instance_SBox_Instance_0_L0), .Z0_f (new_AGEMA_signal_3864), .Z1_t (new_AGEMA_signal_3865), .Z1_f (new_AGEMA_signal_3866) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_0_XOR2_U1 ( .A0_t (LED_128_Instance_addconst_out[1]), .A0_f (new_AGEMA_signal_3639), .A1_t (new_AGEMA_signal_3640), .A1_f (new_AGEMA_signal_3641), .B0_t (LED_128_Instance_addconst_out[0]), .B0_f (new_AGEMA_signal_3636), .B1_t (new_AGEMA_signal_3637), .B1_f (new_AGEMA_signal_3638), .Z0_t (LED_128_Instance_SBox_Instance_0_L1), .Z0_f (new_AGEMA_signal_3867), .Z1_t (new_AGEMA_signal_3868), .Z1_f (new_AGEMA_signal_3869) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_0_XOR3_U1 ( .A0_t (LED_128_Instance_SBox_Instance_0_L1), .A0_f (new_AGEMA_signal_3867), .A1_t (new_AGEMA_signal_3868), .A1_f (new_AGEMA_signal_3869), .B0_t (LED_128_Instance_addroundkey_out[3]), .B0_f (new_AGEMA_signal_3645), .B1_t (new_AGEMA_signal_3646), .B1_f (new_AGEMA_signal_3647), .Z0_t (LED_128_Instance_SBox_Instance_0_L2), .Z0_f (new_AGEMA_signal_4044), .Z1_t (new_AGEMA_signal_4045), .Z1_f (new_AGEMA_signal_4046) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_SBox_Instance_0_XOR16_U1 ( .A0_t (LED_128_Instance_SBox_Instance_0_T0), .A0_f (new_AGEMA_signal_4053), .A1_t (new_AGEMA_signal_4054), .A1_f (new_AGEMA_signal_4055), .B0_t (LED_128_Instance_SBox_Instance_0_L2), .B0_f (new_AGEMA_signal_4044), .B1_t (new_AGEMA_signal_4045), .B1_f (new_AGEMA_signal_4046), .Z0_t (LED_128_Instance_SBox_Instance_0_Q2), .Z0_f (new_AGEMA_signal_4284), .Z1_t (new_AGEMA_signal_4285), .Z1_f (new_AGEMA_signal_4286) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_0_XOR4_U1 ( .A0_t (LED_128_Instance_addroundkey_out[3]), .A0_f (new_AGEMA_signal_3645), .A1_t (new_AGEMA_signal_3646), .A1_f (new_AGEMA_signal_3647), .B0_t (LED_128_Instance_addconst_out[0]), .B0_f (new_AGEMA_signal_3636), .B1_t (new_AGEMA_signal_3637), .B1_f (new_AGEMA_signal_3638), .Z0_t (LED_128_Instance_SBox_Instance_0_L3), .Z0_f (new_AGEMA_signal_3870), .Z1_t (new_AGEMA_signal_3871), .Z1_f (new_AGEMA_signal_3872) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_0_XOR5_U1 ( .A0_t (LED_128_Instance_SBox_Instance_0_L3), .A0_f (new_AGEMA_signal_3870), .A1_t (new_AGEMA_signal_3871), .A1_f (new_AGEMA_signal_3872), .B0_t (LED_128_Instance_SBox_Instance_0_L0), .B0_f (new_AGEMA_signal_3864), .B1_t (new_AGEMA_signal_3865), .B1_f (new_AGEMA_signal_3866), .Z0_t (LED_128_Instance_SBox_Instance_0_Q3), .Z0_f (new_AGEMA_signal_4047), .Z1_t (new_AGEMA_signal_4048), .Z1_f (new_AGEMA_signal_4049) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_0_XOR6_U1 ( .A0_t (LED_128_Instance_addroundkey_out[3]), .A0_f (new_AGEMA_signal_3645), .A1_t (new_AGEMA_signal_3646), .A1_f (new_AGEMA_signal_3647), .B0_t (LED_128_Instance_addconst_out[1]), .B0_f (new_AGEMA_signal_3639), .B1_t (new_AGEMA_signal_3640), .B1_f (new_AGEMA_signal_3641), .Z0_t (LED_128_Instance_SBox_Instance_0_L4), .Z0_f (new_AGEMA_signal_3873), .Z1_t (new_AGEMA_signal_3874), .Z1_f (new_AGEMA_signal_3875) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_0_XOR7_U1 ( .A0_t (LED_128_Instance_SBox_Instance_0_T0), .A0_f (new_AGEMA_signal_4053), .A1_t (new_AGEMA_signal_4054), .A1_f (new_AGEMA_signal_4055), .B0_t (LED_128_Instance_SBox_Instance_0_T2), .B0_f (new_AGEMA_signal_3876), .B1_t (new_AGEMA_signal_3877), .B1_f (new_AGEMA_signal_3878), .Z0_t (LED_128_Instance_SBox_Instance_0_L5), .Z0_f (new_AGEMA_signal_4287), .Z1_t (new_AGEMA_signal_4288), .Z1_f (new_AGEMA_signal_4289) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_SBox_Instance_0_XOR8_U1 ( .A0_t (LED_128_Instance_SBox_Instance_0_L4), .A0_f (new_AGEMA_signal_3873), .A1_t (new_AGEMA_signal_3874), .A1_f (new_AGEMA_signal_3875), .B0_t (LED_128_Instance_SBox_Instance_0_L5), .B0_f (new_AGEMA_signal_4287), .B1_t (new_AGEMA_signal_4288), .B1_f (new_AGEMA_signal_4289), .Z0_t (LED_128_Instance_SBox_Instance_0_Q6), .Z0_f (new_AGEMA_signal_4422), .Z1_t (new_AGEMA_signal_4423), .Z1_f (new_AGEMA_signal_4424) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_0_XOR9_U1 ( .A0_t (LED_128_Instance_SBox_Instance_0_L1), .A0_f (new_AGEMA_signal_3867), .A1_t (new_AGEMA_signal_3868), .A1_f (new_AGEMA_signal_3869), .B0_t (LED_128_Instance_addconst_out[2]), .B0_f (new_AGEMA_signal_3642), .B1_t (new_AGEMA_signal_3643), .B1_f (new_AGEMA_signal_3644), .Z0_t (LED_128_Instance_SBox_Instance_0_Q7), .Z0_f (new_AGEMA_signal_4050), .Z1_t (new_AGEMA_signal_4051), .Z1_f (new_AGEMA_signal_4052) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_0_AND1_U1 ( .A0_t (LED_128_Instance_SBox_Instance_0_L0), .A0_f (new_AGEMA_signal_3864), .A1_t (new_AGEMA_signal_3865), .A1_f (new_AGEMA_signal_3866), .B0_t (LED_128_Instance_addroundkey_out[3]), .B0_f (new_AGEMA_signal_3645), .B1_t (new_AGEMA_signal_3646), .B1_f (new_AGEMA_signal_3647), .Z0_t (LED_128_Instance_SBox_Instance_0_T0), .Z0_f (new_AGEMA_signal_4053), .Z1_t (new_AGEMA_signal_4054), .Z1_f (new_AGEMA_signal_4055) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_0_AND2_U1 ( .A0_t (LED_128_Instance_SBox_Instance_0_Q2), .A0_f (new_AGEMA_signal_4284), .A1_t (new_AGEMA_signal_4285), .A1_f (new_AGEMA_signal_4286), .B0_t (LED_128_Instance_SBox_Instance_0_Q3), .B0_f (new_AGEMA_signal_4047), .B1_t (new_AGEMA_signal_4048), .B1_f (new_AGEMA_signal_4049), .Z0_t (LED_128_Instance_SBox_Instance_0_T1), .Z0_f (new_AGEMA_signal_4425), .Z1_t (new_AGEMA_signal_4426), .Z1_f (new_AGEMA_signal_4427) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_0_AND3_U1 ( .A0_t (LED_128_Instance_addconst_out[1]), .A0_f (new_AGEMA_signal_3639), .A1_t (new_AGEMA_signal_3640), .A1_f (new_AGEMA_signal_3641), .B0_t (LED_128_Instance_addconst_out[2]), .B0_f (new_AGEMA_signal_3642), .B1_t (new_AGEMA_signal_3643), .B1_f (new_AGEMA_signal_3644), .Z0_t (LED_128_Instance_SBox_Instance_0_T2), .Z0_f (new_AGEMA_signal_3876), .Z1_t (new_AGEMA_signal_3877), .Z1_f (new_AGEMA_signal_3878) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_0_AND4_U1 ( .A0_t (LED_128_Instance_SBox_Instance_0_Q6), .A0_f (new_AGEMA_signal_4422), .A1_t (new_AGEMA_signal_4423), .A1_f (new_AGEMA_signal_4424), .B0_t (LED_128_Instance_SBox_Instance_0_Q7), .B0_f (new_AGEMA_signal_4050), .B1_t (new_AGEMA_signal_4051), .B1_f (new_AGEMA_signal_4052), .Z0_t (LED_128_Instance_SBox_Instance_0_T3), .Z0_f (new_AGEMA_signal_4524), .Z1_t (new_AGEMA_signal_4525), .Z1_f (new_AGEMA_signal_4526) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_0_XOR10_U1 ( .A0_t (LED_128_Instance_SBox_Instance_0_L5), .A0_f (new_AGEMA_signal_4287), .A1_t (new_AGEMA_signal_4288), .A1_f (new_AGEMA_signal_4289), .B0_t (LED_128_Instance_SBox_Instance_0_T3), .B0_f (new_AGEMA_signal_4524), .B1_t (new_AGEMA_signal_4525), .B1_f (new_AGEMA_signal_4526), .Z0_t (LED_128_Instance_SBox_Instance_0_L7), .Z0_f (new_AGEMA_signal_4620), .Z1_t (new_AGEMA_signal_4621), .Z1_f (new_AGEMA_signal_4622) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_0_XOR11_U1 ( .A0_t (LED_128_Instance_addconst_out[0]), .A0_f (new_AGEMA_signal_3636), .A1_t (new_AGEMA_signal_3637), .A1_f (new_AGEMA_signal_3638), .B0_t (LED_128_Instance_SBox_Instance_0_L7), .B0_f (new_AGEMA_signal_4620), .B1_t (new_AGEMA_signal_4621), .B1_f (new_AGEMA_signal_4622), .Z0_t (LED_128_Instance_subcells_out[3]), .Z0_f (new_AGEMA_signal_4752), .Z1_t (new_AGEMA_signal_4753), .Z1_f (new_AGEMA_signal_4754) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_0_XOR12_U1 ( .A0_t (LED_128_Instance_SBox_Instance_0_L5), .A0_f (new_AGEMA_signal_4287), .A1_t (new_AGEMA_signal_4288), .A1_f (new_AGEMA_signal_4289), .B0_t (LED_128_Instance_SBox_Instance_0_T1), .B0_f (new_AGEMA_signal_4425), .B1_t (new_AGEMA_signal_4426), .B1_f (new_AGEMA_signal_4427), .Z0_t (LED_128_Instance_SBox_Instance_0_L8), .Z0_f (new_AGEMA_signal_4527), .Z1_t (new_AGEMA_signal_4528), .Z1_f (new_AGEMA_signal_4529) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_0_XOR13_U1 ( .A0_t (LED_128_Instance_SBox_Instance_0_L1), .A0_f (new_AGEMA_signal_3867), .A1_t (new_AGEMA_signal_3868), .A1_f (new_AGEMA_signal_3869), .B0_t (LED_128_Instance_SBox_Instance_0_L8), .B0_f (new_AGEMA_signal_4527), .B1_t (new_AGEMA_signal_4528), .B1_f (new_AGEMA_signal_4529), .Z0_t (LED_128_Instance_subcells_out[2]), .Z0_f (new_AGEMA_signal_4623), .Z1_t (new_AGEMA_signal_4624), .Z1_f (new_AGEMA_signal_4625) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_0_XOR14_U1 ( .A0_t (LED_128_Instance_SBox_Instance_0_L4), .A0_f (new_AGEMA_signal_3873), .A1_t (new_AGEMA_signal_3874), .A1_f (new_AGEMA_signal_3875), .B0_t (LED_128_Instance_SBox_Instance_0_T3), .B0_f (new_AGEMA_signal_4524), .B1_t (new_AGEMA_signal_4525), .B1_f (new_AGEMA_signal_4526), .Z0_t (LED_128_Instance_subcells_out[1]), .Z0_f (new_AGEMA_signal_4626), .Z1_t (new_AGEMA_signal_4627), .Z1_f (new_AGEMA_signal_4628) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_0_XOR15_U1 ( .A0_t (LED_128_Instance_SBox_Instance_0_L3), .A0_f (new_AGEMA_signal_3870), .A1_t (new_AGEMA_signal_3871), .A1_f (new_AGEMA_signal_3872), .B0_t (LED_128_Instance_SBox_Instance_0_T2), .B0_f (new_AGEMA_signal_3876), .B1_t (new_AGEMA_signal_3877), .B1_f (new_AGEMA_signal_3878), .Z0_t (LED_128_Instance_subcells_out[0]), .Z0_f (new_AGEMA_signal_4056), .Z1_t (new_AGEMA_signal_4057), .Z1_f (new_AGEMA_signal_4058) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_1_XOR1_U1 ( .A0_t (LED_128_Instance_addconst_out[6]), .A0_f (new_AGEMA_signal_3834), .A1_t (new_AGEMA_signal_3835), .A1_f (new_AGEMA_signal_3836), .B0_t (LED_128_Instance_addconst_out[5]), .B0_f (new_AGEMA_signal_3861), .B1_t (new_AGEMA_signal_3862), .B1_f (new_AGEMA_signal_3863), .Z0_t (LED_128_Instance_SBox_Instance_1_L0), .Z0_f (new_AGEMA_signal_4059), .Z1_t (new_AGEMA_signal_4060), .Z1_f (new_AGEMA_signal_4061) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_1_XOR2_U1 ( .A0_t (LED_128_Instance_addconst_out[5]), .A0_f (new_AGEMA_signal_3861), .A1_t (new_AGEMA_signal_3862), .A1_f (new_AGEMA_signal_3863), .B0_t (LED_128_Instance_addconst_out[4]), .B0_f (new_AGEMA_signal_3843), .B1_t (new_AGEMA_signal_3844), .B1_f (new_AGEMA_signal_3845), .Z0_t (LED_128_Instance_SBox_Instance_1_L1), .Z0_f (new_AGEMA_signal_4062), .Z1_t (new_AGEMA_signal_4063), .Z1_f (new_AGEMA_signal_4064) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_1_XOR3_U1 ( .A0_t (LED_128_Instance_SBox_Instance_1_L1), .A0_f (new_AGEMA_signal_4062), .A1_t (new_AGEMA_signal_4063), .A1_f (new_AGEMA_signal_4064), .B0_t (LED_128_Instance_addconst_out[7]), .B0_f (new_AGEMA_signal_3657), .B1_t (new_AGEMA_signal_3658), .B1_f (new_AGEMA_signal_3659), .Z0_t (LED_128_Instance_SBox_Instance_1_L2), .Z0_f (new_AGEMA_signal_4290), .Z1_t (new_AGEMA_signal_4291), .Z1_f (new_AGEMA_signal_4292) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_SBox_Instance_1_XOR16_U1 ( .A0_t (LED_128_Instance_SBox_Instance_1_T0), .A0_f (new_AGEMA_signal_4299), .A1_t (new_AGEMA_signal_4300), .A1_f (new_AGEMA_signal_4301), .B0_t (LED_128_Instance_SBox_Instance_1_L2), .B0_f (new_AGEMA_signal_4290), .B1_t (new_AGEMA_signal_4291), .B1_f (new_AGEMA_signal_4292), .Z0_t (LED_128_Instance_SBox_Instance_1_Q2), .Z0_f (new_AGEMA_signal_4428), .Z1_t (new_AGEMA_signal_4429), .Z1_f (new_AGEMA_signal_4430) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_1_XOR4_U1 ( .A0_t (LED_128_Instance_addconst_out[7]), .A0_f (new_AGEMA_signal_3657), .A1_t (new_AGEMA_signal_3658), .A1_f (new_AGEMA_signal_3659), .B0_t (LED_128_Instance_addconst_out[4]), .B0_f (new_AGEMA_signal_3843), .B1_t (new_AGEMA_signal_3844), .B1_f (new_AGEMA_signal_3845), .Z0_t (LED_128_Instance_SBox_Instance_1_L3), .Z0_f (new_AGEMA_signal_4065), .Z1_t (new_AGEMA_signal_4066), .Z1_f (new_AGEMA_signal_4067) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_1_XOR5_U1 ( .A0_t (LED_128_Instance_SBox_Instance_1_L3), .A0_f (new_AGEMA_signal_4065), .A1_t (new_AGEMA_signal_4066), .A1_f (new_AGEMA_signal_4067), .B0_t (LED_128_Instance_SBox_Instance_1_L0), .B0_f (new_AGEMA_signal_4059), .B1_t (new_AGEMA_signal_4060), .B1_f (new_AGEMA_signal_4061), .Z0_t (LED_128_Instance_SBox_Instance_1_Q3), .Z0_f (new_AGEMA_signal_4293), .Z1_t (new_AGEMA_signal_4294), .Z1_f (new_AGEMA_signal_4295) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_1_XOR6_U1 ( .A0_t (LED_128_Instance_addconst_out[7]), .A0_f (new_AGEMA_signal_3657), .A1_t (new_AGEMA_signal_3658), .A1_f (new_AGEMA_signal_3659), .B0_t (LED_128_Instance_addconst_out[5]), .B0_f (new_AGEMA_signal_3861), .B1_t (new_AGEMA_signal_3862), .B1_f (new_AGEMA_signal_3863), .Z0_t (LED_128_Instance_SBox_Instance_1_L4), .Z0_f (new_AGEMA_signal_4068), .Z1_t (new_AGEMA_signal_4069), .Z1_f (new_AGEMA_signal_4070) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_1_XOR7_U1 ( .A0_t (LED_128_Instance_SBox_Instance_1_T0), .A0_f (new_AGEMA_signal_4299), .A1_t (new_AGEMA_signal_4300), .A1_f (new_AGEMA_signal_4301), .B0_t (LED_128_Instance_SBox_Instance_1_T2), .B0_f (new_AGEMA_signal_4071), .B1_t (new_AGEMA_signal_4072), .B1_f (new_AGEMA_signal_4073), .Z0_t (LED_128_Instance_SBox_Instance_1_L5), .Z0_f (new_AGEMA_signal_4431), .Z1_t (new_AGEMA_signal_4432), .Z1_f (new_AGEMA_signal_4433) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_SBox_Instance_1_XOR8_U1 ( .A0_t (LED_128_Instance_SBox_Instance_1_L4), .A0_f (new_AGEMA_signal_4068), .A1_t (new_AGEMA_signal_4069), .A1_f (new_AGEMA_signal_4070), .B0_t (LED_128_Instance_SBox_Instance_1_L5), .B0_f (new_AGEMA_signal_4431), .B1_t (new_AGEMA_signal_4432), .B1_f (new_AGEMA_signal_4433), .Z0_t (LED_128_Instance_SBox_Instance_1_Q6), .Z0_f (new_AGEMA_signal_4530), .Z1_t (new_AGEMA_signal_4531), .Z1_f (new_AGEMA_signal_4532) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_1_XOR9_U1 ( .A0_t (LED_128_Instance_SBox_Instance_1_L1), .A0_f (new_AGEMA_signal_4062), .A1_t (new_AGEMA_signal_4063), .A1_f (new_AGEMA_signal_4064), .B0_t (LED_128_Instance_addconst_out[6]), .B0_f (new_AGEMA_signal_3834), .B1_t (new_AGEMA_signal_3835), .B1_f (new_AGEMA_signal_3836), .Z0_t (LED_128_Instance_SBox_Instance_1_Q7), .Z0_f (new_AGEMA_signal_4296), .Z1_t (new_AGEMA_signal_4297), .Z1_f (new_AGEMA_signal_4298) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_1_AND1_U1 ( .A0_t (LED_128_Instance_SBox_Instance_1_L0), .A0_f (new_AGEMA_signal_4059), .A1_t (new_AGEMA_signal_4060), .A1_f (new_AGEMA_signal_4061), .B0_t (LED_128_Instance_addconst_out[7]), .B0_f (new_AGEMA_signal_3657), .B1_t (new_AGEMA_signal_3658), .B1_f (new_AGEMA_signal_3659), .Z0_t (LED_128_Instance_SBox_Instance_1_T0), .Z0_f (new_AGEMA_signal_4299), .Z1_t (new_AGEMA_signal_4300), .Z1_f (new_AGEMA_signal_4301) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_1_AND2_U1 ( .A0_t (LED_128_Instance_SBox_Instance_1_Q2), .A0_f (new_AGEMA_signal_4428), .A1_t (new_AGEMA_signal_4429), .A1_f (new_AGEMA_signal_4430), .B0_t (LED_128_Instance_SBox_Instance_1_Q3), .B0_f (new_AGEMA_signal_4293), .B1_t (new_AGEMA_signal_4294), .B1_f (new_AGEMA_signal_4295), .Z0_t (LED_128_Instance_SBox_Instance_1_T1), .Z0_f (new_AGEMA_signal_4533), .Z1_t (new_AGEMA_signal_4534), .Z1_f (new_AGEMA_signal_4535) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_1_AND3_U1 ( .A0_t (LED_128_Instance_addconst_out[5]), .A0_f (new_AGEMA_signal_3861), .A1_t (new_AGEMA_signal_3862), .A1_f (new_AGEMA_signal_3863), .B0_t (LED_128_Instance_addconst_out[6]), .B0_f (new_AGEMA_signal_3834), .B1_t (new_AGEMA_signal_3835), .B1_f (new_AGEMA_signal_3836), .Z0_t (LED_128_Instance_SBox_Instance_1_T2), .Z0_f (new_AGEMA_signal_4071), .Z1_t (new_AGEMA_signal_4072), .Z1_f (new_AGEMA_signal_4073) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_1_AND4_U1 ( .A0_t (LED_128_Instance_SBox_Instance_1_Q6), .A0_f (new_AGEMA_signal_4530), .A1_t (new_AGEMA_signal_4531), .A1_f (new_AGEMA_signal_4532), .B0_t (LED_128_Instance_SBox_Instance_1_Q7), .B0_f (new_AGEMA_signal_4296), .B1_t (new_AGEMA_signal_4297), .B1_f (new_AGEMA_signal_4298), .Z0_t (LED_128_Instance_SBox_Instance_1_T3), .Z0_f (new_AGEMA_signal_4629), .Z1_t (new_AGEMA_signal_4630), .Z1_f (new_AGEMA_signal_4631) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_1_XOR10_U1 ( .A0_t (LED_128_Instance_SBox_Instance_1_L5), .A0_f (new_AGEMA_signal_4431), .A1_t (new_AGEMA_signal_4432), .A1_f (new_AGEMA_signal_4433), .B0_t (LED_128_Instance_SBox_Instance_1_T3), .B0_f (new_AGEMA_signal_4629), .B1_t (new_AGEMA_signal_4630), .B1_f (new_AGEMA_signal_4631), .Z0_t (LED_128_Instance_SBox_Instance_1_L7), .Z0_f (new_AGEMA_signal_4755), .Z1_t (new_AGEMA_signal_4756), .Z1_f (new_AGEMA_signal_4757) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_1_XOR11_U1 ( .A0_t (LED_128_Instance_addconst_out[4]), .A0_f (new_AGEMA_signal_3843), .A1_t (new_AGEMA_signal_3844), .A1_f (new_AGEMA_signal_3845), .B0_t (LED_128_Instance_SBox_Instance_1_L7), .B0_f (new_AGEMA_signal_4755), .B1_t (new_AGEMA_signal_4756), .B1_f (new_AGEMA_signal_4757), .Z0_t (LED_128_Instance_subcells_out[7]), .Z0_f (new_AGEMA_signal_4887), .Z1_t (new_AGEMA_signal_4888), .Z1_f (new_AGEMA_signal_4889) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_1_XOR12_U1 ( .A0_t (LED_128_Instance_SBox_Instance_1_L5), .A0_f (new_AGEMA_signal_4431), .A1_t (new_AGEMA_signal_4432), .A1_f (new_AGEMA_signal_4433), .B0_t (LED_128_Instance_SBox_Instance_1_T1), .B0_f (new_AGEMA_signal_4533), .B1_t (new_AGEMA_signal_4534), .B1_f (new_AGEMA_signal_4535), .Z0_t (LED_128_Instance_SBox_Instance_1_L8), .Z0_f (new_AGEMA_signal_4632), .Z1_t (new_AGEMA_signal_4633), .Z1_f (new_AGEMA_signal_4634) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_1_XOR13_U1 ( .A0_t (LED_128_Instance_SBox_Instance_1_L1), .A0_f (new_AGEMA_signal_4062), .A1_t (new_AGEMA_signal_4063), .A1_f (new_AGEMA_signal_4064), .B0_t (LED_128_Instance_SBox_Instance_1_L8), .B0_f (new_AGEMA_signal_4632), .B1_t (new_AGEMA_signal_4633), .B1_f (new_AGEMA_signal_4634), .Z0_t (LED_128_Instance_subcells_out[6]), .Z0_f (new_AGEMA_signal_4758), .Z1_t (new_AGEMA_signal_4759), .Z1_f (new_AGEMA_signal_4760) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_1_XOR14_U1 ( .A0_t (LED_128_Instance_SBox_Instance_1_L4), .A0_f (new_AGEMA_signal_4068), .A1_t (new_AGEMA_signal_4069), .A1_f (new_AGEMA_signal_4070), .B0_t (LED_128_Instance_SBox_Instance_1_T3), .B0_f (new_AGEMA_signal_4629), .B1_t (new_AGEMA_signal_4630), .B1_f (new_AGEMA_signal_4631), .Z0_t (LED_128_Instance_subcells_out[5]), .Z0_f (new_AGEMA_signal_4761), .Z1_t (new_AGEMA_signal_4762), .Z1_f (new_AGEMA_signal_4763) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_1_XOR15_U1 ( .A0_t (LED_128_Instance_SBox_Instance_1_L3), .A0_f (new_AGEMA_signal_4065), .A1_t (new_AGEMA_signal_4066), .A1_f (new_AGEMA_signal_4067), .B0_t (LED_128_Instance_SBox_Instance_1_T2), .B0_f (new_AGEMA_signal_4071), .B1_t (new_AGEMA_signal_4072), .B1_f (new_AGEMA_signal_4073), .Z0_t (LED_128_Instance_subcells_out[4]), .Z0_f (new_AGEMA_signal_4302), .Z1_t (new_AGEMA_signal_4303), .Z1_f (new_AGEMA_signal_4304) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_2_XOR1_U1 ( .A0_t (LED_128_Instance_addconst_out[10]), .A0_f (new_AGEMA_signal_3666), .A1_t (new_AGEMA_signal_3667), .A1_f (new_AGEMA_signal_3668), .B0_t (LED_128_Instance_addconst_out[9]), .B0_f (new_AGEMA_signal_3663), .B1_t (new_AGEMA_signal_3664), .B1_f (new_AGEMA_signal_3665), .Z0_t (LED_128_Instance_SBox_Instance_2_L0), .Z0_f (new_AGEMA_signal_3879), .Z1_t (new_AGEMA_signal_3880), .Z1_f (new_AGEMA_signal_3881) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_2_XOR2_U1 ( .A0_t (LED_128_Instance_addconst_out[9]), .A0_f (new_AGEMA_signal_3663), .A1_t (new_AGEMA_signal_3664), .A1_f (new_AGEMA_signal_3665), .B0_t (LED_128_Instance_addconst_out[8]), .B0_f (new_AGEMA_signal_3660), .B1_t (new_AGEMA_signal_3661), .B1_f (new_AGEMA_signal_3662), .Z0_t (LED_128_Instance_SBox_Instance_2_L1), .Z0_f (new_AGEMA_signal_3882), .Z1_t (new_AGEMA_signal_3883), .Z1_f (new_AGEMA_signal_3884) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_2_XOR3_U1 ( .A0_t (LED_128_Instance_SBox_Instance_2_L1), .A0_f (new_AGEMA_signal_3882), .A1_t (new_AGEMA_signal_3883), .A1_f (new_AGEMA_signal_3884), .B0_t (LED_128_Instance_addconst_out[11]), .B0_f (new_AGEMA_signal_3669), .B1_t (new_AGEMA_signal_3670), .B1_f (new_AGEMA_signal_3671), .Z0_t (LED_128_Instance_SBox_Instance_2_L2), .Z0_f (new_AGEMA_signal_4074), .Z1_t (new_AGEMA_signal_4075), .Z1_f (new_AGEMA_signal_4076) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_SBox_Instance_2_XOR16_U1 ( .A0_t (LED_128_Instance_SBox_Instance_2_T0), .A0_f (new_AGEMA_signal_4083), .A1_t (new_AGEMA_signal_4084), .A1_f (new_AGEMA_signal_4085), .B0_t (LED_128_Instance_SBox_Instance_2_L2), .B0_f (new_AGEMA_signal_4074), .B1_t (new_AGEMA_signal_4075), .B1_f (new_AGEMA_signal_4076), .Z0_t (LED_128_Instance_SBox_Instance_2_Q2), .Z0_f (new_AGEMA_signal_4305), .Z1_t (new_AGEMA_signal_4306), .Z1_f (new_AGEMA_signal_4307) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_2_XOR4_U1 ( .A0_t (LED_128_Instance_addconst_out[11]), .A0_f (new_AGEMA_signal_3669), .A1_t (new_AGEMA_signal_3670), .A1_f (new_AGEMA_signal_3671), .B0_t (LED_128_Instance_addconst_out[8]), .B0_f (new_AGEMA_signal_3660), .B1_t (new_AGEMA_signal_3661), .B1_f (new_AGEMA_signal_3662), .Z0_t (LED_128_Instance_SBox_Instance_2_L3), .Z0_f (new_AGEMA_signal_3885), .Z1_t (new_AGEMA_signal_3886), .Z1_f (new_AGEMA_signal_3887) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_2_XOR5_U1 ( .A0_t (LED_128_Instance_SBox_Instance_2_L3), .A0_f (new_AGEMA_signal_3885), .A1_t (new_AGEMA_signal_3886), .A1_f (new_AGEMA_signal_3887), .B0_t (LED_128_Instance_SBox_Instance_2_L0), .B0_f (new_AGEMA_signal_3879), .B1_t (new_AGEMA_signal_3880), .B1_f (new_AGEMA_signal_3881), .Z0_t (LED_128_Instance_SBox_Instance_2_Q3), .Z0_f (new_AGEMA_signal_4077), .Z1_t (new_AGEMA_signal_4078), .Z1_f (new_AGEMA_signal_4079) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_2_XOR6_U1 ( .A0_t (LED_128_Instance_addconst_out[11]), .A0_f (new_AGEMA_signal_3669), .A1_t (new_AGEMA_signal_3670), .A1_f (new_AGEMA_signal_3671), .B0_t (LED_128_Instance_addconst_out[9]), .B0_f (new_AGEMA_signal_3663), .B1_t (new_AGEMA_signal_3664), .B1_f (new_AGEMA_signal_3665), .Z0_t (LED_128_Instance_SBox_Instance_2_L4), .Z0_f (new_AGEMA_signal_3888), .Z1_t (new_AGEMA_signal_3889), .Z1_f (new_AGEMA_signal_3890) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_2_XOR7_U1 ( .A0_t (LED_128_Instance_SBox_Instance_2_T0), .A0_f (new_AGEMA_signal_4083), .A1_t (new_AGEMA_signal_4084), .A1_f (new_AGEMA_signal_4085), .B0_t (LED_128_Instance_SBox_Instance_2_T2), .B0_f (new_AGEMA_signal_3891), .B1_t (new_AGEMA_signal_3892), .B1_f (new_AGEMA_signal_3893), .Z0_t (LED_128_Instance_SBox_Instance_2_L5), .Z0_f (new_AGEMA_signal_4308), .Z1_t (new_AGEMA_signal_4309), .Z1_f (new_AGEMA_signal_4310) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_SBox_Instance_2_XOR8_U1 ( .A0_t (LED_128_Instance_SBox_Instance_2_L4), .A0_f (new_AGEMA_signal_3888), .A1_t (new_AGEMA_signal_3889), .A1_f (new_AGEMA_signal_3890), .B0_t (LED_128_Instance_SBox_Instance_2_L5), .B0_f (new_AGEMA_signal_4308), .B1_t (new_AGEMA_signal_4309), .B1_f (new_AGEMA_signal_4310), .Z0_t (LED_128_Instance_SBox_Instance_2_Q6), .Z0_f (new_AGEMA_signal_4434), .Z1_t (new_AGEMA_signal_4435), .Z1_f (new_AGEMA_signal_4436) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_2_XOR9_U1 ( .A0_t (LED_128_Instance_SBox_Instance_2_L1), .A0_f (new_AGEMA_signal_3882), .A1_t (new_AGEMA_signal_3883), .A1_f (new_AGEMA_signal_3884), .B0_t (LED_128_Instance_addconst_out[10]), .B0_f (new_AGEMA_signal_3666), .B1_t (new_AGEMA_signal_3667), .B1_f (new_AGEMA_signal_3668), .Z0_t (LED_128_Instance_SBox_Instance_2_Q7), .Z0_f (new_AGEMA_signal_4080), .Z1_t (new_AGEMA_signal_4081), .Z1_f (new_AGEMA_signal_4082) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_2_AND1_U1 ( .A0_t (LED_128_Instance_SBox_Instance_2_L0), .A0_f (new_AGEMA_signal_3879), .A1_t (new_AGEMA_signal_3880), .A1_f (new_AGEMA_signal_3881), .B0_t (LED_128_Instance_addconst_out[11]), .B0_f (new_AGEMA_signal_3669), .B1_t (new_AGEMA_signal_3670), .B1_f (new_AGEMA_signal_3671), .Z0_t (LED_128_Instance_SBox_Instance_2_T0), .Z0_f (new_AGEMA_signal_4083), .Z1_t (new_AGEMA_signal_4084), .Z1_f (new_AGEMA_signal_4085) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_2_AND2_U1 ( .A0_t (LED_128_Instance_SBox_Instance_2_Q2), .A0_f (new_AGEMA_signal_4305), .A1_t (new_AGEMA_signal_4306), .A1_f (new_AGEMA_signal_4307), .B0_t (LED_128_Instance_SBox_Instance_2_Q3), .B0_f (new_AGEMA_signal_4077), .B1_t (new_AGEMA_signal_4078), .B1_f (new_AGEMA_signal_4079), .Z0_t (LED_128_Instance_SBox_Instance_2_T1), .Z0_f (new_AGEMA_signal_4437), .Z1_t (new_AGEMA_signal_4438), .Z1_f (new_AGEMA_signal_4439) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_2_AND3_U1 ( .A0_t (LED_128_Instance_addconst_out[9]), .A0_f (new_AGEMA_signal_3663), .A1_t (new_AGEMA_signal_3664), .A1_f (new_AGEMA_signal_3665), .B0_t (LED_128_Instance_addconst_out[10]), .B0_f (new_AGEMA_signal_3666), .B1_t (new_AGEMA_signal_3667), .B1_f (new_AGEMA_signal_3668), .Z0_t (LED_128_Instance_SBox_Instance_2_T2), .Z0_f (new_AGEMA_signal_3891), .Z1_t (new_AGEMA_signal_3892), .Z1_f (new_AGEMA_signal_3893) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_2_AND4_U1 ( .A0_t (LED_128_Instance_SBox_Instance_2_Q6), .A0_f (new_AGEMA_signal_4434), .A1_t (new_AGEMA_signal_4435), .A1_f (new_AGEMA_signal_4436), .B0_t (LED_128_Instance_SBox_Instance_2_Q7), .B0_f (new_AGEMA_signal_4080), .B1_t (new_AGEMA_signal_4081), .B1_f (new_AGEMA_signal_4082), .Z0_t (LED_128_Instance_SBox_Instance_2_T3), .Z0_f (new_AGEMA_signal_4536), .Z1_t (new_AGEMA_signal_4537), .Z1_f (new_AGEMA_signal_4538) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_2_XOR10_U1 ( .A0_t (LED_128_Instance_SBox_Instance_2_L5), .A0_f (new_AGEMA_signal_4308), .A1_t (new_AGEMA_signal_4309), .A1_f (new_AGEMA_signal_4310), .B0_t (LED_128_Instance_SBox_Instance_2_T3), .B0_f (new_AGEMA_signal_4536), .B1_t (new_AGEMA_signal_4537), .B1_f (new_AGEMA_signal_4538), .Z0_t (LED_128_Instance_SBox_Instance_2_L7), .Z0_f (new_AGEMA_signal_4635), .Z1_t (new_AGEMA_signal_4636), .Z1_f (new_AGEMA_signal_4637) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_2_XOR11_U1 ( .A0_t (LED_128_Instance_addconst_out[8]), .A0_f (new_AGEMA_signal_3660), .A1_t (new_AGEMA_signal_3661), .A1_f (new_AGEMA_signal_3662), .B0_t (LED_128_Instance_SBox_Instance_2_L7), .B0_f (new_AGEMA_signal_4635), .B1_t (new_AGEMA_signal_4636), .B1_f (new_AGEMA_signal_4637), .Z0_t (LED_128_Instance_subcells_out[11]), .Z0_f (new_AGEMA_signal_4764), .Z1_t (new_AGEMA_signal_4765), .Z1_f (new_AGEMA_signal_4766) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_2_XOR12_U1 ( .A0_t (LED_128_Instance_SBox_Instance_2_L5), .A0_f (new_AGEMA_signal_4308), .A1_t (new_AGEMA_signal_4309), .A1_f (new_AGEMA_signal_4310), .B0_t (LED_128_Instance_SBox_Instance_2_T1), .B0_f (new_AGEMA_signal_4437), .B1_t (new_AGEMA_signal_4438), .B1_f (new_AGEMA_signal_4439), .Z0_t (LED_128_Instance_SBox_Instance_2_L8), .Z0_f (new_AGEMA_signal_4539), .Z1_t (new_AGEMA_signal_4540), .Z1_f (new_AGEMA_signal_4541) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_2_XOR13_U1 ( .A0_t (LED_128_Instance_SBox_Instance_2_L1), .A0_f (new_AGEMA_signal_3882), .A1_t (new_AGEMA_signal_3883), .A1_f (new_AGEMA_signal_3884), .B0_t (LED_128_Instance_SBox_Instance_2_L8), .B0_f (new_AGEMA_signal_4539), .B1_t (new_AGEMA_signal_4540), .B1_f (new_AGEMA_signal_4541), .Z0_t (LED_128_Instance_subcells_out[10]), .Z0_f (new_AGEMA_signal_4638), .Z1_t (new_AGEMA_signal_4639), .Z1_f (new_AGEMA_signal_4640) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_2_XOR14_U1 ( .A0_t (LED_128_Instance_SBox_Instance_2_L4), .A0_f (new_AGEMA_signal_3888), .A1_t (new_AGEMA_signal_3889), .A1_f (new_AGEMA_signal_3890), .B0_t (LED_128_Instance_SBox_Instance_2_T3), .B0_f (new_AGEMA_signal_4536), .B1_t (new_AGEMA_signal_4537), .B1_f (new_AGEMA_signal_4538), .Z0_t (LED_128_Instance_subcells_out[9]), .Z0_f (new_AGEMA_signal_4641), .Z1_t (new_AGEMA_signal_4642), .Z1_f (new_AGEMA_signal_4643) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_2_XOR15_U1 ( .A0_t (LED_128_Instance_SBox_Instance_2_L3), .A0_f (new_AGEMA_signal_3885), .A1_t (new_AGEMA_signal_3886), .A1_f (new_AGEMA_signal_3887), .B0_t (LED_128_Instance_SBox_Instance_2_T2), .B0_f (new_AGEMA_signal_3891), .B1_t (new_AGEMA_signal_3892), .B1_f (new_AGEMA_signal_3893), .Z0_t (LED_128_Instance_subcells_out[8]), .Z0_f (new_AGEMA_signal_4086), .Z1_t (new_AGEMA_signal_4087), .Z1_f (new_AGEMA_signal_4088) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_3_XOR1_U1 ( .A0_t (LED_128_Instance_addconst_out[14]), .A0_f (new_AGEMA_signal_3678), .A1_t (new_AGEMA_signal_3679), .A1_f (new_AGEMA_signal_3680), .B0_t (LED_128_Instance_addconst_out[13]), .B0_f (new_AGEMA_signal_3675), .B1_t (new_AGEMA_signal_3676), .B1_f (new_AGEMA_signal_3677), .Z0_t (LED_128_Instance_SBox_Instance_3_L0), .Z0_f (new_AGEMA_signal_3894), .Z1_t (new_AGEMA_signal_3895), .Z1_f (new_AGEMA_signal_3896) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_3_XOR2_U1 ( .A0_t (LED_128_Instance_addconst_out[13]), .A0_f (new_AGEMA_signal_3675), .A1_t (new_AGEMA_signal_3676), .A1_f (new_AGEMA_signal_3677), .B0_t (LED_128_Instance_addconst_out[12]), .B0_f (new_AGEMA_signal_3672), .B1_t (new_AGEMA_signal_3673), .B1_f (new_AGEMA_signal_3674), .Z0_t (LED_128_Instance_SBox_Instance_3_L1), .Z0_f (new_AGEMA_signal_3897), .Z1_t (new_AGEMA_signal_3898), .Z1_f (new_AGEMA_signal_3899) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_3_XOR3_U1 ( .A0_t (LED_128_Instance_SBox_Instance_3_L1), .A0_f (new_AGEMA_signal_3897), .A1_t (new_AGEMA_signal_3898), .A1_f (new_AGEMA_signal_3899), .B0_t (LED_128_Instance_addconst_out[15]), .B0_f (new_AGEMA_signal_3681), .B1_t (new_AGEMA_signal_3682), .B1_f (new_AGEMA_signal_3683), .Z0_t (LED_128_Instance_SBox_Instance_3_L2), .Z0_f (new_AGEMA_signal_4089), .Z1_t (new_AGEMA_signal_4090), .Z1_f (new_AGEMA_signal_4091) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_SBox_Instance_3_XOR16_U1 ( .A0_t (LED_128_Instance_SBox_Instance_3_T0), .A0_f (new_AGEMA_signal_4098), .A1_t (new_AGEMA_signal_4099), .A1_f (new_AGEMA_signal_4100), .B0_t (LED_128_Instance_SBox_Instance_3_L2), .B0_f (new_AGEMA_signal_4089), .B1_t (new_AGEMA_signal_4090), .B1_f (new_AGEMA_signal_4091), .Z0_t (LED_128_Instance_SBox_Instance_3_Q2), .Z0_f (new_AGEMA_signal_4311), .Z1_t (new_AGEMA_signal_4312), .Z1_f (new_AGEMA_signal_4313) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_3_XOR4_U1 ( .A0_t (LED_128_Instance_addconst_out[15]), .A0_f (new_AGEMA_signal_3681), .A1_t (new_AGEMA_signal_3682), .A1_f (new_AGEMA_signal_3683), .B0_t (LED_128_Instance_addconst_out[12]), .B0_f (new_AGEMA_signal_3672), .B1_t (new_AGEMA_signal_3673), .B1_f (new_AGEMA_signal_3674), .Z0_t (LED_128_Instance_SBox_Instance_3_L3), .Z0_f (new_AGEMA_signal_3900), .Z1_t (new_AGEMA_signal_3901), .Z1_f (new_AGEMA_signal_3902) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_3_XOR5_U1 ( .A0_t (LED_128_Instance_SBox_Instance_3_L3), .A0_f (new_AGEMA_signal_3900), .A1_t (new_AGEMA_signal_3901), .A1_f (new_AGEMA_signal_3902), .B0_t (LED_128_Instance_SBox_Instance_3_L0), .B0_f (new_AGEMA_signal_3894), .B1_t (new_AGEMA_signal_3895), .B1_f (new_AGEMA_signal_3896), .Z0_t (LED_128_Instance_SBox_Instance_3_Q3), .Z0_f (new_AGEMA_signal_4092), .Z1_t (new_AGEMA_signal_4093), .Z1_f (new_AGEMA_signal_4094) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_3_XOR6_U1 ( .A0_t (LED_128_Instance_addconst_out[15]), .A0_f (new_AGEMA_signal_3681), .A1_t (new_AGEMA_signal_3682), .A1_f (new_AGEMA_signal_3683), .B0_t (LED_128_Instance_addconst_out[13]), .B0_f (new_AGEMA_signal_3675), .B1_t (new_AGEMA_signal_3676), .B1_f (new_AGEMA_signal_3677), .Z0_t (LED_128_Instance_SBox_Instance_3_L4), .Z0_f (new_AGEMA_signal_3903), .Z1_t (new_AGEMA_signal_3904), .Z1_f (new_AGEMA_signal_3905) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_3_XOR7_U1 ( .A0_t (LED_128_Instance_SBox_Instance_3_T0), .A0_f (new_AGEMA_signal_4098), .A1_t (new_AGEMA_signal_4099), .A1_f (new_AGEMA_signal_4100), .B0_t (LED_128_Instance_SBox_Instance_3_T2), .B0_f (new_AGEMA_signal_3906), .B1_t (new_AGEMA_signal_3907), .B1_f (new_AGEMA_signal_3908), .Z0_t (LED_128_Instance_SBox_Instance_3_L5), .Z0_f (new_AGEMA_signal_4314), .Z1_t (new_AGEMA_signal_4315), .Z1_f (new_AGEMA_signal_4316) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_SBox_Instance_3_XOR8_U1 ( .A0_t (LED_128_Instance_SBox_Instance_3_L4), .A0_f (new_AGEMA_signal_3903), .A1_t (new_AGEMA_signal_3904), .A1_f (new_AGEMA_signal_3905), .B0_t (LED_128_Instance_SBox_Instance_3_L5), .B0_f (new_AGEMA_signal_4314), .B1_t (new_AGEMA_signal_4315), .B1_f (new_AGEMA_signal_4316), .Z0_t (LED_128_Instance_SBox_Instance_3_Q6), .Z0_f (new_AGEMA_signal_4440), .Z1_t (new_AGEMA_signal_4441), .Z1_f (new_AGEMA_signal_4442) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_3_XOR9_U1 ( .A0_t (LED_128_Instance_SBox_Instance_3_L1), .A0_f (new_AGEMA_signal_3897), .A1_t (new_AGEMA_signal_3898), .A1_f (new_AGEMA_signal_3899), .B0_t (LED_128_Instance_addconst_out[14]), .B0_f (new_AGEMA_signal_3678), .B1_t (new_AGEMA_signal_3679), .B1_f (new_AGEMA_signal_3680), .Z0_t (LED_128_Instance_SBox_Instance_3_Q7), .Z0_f (new_AGEMA_signal_4095), .Z1_t (new_AGEMA_signal_4096), .Z1_f (new_AGEMA_signal_4097) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_3_AND1_U1 ( .A0_t (LED_128_Instance_SBox_Instance_3_L0), .A0_f (new_AGEMA_signal_3894), .A1_t (new_AGEMA_signal_3895), .A1_f (new_AGEMA_signal_3896), .B0_t (LED_128_Instance_addconst_out[15]), .B0_f (new_AGEMA_signal_3681), .B1_t (new_AGEMA_signal_3682), .B1_f (new_AGEMA_signal_3683), .Z0_t (LED_128_Instance_SBox_Instance_3_T0), .Z0_f (new_AGEMA_signal_4098), .Z1_t (new_AGEMA_signal_4099), .Z1_f (new_AGEMA_signal_4100) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_3_AND2_U1 ( .A0_t (LED_128_Instance_SBox_Instance_3_Q2), .A0_f (new_AGEMA_signal_4311), .A1_t (new_AGEMA_signal_4312), .A1_f (new_AGEMA_signal_4313), .B0_t (LED_128_Instance_SBox_Instance_3_Q3), .B0_f (new_AGEMA_signal_4092), .B1_t (new_AGEMA_signal_4093), .B1_f (new_AGEMA_signal_4094), .Z0_t (LED_128_Instance_SBox_Instance_3_T1), .Z0_f (new_AGEMA_signal_4443), .Z1_t (new_AGEMA_signal_4444), .Z1_f (new_AGEMA_signal_4445) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_3_AND3_U1 ( .A0_t (LED_128_Instance_addconst_out[13]), .A0_f (new_AGEMA_signal_3675), .A1_t (new_AGEMA_signal_3676), .A1_f (new_AGEMA_signal_3677), .B0_t (LED_128_Instance_addconst_out[14]), .B0_f (new_AGEMA_signal_3678), .B1_t (new_AGEMA_signal_3679), .B1_f (new_AGEMA_signal_3680), .Z0_t (LED_128_Instance_SBox_Instance_3_T2), .Z0_f (new_AGEMA_signal_3906), .Z1_t (new_AGEMA_signal_3907), .Z1_f (new_AGEMA_signal_3908) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_3_AND4_U1 ( .A0_t (LED_128_Instance_SBox_Instance_3_Q6), .A0_f (new_AGEMA_signal_4440), .A1_t (new_AGEMA_signal_4441), .A1_f (new_AGEMA_signal_4442), .B0_t (LED_128_Instance_SBox_Instance_3_Q7), .B0_f (new_AGEMA_signal_4095), .B1_t (new_AGEMA_signal_4096), .B1_f (new_AGEMA_signal_4097), .Z0_t (LED_128_Instance_SBox_Instance_3_T3), .Z0_f (new_AGEMA_signal_4542), .Z1_t (new_AGEMA_signal_4543), .Z1_f (new_AGEMA_signal_4544) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_3_XOR10_U1 ( .A0_t (LED_128_Instance_SBox_Instance_3_L5), .A0_f (new_AGEMA_signal_4314), .A1_t (new_AGEMA_signal_4315), .A1_f (new_AGEMA_signal_4316), .B0_t (LED_128_Instance_SBox_Instance_3_T3), .B0_f (new_AGEMA_signal_4542), .B1_t (new_AGEMA_signal_4543), .B1_f (new_AGEMA_signal_4544), .Z0_t (LED_128_Instance_SBox_Instance_3_L7), .Z0_f (new_AGEMA_signal_4644), .Z1_t (new_AGEMA_signal_4645), .Z1_f (new_AGEMA_signal_4646) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_3_XOR11_U1 ( .A0_t (LED_128_Instance_addconst_out[12]), .A0_f (new_AGEMA_signal_3672), .A1_t (new_AGEMA_signal_3673), .A1_f (new_AGEMA_signal_3674), .B0_t (LED_128_Instance_SBox_Instance_3_L7), .B0_f (new_AGEMA_signal_4644), .B1_t (new_AGEMA_signal_4645), .B1_f (new_AGEMA_signal_4646), .Z0_t (LED_128_Instance_subcells_out[15]), .Z0_f (new_AGEMA_signal_4767), .Z1_t (new_AGEMA_signal_4768), .Z1_f (new_AGEMA_signal_4769) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_3_XOR12_U1 ( .A0_t (LED_128_Instance_SBox_Instance_3_L5), .A0_f (new_AGEMA_signal_4314), .A1_t (new_AGEMA_signal_4315), .A1_f (new_AGEMA_signal_4316), .B0_t (LED_128_Instance_SBox_Instance_3_T1), .B0_f (new_AGEMA_signal_4443), .B1_t (new_AGEMA_signal_4444), .B1_f (new_AGEMA_signal_4445), .Z0_t (LED_128_Instance_SBox_Instance_3_L8), .Z0_f (new_AGEMA_signal_4545), .Z1_t (new_AGEMA_signal_4546), .Z1_f (new_AGEMA_signal_4547) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_3_XOR13_U1 ( .A0_t (LED_128_Instance_SBox_Instance_3_L1), .A0_f (new_AGEMA_signal_3897), .A1_t (new_AGEMA_signal_3898), .A1_f (new_AGEMA_signal_3899), .B0_t (LED_128_Instance_SBox_Instance_3_L8), .B0_f (new_AGEMA_signal_4545), .B1_t (new_AGEMA_signal_4546), .B1_f (new_AGEMA_signal_4547), .Z0_t (LED_128_Instance_subcells_out[14]), .Z0_f (new_AGEMA_signal_4647), .Z1_t (new_AGEMA_signal_4648), .Z1_f (new_AGEMA_signal_4649) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_3_XOR14_U1 ( .A0_t (LED_128_Instance_SBox_Instance_3_L4), .A0_f (new_AGEMA_signal_3903), .A1_t (new_AGEMA_signal_3904), .A1_f (new_AGEMA_signal_3905), .B0_t (LED_128_Instance_SBox_Instance_3_T3), .B0_f (new_AGEMA_signal_4542), .B1_t (new_AGEMA_signal_4543), .B1_f (new_AGEMA_signal_4544), .Z0_t (LED_128_Instance_subcells_out[13]), .Z0_f (new_AGEMA_signal_4650), .Z1_t (new_AGEMA_signal_4651), .Z1_f (new_AGEMA_signal_4652) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_3_XOR15_U1 ( .A0_t (LED_128_Instance_SBox_Instance_3_L3), .A0_f (new_AGEMA_signal_3900), .A1_t (new_AGEMA_signal_3901), .A1_f (new_AGEMA_signal_3902), .B0_t (LED_128_Instance_SBox_Instance_3_T2), .B0_f (new_AGEMA_signal_3906), .B1_t (new_AGEMA_signal_3907), .B1_f (new_AGEMA_signal_3908), .Z0_t (LED_128_Instance_subcells_out[12]), .Z0_f (new_AGEMA_signal_4101), .Z1_t (new_AGEMA_signal_4102), .Z1_f (new_AGEMA_signal_4103) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_4_XOR1_U1 ( .A0_t (LED_128_Instance_addconst_out[18]), .A0_f (new_AGEMA_signal_3690), .A1_t (new_AGEMA_signal_3691), .A1_f (new_AGEMA_signal_3692), .B0_t (LED_128_Instance_addconst_out[17]), .B0_f (new_AGEMA_signal_3687), .B1_t (new_AGEMA_signal_3688), .B1_f (new_AGEMA_signal_3689), .Z0_t (LED_128_Instance_SBox_Instance_4_L0), .Z0_f (new_AGEMA_signal_3909), .Z1_t (new_AGEMA_signal_3910), .Z1_f (new_AGEMA_signal_3911) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_4_XOR2_U1 ( .A0_t (LED_128_Instance_addconst_out[17]), .A0_f (new_AGEMA_signal_3687), .A1_t (new_AGEMA_signal_3688), .A1_f (new_AGEMA_signal_3689), .B0_t (LED_128_Instance_addroundkey_out[16]), .B0_f (new_AGEMA_signal_3684), .B1_t (new_AGEMA_signal_3685), .B1_f (new_AGEMA_signal_3686), .Z0_t (LED_128_Instance_SBox_Instance_4_L1), .Z0_f (new_AGEMA_signal_3912), .Z1_t (new_AGEMA_signal_3913), .Z1_f (new_AGEMA_signal_3914) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_4_XOR3_U1 ( .A0_t (LED_128_Instance_SBox_Instance_4_L1), .A0_f (new_AGEMA_signal_3912), .A1_t (new_AGEMA_signal_3913), .A1_f (new_AGEMA_signal_3914), .B0_t (LED_128_Instance_addroundkey_out[19]), .B0_f (new_AGEMA_signal_3693), .B1_t (new_AGEMA_signal_3694), .B1_f (new_AGEMA_signal_3695), .Z0_t (LED_128_Instance_SBox_Instance_4_L2), .Z0_f (new_AGEMA_signal_4104), .Z1_t (new_AGEMA_signal_4105), .Z1_f (new_AGEMA_signal_4106) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_SBox_Instance_4_XOR16_U1 ( .A0_t (LED_128_Instance_SBox_Instance_4_T0), .A0_f (new_AGEMA_signal_4113), .A1_t (new_AGEMA_signal_4114), .A1_f (new_AGEMA_signal_4115), .B0_t (LED_128_Instance_SBox_Instance_4_L2), .B0_f (new_AGEMA_signal_4104), .B1_t (new_AGEMA_signal_4105), .B1_f (new_AGEMA_signal_4106), .Z0_t (LED_128_Instance_SBox_Instance_4_Q2), .Z0_f (new_AGEMA_signal_4317), .Z1_t (new_AGEMA_signal_4318), .Z1_f (new_AGEMA_signal_4319) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_4_XOR4_U1 ( .A0_t (LED_128_Instance_addroundkey_out[19]), .A0_f (new_AGEMA_signal_3693), .A1_t (new_AGEMA_signal_3694), .A1_f (new_AGEMA_signal_3695), .B0_t (LED_128_Instance_addroundkey_out[16]), .B0_f (new_AGEMA_signal_3684), .B1_t (new_AGEMA_signal_3685), .B1_f (new_AGEMA_signal_3686), .Z0_t (LED_128_Instance_SBox_Instance_4_L3), .Z0_f (new_AGEMA_signal_3915), .Z1_t (new_AGEMA_signal_3916), .Z1_f (new_AGEMA_signal_3917) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_4_XOR5_U1 ( .A0_t (LED_128_Instance_SBox_Instance_4_L3), .A0_f (new_AGEMA_signal_3915), .A1_t (new_AGEMA_signal_3916), .A1_f (new_AGEMA_signal_3917), .B0_t (LED_128_Instance_SBox_Instance_4_L0), .B0_f (new_AGEMA_signal_3909), .B1_t (new_AGEMA_signal_3910), .B1_f (new_AGEMA_signal_3911), .Z0_t (LED_128_Instance_SBox_Instance_4_Q3), .Z0_f (new_AGEMA_signal_4107), .Z1_t (new_AGEMA_signal_4108), .Z1_f (new_AGEMA_signal_4109) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_4_XOR6_U1 ( .A0_t (LED_128_Instance_addroundkey_out[19]), .A0_f (new_AGEMA_signal_3693), .A1_t (new_AGEMA_signal_3694), .A1_f (new_AGEMA_signal_3695), .B0_t (LED_128_Instance_addconst_out[17]), .B0_f (new_AGEMA_signal_3687), .B1_t (new_AGEMA_signal_3688), .B1_f (new_AGEMA_signal_3689), .Z0_t (LED_128_Instance_SBox_Instance_4_L4), .Z0_f (new_AGEMA_signal_3918), .Z1_t (new_AGEMA_signal_3919), .Z1_f (new_AGEMA_signal_3920) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_4_XOR7_U1 ( .A0_t (LED_128_Instance_SBox_Instance_4_T0), .A0_f (new_AGEMA_signal_4113), .A1_t (new_AGEMA_signal_4114), .A1_f (new_AGEMA_signal_4115), .B0_t (LED_128_Instance_SBox_Instance_4_T2), .B0_f (new_AGEMA_signal_3921), .B1_t (new_AGEMA_signal_3922), .B1_f (new_AGEMA_signal_3923), .Z0_t (LED_128_Instance_SBox_Instance_4_L5), .Z0_f (new_AGEMA_signal_4320), .Z1_t (new_AGEMA_signal_4321), .Z1_f (new_AGEMA_signal_4322) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_SBox_Instance_4_XOR8_U1 ( .A0_t (LED_128_Instance_SBox_Instance_4_L4), .A0_f (new_AGEMA_signal_3918), .A1_t (new_AGEMA_signal_3919), .A1_f (new_AGEMA_signal_3920), .B0_t (LED_128_Instance_SBox_Instance_4_L5), .B0_f (new_AGEMA_signal_4320), .B1_t (new_AGEMA_signal_4321), .B1_f (new_AGEMA_signal_4322), .Z0_t (LED_128_Instance_SBox_Instance_4_Q6), .Z0_f (new_AGEMA_signal_4446), .Z1_t (new_AGEMA_signal_4447), .Z1_f (new_AGEMA_signal_4448) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_4_XOR9_U1 ( .A0_t (LED_128_Instance_SBox_Instance_4_L1), .A0_f (new_AGEMA_signal_3912), .A1_t (new_AGEMA_signal_3913), .A1_f (new_AGEMA_signal_3914), .B0_t (LED_128_Instance_addconst_out[18]), .B0_f (new_AGEMA_signal_3690), .B1_t (new_AGEMA_signal_3691), .B1_f (new_AGEMA_signal_3692), .Z0_t (LED_128_Instance_SBox_Instance_4_Q7), .Z0_f (new_AGEMA_signal_4110), .Z1_t (new_AGEMA_signal_4111), .Z1_f (new_AGEMA_signal_4112) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_4_AND1_U1 ( .A0_t (LED_128_Instance_SBox_Instance_4_L0), .A0_f (new_AGEMA_signal_3909), .A1_t (new_AGEMA_signal_3910), .A1_f (new_AGEMA_signal_3911), .B0_t (LED_128_Instance_addroundkey_out[19]), .B0_f (new_AGEMA_signal_3693), .B1_t (new_AGEMA_signal_3694), .B1_f (new_AGEMA_signal_3695), .Z0_t (LED_128_Instance_SBox_Instance_4_T0), .Z0_f (new_AGEMA_signal_4113), .Z1_t (new_AGEMA_signal_4114), .Z1_f (new_AGEMA_signal_4115) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_4_AND2_U1 ( .A0_t (LED_128_Instance_SBox_Instance_4_Q2), .A0_f (new_AGEMA_signal_4317), .A1_t (new_AGEMA_signal_4318), .A1_f (new_AGEMA_signal_4319), .B0_t (LED_128_Instance_SBox_Instance_4_Q3), .B0_f (new_AGEMA_signal_4107), .B1_t (new_AGEMA_signal_4108), .B1_f (new_AGEMA_signal_4109), .Z0_t (LED_128_Instance_SBox_Instance_4_T1), .Z0_f (new_AGEMA_signal_4449), .Z1_t (new_AGEMA_signal_4450), .Z1_f (new_AGEMA_signal_4451) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_4_AND3_U1 ( .A0_t (LED_128_Instance_addconst_out[17]), .A0_f (new_AGEMA_signal_3687), .A1_t (new_AGEMA_signal_3688), .A1_f (new_AGEMA_signal_3689), .B0_t (LED_128_Instance_addconst_out[18]), .B0_f (new_AGEMA_signal_3690), .B1_t (new_AGEMA_signal_3691), .B1_f (new_AGEMA_signal_3692), .Z0_t (LED_128_Instance_SBox_Instance_4_T2), .Z0_f (new_AGEMA_signal_3921), .Z1_t (new_AGEMA_signal_3922), .Z1_f (new_AGEMA_signal_3923) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_4_AND4_U1 ( .A0_t (LED_128_Instance_SBox_Instance_4_Q6), .A0_f (new_AGEMA_signal_4446), .A1_t (new_AGEMA_signal_4447), .A1_f (new_AGEMA_signal_4448), .B0_t (LED_128_Instance_SBox_Instance_4_Q7), .B0_f (new_AGEMA_signal_4110), .B1_t (new_AGEMA_signal_4111), .B1_f (new_AGEMA_signal_4112), .Z0_t (LED_128_Instance_SBox_Instance_4_T3), .Z0_f (new_AGEMA_signal_4548), .Z1_t (new_AGEMA_signal_4549), .Z1_f (new_AGEMA_signal_4550) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_4_XOR10_U1 ( .A0_t (LED_128_Instance_SBox_Instance_4_L5), .A0_f (new_AGEMA_signal_4320), .A1_t (new_AGEMA_signal_4321), .A1_f (new_AGEMA_signal_4322), .B0_t (LED_128_Instance_SBox_Instance_4_T3), .B0_f (new_AGEMA_signal_4548), .B1_t (new_AGEMA_signal_4549), .B1_f (new_AGEMA_signal_4550), .Z0_t (LED_128_Instance_SBox_Instance_4_L7), .Z0_f (new_AGEMA_signal_4653), .Z1_t (new_AGEMA_signal_4654), .Z1_f (new_AGEMA_signal_4655) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_4_XOR11_U1 ( .A0_t (LED_128_Instance_addroundkey_out[16]), .A0_f (new_AGEMA_signal_3684), .A1_t (new_AGEMA_signal_3685), .A1_f (new_AGEMA_signal_3686), .B0_t (LED_128_Instance_SBox_Instance_4_L7), .B0_f (new_AGEMA_signal_4653), .B1_t (new_AGEMA_signal_4654), .B1_f (new_AGEMA_signal_4655), .Z0_t (LED_128_Instance_subcells_out[19]), .Z0_f (new_AGEMA_signal_4770), .Z1_t (new_AGEMA_signal_4771), .Z1_f (new_AGEMA_signal_4772) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_4_XOR12_U1 ( .A0_t (LED_128_Instance_SBox_Instance_4_L5), .A0_f (new_AGEMA_signal_4320), .A1_t (new_AGEMA_signal_4321), .A1_f (new_AGEMA_signal_4322), .B0_t (LED_128_Instance_SBox_Instance_4_T1), .B0_f (new_AGEMA_signal_4449), .B1_t (new_AGEMA_signal_4450), .B1_f (new_AGEMA_signal_4451), .Z0_t (LED_128_Instance_SBox_Instance_4_L8), .Z0_f (new_AGEMA_signal_4551), .Z1_t (new_AGEMA_signal_4552), .Z1_f (new_AGEMA_signal_4553) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_4_XOR13_U1 ( .A0_t (LED_128_Instance_SBox_Instance_4_L1), .A0_f (new_AGEMA_signal_3912), .A1_t (new_AGEMA_signal_3913), .A1_f (new_AGEMA_signal_3914), .B0_t (LED_128_Instance_SBox_Instance_4_L8), .B0_f (new_AGEMA_signal_4551), .B1_t (new_AGEMA_signal_4552), .B1_f (new_AGEMA_signal_4553), .Z0_t (LED_128_Instance_subcells_out[18]), .Z0_f (new_AGEMA_signal_4656), .Z1_t (new_AGEMA_signal_4657), .Z1_f (new_AGEMA_signal_4658) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_4_XOR14_U1 ( .A0_t (LED_128_Instance_SBox_Instance_4_L4), .A0_f (new_AGEMA_signal_3918), .A1_t (new_AGEMA_signal_3919), .A1_f (new_AGEMA_signal_3920), .B0_t (LED_128_Instance_SBox_Instance_4_T3), .B0_f (new_AGEMA_signal_4548), .B1_t (new_AGEMA_signal_4549), .B1_f (new_AGEMA_signal_4550), .Z0_t (LED_128_Instance_subcells_out[17]), .Z0_f (new_AGEMA_signal_4659), .Z1_t (new_AGEMA_signal_4660), .Z1_f (new_AGEMA_signal_4661) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_4_XOR15_U1 ( .A0_t (LED_128_Instance_SBox_Instance_4_L3), .A0_f (new_AGEMA_signal_3915), .A1_t (new_AGEMA_signal_3916), .A1_f (new_AGEMA_signal_3917), .B0_t (LED_128_Instance_SBox_Instance_4_T2), .B0_f (new_AGEMA_signal_3921), .B1_t (new_AGEMA_signal_3922), .B1_f (new_AGEMA_signal_3923), .Z0_t (LED_128_Instance_subcells_out[16]), .Z0_f (new_AGEMA_signal_4116), .Z1_t (new_AGEMA_signal_4117), .Z1_f (new_AGEMA_signal_4118) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_5_XOR1_U1 ( .A0_t (LED_128_Instance_addconst_out[22]), .A0_f (new_AGEMA_signal_3837), .A1_t (new_AGEMA_signal_3838), .A1_f (new_AGEMA_signal_3839), .B0_t (LED_128_Instance_addconst_out[21]), .B0_f (new_AGEMA_signal_3855), .B1_t (new_AGEMA_signal_3856), .B1_f (new_AGEMA_signal_3857), .Z0_t (LED_128_Instance_SBox_Instance_5_L0), .Z0_f (new_AGEMA_signal_4119), .Z1_t (new_AGEMA_signal_4120), .Z1_f (new_AGEMA_signal_4121) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_5_XOR2_U1 ( .A0_t (LED_128_Instance_addconst_out[21]), .A0_f (new_AGEMA_signal_3855), .A1_t (new_AGEMA_signal_3856), .A1_f (new_AGEMA_signal_3857), .B0_t (LED_128_Instance_addconst_out[20]), .B0_f (new_AGEMA_signal_3849), .B1_t (new_AGEMA_signal_3850), .B1_f (new_AGEMA_signal_3851), .Z0_t (LED_128_Instance_SBox_Instance_5_L1), .Z0_f (new_AGEMA_signal_4122), .Z1_t (new_AGEMA_signal_4123), .Z1_f (new_AGEMA_signal_4124) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_5_XOR3_U1 ( .A0_t (LED_128_Instance_SBox_Instance_5_L1), .A0_f (new_AGEMA_signal_4122), .A1_t (new_AGEMA_signal_4123), .A1_f (new_AGEMA_signal_4124), .B0_t (LED_128_Instance_addconst_out[23]), .B0_f (new_AGEMA_signal_3705), .B1_t (new_AGEMA_signal_3706), .B1_f (new_AGEMA_signal_3707), .Z0_t (LED_128_Instance_SBox_Instance_5_L2), .Z0_f (new_AGEMA_signal_4323), .Z1_t (new_AGEMA_signal_4324), .Z1_f (new_AGEMA_signal_4325) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_SBox_Instance_5_XOR16_U1 ( .A0_t (LED_128_Instance_SBox_Instance_5_T0), .A0_f (new_AGEMA_signal_4332), .A1_t (new_AGEMA_signal_4333), .A1_f (new_AGEMA_signal_4334), .B0_t (LED_128_Instance_SBox_Instance_5_L2), .B0_f (new_AGEMA_signal_4323), .B1_t (new_AGEMA_signal_4324), .B1_f (new_AGEMA_signal_4325), .Z0_t (LED_128_Instance_SBox_Instance_5_Q2), .Z0_f (new_AGEMA_signal_4452), .Z1_t (new_AGEMA_signal_4453), .Z1_f (new_AGEMA_signal_4454) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_5_XOR4_U1 ( .A0_t (LED_128_Instance_addconst_out[23]), .A0_f (new_AGEMA_signal_3705), .A1_t (new_AGEMA_signal_3706), .A1_f (new_AGEMA_signal_3707), .B0_t (LED_128_Instance_addconst_out[20]), .B0_f (new_AGEMA_signal_3849), .B1_t (new_AGEMA_signal_3850), .B1_f (new_AGEMA_signal_3851), .Z0_t (LED_128_Instance_SBox_Instance_5_L3), .Z0_f (new_AGEMA_signal_4125), .Z1_t (new_AGEMA_signal_4126), .Z1_f (new_AGEMA_signal_4127) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_5_XOR5_U1 ( .A0_t (LED_128_Instance_SBox_Instance_5_L3), .A0_f (new_AGEMA_signal_4125), .A1_t (new_AGEMA_signal_4126), .A1_f (new_AGEMA_signal_4127), .B0_t (LED_128_Instance_SBox_Instance_5_L0), .B0_f (new_AGEMA_signal_4119), .B1_t (new_AGEMA_signal_4120), .B1_f (new_AGEMA_signal_4121), .Z0_t (LED_128_Instance_SBox_Instance_5_Q3), .Z0_f (new_AGEMA_signal_4326), .Z1_t (new_AGEMA_signal_4327), .Z1_f (new_AGEMA_signal_4328) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_5_XOR6_U1 ( .A0_t (LED_128_Instance_addconst_out[23]), .A0_f (new_AGEMA_signal_3705), .A1_t (new_AGEMA_signal_3706), .A1_f (new_AGEMA_signal_3707), .B0_t (LED_128_Instance_addconst_out[21]), .B0_f (new_AGEMA_signal_3855), .B1_t (new_AGEMA_signal_3856), .B1_f (new_AGEMA_signal_3857), .Z0_t (LED_128_Instance_SBox_Instance_5_L4), .Z0_f (new_AGEMA_signal_4128), .Z1_t (new_AGEMA_signal_4129), .Z1_f (new_AGEMA_signal_4130) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_5_XOR7_U1 ( .A0_t (LED_128_Instance_SBox_Instance_5_T0), .A0_f (new_AGEMA_signal_4332), .A1_t (new_AGEMA_signal_4333), .A1_f (new_AGEMA_signal_4334), .B0_t (LED_128_Instance_SBox_Instance_5_T2), .B0_f (new_AGEMA_signal_4131), .B1_t (new_AGEMA_signal_4132), .B1_f (new_AGEMA_signal_4133), .Z0_t (LED_128_Instance_SBox_Instance_5_L5), .Z0_f (new_AGEMA_signal_4455), .Z1_t (new_AGEMA_signal_4456), .Z1_f (new_AGEMA_signal_4457) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_SBox_Instance_5_XOR8_U1 ( .A0_t (LED_128_Instance_SBox_Instance_5_L4), .A0_f (new_AGEMA_signal_4128), .A1_t (new_AGEMA_signal_4129), .A1_f (new_AGEMA_signal_4130), .B0_t (LED_128_Instance_SBox_Instance_5_L5), .B0_f (new_AGEMA_signal_4455), .B1_t (new_AGEMA_signal_4456), .B1_f (new_AGEMA_signal_4457), .Z0_t (LED_128_Instance_SBox_Instance_5_Q6), .Z0_f (new_AGEMA_signal_4554), .Z1_t (new_AGEMA_signal_4555), .Z1_f (new_AGEMA_signal_4556) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_5_XOR9_U1 ( .A0_t (LED_128_Instance_SBox_Instance_5_L1), .A0_f (new_AGEMA_signal_4122), .A1_t (new_AGEMA_signal_4123), .A1_f (new_AGEMA_signal_4124), .B0_t (LED_128_Instance_addconst_out[22]), .B0_f (new_AGEMA_signal_3837), .B1_t (new_AGEMA_signal_3838), .B1_f (new_AGEMA_signal_3839), .Z0_t (LED_128_Instance_SBox_Instance_5_Q7), .Z0_f (new_AGEMA_signal_4329), .Z1_t (new_AGEMA_signal_4330), .Z1_f (new_AGEMA_signal_4331) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_5_AND1_U1 ( .A0_t (LED_128_Instance_SBox_Instance_5_L0), .A0_f (new_AGEMA_signal_4119), .A1_t (new_AGEMA_signal_4120), .A1_f (new_AGEMA_signal_4121), .B0_t (LED_128_Instance_addconst_out[23]), .B0_f (new_AGEMA_signal_3705), .B1_t (new_AGEMA_signal_3706), .B1_f (new_AGEMA_signal_3707), .Z0_t (LED_128_Instance_SBox_Instance_5_T0), .Z0_f (new_AGEMA_signal_4332), .Z1_t (new_AGEMA_signal_4333), .Z1_f (new_AGEMA_signal_4334) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_5_AND2_U1 ( .A0_t (LED_128_Instance_SBox_Instance_5_Q2), .A0_f (new_AGEMA_signal_4452), .A1_t (new_AGEMA_signal_4453), .A1_f (new_AGEMA_signal_4454), .B0_t (LED_128_Instance_SBox_Instance_5_Q3), .B0_f (new_AGEMA_signal_4326), .B1_t (new_AGEMA_signal_4327), .B1_f (new_AGEMA_signal_4328), .Z0_t (LED_128_Instance_SBox_Instance_5_T1), .Z0_f (new_AGEMA_signal_4557), .Z1_t (new_AGEMA_signal_4558), .Z1_f (new_AGEMA_signal_4559) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_5_AND3_U1 ( .A0_t (LED_128_Instance_addconst_out[21]), .A0_f (new_AGEMA_signal_3855), .A1_t (new_AGEMA_signal_3856), .A1_f (new_AGEMA_signal_3857), .B0_t (LED_128_Instance_addconst_out[22]), .B0_f (new_AGEMA_signal_3837), .B1_t (new_AGEMA_signal_3838), .B1_f (new_AGEMA_signal_3839), .Z0_t (LED_128_Instance_SBox_Instance_5_T2), .Z0_f (new_AGEMA_signal_4131), .Z1_t (new_AGEMA_signal_4132), .Z1_f (new_AGEMA_signal_4133) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_5_AND4_U1 ( .A0_t (LED_128_Instance_SBox_Instance_5_Q6), .A0_f (new_AGEMA_signal_4554), .A1_t (new_AGEMA_signal_4555), .A1_f (new_AGEMA_signal_4556), .B0_t (LED_128_Instance_SBox_Instance_5_Q7), .B0_f (new_AGEMA_signal_4329), .B1_t (new_AGEMA_signal_4330), .B1_f (new_AGEMA_signal_4331), .Z0_t (LED_128_Instance_SBox_Instance_5_T3), .Z0_f (new_AGEMA_signal_4662), .Z1_t (new_AGEMA_signal_4663), .Z1_f (new_AGEMA_signal_4664) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_5_XOR10_U1 ( .A0_t (LED_128_Instance_SBox_Instance_5_L5), .A0_f (new_AGEMA_signal_4455), .A1_t (new_AGEMA_signal_4456), .A1_f (new_AGEMA_signal_4457), .B0_t (LED_128_Instance_SBox_Instance_5_T3), .B0_f (new_AGEMA_signal_4662), .B1_t (new_AGEMA_signal_4663), .B1_f (new_AGEMA_signal_4664), .Z0_t (LED_128_Instance_SBox_Instance_5_L7), .Z0_f (new_AGEMA_signal_4773), .Z1_t (new_AGEMA_signal_4774), .Z1_f (new_AGEMA_signal_4775) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_5_XOR11_U1 ( .A0_t (LED_128_Instance_addconst_out[20]), .A0_f (new_AGEMA_signal_3849), .A1_t (new_AGEMA_signal_3850), .A1_f (new_AGEMA_signal_3851), .B0_t (LED_128_Instance_SBox_Instance_5_L7), .B0_f (new_AGEMA_signal_4773), .B1_t (new_AGEMA_signal_4774), .B1_f (new_AGEMA_signal_4775), .Z0_t (LED_128_Instance_subcells_out[23]), .Z0_f (new_AGEMA_signal_4890), .Z1_t (new_AGEMA_signal_4891), .Z1_f (new_AGEMA_signal_4892) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_5_XOR12_U1 ( .A0_t (LED_128_Instance_SBox_Instance_5_L5), .A0_f (new_AGEMA_signal_4455), .A1_t (new_AGEMA_signal_4456), .A1_f (new_AGEMA_signal_4457), .B0_t (LED_128_Instance_SBox_Instance_5_T1), .B0_f (new_AGEMA_signal_4557), .B1_t (new_AGEMA_signal_4558), .B1_f (new_AGEMA_signal_4559), .Z0_t (LED_128_Instance_SBox_Instance_5_L8), .Z0_f (new_AGEMA_signal_4665), .Z1_t (new_AGEMA_signal_4666), .Z1_f (new_AGEMA_signal_4667) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_5_XOR13_U1 ( .A0_t (LED_128_Instance_SBox_Instance_5_L1), .A0_f (new_AGEMA_signal_4122), .A1_t (new_AGEMA_signal_4123), .A1_f (new_AGEMA_signal_4124), .B0_t (LED_128_Instance_SBox_Instance_5_L8), .B0_f (new_AGEMA_signal_4665), .B1_t (new_AGEMA_signal_4666), .B1_f (new_AGEMA_signal_4667), .Z0_t (LED_128_Instance_subcells_out[22]), .Z0_f (new_AGEMA_signal_4776), .Z1_t (new_AGEMA_signal_4777), .Z1_f (new_AGEMA_signal_4778) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_5_XOR14_U1 ( .A0_t (LED_128_Instance_SBox_Instance_5_L4), .A0_f (new_AGEMA_signal_4128), .A1_t (new_AGEMA_signal_4129), .A1_f (new_AGEMA_signal_4130), .B0_t (LED_128_Instance_SBox_Instance_5_T3), .B0_f (new_AGEMA_signal_4662), .B1_t (new_AGEMA_signal_4663), .B1_f (new_AGEMA_signal_4664), .Z0_t (LED_128_Instance_subcells_out[21]), .Z0_f (new_AGEMA_signal_4779), .Z1_t (new_AGEMA_signal_4780), .Z1_f (new_AGEMA_signal_4781) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_5_XOR15_U1 ( .A0_t (LED_128_Instance_SBox_Instance_5_L3), .A0_f (new_AGEMA_signal_4125), .A1_t (new_AGEMA_signal_4126), .A1_f (new_AGEMA_signal_4127), .B0_t (LED_128_Instance_SBox_Instance_5_T2), .B0_f (new_AGEMA_signal_4131), .B1_t (new_AGEMA_signal_4132), .B1_f (new_AGEMA_signal_4133), .Z0_t (LED_128_Instance_subcells_out[20]), .Z0_f (new_AGEMA_signal_4335), .Z1_t (new_AGEMA_signal_4336), .Z1_f (new_AGEMA_signal_4337) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_6_XOR1_U1 ( .A0_t (LED_128_Instance_addconst_out[26]), .A0_f (new_AGEMA_signal_3714), .A1_t (new_AGEMA_signal_3715), .A1_f (new_AGEMA_signal_3716), .B0_t (LED_128_Instance_addconst_out[25]), .B0_f (new_AGEMA_signal_3711), .B1_t (new_AGEMA_signal_3712), .B1_f (new_AGEMA_signal_3713), .Z0_t (LED_128_Instance_SBox_Instance_6_L0), .Z0_f (new_AGEMA_signal_3924), .Z1_t (new_AGEMA_signal_3925), .Z1_f (new_AGEMA_signal_3926) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_6_XOR2_U1 ( .A0_t (LED_128_Instance_addconst_out[25]), .A0_f (new_AGEMA_signal_3711), .A1_t (new_AGEMA_signal_3712), .A1_f (new_AGEMA_signal_3713), .B0_t (LED_128_Instance_addconst_out[24]), .B0_f (new_AGEMA_signal_3708), .B1_t (new_AGEMA_signal_3709), .B1_f (new_AGEMA_signal_3710), .Z0_t (LED_128_Instance_SBox_Instance_6_L1), .Z0_f (new_AGEMA_signal_3927), .Z1_t (new_AGEMA_signal_3928), .Z1_f (new_AGEMA_signal_3929) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_6_XOR3_U1 ( .A0_t (LED_128_Instance_SBox_Instance_6_L1), .A0_f (new_AGEMA_signal_3927), .A1_t (new_AGEMA_signal_3928), .A1_f (new_AGEMA_signal_3929), .B0_t (LED_128_Instance_addconst_out[27]), .B0_f (new_AGEMA_signal_3717), .B1_t (new_AGEMA_signal_3718), .B1_f (new_AGEMA_signal_3719), .Z0_t (LED_128_Instance_SBox_Instance_6_L2), .Z0_f (new_AGEMA_signal_4134), .Z1_t (new_AGEMA_signal_4135), .Z1_f (new_AGEMA_signal_4136) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_SBox_Instance_6_XOR16_U1 ( .A0_t (LED_128_Instance_SBox_Instance_6_T0), .A0_f (new_AGEMA_signal_4143), .A1_t (new_AGEMA_signal_4144), .A1_f (new_AGEMA_signal_4145), .B0_t (LED_128_Instance_SBox_Instance_6_L2), .B0_f (new_AGEMA_signal_4134), .B1_t (new_AGEMA_signal_4135), .B1_f (new_AGEMA_signal_4136), .Z0_t (LED_128_Instance_SBox_Instance_6_Q2), .Z0_f (new_AGEMA_signal_4338), .Z1_t (new_AGEMA_signal_4339), .Z1_f (new_AGEMA_signal_4340) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_6_XOR4_U1 ( .A0_t (LED_128_Instance_addconst_out[27]), .A0_f (new_AGEMA_signal_3717), .A1_t (new_AGEMA_signal_3718), .A1_f (new_AGEMA_signal_3719), .B0_t (LED_128_Instance_addconst_out[24]), .B0_f (new_AGEMA_signal_3708), .B1_t (new_AGEMA_signal_3709), .B1_f (new_AGEMA_signal_3710), .Z0_t (LED_128_Instance_SBox_Instance_6_L3), .Z0_f (new_AGEMA_signal_3930), .Z1_t (new_AGEMA_signal_3931), .Z1_f (new_AGEMA_signal_3932) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_6_XOR5_U1 ( .A0_t (LED_128_Instance_SBox_Instance_6_L3), .A0_f (new_AGEMA_signal_3930), .A1_t (new_AGEMA_signal_3931), .A1_f (new_AGEMA_signal_3932), .B0_t (LED_128_Instance_SBox_Instance_6_L0), .B0_f (new_AGEMA_signal_3924), .B1_t (new_AGEMA_signal_3925), .B1_f (new_AGEMA_signal_3926), .Z0_t (LED_128_Instance_SBox_Instance_6_Q3), .Z0_f (new_AGEMA_signal_4137), .Z1_t (new_AGEMA_signal_4138), .Z1_f (new_AGEMA_signal_4139) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_6_XOR6_U1 ( .A0_t (LED_128_Instance_addconst_out[27]), .A0_f (new_AGEMA_signal_3717), .A1_t (new_AGEMA_signal_3718), .A1_f (new_AGEMA_signal_3719), .B0_t (LED_128_Instance_addconst_out[25]), .B0_f (new_AGEMA_signal_3711), .B1_t (new_AGEMA_signal_3712), .B1_f (new_AGEMA_signal_3713), .Z0_t (LED_128_Instance_SBox_Instance_6_L4), .Z0_f (new_AGEMA_signal_3933), .Z1_t (new_AGEMA_signal_3934), .Z1_f (new_AGEMA_signal_3935) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_6_XOR7_U1 ( .A0_t (LED_128_Instance_SBox_Instance_6_T0), .A0_f (new_AGEMA_signal_4143), .A1_t (new_AGEMA_signal_4144), .A1_f (new_AGEMA_signal_4145), .B0_t (LED_128_Instance_SBox_Instance_6_T2), .B0_f (new_AGEMA_signal_3936), .B1_t (new_AGEMA_signal_3937), .B1_f (new_AGEMA_signal_3938), .Z0_t (LED_128_Instance_SBox_Instance_6_L5), .Z0_f (new_AGEMA_signal_4341), .Z1_t (new_AGEMA_signal_4342), .Z1_f (new_AGEMA_signal_4343) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_SBox_Instance_6_XOR8_U1 ( .A0_t (LED_128_Instance_SBox_Instance_6_L4), .A0_f (new_AGEMA_signal_3933), .A1_t (new_AGEMA_signal_3934), .A1_f (new_AGEMA_signal_3935), .B0_t (LED_128_Instance_SBox_Instance_6_L5), .B0_f (new_AGEMA_signal_4341), .B1_t (new_AGEMA_signal_4342), .B1_f (new_AGEMA_signal_4343), .Z0_t (LED_128_Instance_SBox_Instance_6_Q6), .Z0_f (new_AGEMA_signal_4458), .Z1_t (new_AGEMA_signal_4459), .Z1_f (new_AGEMA_signal_4460) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_6_XOR9_U1 ( .A0_t (LED_128_Instance_SBox_Instance_6_L1), .A0_f (new_AGEMA_signal_3927), .A1_t (new_AGEMA_signal_3928), .A1_f (new_AGEMA_signal_3929), .B0_t (LED_128_Instance_addconst_out[26]), .B0_f (new_AGEMA_signal_3714), .B1_t (new_AGEMA_signal_3715), .B1_f (new_AGEMA_signal_3716), .Z0_t (LED_128_Instance_SBox_Instance_6_Q7), .Z0_f (new_AGEMA_signal_4140), .Z1_t (new_AGEMA_signal_4141), .Z1_f (new_AGEMA_signal_4142) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_6_AND1_U1 ( .A0_t (LED_128_Instance_SBox_Instance_6_L0), .A0_f (new_AGEMA_signal_3924), .A1_t (new_AGEMA_signal_3925), .A1_f (new_AGEMA_signal_3926), .B0_t (LED_128_Instance_addconst_out[27]), .B0_f (new_AGEMA_signal_3717), .B1_t (new_AGEMA_signal_3718), .B1_f (new_AGEMA_signal_3719), .Z0_t (LED_128_Instance_SBox_Instance_6_T0), .Z0_f (new_AGEMA_signal_4143), .Z1_t (new_AGEMA_signal_4144), .Z1_f (new_AGEMA_signal_4145) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_6_AND2_U1 ( .A0_t (LED_128_Instance_SBox_Instance_6_Q2), .A0_f (new_AGEMA_signal_4338), .A1_t (new_AGEMA_signal_4339), .A1_f (new_AGEMA_signal_4340), .B0_t (LED_128_Instance_SBox_Instance_6_Q3), .B0_f (new_AGEMA_signal_4137), .B1_t (new_AGEMA_signal_4138), .B1_f (new_AGEMA_signal_4139), .Z0_t (LED_128_Instance_SBox_Instance_6_T1), .Z0_f (new_AGEMA_signal_4461), .Z1_t (new_AGEMA_signal_4462), .Z1_f (new_AGEMA_signal_4463) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_6_AND3_U1 ( .A0_t (LED_128_Instance_addconst_out[25]), .A0_f (new_AGEMA_signal_3711), .A1_t (new_AGEMA_signal_3712), .A1_f (new_AGEMA_signal_3713), .B0_t (LED_128_Instance_addconst_out[26]), .B0_f (new_AGEMA_signal_3714), .B1_t (new_AGEMA_signal_3715), .B1_f (new_AGEMA_signal_3716), .Z0_t (LED_128_Instance_SBox_Instance_6_T2), .Z0_f (new_AGEMA_signal_3936), .Z1_t (new_AGEMA_signal_3937), .Z1_f (new_AGEMA_signal_3938) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_6_AND4_U1 ( .A0_t (LED_128_Instance_SBox_Instance_6_Q6), .A0_f (new_AGEMA_signal_4458), .A1_t (new_AGEMA_signal_4459), .A1_f (new_AGEMA_signal_4460), .B0_t (LED_128_Instance_SBox_Instance_6_Q7), .B0_f (new_AGEMA_signal_4140), .B1_t (new_AGEMA_signal_4141), .B1_f (new_AGEMA_signal_4142), .Z0_t (LED_128_Instance_SBox_Instance_6_T3), .Z0_f (new_AGEMA_signal_4560), .Z1_t (new_AGEMA_signal_4561), .Z1_f (new_AGEMA_signal_4562) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_6_XOR10_U1 ( .A0_t (LED_128_Instance_SBox_Instance_6_L5), .A0_f (new_AGEMA_signal_4341), .A1_t (new_AGEMA_signal_4342), .A1_f (new_AGEMA_signal_4343), .B0_t (LED_128_Instance_SBox_Instance_6_T3), .B0_f (new_AGEMA_signal_4560), .B1_t (new_AGEMA_signal_4561), .B1_f (new_AGEMA_signal_4562), .Z0_t (LED_128_Instance_SBox_Instance_6_L7), .Z0_f (new_AGEMA_signal_4668), .Z1_t (new_AGEMA_signal_4669), .Z1_f (new_AGEMA_signal_4670) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_6_XOR11_U1 ( .A0_t (LED_128_Instance_addconst_out[24]), .A0_f (new_AGEMA_signal_3708), .A1_t (new_AGEMA_signal_3709), .A1_f (new_AGEMA_signal_3710), .B0_t (LED_128_Instance_SBox_Instance_6_L7), .B0_f (new_AGEMA_signal_4668), .B1_t (new_AGEMA_signal_4669), .B1_f (new_AGEMA_signal_4670), .Z0_t (LED_128_Instance_subcells_out[27]), .Z0_f (new_AGEMA_signal_4782), .Z1_t (new_AGEMA_signal_4783), .Z1_f (new_AGEMA_signal_4784) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_6_XOR12_U1 ( .A0_t (LED_128_Instance_SBox_Instance_6_L5), .A0_f (new_AGEMA_signal_4341), .A1_t (new_AGEMA_signal_4342), .A1_f (new_AGEMA_signal_4343), .B0_t (LED_128_Instance_SBox_Instance_6_T1), .B0_f (new_AGEMA_signal_4461), .B1_t (new_AGEMA_signal_4462), .B1_f (new_AGEMA_signal_4463), .Z0_t (LED_128_Instance_SBox_Instance_6_L8), .Z0_f (new_AGEMA_signal_4563), .Z1_t (new_AGEMA_signal_4564), .Z1_f (new_AGEMA_signal_4565) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_6_XOR13_U1 ( .A0_t (LED_128_Instance_SBox_Instance_6_L1), .A0_f (new_AGEMA_signal_3927), .A1_t (new_AGEMA_signal_3928), .A1_f (new_AGEMA_signal_3929), .B0_t (LED_128_Instance_SBox_Instance_6_L8), .B0_f (new_AGEMA_signal_4563), .B1_t (new_AGEMA_signal_4564), .B1_f (new_AGEMA_signal_4565), .Z0_t (LED_128_Instance_subcells_out[26]), .Z0_f (new_AGEMA_signal_4671), .Z1_t (new_AGEMA_signal_4672), .Z1_f (new_AGEMA_signal_4673) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_6_XOR14_U1 ( .A0_t (LED_128_Instance_SBox_Instance_6_L4), .A0_f (new_AGEMA_signal_3933), .A1_t (new_AGEMA_signal_3934), .A1_f (new_AGEMA_signal_3935), .B0_t (LED_128_Instance_SBox_Instance_6_T3), .B0_f (new_AGEMA_signal_4560), .B1_t (new_AGEMA_signal_4561), .B1_f (new_AGEMA_signal_4562), .Z0_t (LED_128_Instance_subcells_out[25]), .Z0_f (new_AGEMA_signal_4674), .Z1_t (new_AGEMA_signal_4675), .Z1_f (new_AGEMA_signal_4676) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_6_XOR15_U1 ( .A0_t (LED_128_Instance_SBox_Instance_6_L3), .A0_f (new_AGEMA_signal_3930), .A1_t (new_AGEMA_signal_3931), .A1_f (new_AGEMA_signal_3932), .B0_t (LED_128_Instance_SBox_Instance_6_T2), .B0_f (new_AGEMA_signal_3936), .B1_t (new_AGEMA_signal_3937), .B1_f (new_AGEMA_signal_3938), .Z0_t (LED_128_Instance_subcells_out[24]), .Z0_f (new_AGEMA_signal_4146), .Z1_t (new_AGEMA_signal_4147), .Z1_f (new_AGEMA_signal_4148) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_7_XOR1_U1 ( .A0_t (LED_128_Instance_addconst_out[30]), .A0_f (new_AGEMA_signal_3726), .A1_t (new_AGEMA_signal_3727), .A1_f (new_AGEMA_signal_3728), .B0_t (LED_128_Instance_addconst_out[29]), .B0_f (new_AGEMA_signal_3723), .B1_t (new_AGEMA_signal_3724), .B1_f (new_AGEMA_signal_3725), .Z0_t (LED_128_Instance_SBox_Instance_7_L0), .Z0_f (new_AGEMA_signal_3939), .Z1_t (new_AGEMA_signal_3940), .Z1_f (new_AGEMA_signal_3941) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_7_XOR2_U1 ( .A0_t (LED_128_Instance_addconst_out[29]), .A0_f (new_AGEMA_signal_3723), .A1_t (new_AGEMA_signal_3724), .A1_f (new_AGEMA_signal_3725), .B0_t (LED_128_Instance_addconst_out[28]), .B0_f (new_AGEMA_signal_3720), .B1_t (new_AGEMA_signal_3721), .B1_f (new_AGEMA_signal_3722), .Z0_t (LED_128_Instance_SBox_Instance_7_L1), .Z0_f (new_AGEMA_signal_3942), .Z1_t (new_AGEMA_signal_3943), .Z1_f (new_AGEMA_signal_3944) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_7_XOR3_U1 ( .A0_t (LED_128_Instance_SBox_Instance_7_L1), .A0_f (new_AGEMA_signal_3942), .A1_t (new_AGEMA_signal_3943), .A1_f (new_AGEMA_signal_3944), .B0_t (LED_128_Instance_addconst_out[31]), .B0_f (new_AGEMA_signal_3729), .B1_t (new_AGEMA_signal_3730), .B1_f (new_AGEMA_signal_3731), .Z0_t (LED_128_Instance_SBox_Instance_7_L2), .Z0_f (new_AGEMA_signal_4149), .Z1_t (new_AGEMA_signal_4150), .Z1_f (new_AGEMA_signal_4151) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_SBox_Instance_7_XOR16_U1 ( .A0_t (LED_128_Instance_SBox_Instance_7_T0), .A0_f (new_AGEMA_signal_4158), .A1_t (new_AGEMA_signal_4159), .A1_f (new_AGEMA_signal_4160), .B0_t (LED_128_Instance_SBox_Instance_7_L2), .B0_f (new_AGEMA_signal_4149), .B1_t (new_AGEMA_signal_4150), .B1_f (new_AGEMA_signal_4151), .Z0_t (LED_128_Instance_SBox_Instance_7_Q2), .Z0_f (new_AGEMA_signal_4344), .Z1_t (new_AGEMA_signal_4345), .Z1_f (new_AGEMA_signal_4346) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_7_XOR4_U1 ( .A0_t (LED_128_Instance_addconst_out[31]), .A0_f (new_AGEMA_signal_3729), .A1_t (new_AGEMA_signal_3730), .A1_f (new_AGEMA_signal_3731), .B0_t (LED_128_Instance_addconst_out[28]), .B0_f (new_AGEMA_signal_3720), .B1_t (new_AGEMA_signal_3721), .B1_f (new_AGEMA_signal_3722), .Z0_t (LED_128_Instance_SBox_Instance_7_L3), .Z0_f (new_AGEMA_signal_3945), .Z1_t (new_AGEMA_signal_3946), .Z1_f (new_AGEMA_signal_3947) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_7_XOR5_U1 ( .A0_t (LED_128_Instance_SBox_Instance_7_L3), .A0_f (new_AGEMA_signal_3945), .A1_t (new_AGEMA_signal_3946), .A1_f (new_AGEMA_signal_3947), .B0_t (LED_128_Instance_SBox_Instance_7_L0), .B0_f (new_AGEMA_signal_3939), .B1_t (new_AGEMA_signal_3940), .B1_f (new_AGEMA_signal_3941), .Z0_t (LED_128_Instance_SBox_Instance_7_Q3), .Z0_f (new_AGEMA_signal_4152), .Z1_t (new_AGEMA_signal_4153), .Z1_f (new_AGEMA_signal_4154) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_7_XOR6_U1 ( .A0_t (LED_128_Instance_addconst_out[31]), .A0_f (new_AGEMA_signal_3729), .A1_t (new_AGEMA_signal_3730), .A1_f (new_AGEMA_signal_3731), .B0_t (LED_128_Instance_addconst_out[29]), .B0_f (new_AGEMA_signal_3723), .B1_t (new_AGEMA_signal_3724), .B1_f (new_AGEMA_signal_3725), .Z0_t (LED_128_Instance_SBox_Instance_7_L4), .Z0_f (new_AGEMA_signal_3948), .Z1_t (new_AGEMA_signal_3949), .Z1_f (new_AGEMA_signal_3950) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_7_XOR7_U1 ( .A0_t (LED_128_Instance_SBox_Instance_7_T0), .A0_f (new_AGEMA_signal_4158), .A1_t (new_AGEMA_signal_4159), .A1_f (new_AGEMA_signal_4160), .B0_t (LED_128_Instance_SBox_Instance_7_T2), .B0_f (new_AGEMA_signal_3951), .B1_t (new_AGEMA_signal_3952), .B1_f (new_AGEMA_signal_3953), .Z0_t (LED_128_Instance_SBox_Instance_7_L5), .Z0_f (new_AGEMA_signal_4347), .Z1_t (new_AGEMA_signal_4348), .Z1_f (new_AGEMA_signal_4349) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_SBox_Instance_7_XOR8_U1 ( .A0_t (LED_128_Instance_SBox_Instance_7_L4), .A0_f (new_AGEMA_signal_3948), .A1_t (new_AGEMA_signal_3949), .A1_f (new_AGEMA_signal_3950), .B0_t (LED_128_Instance_SBox_Instance_7_L5), .B0_f (new_AGEMA_signal_4347), .B1_t (new_AGEMA_signal_4348), .B1_f (new_AGEMA_signal_4349), .Z0_t (LED_128_Instance_SBox_Instance_7_Q6), .Z0_f (new_AGEMA_signal_4464), .Z1_t (new_AGEMA_signal_4465), .Z1_f (new_AGEMA_signal_4466) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_7_XOR9_U1 ( .A0_t (LED_128_Instance_SBox_Instance_7_L1), .A0_f (new_AGEMA_signal_3942), .A1_t (new_AGEMA_signal_3943), .A1_f (new_AGEMA_signal_3944), .B0_t (LED_128_Instance_addconst_out[30]), .B0_f (new_AGEMA_signal_3726), .B1_t (new_AGEMA_signal_3727), .B1_f (new_AGEMA_signal_3728), .Z0_t (LED_128_Instance_SBox_Instance_7_Q7), .Z0_f (new_AGEMA_signal_4155), .Z1_t (new_AGEMA_signal_4156), .Z1_f (new_AGEMA_signal_4157) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_7_AND1_U1 ( .A0_t (LED_128_Instance_SBox_Instance_7_L0), .A0_f (new_AGEMA_signal_3939), .A1_t (new_AGEMA_signal_3940), .A1_f (new_AGEMA_signal_3941), .B0_t (LED_128_Instance_addconst_out[31]), .B0_f (new_AGEMA_signal_3729), .B1_t (new_AGEMA_signal_3730), .B1_f (new_AGEMA_signal_3731), .Z0_t (LED_128_Instance_SBox_Instance_7_T0), .Z0_f (new_AGEMA_signal_4158), .Z1_t (new_AGEMA_signal_4159), .Z1_f (new_AGEMA_signal_4160) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_7_AND2_U1 ( .A0_t (LED_128_Instance_SBox_Instance_7_Q2), .A0_f (new_AGEMA_signal_4344), .A1_t (new_AGEMA_signal_4345), .A1_f (new_AGEMA_signal_4346), .B0_t (LED_128_Instance_SBox_Instance_7_Q3), .B0_f (new_AGEMA_signal_4152), .B1_t (new_AGEMA_signal_4153), .B1_f (new_AGEMA_signal_4154), .Z0_t (LED_128_Instance_SBox_Instance_7_T1), .Z0_f (new_AGEMA_signal_4467), .Z1_t (new_AGEMA_signal_4468), .Z1_f (new_AGEMA_signal_4469) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_7_AND3_U1 ( .A0_t (LED_128_Instance_addconst_out[29]), .A0_f (new_AGEMA_signal_3723), .A1_t (new_AGEMA_signal_3724), .A1_f (new_AGEMA_signal_3725), .B0_t (LED_128_Instance_addconst_out[30]), .B0_f (new_AGEMA_signal_3726), .B1_t (new_AGEMA_signal_3727), .B1_f (new_AGEMA_signal_3728), .Z0_t (LED_128_Instance_SBox_Instance_7_T2), .Z0_f (new_AGEMA_signal_3951), .Z1_t (new_AGEMA_signal_3952), .Z1_f (new_AGEMA_signal_3953) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_7_AND4_U1 ( .A0_t (LED_128_Instance_SBox_Instance_7_Q6), .A0_f (new_AGEMA_signal_4464), .A1_t (new_AGEMA_signal_4465), .A1_f (new_AGEMA_signal_4466), .B0_t (LED_128_Instance_SBox_Instance_7_Q7), .B0_f (new_AGEMA_signal_4155), .B1_t (new_AGEMA_signal_4156), .B1_f (new_AGEMA_signal_4157), .Z0_t (LED_128_Instance_SBox_Instance_7_T3), .Z0_f (new_AGEMA_signal_4566), .Z1_t (new_AGEMA_signal_4567), .Z1_f (new_AGEMA_signal_4568) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_7_XOR10_U1 ( .A0_t (LED_128_Instance_SBox_Instance_7_L5), .A0_f (new_AGEMA_signal_4347), .A1_t (new_AGEMA_signal_4348), .A1_f (new_AGEMA_signal_4349), .B0_t (LED_128_Instance_SBox_Instance_7_T3), .B0_f (new_AGEMA_signal_4566), .B1_t (new_AGEMA_signal_4567), .B1_f (new_AGEMA_signal_4568), .Z0_t (LED_128_Instance_SBox_Instance_7_L7), .Z0_f (new_AGEMA_signal_4677), .Z1_t (new_AGEMA_signal_4678), .Z1_f (new_AGEMA_signal_4679) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_7_XOR11_U1 ( .A0_t (LED_128_Instance_addconst_out[28]), .A0_f (new_AGEMA_signal_3720), .A1_t (new_AGEMA_signal_3721), .A1_f (new_AGEMA_signal_3722), .B0_t (LED_128_Instance_SBox_Instance_7_L7), .B0_f (new_AGEMA_signal_4677), .B1_t (new_AGEMA_signal_4678), .B1_f (new_AGEMA_signal_4679), .Z0_t (LED_128_Instance_subcells_out[31]), .Z0_f (new_AGEMA_signal_4785), .Z1_t (new_AGEMA_signal_4786), .Z1_f (new_AGEMA_signal_4787) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_7_XOR12_U1 ( .A0_t (LED_128_Instance_SBox_Instance_7_L5), .A0_f (new_AGEMA_signal_4347), .A1_t (new_AGEMA_signal_4348), .A1_f (new_AGEMA_signal_4349), .B0_t (LED_128_Instance_SBox_Instance_7_T1), .B0_f (new_AGEMA_signal_4467), .B1_t (new_AGEMA_signal_4468), .B1_f (new_AGEMA_signal_4469), .Z0_t (LED_128_Instance_SBox_Instance_7_L8), .Z0_f (new_AGEMA_signal_4569), .Z1_t (new_AGEMA_signal_4570), .Z1_f (new_AGEMA_signal_4571) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_7_XOR13_U1 ( .A0_t (LED_128_Instance_SBox_Instance_7_L1), .A0_f (new_AGEMA_signal_3942), .A1_t (new_AGEMA_signal_3943), .A1_f (new_AGEMA_signal_3944), .B0_t (LED_128_Instance_SBox_Instance_7_L8), .B0_f (new_AGEMA_signal_4569), .B1_t (new_AGEMA_signal_4570), .B1_f (new_AGEMA_signal_4571), .Z0_t (LED_128_Instance_subcells_out[30]), .Z0_f (new_AGEMA_signal_4680), .Z1_t (new_AGEMA_signal_4681), .Z1_f (new_AGEMA_signal_4682) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_7_XOR14_U1 ( .A0_t (LED_128_Instance_SBox_Instance_7_L4), .A0_f (new_AGEMA_signal_3948), .A1_t (new_AGEMA_signal_3949), .A1_f (new_AGEMA_signal_3950), .B0_t (LED_128_Instance_SBox_Instance_7_T3), .B0_f (new_AGEMA_signal_4566), .B1_t (new_AGEMA_signal_4567), .B1_f (new_AGEMA_signal_4568), .Z0_t (LED_128_Instance_subcells_out[29]), .Z0_f (new_AGEMA_signal_4683), .Z1_t (new_AGEMA_signal_4684), .Z1_f (new_AGEMA_signal_4685) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_7_XOR15_U1 ( .A0_t (LED_128_Instance_SBox_Instance_7_L3), .A0_f (new_AGEMA_signal_3945), .A1_t (new_AGEMA_signal_3946), .A1_f (new_AGEMA_signal_3947), .B0_t (LED_128_Instance_SBox_Instance_7_T2), .B0_f (new_AGEMA_signal_3951), .B1_t (new_AGEMA_signal_3952), .B1_f (new_AGEMA_signal_3953), .Z0_t (LED_128_Instance_subcells_out[28]), .Z0_f (new_AGEMA_signal_4161), .Z1_t (new_AGEMA_signal_4162), .Z1_f (new_AGEMA_signal_4163) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_8_XOR1_U1 ( .A0_t (LED_128_Instance_addconst_out[34]), .A0_f (new_AGEMA_signal_3738), .A1_t (new_AGEMA_signal_3739), .A1_f (new_AGEMA_signal_3740), .B0_t (LED_128_Instance_addroundkey_out[33]), .B0_f (new_AGEMA_signal_3735), .B1_t (new_AGEMA_signal_3736), .B1_f (new_AGEMA_signal_3737), .Z0_t (LED_128_Instance_SBox_Instance_8_L0), .Z0_f (new_AGEMA_signal_3954), .Z1_t (new_AGEMA_signal_3955), .Z1_f (new_AGEMA_signal_3956) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_8_XOR2_U1 ( .A0_t (LED_128_Instance_addroundkey_out[33]), .A0_f (new_AGEMA_signal_3735), .A1_t (new_AGEMA_signal_3736), .A1_f (new_AGEMA_signal_3737), .B0_t (LED_128_Instance_addconst_out[32]), .B0_f (new_AGEMA_signal_3732), .B1_t (new_AGEMA_signal_3733), .B1_f (new_AGEMA_signal_3734), .Z0_t (LED_128_Instance_SBox_Instance_8_L1), .Z0_f (new_AGEMA_signal_3957), .Z1_t (new_AGEMA_signal_3958), .Z1_f (new_AGEMA_signal_3959) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_8_XOR3_U1 ( .A0_t (LED_128_Instance_SBox_Instance_8_L1), .A0_f (new_AGEMA_signal_3957), .A1_t (new_AGEMA_signal_3958), .A1_f (new_AGEMA_signal_3959), .B0_t (LED_128_Instance_addconst_out[35]), .B0_f (new_AGEMA_signal_3741), .B1_t (new_AGEMA_signal_3742), .B1_f (new_AGEMA_signal_3743), .Z0_t (LED_128_Instance_SBox_Instance_8_L2), .Z0_f (new_AGEMA_signal_4164), .Z1_t (new_AGEMA_signal_4165), .Z1_f (new_AGEMA_signal_4166) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_SBox_Instance_8_XOR16_U1 ( .A0_t (LED_128_Instance_SBox_Instance_8_T0), .A0_f (new_AGEMA_signal_4173), .A1_t (new_AGEMA_signal_4174), .A1_f (new_AGEMA_signal_4175), .B0_t (LED_128_Instance_SBox_Instance_8_L2), .B0_f (new_AGEMA_signal_4164), .B1_t (new_AGEMA_signal_4165), .B1_f (new_AGEMA_signal_4166), .Z0_t (LED_128_Instance_SBox_Instance_8_Q2), .Z0_f (new_AGEMA_signal_4350), .Z1_t (new_AGEMA_signal_4351), .Z1_f (new_AGEMA_signal_4352) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_8_XOR4_U1 ( .A0_t (LED_128_Instance_addconst_out[35]), .A0_f (new_AGEMA_signal_3741), .A1_t (new_AGEMA_signal_3742), .A1_f (new_AGEMA_signal_3743), .B0_t (LED_128_Instance_addconst_out[32]), .B0_f (new_AGEMA_signal_3732), .B1_t (new_AGEMA_signal_3733), .B1_f (new_AGEMA_signal_3734), .Z0_t (LED_128_Instance_SBox_Instance_8_L3), .Z0_f (new_AGEMA_signal_3960), .Z1_t (new_AGEMA_signal_3961), .Z1_f (new_AGEMA_signal_3962) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_8_XOR5_U1 ( .A0_t (LED_128_Instance_SBox_Instance_8_L3), .A0_f (new_AGEMA_signal_3960), .A1_t (new_AGEMA_signal_3961), .A1_f (new_AGEMA_signal_3962), .B0_t (LED_128_Instance_SBox_Instance_8_L0), .B0_f (new_AGEMA_signal_3954), .B1_t (new_AGEMA_signal_3955), .B1_f (new_AGEMA_signal_3956), .Z0_t (LED_128_Instance_SBox_Instance_8_Q3), .Z0_f (new_AGEMA_signal_4167), .Z1_t (new_AGEMA_signal_4168), .Z1_f (new_AGEMA_signal_4169) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_8_XOR6_U1 ( .A0_t (LED_128_Instance_addconst_out[35]), .A0_f (new_AGEMA_signal_3741), .A1_t (new_AGEMA_signal_3742), .A1_f (new_AGEMA_signal_3743), .B0_t (LED_128_Instance_addroundkey_out[33]), .B0_f (new_AGEMA_signal_3735), .B1_t (new_AGEMA_signal_3736), .B1_f (new_AGEMA_signal_3737), .Z0_t (LED_128_Instance_SBox_Instance_8_L4), .Z0_f (new_AGEMA_signal_3963), .Z1_t (new_AGEMA_signal_3964), .Z1_f (new_AGEMA_signal_3965) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_8_XOR7_U1 ( .A0_t (LED_128_Instance_SBox_Instance_8_T0), .A0_f (new_AGEMA_signal_4173), .A1_t (new_AGEMA_signal_4174), .A1_f (new_AGEMA_signal_4175), .B0_t (LED_128_Instance_SBox_Instance_8_T2), .B0_f (new_AGEMA_signal_3966), .B1_t (new_AGEMA_signal_3967), .B1_f (new_AGEMA_signal_3968), .Z0_t (LED_128_Instance_SBox_Instance_8_L5), .Z0_f (new_AGEMA_signal_4353), .Z1_t (new_AGEMA_signal_4354), .Z1_f (new_AGEMA_signal_4355) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_SBox_Instance_8_XOR8_U1 ( .A0_t (LED_128_Instance_SBox_Instance_8_L4), .A0_f (new_AGEMA_signal_3963), .A1_t (new_AGEMA_signal_3964), .A1_f (new_AGEMA_signal_3965), .B0_t (LED_128_Instance_SBox_Instance_8_L5), .B0_f (new_AGEMA_signal_4353), .B1_t (new_AGEMA_signal_4354), .B1_f (new_AGEMA_signal_4355), .Z0_t (LED_128_Instance_SBox_Instance_8_Q6), .Z0_f (new_AGEMA_signal_4470), .Z1_t (new_AGEMA_signal_4471), .Z1_f (new_AGEMA_signal_4472) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_8_XOR9_U1 ( .A0_t (LED_128_Instance_SBox_Instance_8_L1), .A0_f (new_AGEMA_signal_3957), .A1_t (new_AGEMA_signal_3958), .A1_f (new_AGEMA_signal_3959), .B0_t (LED_128_Instance_addconst_out[34]), .B0_f (new_AGEMA_signal_3738), .B1_t (new_AGEMA_signal_3739), .B1_f (new_AGEMA_signal_3740), .Z0_t (LED_128_Instance_SBox_Instance_8_Q7), .Z0_f (new_AGEMA_signal_4170), .Z1_t (new_AGEMA_signal_4171), .Z1_f (new_AGEMA_signal_4172) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_8_AND1_U1 ( .A0_t (LED_128_Instance_SBox_Instance_8_L0), .A0_f (new_AGEMA_signal_3954), .A1_t (new_AGEMA_signal_3955), .A1_f (new_AGEMA_signal_3956), .B0_t (LED_128_Instance_addconst_out[35]), .B0_f (new_AGEMA_signal_3741), .B1_t (new_AGEMA_signal_3742), .B1_f (new_AGEMA_signal_3743), .Z0_t (LED_128_Instance_SBox_Instance_8_T0), .Z0_f (new_AGEMA_signal_4173), .Z1_t (new_AGEMA_signal_4174), .Z1_f (new_AGEMA_signal_4175) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_8_AND2_U1 ( .A0_t (LED_128_Instance_SBox_Instance_8_Q2), .A0_f (new_AGEMA_signal_4350), .A1_t (new_AGEMA_signal_4351), .A1_f (new_AGEMA_signal_4352), .B0_t (LED_128_Instance_SBox_Instance_8_Q3), .B0_f (new_AGEMA_signal_4167), .B1_t (new_AGEMA_signal_4168), .B1_f (new_AGEMA_signal_4169), .Z0_t (LED_128_Instance_SBox_Instance_8_T1), .Z0_f (new_AGEMA_signal_4473), .Z1_t (new_AGEMA_signal_4474), .Z1_f (new_AGEMA_signal_4475) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_8_AND3_U1 ( .A0_t (LED_128_Instance_addroundkey_out[33]), .A0_f (new_AGEMA_signal_3735), .A1_t (new_AGEMA_signal_3736), .A1_f (new_AGEMA_signal_3737), .B0_t (LED_128_Instance_addconst_out[34]), .B0_f (new_AGEMA_signal_3738), .B1_t (new_AGEMA_signal_3739), .B1_f (new_AGEMA_signal_3740), .Z0_t (LED_128_Instance_SBox_Instance_8_T2), .Z0_f (new_AGEMA_signal_3966), .Z1_t (new_AGEMA_signal_3967), .Z1_f (new_AGEMA_signal_3968) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_8_AND4_U1 ( .A0_t (LED_128_Instance_SBox_Instance_8_Q6), .A0_f (new_AGEMA_signal_4470), .A1_t (new_AGEMA_signal_4471), .A1_f (new_AGEMA_signal_4472), .B0_t (LED_128_Instance_SBox_Instance_8_Q7), .B0_f (new_AGEMA_signal_4170), .B1_t (new_AGEMA_signal_4171), .B1_f (new_AGEMA_signal_4172), .Z0_t (LED_128_Instance_SBox_Instance_8_T3), .Z0_f (new_AGEMA_signal_4572), .Z1_t (new_AGEMA_signal_4573), .Z1_f (new_AGEMA_signal_4574) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_8_XOR10_U1 ( .A0_t (LED_128_Instance_SBox_Instance_8_L5), .A0_f (new_AGEMA_signal_4353), .A1_t (new_AGEMA_signal_4354), .A1_f (new_AGEMA_signal_4355), .B0_t (LED_128_Instance_SBox_Instance_8_T3), .B0_f (new_AGEMA_signal_4572), .B1_t (new_AGEMA_signal_4573), .B1_f (new_AGEMA_signal_4574), .Z0_t (LED_128_Instance_SBox_Instance_8_L7), .Z0_f (new_AGEMA_signal_4686), .Z1_t (new_AGEMA_signal_4687), .Z1_f (new_AGEMA_signal_4688) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_8_XOR11_U1 ( .A0_t (LED_128_Instance_addconst_out[32]), .A0_f (new_AGEMA_signal_3732), .A1_t (new_AGEMA_signal_3733), .A1_f (new_AGEMA_signal_3734), .B0_t (LED_128_Instance_SBox_Instance_8_L7), .B0_f (new_AGEMA_signal_4686), .B1_t (new_AGEMA_signal_4687), .B1_f (new_AGEMA_signal_4688), .Z0_t (LED_128_Instance_subcells_out[35]), .Z0_f (new_AGEMA_signal_4788), .Z1_t (new_AGEMA_signal_4789), .Z1_f (new_AGEMA_signal_4790) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_8_XOR12_U1 ( .A0_t (LED_128_Instance_SBox_Instance_8_L5), .A0_f (new_AGEMA_signal_4353), .A1_t (new_AGEMA_signal_4354), .A1_f (new_AGEMA_signal_4355), .B0_t (LED_128_Instance_SBox_Instance_8_T1), .B0_f (new_AGEMA_signal_4473), .B1_t (new_AGEMA_signal_4474), .B1_f (new_AGEMA_signal_4475), .Z0_t (LED_128_Instance_SBox_Instance_8_L8), .Z0_f (new_AGEMA_signal_4575), .Z1_t (new_AGEMA_signal_4576), .Z1_f (new_AGEMA_signal_4577) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_8_XOR13_U1 ( .A0_t (LED_128_Instance_SBox_Instance_8_L1), .A0_f (new_AGEMA_signal_3957), .A1_t (new_AGEMA_signal_3958), .A1_f (new_AGEMA_signal_3959), .B0_t (LED_128_Instance_SBox_Instance_8_L8), .B0_f (new_AGEMA_signal_4575), .B1_t (new_AGEMA_signal_4576), .B1_f (new_AGEMA_signal_4577), .Z0_t (LED_128_Instance_subcells_out[34]), .Z0_f (new_AGEMA_signal_4689), .Z1_t (new_AGEMA_signal_4690), .Z1_f (new_AGEMA_signal_4691) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_8_XOR14_U1 ( .A0_t (LED_128_Instance_SBox_Instance_8_L4), .A0_f (new_AGEMA_signal_3963), .A1_t (new_AGEMA_signal_3964), .A1_f (new_AGEMA_signal_3965), .B0_t (LED_128_Instance_SBox_Instance_8_T3), .B0_f (new_AGEMA_signal_4572), .B1_t (new_AGEMA_signal_4573), .B1_f (new_AGEMA_signal_4574), .Z0_t (LED_128_Instance_subcells_out[33]), .Z0_f (new_AGEMA_signal_4692), .Z1_t (new_AGEMA_signal_4693), .Z1_f (new_AGEMA_signal_4694) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_8_XOR15_U1 ( .A0_t (LED_128_Instance_SBox_Instance_8_L3), .A0_f (new_AGEMA_signal_3960), .A1_t (new_AGEMA_signal_3961), .A1_f (new_AGEMA_signal_3962), .B0_t (LED_128_Instance_SBox_Instance_8_T2), .B0_f (new_AGEMA_signal_3966), .B1_t (new_AGEMA_signal_3967), .B1_f (new_AGEMA_signal_3968), .Z0_t (LED_128_Instance_subcells_out[32]), .Z0_f (new_AGEMA_signal_4176), .Z1_t (new_AGEMA_signal_4177), .Z1_f (new_AGEMA_signal_4178) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_9_XOR1_U1 ( .A0_t (LED_128_Instance_addconst_out[38]), .A0_f (new_AGEMA_signal_3831), .A1_t (new_AGEMA_signal_3832), .A1_f (new_AGEMA_signal_3833), .B0_t (LED_128_Instance_addconst_out[37]), .B0_f (new_AGEMA_signal_3858), .B1_t (new_AGEMA_signal_3859), .B1_f (new_AGEMA_signal_3860), .Z0_t (LED_128_Instance_SBox_Instance_9_L0), .Z0_f (new_AGEMA_signal_4179), .Z1_t (new_AGEMA_signal_4180), .Z1_f (new_AGEMA_signal_4181) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_9_XOR2_U1 ( .A0_t (LED_128_Instance_addconst_out[37]), .A0_f (new_AGEMA_signal_3858), .A1_t (new_AGEMA_signal_3859), .A1_f (new_AGEMA_signal_3860), .B0_t (LED_128_Instance_addconst_out[36]), .B0_f (new_AGEMA_signal_3840), .B1_t (new_AGEMA_signal_3841), .B1_f (new_AGEMA_signal_3842), .Z0_t (LED_128_Instance_SBox_Instance_9_L1), .Z0_f (new_AGEMA_signal_4182), .Z1_t (new_AGEMA_signal_4183), .Z1_f (new_AGEMA_signal_4184) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_9_XOR3_U1 ( .A0_t (LED_128_Instance_SBox_Instance_9_L1), .A0_f (new_AGEMA_signal_4182), .A1_t (new_AGEMA_signal_4183), .A1_f (new_AGEMA_signal_4184), .B0_t (LED_128_Instance_addconst_out[39]), .B0_f (new_AGEMA_signal_3753), .B1_t (new_AGEMA_signal_3754), .B1_f (new_AGEMA_signal_3755), .Z0_t (LED_128_Instance_SBox_Instance_9_L2), .Z0_f (new_AGEMA_signal_4356), .Z1_t (new_AGEMA_signal_4357), .Z1_f (new_AGEMA_signal_4358) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_SBox_Instance_9_XOR16_U1 ( .A0_t (LED_128_Instance_SBox_Instance_9_T0), .A0_f (new_AGEMA_signal_4365), .A1_t (new_AGEMA_signal_4366), .A1_f (new_AGEMA_signal_4367), .B0_t (LED_128_Instance_SBox_Instance_9_L2), .B0_f (new_AGEMA_signal_4356), .B1_t (new_AGEMA_signal_4357), .B1_f (new_AGEMA_signal_4358), .Z0_t (LED_128_Instance_SBox_Instance_9_Q2), .Z0_f (new_AGEMA_signal_4476), .Z1_t (new_AGEMA_signal_4477), .Z1_f (new_AGEMA_signal_4478) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_9_XOR4_U1 ( .A0_t (LED_128_Instance_addconst_out[39]), .A0_f (new_AGEMA_signal_3753), .A1_t (new_AGEMA_signal_3754), .A1_f (new_AGEMA_signal_3755), .B0_t (LED_128_Instance_addconst_out[36]), .B0_f (new_AGEMA_signal_3840), .B1_t (new_AGEMA_signal_3841), .B1_f (new_AGEMA_signal_3842), .Z0_t (LED_128_Instance_SBox_Instance_9_L3), .Z0_f (new_AGEMA_signal_4185), .Z1_t (new_AGEMA_signal_4186), .Z1_f (new_AGEMA_signal_4187) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_9_XOR5_U1 ( .A0_t (LED_128_Instance_SBox_Instance_9_L3), .A0_f (new_AGEMA_signal_4185), .A1_t (new_AGEMA_signal_4186), .A1_f (new_AGEMA_signal_4187), .B0_t (LED_128_Instance_SBox_Instance_9_L0), .B0_f (new_AGEMA_signal_4179), .B1_t (new_AGEMA_signal_4180), .B1_f (new_AGEMA_signal_4181), .Z0_t (LED_128_Instance_SBox_Instance_9_Q3), .Z0_f (new_AGEMA_signal_4359), .Z1_t (new_AGEMA_signal_4360), .Z1_f (new_AGEMA_signal_4361) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_9_XOR6_U1 ( .A0_t (LED_128_Instance_addconst_out[39]), .A0_f (new_AGEMA_signal_3753), .A1_t (new_AGEMA_signal_3754), .A1_f (new_AGEMA_signal_3755), .B0_t (LED_128_Instance_addconst_out[37]), .B0_f (new_AGEMA_signal_3858), .B1_t (new_AGEMA_signal_3859), .B1_f (new_AGEMA_signal_3860), .Z0_t (LED_128_Instance_SBox_Instance_9_L4), .Z0_f (new_AGEMA_signal_4188), .Z1_t (new_AGEMA_signal_4189), .Z1_f (new_AGEMA_signal_4190) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_9_XOR7_U1 ( .A0_t (LED_128_Instance_SBox_Instance_9_T0), .A0_f (new_AGEMA_signal_4365), .A1_t (new_AGEMA_signal_4366), .A1_f (new_AGEMA_signal_4367), .B0_t (LED_128_Instance_SBox_Instance_9_T2), .B0_f (new_AGEMA_signal_4191), .B1_t (new_AGEMA_signal_4192), .B1_f (new_AGEMA_signal_4193), .Z0_t (LED_128_Instance_SBox_Instance_9_L5), .Z0_f (new_AGEMA_signal_4479), .Z1_t (new_AGEMA_signal_4480), .Z1_f (new_AGEMA_signal_4481) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_SBox_Instance_9_XOR8_U1 ( .A0_t (LED_128_Instance_SBox_Instance_9_L4), .A0_f (new_AGEMA_signal_4188), .A1_t (new_AGEMA_signal_4189), .A1_f (new_AGEMA_signal_4190), .B0_t (LED_128_Instance_SBox_Instance_9_L5), .B0_f (new_AGEMA_signal_4479), .B1_t (new_AGEMA_signal_4480), .B1_f (new_AGEMA_signal_4481), .Z0_t (LED_128_Instance_SBox_Instance_9_Q6), .Z0_f (new_AGEMA_signal_4578), .Z1_t (new_AGEMA_signal_4579), .Z1_f (new_AGEMA_signal_4580) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_9_XOR9_U1 ( .A0_t (LED_128_Instance_SBox_Instance_9_L1), .A0_f (new_AGEMA_signal_4182), .A1_t (new_AGEMA_signal_4183), .A1_f (new_AGEMA_signal_4184), .B0_t (LED_128_Instance_addconst_out[38]), .B0_f (new_AGEMA_signal_3831), .B1_t (new_AGEMA_signal_3832), .B1_f (new_AGEMA_signal_3833), .Z0_t (LED_128_Instance_SBox_Instance_9_Q7), .Z0_f (new_AGEMA_signal_4362), .Z1_t (new_AGEMA_signal_4363), .Z1_f (new_AGEMA_signal_4364) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_9_AND1_U1 ( .A0_t (LED_128_Instance_SBox_Instance_9_L0), .A0_f (new_AGEMA_signal_4179), .A1_t (new_AGEMA_signal_4180), .A1_f (new_AGEMA_signal_4181), .B0_t (LED_128_Instance_addconst_out[39]), .B0_f (new_AGEMA_signal_3753), .B1_t (new_AGEMA_signal_3754), .B1_f (new_AGEMA_signal_3755), .Z0_t (LED_128_Instance_SBox_Instance_9_T0), .Z0_f (new_AGEMA_signal_4365), .Z1_t (new_AGEMA_signal_4366), .Z1_f (new_AGEMA_signal_4367) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_9_AND2_U1 ( .A0_t (LED_128_Instance_SBox_Instance_9_Q2), .A0_f (new_AGEMA_signal_4476), .A1_t (new_AGEMA_signal_4477), .A1_f (new_AGEMA_signal_4478), .B0_t (LED_128_Instance_SBox_Instance_9_Q3), .B0_f (new_AGEMA_signal_4359), .B1_t (new_AGEMA_signal_4360), .B1_f (new_AGEMA_signal_4361), .Z0_t (LED_128_Instance_SBox_Instance_9_T1), .Z0_f (new_AGEMA_signal_4581), .Z1_t (new_AGEMA_signal_4582), .Z1_f (new_AGEMA_signal_4583) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_9_AND3_U1 ( .A0_t (LED_128_Instance_addconst_out[37]), .A0_f (new_AGEMA_signal_3858), .A1_t (new_AGEMA_signal_3859), .A1_f (new_AGEMA_signal_3860), .B0_t (LED_128_Instance_addconst_out[38]), .B0_f (new_AGEMA_signal_3831), .B1_t (new_AGEMA_signal_3832), .B1_f (new_AGEMA_signal_3833), .Z0_t (LED_128_Instance_SBox_Instance_9_T2), .Z0_f (new_AGEMA_signal_4191), .Z1_t (new_AGEMA_signal_4192), .Z1_f (new_AGEMA_signal_4193) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_9_AND4_U1 ( .A0_t (LED_128_Instance_SBox_Instance_9_Q6), .A0_f (new_AGEMA_signal_4578), .A1_t (new_AGEMA_signal_4579), .A1_f (new_AGEMA_signal_4580), .B0_t (LED_128_Instance_SBox_Instance_9_Q7), .B0_f (new_AGEMA_signal_4362), .B1_t (new_AGEMA_signal_4363), .B1_f (new_AGEMA_signal_4364), .Z0_t (LED_128_Instance_SBox_Instance_9_T3), .Z0_f (new_AGEMA_signal_4695), .Z1_t (new_AGEMA_signal_4696), .Z1_f (new_AGEMA_signal_4697) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_9_XOR10_U1 ( .A0_t (LED_128_Instance_SBox_Instance_9_L5), .A0_f (new_AGEMA_signal_4479), .A1_t (new_AGEMA_signal_4480), .A1_f (new_AGEMA_signal_4481), .B0_t (LED_128_Instance_SBox_Instance_9_T3), .B0_f (new_AGEMA_signal_4695), .B1_t (new_AGEMA_signal_4696), .B1_f (new_AGEMA_signal_4697), .Z0_t (LED_128_Instance_SBox_Instance_9_L7), .Z0_f (new_AGEMA_signal_4791), .Z1_t (new_AGEMA_signal_4792), .Z1_f (new_AGEMA_signal_4793) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_9_XOR11_U1 ( .A0_t (LED_128_Instance_addconst_out[36]), .A0_f (new_AGEMA_signal_3840), .A1_t (new_AGEMA_signal_3841), .A1_f (new_AGEMA_signal_3842), .B0_t (LED_128_Instance_SBox_Instance_9_L7), .B0_f (new_AGEMA_signal_4791), .B1_t (new_AGEMA_signal_4792), .B1_f (new_AGEMA_signal_4793), .Z0_t (LED_128_Instance_subcells_out[39]), .Z0_f (new_AGEMA_signal_4893), .Z1_t (new_AGEMA_signal_4894), .Z1_f (new_AGEMA_signal_4895) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_9_XOR12_U1 ( .A0_t (LED_128_Instance_SBox_Instance_9_L5), .A0_f (new_AGEMA_signal_4479), .A1_t (new_AGEMA_signal_4480), .A1_f (new_AGEMA_signal_4481), .B0_t (LED_128_Instance_SBox_Instance_9_T1), .B0_f (new_AGEMA_signal_4581), .B1_t (new_AGEMA_signal_4582), .B1_f (new_AGEMA_signal_4583), .Z0_t (LED_128_Instance_SBox_Instance_9_L8), .Z0_f (new_AGEMA_signal_4698), .Z1_t (new_AGEMA_signal_4699), .Z1_f (new_AGEMA_signal_4700) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_9_XOR13_U1 ( .A0_t (LED_128_Instance_SBox_Instance_9_L1), .A0_f (new_AGEMA_signal_4182), .A1_t (new_AGEMA_signal_4183), .A1_f (new_AGEMA_signal_4184), .B0_t (LED_128_Instance_SBox_Instance_9_L8), .B0_f (new_AGEMA_signal_4698), .B1_t (new_AGEMA_signal_4699), .B1_f (new_AGEMA_signal_4700), .Z0_t (LED_128_Instance_subcells_out[38]), .Z0_f (new_AGEMA_signal_4794), .Z1_t (new_AGEMA_signal_4795), .Z1_f (new_AGEMA_signal_4796) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_9_XOR14_U1 ( .A0_t (LED_128_Instance_SBox_Instance_9_L4), .A0_f (new_AGEMA_signal_4188), .A1_t (new_AGEMA_signal_4189), .A1_f (new_AGEMA_signal_4190), .B0_t (LED_128_Instance_SBox_Instance_9_T3), .B0_f (new_AGEMA_signal_4695), .B1_t (new_AGEMA_signal_4696), .B1_f (new_AGEMA_signal_4697), .Z0_t (LED_128_Instance_subcells_out[37]), .Z0_f (new_AGEMA_signal_4797), .Z1_t (new_AGEMA_signal_4798), .Z1_f (new_AGEMA_signal_4799) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_9_XOR15_U1 ( .A0_t (LED_128_Instance_SBox_Instance_9_L3), .A0_f (new_AGEMA_signal_4185), .A1_t (new_AGEMA_signal_4186), .A1_f (new_AGEMA_signal_4187), .B0_t (LED_128_Instance_SBox_Instance_9_T2), .B0_f (new_AGEMA_signal_4191), .B1_t (new_AGEMA_signal_4192), .B1_f (new_AGEMA_signal_4193), .Z0_t (LED_128_Instance_subcells_out[36]), .Z0_f (new_AGEMA_signal_4368), .Z1_t (new_AGEMA_signal_4369), .Z1_f (new_AGEMA_signal_4370) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_10_XOR1_U1 ( .A0_t (LED_128_Instance_addconst_out[42]), .A0_f (new_AGEMA_signal_3762), .A1_t (new_AGEMA_signal_3763), .A1_f (new_AGEMA_signal_3764), .B0_t (LED_128_Instance_addconst_out[41]), .B0_f (new_AGEMA_signal_3759), .B1_t (new_AGEMA_signal_3760), .B1_f (new_AGEMA_signal_3761), .Z0_t (LED_128_Instance_SBox_Instance_10_L0), .Z0_f (new_AGEMA_signal_3969), .Z1_t (new_AGEMA_signal_3970), .Z1_f (new_AGEMA_signal_3971) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_10_XOR2_U1 ( .A0_t (LED_128_Instance_addconst_out[41]), .A0_f (new_AGEMA_signal_3759), .A1_t (new_AGEMA_signal_3760), .A1_f (new_AGEMA_signal_3761), .B0_t (LED_128_Instance_addconst_out[40]), .B0_f (new_AGEMA_signal_3756), .B1_t (new_AGEMA_signal_3757), .B1_f (new_AGEMA_signal_3758), .Z0_t (LED_128_Instance_SBox_Instance_10_L1), .Z0_f (new_AGEMA_signal_3972), .Z1_t (new_AGEMA_signal_3973), .Z1_f (new_AGEMA_signal_3974) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_10_XOR3_U1 ( .A0_t (LED_128_Instance_SBox_Instance_10_L1), .A0_f (new_AGEMA_signal_3972), .A1_t (new_AGEMA_signal_3973), .A1_f (new_AGEMA_signal_3974), .B0_t (LED_128_Instance_addconst_out[43]), .B0_f (new_AGEMA_signal_3765), .B1_t (new_AGEMA_signal_3766), .B1_f (new_AGEMA_signal_3767), .Z0_t (LED_128_Instance_SBox_Instance_10_L2), .Z0_f (new_AGEMA_signal_4194), .Z1_t (new_AGEMA_signal_4195), .Z1_f (new_AGEMA_signal_4196) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_SBox_Instance_10_XOR16_U1 ( .A0_t (LED_128_Instance_SBox_Instance_10_T0), .A0_f (new_AGEMA_signal_4203), .A1_t (new_AGEMA_signal_4204), .A1_f (new_AGEMA_signal_4205), .B0_t (LED_128_Instance_SBox_Instance_10_L2), .B0_f (new_AGEMA_signal_4194), .B1_t (new_AGEMA_signal_4195), .B1_f (new_AGEMA_signal_4196), .Z0_t (LED_128_Instance_SBox_Instance_10_Q2), .Z0_f (new_AGEMA_signal_4371), .Z1_t (new_AGEMA_signal_4372), .Z1_f (new_AGEMA_signal_4373) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_10_XOR4_U1 ( .A0_t (LED_128_Instance_addconst_out[43]), .A0_f (new_AGEMA_signal_3765), .A1_t (new_AGEMA_signal_3766), .A1_f (new_AGEMA_signal_3767), .B0_t (LED_128_Instance_addconst_out[40]), .B0_f (new_AGEMA_signal_3756), .B1_t (new_AGEMA_signal_3757), .B1_f (new_AGEMA_signal_3758), .Z0_t (LED_128_Instance_SBox_Instance_10_L3), .Z0_f (new_AGEMA_signal_3975), .Z1_t (new_AGEMA_signal_3976), .Z1_f (new_AGEMA_signal_3977) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_10_XOR5_U1 ( .A0_t (LED_128_Instance_SBox_Instance_10_L3), .A0_f (new_AGEMA_signal_3975), .A1_t (new_AGEMA_signal_3976), .A1_f (new_AGEMA_signal_3977), .B0_t (LED_128_Instance_SBox_Instance_10_L0), .B0_f (new_AGEMA_signal_3969), .B1_t (new_AGEMA_signal_3970), .B1_f (new_AGEMA_signal_3971), .Z0_t (LED_128_Instance_SBox_Instance_10_Q3), .Z0_f (new_AGEMA_signal_4197), .Z1_t (new_AGEMA_signal_4198), .Z1_f (new_AGEMA_signal_4199) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_10_XOR6_U1 ( .A0_t (LED_128_Instance_addconst_out[43]), .A0_f (new_AGEMA_signal_3765), .A1_t (new_AGEMA_signal_3766), .A1_f (new_AGEMA_signal_3767), .B0_t (LED_128_Instance_addconst_out[41]), .B0_f (new_AGEMA_signal_3759), .B1_t (new_AGEMA_signal_3760), .B1_f (new_AGEMA_signal_3761), .Z0_t (LED_128_Instance_SBox_Instance_10_L4), .Z0_f (new_AGEMA_signal_3978), .Z1_t (new_AGEMA_signal_3979), .Z1_f (new_AGEMA_signal_3980) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_10_XOR7_U1 ( .A0_t (LED_128_Instance_SBox_Instance_10_T0), .A0_f (new_AGEMA_signal_4203), .A1_t (new_AGEMA_signal_4204), .A1_f (new_AGEMA_signal_4205), .B0_t (LED_128_Instance_SBox_Instance_10_T2), .B0_f (new_AGEMA_signal_3981), .B1_t (new_AGEMA_signal_3982), .B1_f (new_AGEMA_signal_3983), .Z0_t (LED_128_Instance_SBox_Instance_10_L5), .Z0_f (new_AGEMA_signal_4374), .Z1_t (new_AGEMA_signal_4375), .Z1_f (new_AGEMA_signal_4376) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_SBox_Instance_10_XOR8_U1 ( .A0_t (LED_128_Instance_SBox_Instance_10_L4), .A0_f (new_AGEMA_signal_3978), .A1_t (new_AGEMA_signal_3979), .A1_f (new_AGEMA_signal_3980), .B0_t (LED_128_Instance_SBox_Instance_10_L5), .B0_f (new_AGEMA_signal_4374), .B1_t (new_AGEMA_signal_4375), .B1_f (new_AGEMA_signal_4376), .Z0_t (LED_128_Instance_SBox_Instance_10_Q6), .Z0_f (new_AGEMA_signal_4482), .Z1_t (new_AGEMA_signal_4483), .Z1_f (new_AGEMA_signal_4484) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_10_XOR9_U1 ( .A0_t (LED_128_Instance_SBox_Instance_10_L1), .A0_f (new_AGEMA_signal_3972), .A1_t (new_AGEMA_signal_3973), .A1_f (new_AGEMA_signal_3974), .B0_t (LED_128_Instance_addconst_out[42]), .B0_f (new_AGEMA_signal_3762), .B1_t (new_AGEMA_signal_3763), .B1_f (new_AGEMA_signal_3764), .Z0_t (LED_128_Instance_SBox_Instance_10_Q7), .Z0_f (new_AGEMA_signal_4200), .Z1_t (new_AGEMA_signal_4201), .Z1_f (new_AGEMA_signal_4202) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_10_AND1_U1 ( .A0_t (LED_128_Instance_SBox_Instance_10_L0), .A0_f (new_AGEMA_signal_3969), .A1_t (new_AGEMA_signal_3970), .A1_f (new_AGEMA_signal_3971), .B0_t (LED_128_Instance_addconst_out[43]), .B0_f (new_AGEMA_signal_3765), .B1_t (new_AGEMA_signal_3766), .B1_f (new_AGEMA_signal_3767), .Z0_t (LED_128_Instance_SBox_Instance_10_T0), .Z0_f (new_AGEMA_signal_4203), .Z1_t (new_AGEMA_signal_4204), .Z1_f (new_AGEMA_signal_4205) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_10_AND2_U1 ( .A0_t (LED_128_Instance_SBox_Instance_10_Q2), .A0_f (new_AGEMA_signal_4371), .A1_t (new_AGEMA_signal_4372), .A1_f (new_AGEMA_signal_4373), .B0_t (LED_128_Instance_SBox_Instance_10_Q3), .B0_f (new_AGEMA_signal_4197), .B1_t (new_AGEMA_signal_4198), .B1_f (new_AGEMA_signal_4199), .Z0_t (LED_128_Instance_SBox_Instance_10_T1), .Z0_f (new_AGEMA_signal_4485), .Z1_t (new_AGEMA_signal_4486), .Z1_f (new_AGEMA_signal_4487) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_10_AND3_U1 ( .A0_t (LED_128_Instance_addconst_out[41]), .A0_f (new_AGEMA_signal_3759), .A1_t (new_AGEMA_signal_3760), .A1_f (new_AGEMA_signal_3761), .B0_t (LED_128_Instance_addconst_out[42]), .B0_f (new_AGEMA_signal_3762), .B1_t (new_AGEMA_signal_3763), .B1_f (new_AGEMA_signal_3764), .Z0_t (LED_128_Instance_SBox_Instance_10_T2), .Z0_f (new_AGEMA_signal_3981), .Z1_t (new_AGEMA_signal_3982), .Z1_f (new_AGEMA_signal_3983) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_10_AND4_U1 ( .A0_t (LED_128_Instance_SBox_Instance_10_Q6), .A0_f (new_AGEMA_signal_4482), .A1_t (new_AGEMA_signal_4483), .A1_f (new_AGEMA_signal_4484), .B0_t (LED_128_Instance_SBox_Instance_10_Q7), .B0_f (new_AGEMA_signal_4200), .B1_t (new_AGEMA_signal_4201), .B1_f (new_AGEMA_signal_4202), .Z0_t (LED_128_Instance_SBox_Instance_10_T3), .Z0_f (new_AGEMA_signal_4584), .Z1_t (new_AGEMA_signal_4585), .Z1_f (new_AGEMA_signal_4586) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_10_XOR10_U1 ( .A0_t (LED_128_Instance_SBox_Instance_10_L5), .A0_f (new_AGEMA_signal_4374), .A1_t (new_AGEMA_signal_4375), .A1_f (new_AGEMA_signal_4376), .B0_t (LED_128_Instance_SBox_Instance_10_T3), .B0_f (new_AGEMA_signal_4584), .B1_t (new_AGEMA_signal_4585), .B1_f (new_AGEMA_signal_4586), .Z0_t (LED_128_Instance_SBox_Instance_10_L7), .Z0_f (new_AGEMA_signal_4701), .Z1_t (new_AGEMA_signal_4702), .Z1_f (new_AGEMA_signal_4703) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_10_XOR11_U1 ( .A0_t (LED_128_Instance_addconst_out[40]), .A0_f (new_AGEMA_signal_3756), .A1_t (new_AGEMA_signal_3757), .A1_f (new_AGEMA_signal_3758), .B0_t (LED_128_Instance_SBox_Instance_10_L7), .B0_f (new_AGEMA_signal_4701), .B1_t (new_AGEMA_signal_4702), .B1_f (new_AGEMA_signal_4703), .Z0_t (LED_128_Instance_subcells_out[43]), .Z0_f (new_AGEMA_signal_4800), .Z1_t (new_AGEMA_signal_4801), .Z1_f (new_AGEMA_signal_4802) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_10_XOR12_U1 ( .A0_t (LED_128_Instance_SBox_Instance_10_L5), .A0_f (new_AGEMA_signal_4374), .A1_t (new_AGEMA_signal_4375), .A1_f (new_AGEMA_signal_4376), .B0_t (LED_128_Instance_SBox_Instance_10_T1), .B0_f (new_AGEMA_signal_4485), .B1_t (new_AGEMA_signal_4486), .B1_f (new_AGEMA_signal_4487), .Z0_t (LED_128_Instance_SBox_Instance_10_L8), .Z0_f (new_AGEMA_signal_4587), .Z1_t (new_AGEMA_signal_4588), .Z1_f (new_AGEMA_signal_4589) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_10_XOR13_U1 ( .A0_t (LED_128_Instance_SBox_Instance_10_L1), .A0_f (new_AGEMA_signal_3972), .A1_t (new_AGEMA_signal_3973), .A1_f (new_AGEMA_signal_3974), .B0_t (LED_128_Instance_SBox_Instance_10_L8), .B0_f (new_AGEMA_signal_4587), .B1_t (new_AGEMA_signal_4588), .B1_f (new_AGEMA_signal_4589), .Z0_t (LED_128_Instance_subcells_out[42]), .Z0_f (new_AGEMA_signal_4704), .Z1_t (new_AGEMA_signal_4705), .Z1_f (new_AGEMA_signal_4706) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_10_XOR14_U1 ( .A0_t (LED_128_Instance_SBox_Instance_10_L4), .A0_f (new_AGEMA_signal_3978), .A1_t (new_AGEMA_signal_3979), .A1_f (new_AGEMA_signal_3980), .B0_t (LED_128_Instance_SBox_Instance_10_T3), .B0_f (new_AGEMA_signal_4584), .B1_t (new_AGEMA_signal_4585), .B1_f (new_AGEMA_signal_4586), .Z0_t (LED_128_Instance_subcells_out[41]), .Z0_f (new_AGEMA_signal_4707), .Z1_t (new_AGEMA_signal_4708), .Z1_f (new_AGEMA_signal_4709) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_10_XOR15_U1 ( .A0_t (LED_128_Instance_SBox_Instance_10_L3), .A0_f (new_AGEMA_signal_3975), .A1_t (new_AGEMA_signal_3976), .A1_f (new_AGEMA_signal_3977), .B0_t (LED_128_Instance_SBox_Instance_10_T2), .B0_f (new_AGEMA_signal_3981), .B1_t (new_AGEMA_signal_3982), .B1_f (new_AGEMA_signal_3983), .Z0_t (LED_128_Instance_subcells_out[40]), .Z0_f (new_AGEMA_signal_4206), .Z1_t (new_AGEMA_signal_4207), .Z1_f (new_AGEMA_signal_4208) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_11_XOR1_U1 ( .A0_t (LED_128_Instance_addconst_out[46]), .A0_f (new_AGEMA_signal_3774), .A1_t (new_AGEMA_signal_3775), .A1_f (new_AGEMA_signal_3776), .B0_t (LED_128_Instance_addconst_out[45]), .B0_f (new_AGEMA_signal_3771), .B1_t (new_AGEMA_signal_3772), .B1_f (new_AGEMA_signal_3773), .Z0_t (LED_128_Instance_SBox_Instance_11_L0), .Z0_f (new_AGEMA_signal_3984), .Z1_t (new_AGEMA_signal_3985), .Z1_f (new_AGEMA_signal_3986) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_11_XOR2_U1 ( .A0_t (LED_128_Instance_addconst_out[45]), .A0_f (new_AGEMA_signal_3771), .A1_t (new_AGEMA_signal_3772), .A1_f (new_AGEMA_signal_3773), .B0_t (LED_128_Instance_addconst_out[44]), .B0_f (new_AGEMA_signal_3768), .B1_t (new_AGEMA_signal_3769), .B1_f (new_AGEMA_signal_3770), .Z0_t (LED_128_Instance_SBox_Instance_11_L1), .Z0_f (new_AGEMA_signal_3987), .Z1_t (new_AGEMA_signal_3988), .Z1_f (new_AGEMA_signal_3989) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_11_XOR3_U1 ( .A0_t (LED_128_Instance_SBox_Instance_11_L1), .A0_f (new_AGEMA_signal_3987), .A1_t (new_AGEMA_signal_3988), .A1_f (new_AGEMA_signal_3989), .B0_t (LED_128_Instance_addconst_out[47]), .B0_f (new_AGEMA_signal_3777), .B1_t (new_AGEMA_signal_3778), .B1_f (new_AGEMA_signal_3779), .Z0_t (LED_128_Instance_SBox_Instance_11_L2), .Z0_f (new_AGEMA_signal_4209), .Z1_t (new_AGEMA_signal_4210), .Z1_f (new_AGEMA_signal_4211) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_SBox_Instance_11_XOR16_U1 ( .A0_t (LED_128_Instance_SBox_Instance_11_T0), .A0_f (new_AGEMA_signal_4218), .A1_t (new_AGEMA_signal_4219), .A1_f (new_AGEMA_signal_4220), .B0_t (LED_128_Instance_SBox_Instance_11_L2), .B0_f (new_AGEMA_signal_4209), .B1_t (new_AGEMA_signal_4210), .B1_f (new_AGEMA_signal_4211), .Z0_t (LED_128_Instance_SBox_Instance_11_Q2), .Z0_f (new_AGEMA_signal_4377), .Z1_t (new_AGEMA_signal_4378), .Z1_f (new_AGEMA_signal_4379) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_11_XOR4_U1 ( .A0_t (LED_128_Instance_addconst_out[47]), .A0_f (new_AGEMA_signal_3777), .A1_t (new_AGEMA_signal_3778), .A1_f (new_AGEMA_signal_3779), .B0_t (LED_128_Instance_addconst_out[44]), .B0_f (new_AGEMA_signal_3768), .B1_t (new_AGEMA_signal_3769), .B1_f (new_AGEMA_signal_3770), .Z0_t (LED_128_Instance_SBox_Instance_11_L3), .Z0_f (new_AGEMA_signal_3990), .Z1_t (new_AGEMA_signal_3991), .Z1_f (new_AGEMA_signal_3992) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_11_XOR5_U1 ( .A0_t (LED_128_Instance_SBox_Instance_11_L3), .A0_f (new_AGEMA_signal_3990), .A1_t (new_AGEMA_signal_3991), .A1_f (new_AGEMA_signal_3992), .B0_t (LED_128_Instance_SBox_Instance_11_L0), .B0_f (new_AGEMA_signal_3984), .B1_t (new_AGEMA_signal_3985), .B1_f (new_AGEMA_signal_3986), .Z0_t (LED_128_Instance_SBox_Instance_11_Q3), .Z0_f (new_AGEMA_signal_4212), .Z1_t (new_AGEMA_signal_4213), .Z1_f (new_AGEMA_signal_4214) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_11_XOR6_U1 ( .A0_t (LED_128_Instance_addconst_out[47]), .A0_f (new_AGEMA_signal_3777), .A1_t (new_AGEMA_signal_3778), .A1_f (new_AGEMA_signal_3779), .B0_t (LED_128_Instance_addconst_out[45]), .B0_f (new_AGEMA_signal_3771), .B1_t (new_AGEMA_signal_3772), .B1_f (new_AGEMA_signal_3773), .Z0_t (LED_128_Instance_SBox_Instance_11_L4), .Z0_f (new_AGEMA_signal_3993), .Z1_t (new_AGEMA_signal_3994), .Z1_f (new_AGEMA_signal_3995) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_11_XOR7_U1 ( .A0_t (LED_128_Instance_SBox_Instance_11_T0), .A0_f (new_AGEMA_signal_4218), .A1_t (new_AGEMA_signal_4219), .A1_f (new_AGEMA_signal_4220), .B0_t (LED_128_Instance_SBox_Instance_11_T2), .B0_f (new_AGEMA_signal_3996), .B1_t (new_AGEMA_signal_3997), .B1_f (new_AGEMA_signal_3998), .Z0_t (LED_128_Instance_SBox_Instance_11_L5), .Z0_f (new_AGEMA_signal_4380), .Z1_t (new_AGEMA_signal_4381), .Z1_f (new_AGEMA_signal_4382) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_SBox_Instance_11_XOR8_U1 ( .A0_t (LED_128_Instance_SBox_Instance_11_L4), .A0_f (new_AGEMA_signal_3993), .A1_t (new_AGEMA_signal_3994), .A1_f (new_AGEMA_signal_3995), .B0_t (LED_128_Instance_SBox_Instance_11_L5), .B0_f (new_AGEMA_signal_4380), .B1_t (new_AGEMA_signal_4381), .B1_f (new_AGEMA_signal_4382), .Z0_t (LED_128_Instance_SBox_Instance_11_Q6), .Z0_f (new_AGEMA_signal_4488), .Z1_t (new_AGEMA_signal_4489), .Z1_f (new_AGEMA_signal_4490) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_11_XOR9_U1 ( .A0_t (LED_128_Instance_SBox_Instance_11_L1), .A0_f (new_AGEMA_signal_3987), .A1_t (new_AGEMA_signal_3988), .A1_f (new_AGEMA_signal_3989), .B0_t (LED_128_Instance_addconst_out[46]), .B0_f (new_AGEMA_signal_3774), .B1_t (new_AGEMA_signal_3775), .B1_f (new_AGEMA_signal_3776), .Z0_t (LED_128_Instance_SBox_Instance_11_Q7), .Z0_f (new_AGEMA_signal_4215), .Z1_t (new_AGEMA_signal_4216), .Z1_f (new_AGEMA_signal_4217) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_11_AND1_U1 ( .A0_t (LED_128_Instance_SBox_Instance_11_L0), .A0_f (new_AGEMA_signal_3984), .A1_t (new_AGEMA_signal_3985), .A1_f (new_AGEMA_signal_3986), .B0_t (LED_128_Instance_addconst_out[47]), .B0_f (new_AGEMA_signal_3777), .B1_t (new_AGEMA_signal_3778), .B1_f (new_AGEMA_signal_3779), .Z0_t (LED_128_Instance_SBox_Instance_11_T0), .Z0_f (new_AGEMA_signal_4218), .Z1_t (new_AGEMA_signal_4219), .Z1_f (new_AGEMA_signal_4220) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_11_AND2_U1 ( .A0_t (LED_128_Instance_SBox_Instance_11_Q2), .A0_f (new_AGEMA_signal_4377), .A1_t (new_AGEMA_signal_4378), .A1_f (new_AGEMA_signal_4379), .B0_t (LED_128_Instance_SBox_Instance_11_Q3), .B0_f (new_AGEMA_signal_4212), .B1_t (new_AGEMA_signal_4213), .B1_f (new_AGEMA_signal_4214), .Z0_t (LED_128_Instance_SBox_Instance_11_T1), .Z0_f (new_AGEMA_signal_4491), .Z1_t (new_AGEMA_signal_4492), .Z1_f (new_AGEMA_signal_4493) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_11_AND3_U1 ( .A0_t (LED_128_Instance_addconst_out[45]), .A0_f (new_AGEMA_signal_3771), .A1_t (new_AGEMA_signal_3772), .A1_f (new_AGEMA_signal_3773), .B0_t (LED_128_Instance_addconst_out[46]), .B0_f (new_AGEMA_signal_3774), .B1_t (new_AGEMA_signal_3775), .B1_f (new_AGEMA_signal_3776), .Z0_t (LED_128_Instance_SBox_Instance_11_T2), .Z0_f (new_AGEMA_signal_3996), .Z1_t (new_AGEMA_signal_3997), .Z1_f (new_AGEMA_signal_3998) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_11_AND4_U1 ( .A0_t (LED_128_Instance_SBox_Instance_11_Q6), .A0_f (new_AGEMA_signal_4488), .A1_t (new_AGEMA_signal_4489), .A1_f (new_AGEMA_signal_4490), .B0_t (LED_128_Instance_SBox_Instance_11_Q7), .B0_f (new_AGEMA_signal_4215), .B1_t (new_AGEMA_signal_4216), .B1_f (new_AGEMA_signal_4217), .Z0_t (LED_128_Instance_SBox_Instance_11_T3), .Z0_f (new_AGEMA_signal_4590), .Z1_t (new_AGEMA_signal_4591), .Z1_f (new_AGEMA_signal_4592) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_11_XOR10_U1 ( .A0_t (LED_128_Instance_SBox_Instance_11_L5), .A0_f (new_AGEMA_signal_4380), .A1_t (new_AGEMA_signal_4381), .A1_f (new_AGEMA_signal_4382), .B0_t (LED_128_Instance_SBox_Instance_11_T3), .B0_f (new_AGEMA_signal_4590), .B1_t (new_AGEMA_signal_4591), .B1_f (new_AGEMA_signal_4592), .Z0_t (LED_128_Instance_SBox_Instance_11_L7), .Z0_f (new_AGEMA_signal_4710), .Z1_t (new_AGEMA_signal_4711), .Z1_f (new_AGEMA_signal_4712) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_11_XOR11_U1 ( .A0_t (LED_128_Instance_addconst_out[44]), .A0_f (new_AGEMA_signal_3768), .A1_t (new_AGEMA_signal_3769), .A1_f (new_AGEMA_signal_3770), .B0_t (LED_128_Instance_SBox_Instance_11_L7), .B0_f (new_AGEMA_signal_4710), .B1_t (new_AGEMA_signal_4711), .B1_f (new_AGEMA_signal_4712), .Z0_t (LED_128_Instance_subcells_out[47]), .Z0_f (new_AGEMA_signal_4803), .Z1_t (new_AGEMA_signal_4804), .Z1_f (new_AGEMA_signal_4805) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_11_XOR12_U1 ( .A0_t (LED_128_Instance_SBox_Instance_11_L5), .A0_f (new_AGEMA_signal_4380), .A1_t (new_AGEMA_signal_4381), .A1_f (new_AGEMA_signal_4382), .B0_t (LED_128_Instance_SBox_Instance_11_T1), .B0_f (new_AGEMA_signal_4491), .B1_t (new_AGEMA_signal_4492), .B1_f (new_AGEMA_signal_4493), .Z0_t (LED_128_Instance_SBox_Instance_11_L8), .Z0_f (new_AGEMA_signal_4593), .Z1_t (new_AGEMA_signal_4594), .Z1_f (new_AGEMA_signal_4595) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_11_XOR13_U1 ( .A0_t (LED_128_Instance_SBox_Instance_11_L1), .A0_f (new_AGEMA_signal_3987), .A1_t (new_AGEMA_signal_3988), .A1_f (new_AGEMA_signal_3989), .B0_t (LED_128_Instance_SBox_Instance_11_L8), .B0_f (new_AGEMA_signal_4593), .B1_t (new_AGEMA_signal_4594), .B1_f (new_AGEMA_signal_4595), .Z0_t (LED_128_Instance_subcells_out[46]), .Z0_f (new_AGEMA_signal_4713), .Z1_t (new_AGEMA_signal_4714), .Z1_f (new_AGEMA_signal_4715) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_11_XOR14_U1 ( .A0_t (LED_128_Instance_SBox_Instance_11_L4), .A0_f (new_AGEMA_signal_3993), .A1_t (new_AGEMA_signal_3994), .A1_f (new_AGEMA_signal_3995), .B0_t (LED_128_Instance_SBox_Instance_11_T3), .B0_f (new_AGEMA_signal_4590), .B1_t (new_AGEMA_signal_4591), .B1_f (new_AGEMA_signal_4592), .Z0_t (LED_128_Instance_subcells_out[45]), .Z0_f (new_AGEMA_signal_4716), .Z1_t (new_AGEMA_signal_4717), .Z1_f (new_AGEMA_signal_4718) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_11_XOR15_U1 ( .A0_t (LED_128_Instance_SBox_Instance_11_L3), .A0_f (new_AGEMA_signal_3990), .A1_t (new_AGEMA_signal_3991), .A1_f (new_AGEMA_signal_3992), .B0_t (LED_128_Instance_SBox_Instance_11_T2), .B0_f (new_AGEMA_signal_3996), .B1_t (new_AGEMA_signal_3997), .B1_f (new_AGEMA_signal_3998), .Z0_t (LED_128_Instance_subcells_out[44]), .Z0_f (new_AGEMA_signal_4221), .Z1_t (new_AGEMA_signal_4222), .Z1_f (new_AGEMA_signal_4223) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_12_XOR1_U1 ( .A0_t (LED_128_Instance_addconst_out[50]), .A0_f (new_AGEMA_signal_3786), .A1_t (new_AGEMA_signal_3787), .A1_f (new_AGEMA_signal_3788), .B0_t (LED_128_Instance_addroundkey_out[49]), .B0_f (new_AGEMA_signal_3783), .B1_t (new_AGEMA_signal_3784), .B1_f (new_AGEMA_signal_3785), .Z0_t (LED_128_Instance_SBox_Instance_12_L0), .Z0_f (new_AGEMA_signal_3999), .Z1_t (new_AGEMA_signal_4000), .Z1_f (new_AGEMA_signal_4001) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_12_XOR2_U1 ( .A0_t (LED_128_Instance_addroundkey_out[49]), .A0_f (new_AGEMA_signal_3783), .A1_t (new_AGEMA_signal_3784), .A1_f (new_AGEMA_signal_3785), .B0_t (LED_128_Instance_addroundkey_out[48]), .B0_f (new_AGEMA_signal_3780), .B1_t (new_AGEMA_signal_3781), .B1_f (new_AGEMA_signal_3782), .Z0_t (LED_128_Instance_SBox_Instance_12_L1), .Z0_f (new_AGEMA_signal_4002), .Z1_t (new_AGEMA_signal_4003), .Z1_f (new_AGEMA_signal_4004) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_12_XOR3_U1 ( .A0_t (LED_128_Instance_SBox_Instance_12_L1), .A0_f (new_AGEMA_signal_4002), .A1_t (new_AGEMA_signal_4003), .A1_f (new_AGEMA_signal_4004), .B0_t (LED_128_Instance_addconst_out[51]), .B0_f (new_AGEMA_signal_3789), .B1_t (new_AGEMA_signal_3790), .B1_f (new_AGEMA_signal_3791), .Z0_t (LED_128_Instance_SBox_Instance_12_L2), .Z0_f (new_AGEMA_signal_4224), .Z1_t (new_AGEMA_signal_4225), .Z1_f (new_AGEMA_signal_4226) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_SBox_Instance_12_XOR16_U1 ( .A0_t (LED_128_Instance_SBox_Instance_12_T0), .A0_f (new_AGEMA_signal_4233), .A1_t (new_AGEMA_signal_4234), .A1_f (new_AGEMA_signal_4235), .B0_t (LED_128_Instance_SBox_Instance_12_L2), .B0_f (new_AGEMA_signal_4224), .B1_t (new_AGEMA_signal_4225), .B1_f (new_AGEMA_signal_4226), .Z0_t (LED_128_Instance_SBox_Instance_12_Q2), .Z0_f (new_AGEMA_signal_4383), .Z1_t (new_AGEMA_signal_4384), .Z1_f (new_AGEMA_signal_4385) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_12_XOR4_U1 ( .A0_t (LED_128_Instance_addconst_out[51]), .A0_f (new_AGEMA_signal_3789), .A1_t (new_AGEMA_signal_3790), .A1_f (new_AGEMA_signal_3791), .B0_t (LED_128_Instance_addroundkey_out[48]), .B0_f (new_AGEMA_signal_3780), .B1_t (new_AGEMA_signal_3781), .B1_f (new_AGEMA_signal_3782), .Z0_t (LED_128_Instance_SBox_Instance_12_L3), .Z0_f (new_AGEMA_signal_4005), .Z1_t (new_AGEMA_signal_4006), .Z1_f (new_AGEMA_signal_4007) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_12_XOR5_U1 ( .A0_t (LED_128_Instance_SBox_Instance_12_L3), .A0_f (new_AGEMA_signal_4005), .A1_t (new_AGEMA_signal_4006), .A1_f (new_AGEMA_signal_4007), .B0_t (LED_128_Instance_SBox_Instance_12_L0), .B0_f (new_AGEMA_signal_3999), .B1_t (new_AGEMA_signal_4000), .B1_f (new_AGEMA_signal_4001), .Z0_t (LED_128_Instance_SBox_Instance_12_Q3), .Z0_f (new_AGEMA_signal_4227), .Z1_t (new_AGEMA_signal_4228), .Z1_f (new_AGEMA_signal_4229) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_12_XOR6_U1 ( .A0_t (LED_128_Instance_addconst_out[51]), .A0_f (new_AGEMA_signal_3789), .A1_t (new_AGEMA_signal_3790), .A1_f (new_AGEMA_signal_3791), .B0_t (LED_128_Instance_addroundkey_out[49]), .B0_f (new_AGEMA_signal_3783), .B1_t (new_AGEMA_signal_3784), .B1_f (new_AGEMA_signal_3785), .Z0_t (LED_128_Instance_SBox_Instance_12_L4), .Z0_f (new_AGEMA_signal_4008), .Z1_t (new_AGEMA_signal_4009), .Z1_f (new_AGEMA_signal_4010) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_12_XOR7_U1 ( .A0_t (LED_128_Instance_SBox_Instance_12_T0), .A0_f (new_AGEMA_signal_4233), .A1_t (new_AGEMA_signal_4234), .A1_f (new_AGEMA_signal_4235), .B0_t (LED_128_Instance_SBox_Instance_12_T2), .B0_f (new_AGEMA_signal_4011), .B1_t (new_AGEMA_signal_4012), .B1_f (new_AGEMA_signal_4013), .Z0_t (LED_128_Instance_SBox_Instance_12_L5), .Z0_f (new_AGEMA_signal_4386), .Z1_t (new_AGEMA_signal_4387), .Z1_f (new_AGEMA_signal_4388) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_SBox_Instance_12_XOR8_U1 ( .A0_t (LED_128_Instance_SBox_Instance_12_L4), .A0_f (new_AGEMA_signal_4008), .A1_t (new_AGEMA_signal_4009), .A1_f (new_AGEMA_signal_4010), .B0_t (LED_128_Instance_SBox_Instance_12_L5), .B0_f (new_AGEMA_signal_4386), .B1_t (new_AGEMA_signal_4387), .B1_f (new_AGEMA_signal_4388), .Z0_t (LED_128_Instance_SBox_Instance_12_Q6), .Z0_f (new_AGEMA_signal_4494), .Z1_t (new_AGEMA_signal_4495), .Z1_f (new_AGEMA_signal_4496) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_12_XOR9_U1 ( .A0_t (LED_128_Instance_SBox_Instance_12_L1), .A0_f (new_AGEMA_signal_4002), .A1_t (new_AGEMA_signal_4003), .A1_f (new_AGEMA_signal_4004), .B0_t (LED_128_Instance_addconst_out[50]), .B0_f (new_AGEMA_signal_3786), .B1_t (new_AGEMA_signal_3787), .B1_f (new_AGEMA_signal_3788), .Z0_t (LED_128_Instance_SBox_Instance_12_Q7), .Z0_f (new_AGEMA_signal_4230), .Z1_t (new_AGEMA_signal_4231), .Z1_f (new_AGEMA_signal_4232) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_12_AND1_U1 ( .A0_t (LED_128_Instance_SBox_Instance_12_L0), .A0_f (new_AGEMA_signal_3999), .A1_t (new_AGEMA_signal_4000), .A1_f (new_AGEMA_signal_4001), .B0_t (LED_128_Instance_addconst_out[51]), .B0_f (new_AGEMA_signal_3789), .B1_t (new_AGEMA_signal_3790), .B1_f (new_AGEMA_signal_3791), .Z0_t (LED_128_Instance_SBox_Instance_12_T0), .Z0_f (new_AGEMA_signal_4233), .Z1_t (new_AGEMA_signal_4234), .Z1_f (new_AGEMA_signal_4235) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_12_AND2_U1 ( .A0_t (LED_128_Instance_SBox_Instance_12_Q2), .A0_f (new_AGEMA_signal_4383), .A1_t (new_AGEMA_signal_4384), .A1_f (new_AGEMA_signal_4385), .B0_t (LED_128_Instance_SBox_Instance_12_Q3), .B0_f (new_AGEMA_signal_4227), .B1_t (new_AGEMA_signal_4228), .B1_f (new_AGEMA_signal_4229), .Z0_t (LED_128_Instance_SBox_Instance_12_T1), .Z0_f (new_AGEMA_signal_4497), .Z1_t (new_AGEMA_signal_4498), .Z1_f (new_AGEMA_signal_4499) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_12_AND3_U1 ( .A0_t (LED_128_Instance_addroundkey_out[49]), .A0_f (new_AGEMA_signal_3783), .A1_t (new_AGEMA_signal_3784), .A1_f (new_AGEMA_signal_3785), .B0_t (LED_128_Instance_addconst_out[50]), .B0_f (new_AGEMA_signal_3786), .B1_t (new_AGEMA_signal_3787), .B1_f (new_AGEMA_signal_3788), .Z0_t (LED_128_Instance_SBox_Instance_12_T2), .Z0_f (new_AGEMA_signal_4011), .Z1_t (new_AGEMA_signal_4012), .Z1_f (new_AGEMA_signal_4013) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_12_AND4_U1 ( .A0_t (LED_128_Instance_SBox_Instance_12_Q6), .A0_f (new_AGEMA_signal_4494), .A1_t (new_AGEMA_signal_4495), .A1_f (new_AGEMA_signal_4496), .B0_t (LED_128_Instance_SBox_Instance_12_Q7), .B0_f (new_AGEMA_signal_4230), .B1_t (new_AGEMA_signal_4231), .B1_f (new_AGEMA_signal_4232), .Z0_t (LED_128_Instance_SBox_Instance_12_T3), .Z0_f (new_AGEMA_signal_4596), .Z1_t (new_AGEMA_signal_4597), .Z1_f (new_AGEMA_signal_4598) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_12_XOR10_U1 ( .A0_t (LED_128_Instance_SBox_Instance_12_L5), .A0_f (new_AGEMA_signal_4386), .A1_t (new_AGEMA_signal_4387), .A1_f (new_AGEMA_signal_4388), .B0_t (LED_128_Instance_SBox_Instance_12_T3), .B0_f (new_AGEMA_signal_4596), .B1_t (new_AGEMA_signal_4597), .B1_f (new_AGEMA_signal_4598), .Z0_t (LED_128_Instance_SBox_Instance_12_L7), .Z0_f (new_AGEMA_signal_4719), .Z1_t (new_AGEMA_signal_4720), .Z1_f (new_AGEMA_signal_4721) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_12_XOR11_U1 ( .A0_t (LED_128_Instance_addroundkey_out[48]), .A0_f (new_AGEMA_signal_3780), .A1_t (new_AGEMA_signal_3781), .A1_f (new_AGEMA_signal_3782), .B0_t (LED_128_Instance_SBox_Instance_12_L7), .B0_f (new_AGEMA_signal_4719), .B1_t (new_AGEMA_signal_4720), .B1_f (new_AGEMA_signal_4721), .Z0_t (LED_128_Instance_subcells_out[51]), .Z0_f (new_AGEMA_signal_4806), .Z1_t (new_AGEMA_signal_4807), .Z1_f (new_AGEMA_signal_4808) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_12_XOR12_U1 ( .A0_t (LED_128_Instance_SBox_Instance_12_L5), .A0_f (new_AGEMA_signal_4386), .A1_t (new_AGEMA_signal_4387), .A1_f (new_AGEMA_signal_4388), .B0_t (LED_128_Instance_SBox_Instance_12_T1), .B0_f (new_AGEMA_signal_4497), .B1_t (new_AGEMA_signal_4498), .B1_f (new_AGEMA_signal_4499), .Z0_t (LED_128_Instance_SBox_Instance_12_L8), .Z0_f (new_AGEMA_signal_4599), .Z1_t (new_AGEMA_signal_4600), .Z1_f (new_AGEMA_signal_4601) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_12_XOR13_U1 ( .A0_t (LED_128_Instance_SBox_Instance_12_L1), .A0_f (new_AGEMA_signal_4002), .A1_t (new_AGEMA_signal_4003), .A1_f (new_AGEMA_signal_4004), .B0_t (LED_128_Instance_SBox_Instance_12_L8), .B0_f (new_AGEMA_signal_4599), .B1_t (new_AGEMA_signal_4600), .B1_f (new_AGEMA_signal_4601), .Z0_t (LED_128_Instance_subcells_out[50]), .Z0_f (new_AGEMA_signal_4722), .Z1_t (new_AGEMA_signal_4723), .Z1_f (new_AGEMA_signal_4724) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_12_XOR14_U1 ( .A0_t (LED_128_Instance_SBox_Instance_12_L4), .A0_f (new_AGEMA_signal_4008), .A1_t (new_AGEMA_signal_4009), .A1_f (new_AGEMA_signal_4010), .B0_t (LED_128_Instance_SBox_Instance_12_T3), .B0_f (new_AGEMA_signal_4596), .B1_t (new_AGEMA_signal_4597), .B1_f (new_AGEMA_signal_4598), .Z0_t (LED_128_Instance_subcells_out[49]), .Z0_f (new_AGEMA_signal_4725), .Z1_t (new_AGEMA_signal_4726), .Z1_f (new_AGEMA_signal_4727) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_12_XOR15_U1 ( .A0_t (LED_128_Instance_SBox_Instance_12_L3), .A0_f (new_AGEMA_signal_4005), .A1_t (new_AGEMA_signal_4006), .A1_f (new_AGEMA_signal_4007), .B0_t (LED_128_Instance_SBox_Instance_12_T2), .B0_f (new_AGEMA_signal_4011), .B1_t (new_AGEMA_signal_4012), .B1_f (new_AGEMA_signal_4013), .Z0_t (LED_128_Instance_subcells_out[48]), .Z0_f (new_AGEMA_signal_4236), .Z1_t (new_AGEMA_signal_4237), .Z1_f (new_AGEMA_signal_4238) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_13_XOR1_U1 ( .A0_t (LED_128_Instance_addconst_out[54]), .A0_f (new_AGEMA_signal_3828), .A1_t (new_AGEMA_signal_3829), .A1_f (new_AGEMA_signal_3830), .B0_t (LED_128_Instance_addconst_out[53]), .B0_f (new_AGEMA_signal_3852), .B1_t (new_AGEMA_signal_3853), .B1_f (new_AGEMA_signal_3854), .Z0_t (LED_128_Instance_SBox_Instance_13_L0), .Z0_f (new_AGEMA_signal_4239), .Z1_t (new_AGEMA_signal_4240), .Z1_f (new_AGEMA_signal_4241) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_13_XOR2_U1 ( .A0_t (LED_128_Instance_addconst_out[53]), .A0_f (new_AGEMA_signal_3852), .A1_t (new_AGEMA_signal_3853), .A1_f (new_AGEMA_signal_3854), .B0_t (LED_128_Instance_addconst_out[52]), .B0_f (new_AGEMA_signal_3846), .B1_t (new_AGEMA_signal_3847), .B1_f (new_AGEMA_signal_3848), .Z0_t (LED_128_Instance_SBox_Instance_13_L1), .Z0_f (new_AGEMA_signal_4242), .Z1_t (new_AGEMA_signal_4243), .Z1_f (new_AGEMA_signal_4244) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_13_XOR3_U1 ( .A0_t (LED_128_Instance_SBox_Instance_13_L1), .A0_f (new_AGEMA_signal_4242), .A1_t (new_AGEMA_signal_4243), .A1_f (new_AGEMA_signal_4244), .B0_t (LED_128_Instance_addconst_out[55]), .B0_f (new_AGEMA_signal_3801), .B1_t (new_AGEMA_signal_3802), .B1_f (new_AGEMA_signal_3803), .Z0_t (LED_128_Instance_SBox_Instance_13_L2), .Z0_f (new_AGEMA_signal_4389), .Z1_t (new_AGEMA_signal_4390), .Z1_f (new_AGEMA_signal_4391) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_SBox_Instance_13_XOR16_U1 ( .A0_t (LED_128_Instance_SBox_Instance_13_T0), .A0_f (new_AGEMA_signal_4398), .A1_t (new_AGEMA_signal_4399), .A1_f (new_AGEMA_signal_4400), .B0_t (LED_128_Instance_SBox_Instance_13_L2), .B0_f (new_AGEMA_signal_4389), .B1_t (new_AGEMA_signal_4390), .B1_f (new_AGEMA_signal_4391), .Z0_t (LED_128_Instance_SBox_Instance_13_Q2), .Z0_f (new_AGEMA_signal_4500), .Z1_t (new_AGEMA_signal_4501), .Z1_f (new_AGEMA_signal_4502) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_13_XOR4_U1 ( .A0_t (LED_128_Instance_addconst_out[55]), .A0_f (new_AGEMA_signal_3801), .A1_t (new_AGEMA_signal_3802), .A1_f (new_AGEMA_signal_3803), .B0_t (LED_128_Instance_addconst_out[52]), .B0_f (new_AGEMA_signal_3846), .B1_t (new_AGEMA_signal_3847), .B1_f (new_AGEMA_signal_3848), .Z0_t (LED_128_Instance_SBox_Instance_13_L3), .Z0_f (new_AGEMA_signal_4245), .Z1_t (new_AGEMA_signal_4246), .Z1_f (new_AGEMA_signal_4247) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_13_XOR5_U1 ( .A0_t (LED_128_Instance_SBox_Instance_13_L3), .A0_f (new_AGEMA_signal_4245), .A1_t (new_AGEMA_signal_4246), .A1_f (new_AGEMA_signal_4247), .B0_t (LED_128_Instance_SBox_Instance_13_L0), .B0_f (new_AGEMA_signal_4239), .B1_t (new_AGEMA_signal_4240), .B1_f (new_AGEMA_signal_4241), .Z0_t (LED_128_Instance_SBox_Instance_13_Q3), .Z0_f (new_AGEMA_signal_4392), .Z1_t (new_AGEMA_signal_4393), .Z1_f (new_AGEMA_signal_4394) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_13_XOR6_U1 ( .A0_t (LED_128_Instance_addconst_out[55]), .A0_f (new_AGEMA_signal_3801), .A1_t (new_AGEMA_signal_3802), .A1_f (new_AGEMA_signal_3803), .B0_t (LED_128_Instance_addconst_out[53]), .B0_f (new_AGEMA_signal_3852), .B1_t (new_AGEMA_signal_3853), .B1_f (new_AGEMA_signal_3854), .Z0_t (LED_128_Instance_SBox_Instance_13_L4), .Z0_f (new_AGEMA_signal_4248), .Z1_t (new_AGEMA_signal_4249), .Z1_f (new_AGEMA_signal_4250) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_13_XOR7_U1 ( .A0_t (LED_128_Instance_SBox_Instance_13_T0), .A0_f (new_AGEMA_signal_4398), .A1_t (new_AGEMA_signal_4399), .A1_f (new_AGEMA_signal_4400), .B0_t (LED_128_Instance_SBox_Instance_13_T2), .B0_f (new_AGEMA_signal_4251), .B1_t (new_AGEMA_signal_4252), .B1_f (new_AGEMA_signal_4253), .Z0_t (LED_128_Instance_SBox_Instance_13_L5), .Z0_f (new_AGEMA_signal_4503), .Z1_t (new_AGEMA_signal_4504), .Z1_f (new_AGEMA_signal_4505) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_SBox_Instance_13_XOR8_U1 ( .A0_t (LED_128_Instance_SBox_Instance_13_L4), .A0_f (new_AGEMA_signal_4248), .A1_t (new_AGEMA_signal_4249), .A1_f (new_AGEMA_signal_4250), .B0_t (LED_128_Instance_SBox_Instance_13_L5), .B0_f (new_AGEMA_signal_4503), .B1_t (new_AGEMA_signal_4504), .B1_f (new_AGEMA_signal_4505), .Z0_t (LED_128_Instance_SBox_Instance_13_Q6), .Z0_f (new_AGEMA_signal_4602), .Z1_t (new_AGEMA_signal_4603), .Z1_f (new_AGEMA_signal_4604) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_13_XOR9_U1 ( .A0_t (LED_128_Instance_SBox_Instance_13_L1), .A0_f (new_AGEMA_signal_4242), .A1_t (new_AGEMA_signal_4243), .A1_f (new_AGEMA_signal_4244), .B0_t (LED_128_Instance_addconst_out[54]), .B0_f (new_AGEMA_signal_3828), .B1_t (new_AGEMA_signal_3829), .B1_f (new_AGEMA_signal_3830), .Z0_t (LED_128_Instance_SBox_Instance_13_Q7), .Z0_f (new_AGEMA_signal_4395), .Z1_t (new_AGEMA_signal_4396), .Z1_f (new_AGEMA_signal_4397) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_13_AND1_U1 ( .A0_t (LED_128_Instance_SBox_Instance_13_L0), .A0_f (new_AGEMA_signal_4239), .A1_t (new_AGEMA_signal_4240), .A1_f (new_AGEMA_signal_4241), .B0_t (LED_128_Instance_addconst_out[55]), .B0_f (new_AGEMA_signal_3801), .B1_t (new_AGEMA_signal_3802), .B1_f (new_AGEMA_signal_3803), .Z0_t (LED_128_Instance_SBox_Instance_13_T0), .Z0_f (new_AGEMA_signal_4398), .Z1_t (new_AGEMA_signal_4399), .Z1_f (new_AGEMA_signal_4400) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_13_AND2_U1 ( .A0_t (LED_128_Instance_SBox_Instance_13_Q2), .A0_f (new_AGEMA_signal_4500), .A1_t (new_AGEMA_signal_4501), .A1_f (new_AGEMA_signal_4502), .B0_t (LED_128_Instance_SBox_Instance_13_Q3), .B0_f (new_AGEMA_signal_4392), .B1_t (new_AGEMA_signal_4393), .B1_f (new_AGEMA_signal_4394), .Z0_t (LED_128_Instance_SBox_Instance_13_T1), .Z0_f (new_AGEMA_signal_4605), .Z1_t (new_AGEMA_signal_4606), .Z1_f (new_AGEMA_signal_4607) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_13_AND3_U1 ( .A0_t (LED_128_Instance_addconst_out[53]), .A0_f (new_AGEMA_signal_3852), .A1_t (new_AGEMA_signal_3853), .A1_f (new_AGEMA_signal_3854), .B0_t (LED_128_Instance_addconst_out[54]), .B0_f (new_AGEMA_signal_3828), .B1_t (new_AGEMA_signal_3829), .B1_f (new_AGEMA_signal_3830), .Z0_t (LED_128_Instance_SBox_Instance_13_T2), .Z0_f (new_AGEMA_signal_4251), .Z1_t (new_AGEMA_signal_4252), .Z1_f (new_AGEMA_signal_4253) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_13_AND4_U1 ( .A0_t (LED_128_Instance_SBox_Instance_13_Q6), .A0_f (new_AGEMA_signal_4602), .A1_t (new_AGEMA_signal_4603), .A1_f (new_AGEMA_signal_4604), .B0_t (LED_128_Instance_SBox_Instance_13_Q7), .B0_f (new_AGEMA_signal_4395), .B1_t (new_AGEMA_signal_4396), .B1_f (new_AGEMA_signal_4397), .Z0_t (LED_128_Instance_SBox_Instance_13_T3), .Z0_f (new_AGEMA_signal_4728), .Z1_t (new_AGEMA_signal_4729), .Z1_f (new_AGEMA_signal_4730) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_13_XOR10_U1 ( .A0_t (LED_128_Instance_SBox_Instance_13_L5), .A0_f (new_AGEMA_signal_4503), .A1_t (new_AGEMA_signal_4504), .A1_f (new_AGEMA_signal_4505), .B0_t (LED_128_Instance_SBox_Instance_13_T3), .B0_f (new_AGEMA_signal_4728), .B1_t (new_AGEMA_signal_4729), .B1_f (new_AGEMA_signal_4730), .Z0_t (LED_128_Instance_SBox_Instance_13_L7), .Z0_f (new_AGEMA_signal_4809), .Z1_t (new_AGEMA_signal_4810), .Z1_f (new_AGEMA_signal_4811) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_13_XOR11_U1 ( .A0_t (LED_128_Instance_addconst_out[52]), .A0_f (new_AGEMA_signal_3846), .A1_t (new_AGEMA_signal_3847), .A1_f (new_AGEMA_signal_3848), .B0_t (LED_128_Instance_SBox_Instance_13_L7), .B0_f (new_AGEMA_signal_4809), .B1_t (new_AGEMA_signal_4810), .B1_f (new_AGEMA_signal_4811), .Z0_t (LED_128_Instance_subcells_out[55]), .Z0_f (new_AGEMA_signal_4896), .Z1_t (new_AGEMA_signal_4897), .Z1_f (new_AGEMA_signal_4898) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_13_XOR12_U1 ( .A0_t (LED_128_Instance_SBox_Instance_13_L5), .A0_f (new_AGEMA_signal_4503), .A1_t (new_AGEMA_signal_4504), .A1_f (new_AGEMA_signal_4505), .B0_t (LED_128_Instance_SBox_Instance_13_T1), .B0_f (new_AGEMA_signal_4605), .B1_t (new_AGEMA_signal_4606), .B1_f (new_AGEMA_signal_4607), .Z0_t (LED_128_Instance_SBox_Instance_13_L8), .Z0_f (new_AGEMA_signal_4731), .Z1_t (new_AGEMA_signal_4732), .Z1_f (new_AGEMA_signal_4733) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_13_XOR13_U1 ( .A0_t (LED_128_Instance_SBox_Instance_13_L1), .A0_f (new_AGEMA_signal_4242), .A1_t (new_AGEMA_signal_4243), .A1_f (new_AGEMA_signal_4244), .B0_t (LED_128_Instance_SBox_Instance_13_L8), .B0_f (new_AGEMA_signal_4731), .B1_t (new_AGEMA_signal_4732), .B1_f (new_AGEMA_signal_4733), .Z0_t (LED_128_Instance_subcells_out[54]), .Z0_f (new_AGEMA_signal_4812), .Z1_t (new_AGEMA_signal_4813), .Z1_f (new_AGEMA_signal_4814) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_13_XOR14_U1 ( .A0_t (LED_128_Instance_SBox_Instance_13_L4), .A0_f (new_AGEMA_signal_4248), .A1_t (new_AGEMA_signal_4249), .A1_f (new_AGEMA_signal_4250), .B0_t (LED_128_Instance_SBox_Instance_13_T3), .B0_f (new_AGEMA_signal_4728), .B1_t (new_AGEMA_signal_4729), .B1_f (new_AGEMA_signal_4730), .Z0_t (LED_128_Instance_subcells_out[53]), .Z0_f (new_AGEMA_signal_4815), .Z1_t (new_AGEMA_signal_4816), .Z1_f (new_AGEMA_signal_4817) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_13_XOR15_U1 ( .A0_t (LED_128_Instance_SBox_Instance_13_L3), .A0_f (new_AGEMA_signal_4245), .A1_t (new_AGEMA_signal_4246), .A1_f (new_AGEMA_signal_4247), .B0_t (LED_128_Instance_SBox_Instance_13_T2), .B0_f (new_AGEMA_signal_4251), .B1_t (new_AGEMA_signal_4252), .B1_f (new_AGEMA_signal_4253), .Z0_t (LED_128_Instance_subcells_out[52]), .Z0_f (new_AGEMA_signal_4401), .Z1_t (new_AGEMA_signal_4402), .Z1_f (new_AGEMA_signal_4403) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_14_XOR1_U1 ( .A0_t (LED_128_Instance_addconst_out[58]), .A0_f (new_AGEMA_signal_3810), .A1_t (new_AGEMA_signal_3811), .A1_f (new_AGEMA_signal_3812), .B0_t (LED_128_Instance_addconst_out[57]), .B0_f (new_AGEMA_signal_3807), .B1_t (new_AGEMA_signal_3808), .B1_f (new_AGEMA_signal_3809), .Z0_t (LED_128_Instance_SBox_Instance_14_L0), .Z0_f (new_AGEMA_signal_4014), .Z1_t (new_AGEMA_signal_4015), .Z1_f (new_AGEMA_signal_4016) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_14_XOR2_U1 ( .A0_t (LED_128_Instance_addconst_out[57]), .A0_f (new_AGEMA_signal_3807), .A1_t (new_AGEMA_signal_3808), .A1_f (new_AGEMA_signal_3809), .B0_t (LED_128_Instance_addconst_out[56]), .B0_f (new_AGEMA_signal_3804), .B1_t (new_AGEMA_signal_3805), .B1_f (new_AGEMA_signal_3806), .Z0_t (LED_128_Instance_SBox_Instance_14_L1), .Z0_f (new_AGEMA_signal_4017), .Z1_t (new_AGEMA_signal_4018), .Z1_f (new_AGEMA_signal_4019) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_14_XOR3_U1 ( .A0_t (LED_128_Instance_SBox_Instance_14_L1), .A0_f (new_AGEMA_signal_4017), .A1_t (new_AGEMA_signal_4018), .A1_f (new_AGEMA_signal_4019), .B0_t (LED_128_Instance_addconst_out[59]), .B0_f (new_AGEMA_signal_3813), .B1_t (new_AGEMA_signal_3814), .B1_f (new_AGEMA_signal_3815), .Z0_t (LED_128_Instance_SBox_Instance_14_L2), .Z0_f (new_AGEMA_signal_4254), .Z1_t (new_AGEMA_signal_4255), .Z1_f (new_AGEMA_signal_4256) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_SBox_Instance_14_XOR16_U1 ( .A0_t (LED_128_Instance_SBox_Instance_14_T0), .A0_f (new_AGEMA_signal_4263), .A1_t (new_AGEMA_signal_4264), .A1_f (new_AGEMA_signal_4265), .B0_t (LED_128_Instance_SBox_Instance_14_L2), .B0_f (new_AGEMA_signal_4254), .B1_t (new_AGEMA_signal_4255), .B1_f (new_AGEMA_signal_4256), .Z0_t (LED_128_Instance_SBox_Instance_14_Q2), .Z0_f (new_AGEMA_signal_4404), .Z1_t (new_AGEMA_signal_4405), .Z1_f (new_AGEMA_signal_4406) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_14_XOR4_U1 ( .A0_t (LED_128_Instance_addconst_out[59]), .A0_f (new_AGEMA_signal_3813), .A1_t (new_AGEMA_signal_3814), .A1_f (new_AGEMA_signal_3815), .B0_t (LED_128_Instance_addconst_out[56]), .B0_f (new_AGEMA_signal_3804), .B1_t (new_AGEMA_signal_3805), .B1_f (new_AGEMA_signal_3806), .Z0_t (LED_128_Instance_SBox_Instance_14_L3), .Z0_f (new_AGEMA_signal_4020), .Z1_t (new_AGEMA_signal_4021), .Z1_f (new_AGEMA_signal_4022) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_14_XOR5_U1 ( .A0_t (LED_128_Instance_SBox_Instance_14_L3), .A0_f (new_AGEMA_signal_4020), .A1_t (new_AGEMA_signal_4021), .A1_f (new_AGEMA_signal_4022), .B0_t (LED_128_Instance_SBox_Instance_14_L0), .B0_f (new_AGEMA_signal_4014), .B1_t (new_AGEMA_signal_4015), .B1_f (new_AGEMA_signal_4016), .Z0_t (LED_128_Instance_SBox_Instance_14_Q3), .Z0_f (new_AGEMA_signal_4257), .Z1_t (new_AGEMA_signal_4258), .Z1_f (new_AGEMA_signal_4259) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_14_XOR6_U1 ( .A0_t (LED_128_Instance_addconst_out[59]), .A0_f (new_AGEMA_signal_3813), .A1_t (new_AGEMA_signal_3814), .A1_f (new_AGEMA_signal_3815), .B0_t (LED_128_Instance_addconst_out[57]), .B0_f (new_AGEMA_signal_3807), .B1_t (new_AGEMA_signal_3808), .B1_f (new_AGEMA_signal_3809), .Z0_t (LED_128_Instance_SBox_Instance_14_L4), .Z0_f (new_AGEMA_signal_4023), .Z1_t (new_AGEMA_signal_4024), .Z1_f (new_AGEMA_signal_4025) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_14_XOR7_U1 ( .A0_t (LED_128_Instance_SBox_Instance_14_T0), .A0_f (new_AGEMA_signal_4263), .A1_t (new_AGEMA_signal_4264), .A1_f (new_AGEMA_signal_4265), .B0_t (LED_128_Instance_SBox_Instance_14_T2), .B0_f (new_AGEMA_signal_4026), .B1_t (new_AGEMA_signal_4027), .B1_f (new_AGEMA_signal_4028), .Z0_t (LED_128_Instance_SBox_Instance_14_L5), .Z0_f (new_AGEMA_signal_4407), .Z1_t (new_AGEMA_signal_4408), .Z1_f (new_AGEMA_signal_4409) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_SBox_Instance_14_XOR8_U1 ( .A0_t (LED_128_Instance_SBox_Instance_14_L4), .A0_f (new_AGEMA_signal_4023), .A1_t (new_AGEMA_signal_4024), .A1_f (new_AGEMA_signal_4025), .B0_t (LED_128_Instance_SBox_Instance_14_L5), .B0_f (new_AGEMA_signal_4407), .B1_t (new_AGEMA_signal_4408), .B1_f (new_AGEMA_signal_4409), .Z0_t (LED_128_Instance_SBox_Instance_14_Q6), .Z0_f (new_AGEMA_signal_4506), .Z1_t (new_AGEMA_signal_4507), .Z1_f (new_AGEMA_signal_4508) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_14_XOR9_U1 ( .A0_t (LED_128_Instance_SBox_Instance_14_L1), .A0_f (new_AGEMA_signal_4017), .A1_t (new_AGEMA_signal_4018), .A1_f (new_AGEMA_signal_4019), .B0_t (LED_128_Instance_addconst_out[58]), .B0_f (new_AGEMA_signal_3810), .B1_t (new_AGEMA_signal_3811), .B1_f (new_AGEMA_signal_3812), .Z0_t (LED_128_Instance_SBox_Instance_14_Q7), .Z0_f (new_AGEMA_signal_4260), .Z1_t (new_AGEMA_signal_4261), .Z1_f (new_AGEMA_signal_4262) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_14_AND1_U1 ( .A0_t (LED_128_Instance_SBox_Instance_14_L0), .A0_f (new_AGEMA_signal_4014), .A1_t (new_AGEMA_signal_4015), .A1_f (new_AGEMA_signal_4016), .B0_t (LED_128_Instance_addconst_out[59]), .B0_f (new_AGEMA_signal_3813), .B1_t (new_AGEMA_signal_3814), .B1_f (new_AGEMA_signal_3815), .Z0_t (LED_128_Instance_SBox_Instance_14_T0), .Z0_f (new_AGEMA_signal_4263), .Z1_t (new_AGEMA_signal_4264), .Z1_f (new_AGEMA_signal_4265) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_14_AND2_U1 ( .A0_t (LED_128_Instance_SBox_Instance_14_Q2), .A0_f (new_AGEMA_signal_4404), .A1_t (new_AGEMA_signal_4405), .A1_f (new_AGEMA_signal_4406), .B0_t (LED_128_Instance_SBox_Instance_14_Q3), .B0_f (new_AGEMA_signal_4257), .B1_t (new_AGEMA_signal_4258), .B1_f (new_AGEMA_signal_4259), .Z0_t (LED_128_Instance_SBox_Instance_14_T1), .Z0_f (new_AGEMA_signal_4509), .Z1_t (new_AGEMA_signal_4510), .Z1_f (new_AGEMA_signal_4511) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_14_AND3_U1 ( .A0_t (LED_128_Instance_addconst_out[57]), .A0_f (new_AGEMA_signal_3807), .A1_t (new_AGEMA_signal_3808), .A1_f (new_AGEMA_signal_3809), .B0_t (LED_128_Instance_addconst_out[58]), .B0_f (new_AGEMA_signal_3810), .B1_t (new_AGEMA_signal_3811), .B1_f (new_AGEMA_signal_3812), .Z0_t (LED_128_Instance_SBox_Instance_14_T2), .Z0_f (new_AGEMA_signal_4026), .Z1_t (new_AGEMA_signal_4027), .Z1_f (new_AGEMA_signal_4028) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_14_AND4_U1 ( .A0_t (LED_128_Instance_SBox_Instance_14_Q6), .A0_f (new_AGEMA_signal_4506), .A1_t (new_AGEMA_signal_4507), .A1_f (new_AGEMA_signal_4508), .B0_t (LED_128_Instance_SBox_Instance_14_Q7), .B0_f (new_AGEMA_signal_4260), .B1_t (new_AGEMA_signal_4261), .B1_f (new_AGEMA_signal_4262), .Z0_t (LED_128_Instance_SBox_Instance_14_T3), .Z0_f (new_AGEMA_signal_4608), .Z1_t (new_AGEMA_signal_4609), .Z1_f (new_AGEMA_signal_4610) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_14_XOR10_U1 ( .A0_t (LED_128_Instance_SBox_Instance_14_L5), .A0_f (new_AGEMA_signal_4407), .A1_t (new_AGEMA_signal_4408), .A1_f (new_AGEMA_signal_4409), .B0_t (LED_128_Instance_SBox_Instance_14_T3), .B0_f (new_AGEMA_signal_4608), .B1_t (new_AGEMA_signal_4609), .B1_f (new_AGEMA_signal_4610), .Z0_t (LED_128_Instance_SBox_Instance_14_L7), .Z0_f (new_AGEMA_signal_4734), .Z1_t (new_AGEMA_signal_4735), .Z1_f (new_AGEMA_signal_4736) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_14_XOR11_U1 ( .A0_t (LED_128_Instance_addconst_out[56]), .A0_f (new_AGEMA_signal_3804), .A1_t (new_AGEMA_signal_3805), .A1_f (new_AGEMA_signal_3806), .B0_t (LED_128_Instance_SBox_Instance_14_L7), .B0_f (new_AGEMA_signal_4734), .B1_t (new_AGEMA_signal_4735), .B1_f (new_AGEMA_signal_4736), .Z0_t (LED_128_Instance_subcells_out[59]), .Z0_f (new_AGEMA_signal_4818), .Z1_t (new_AGEMA_signal_4819), .Z1_f (new_AGEMA_signal_4820) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_14_XOR12_U1 ( .A0_t (LED_128_Instance_SBox_Instance_14_L5), .A0_f (new_AGEMA_signal_4407), .A1_t (new_AGEMA_signal_4408), .A1_f (new_AGEMA_signal_4409), .B0_t (LED_128_Instance_SBox_Instance_14_T1), .B0_f (new_AGEMA_signal_4509), .B1_t (new_AGEMA_signal_4510), .B1_f (new_AGEMA_signal_4511), .Z0_t (LED_128_Instance_SBox_Instance_14_L8), .Z0_f (new_AGEMA_signal_4611), .Z1_t (new_AGEMA_signal_4612), .Z1_f (new_AGEMA_signal_4613) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_14_XOR13_U1 ( .A0_t (LED_128_Instance_SBox_Instance_14_L1), .A0_f (new_AGEMA_signal_4017), .A1_t (new_AGEMA_signal_4018), .A1_f (new_AGEMA_signal_4019), .B0_t (LED_128_Instance_SBox_Instance_14_L8), .B0_f (new_AGEMA_signal_4611), .B1_t (new_AGEMA_signal_4612), .B1_f (new_AGEMA_signal_4613), .Z0_t (LED_128_Instance_subcells_out[58]), .Z0_f (new_AGEMA_signal_4737), .Z1_t (new_AGEMA_signal_4738), .Z1_f (new_AGEMA_signal_4739) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_14_XOR14_U1 ( .A0_t (LED_128_Instance_SBox_Instance_14_L4), .A0_f (new_AGEMA_signal_4023), .A1_t (new_AGEMA_signal_4024), .A1_f (new_AGEMA_signal_4025), .B0_t (LED_128_Instance_SBox_Instance_14_T3), .B0_f (new_AGEMA_signal_4608), .B1_t (new_AGEMA_signal_4609), .B1_f (new_AGEMA_signal_4610), .Z0_t (LED_128_Instance_subcells_out[57]), .Z0_f (new_AGEMA_signal_4740), .Z1_t (new_AGEMA_signal_4741), .Z1_f (new_AGEMA_signal_4742) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_14_XOR15_U1 ( .A0_t (LED_128_Instance_SBox_Instance_14_L3), .A0_f (new_AGEMA_signal_4020), .A1_t (new_AGEMA_signal_4021), .A1_f (new_AGEMA_signal_4022), .B0_t (LED_128_Instance_SBox_Instance_14_T2), .B0_f (new_AGEMA_signal_4026), .B1_t (new_AGEMA_signal_4027), .B1_f (new_AGEMA_signal_4028), .Z0_t (LED_128_Instance_subcells_out[56]), .Z0_f (new_AGEMA_signal_4266), .Z1_t (new_AGEMA_signal_4267), .Z1_f (new_AGEMA_signal_4268) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_15_XOR1_U1 ( .A0_t (LED_128_Instance_addconst_out[62]), .A0_f (new_AGEMA_signal_3822), .A1_t (new_AGEMA_signal_3823), .A1_f (new_AGEMA_signal_3824), .B0_t (LED_128_Instance_addconst_out[61]), .B0_f (new_AGEMA_signal_3819), .B1_t (new_AGEMA_signal_3820), .B1_f (new_AGEMA_signal_3821), .Z0_t (LED_128_Instance_SBox_Instance_15_L0), .Z0_f (new_AGEMA_signal_4029), .Z1_t (new_AGEMA_signal_4030), .Z1_f (new_AGEMA_signal_4031) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_15_XOR2_U1 ( .A0_t (LED_128_Instance_addconst_out[61]), .A0_f (new_AGEMA_signal_3819), .A1_t (new_AGEMA_signal_3820), .A1_f (new_AGEMA_signal_3821), .B0_t (LED_128_Instance_addconst_out[60]), .B0_f (new_AGEMA_signal_3816), .B1_t (new_AGEMA_signal_3817), .B1_f (new_AGEMA_signal_3818), .Z0_t (LED_128_Instance_SBox_Instance_15_L1), .Z0_f (new_AGEMA_signal_4032), .Z1_t (new_AGEMA_signal_4033), .Z1_f (new_AGEMA_signal_4034) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_15_XOR3_U1 ( .A0_t (LED_128_Instance_SBox_Instance_15_L1), .A0_f (new_AGEMA_signal_4032), .A1_t (new_AGEMA_signal_4033), .A1_f (new_AGEMA_signal_4034), .B0_t (LED_128_Instance_addconst_out[63]), .B0_f (new_AGEMA_signal_3825), .B1_t (new_AGEMA_signal_3826), .B1_f (new_AGEMA_signal_3827), .Z0_t (LED_128_Instance_SBox_Instance_15_L2), .Z0_f (new_AGEMA_signal_4269), .Z1_t (new_AGEMA_signal_4270), .Z1_f (new_AGEMA_signal_4271) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_SBox_Instance_15_XOR16_U1 ( .A0_t (LED_128_Instance_SBox_Instance_15_T0), .A0_f (new_AGEMA_signal_4278), .A1_t (new_AGEMA_signal_4279), .A1_f (new_AGEMA_signal_4280), .B0_t (LED_128_Instance_SBox_Instance_15_L2), .B0_f (new_AGEMA_signal_4269), .B1_t (new_AGEMA_signal_4270), .B1_f (new_AGEMA_signal_4271), .Z0_t (LED_128_Instance_SBox_Instance_15_Q2), .Z0_f (new_AGEMA_signal_4410), .Z1_t (new_AGEMA_signal_4411), .Z1_f (new_AGEMA_signal_4412) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_15_XOR4_U1 ( .A0_t (LED_128_Instance_addconst_out[63]), .A0_f (new_AGEMA_signal_3825), .A1_t (new_AGEMA_signal_3826), .A1_f (new_AGEMA_signal_3827), .B0_t (LED_128_Instance_addconst_out[60]), .B0_f (new_AGEMA_signal_3816), .B1_t (new_AGEMA_signal_3817), .B1_f (new_AGEMA_signal_3818), .Z0_t (LED_128_Instance_SBox_Instance_15_L3), .Z0_f (new_AGEMA_signal_4035), .Z1_t (new_AGEMA_signal_4036), .Z1_f (new_AGEMA_signal_4037) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_15_XOR5_U1 ( .A0_t (LED_128_Instance_SBox_Instance_15_L3), .A0_f (new_AGEMA_signal_4035), .A1_t (new_AGEMA_signal_4036), .A1_f (new_AGEMA_signal_4037), .B0_t (LED_128_Instance_SBox_Instance_15_L0), .B0_f (new_AGEMA_signal_4029), .B1_t (new_AGEMA_signal_4030), .B1_f (new_AGEMA_signal_4031), .Z0_t (LED_128_Instance_SBox_Instance_15_Q3), .Z0_f (new_AGEMA_signal_4272), .Z1_t (new_AGEMA_signal_4273), .Z1_f (new_AGEMA_signal_4274) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_15_XOR6_U1 ( .A0_t (LED_128_Instance_addconst_out[63]), .A0_f (new_AGEMA_signal_3825), .A1_t (new_AGEMA_signal_3826), .A1_f (new_AGEMA_signal_3827), .B0_t (LED_128_Instance_addconst_out[61]), .B0_f (new_AGEMA_signal_3819), .B1_t (new_AGEMA_signal_3820), .B1_f (new_AGEMA_signal_3821), .Z0_t (LED_128_Instance_SBox_Instance_15_L4), .Z0_f (new_AGEMA_signal_4038), .Z1_t (new_AGEMA_signal_4039), .Z1_f (new_AGEMA_signal_4040) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_15_XOR7_U1 ( .A0_t (LED_128_Instance_SBox_Instance_15_T0), .A0_f (new_AGEMA_signal_4278), .A1_t (new_AGEMA_signal_4279), .A1_f (new_AGEMA_signal_4280), .B0_t (LED_128_Instance_SBox_Instance_15_T2), .B0_f (new_AGEMA_signal_4041), .B1_t (new_AGEMA_signal_4042), .B1_f (new_AGEMA_signal_4043), .Z0_t (LED_128_Instance_SBox_Instance_15_L5), .Z0_f (new_AGEMA_signal_4413), .Z1_t (new_AGEMA_signal_4414), .Z1_f (new_AGEMA_signal_4415) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_SBox_Instance_15_XOR8_U1 ( .A0_t (LED_128_Instance_SBox_Instance_15_L4), .A0_f (new_AGEMA_signal_4038), .A1_t (new_AGEMA_signal_4039), .A1_f (new_AGEMA_signal_4040), .B0_t (LED_128_Instance_SBox_Instance_15_L5), .B0_f (new_AGEMA_signal_4413), .B1_t (new_AGEMA_signal_4414), .B1_f (new_AGEMA_signal_4415), .Z0_t (LED_128_Instance_SBox_Instance_15_Q6), .Z0_f (new_AGEMA_signal_4512), .Z1_t (new_AGEMA_signal_4513), .Z1_f (new_AGEMA_signal_4514) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_15_XOR9_U1 ( .A0_t (LED_128_Instance_SBox_Instance_15_L1), .A0_f (new_AGEMA_signal_4032), .A1_t (new_AGEMA_signal_4033), .A1_f (new_AGEMA_signal_4034), .B0_t (LED_128_Instance_addconst_out[62]), .B0_f (new_AGEMA_signal_3822), .B1_t (new_AGEMA_signal_3823), .B1_f (new_AGEMA_signal_3824), .Z0_t (LED_128_Instance_SBox_Instance_15_Q7), .Z0_f (new_AGEMA_signal_4275), .Z1_t (new_AGEMA_signal_4276), .Z1_f (new_AGEMA_signal_4277) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_15_AND1_U1 ( .A0_t (LED_128_Instance_SBox_Instance_15_L0), .A0_f (new_AGEMA_signal_4029), .A1_t (new_AGEMA_signal_4030), .A1_f (new_AGEMA_signal_4031), .B0_t (LED_128_Instance_addconst_out[63]), .B0_f (new_AGEMA_signal_3825), .B1_t (new_AGEMA_signal_3826), .B1_f (new_AGEMA_signal_3827), .Z0_t (LED_128_Instance_SBox_Instance_15_T0), .Z0_f (new_AGEMA_signal_4278), .Z1_t (new_AGEMA_signal_4279), .Z1_f (new_AGEMA_signal_4280) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_15_AND2_U1 ( .A0_t (LED_128_Instance_SBox_Instance_15_Q2), .A0_f (new_AGEMA_signal_4410), .A1_t (new_AGEMA_signal_4411), .A1_f (new_AGEMA_signal_4412), .B0_t (LED_128_Instance_SBox_Instance_15_Q3), .B0_f (new_AGEMA_signal_4272), .B1_t (new_AGEMA_signal_4273), .B1_f (new_AGEMA_signal_4274), .Z0_t (LED_128_Instance_SBox_Instance_15_T1), .Z0_f (new_AGEMA_signal_4515), .Z1_t (new_AGEMA_signal_4516), .Z1_f (new_AGEMA_signal_4517) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_15_AND3_U1 ( .A0_t (LED_128_Instance_addconst_out[61]), .A0_f (new_AGEMA_signal_3819), .A1_t (new_AGEMA_signal_3820), .A1_f (new_AGEMA_signal_3821), .B0_t (LED_128_Instance_addconst_out[62]), .B0_f (new_AGEMA_signal_3822), .B1_t (new_AGEMA_signal_3823), .B1_f (new_AGEMA_signal_3824), .Z0_t (LED_128_Instance_SBox_Instance_15_T2), .Z0_f (new_AGEMA_signal_4041), .Z1_t (new_AGEMA_signal_4042), .Z1_f (new_AGEMA_signal_4043) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_15_AND4_U1 ( .A0_t (LED_128_Instance_SBox_Instance_15_Q6), .A0_f (new_AGEMA_signal_4512), .A1_t (new_AGEMA_signal_4513), .A1_f (new_AGEMA_signal_4514), .B0_t (LED_128_Instance_SBox_Instance_15_Q7), .B0_f (new_AGEMA_signal_4275), .B1_t (new_AGEMA_signal_4276), .B1_f (new_AGEMA_signal_4277), .Z0_t (LED_128_Instance_SBox_Instance_15_T3), .Z0_f (new_AGEMA_signal_4614), .Z1_t (new_AGEMA_signal_4615), .Z1_f (new_AGEMA_signal_4616) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_15_XOR10_U1 ( .A0_t (LED_128_Instance_SBox_Instance_15_L5), .A0_f (new_AGEMA_signal_4413), .A1_t (new_AGEMA_signal_4414), .A1_f (new_AGEMA_signal_4415), .B0_t (LED_128_Instance_SBox_Instance_15_T3), .B0_f (new_AGEMA_signal_4614), .B1_t (new_AGEMA_signal_4615), .B1_f (new_AGEMA_signal_4616), .Z0_t (LED_128_Instance_SBox_Instance_15_L7), .Z0_f (new_AGEMA_signal_4743), .Z1_t (new_AGEMA_signal_4744), .Z1_f (new_AGEMA_signal_4745) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_15_XOR11_U1 ( .A0_t (LED_128_Instance_addconst_out[60]), .A0_f (new_AGEMA_signal_3816), .A1_t (new_AGEMA_signal_3817), .A1_f (new_AGEMA_signal_3818), .B0_t (LED_128_Instance_SBox_Instance_15_L7), .B0_f (new_AGEMA_signal_4743), .B1_t (new_AGEMA_signal_4744), .B1_f (new_AGEMA_signal_4745), .Z0_t (LED_128_Instance_subcells_out[63]), .Z0_f (new_AGEMA_signal_4821), .Z1_t (new_AGEMA_signal_4822), .Z1_f (new_AGEMA_signal_4823) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_15_XOR12_U1 ( .A0_t (LED_128_Instance_SBox_Instance_15_L5), .A0_f (new_AGEMA_signal_4413), .A1_t (new_AGEMA_signal_4414), .A1_f (new_AGEMA_signal_4415), .B0_t (LED_128_Instance_SBox_Instance_15_T1), .B0_f (new_AGEMA_signal_4515), .B1_t (new_AGEMA_signal_4516), .B1_f (new_AGEMA_signal_4517), .Z0_t (LED_128_Instance_SBox_Instance_15_L8), .Z0_f (new_AGEMA_signal_4617), .Z1_t (new_AGEMA_signal_4618), .Z1_f (new_AGEMA_signal_4619) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_15_XOR13_U1 ( .A0_t (LED_128_Instance_SBox_Instance_15_L1), .A0_f (new_AGEMA_signal_4032), .A1_t (new_AGEMA_signal_4033), .A1_f (new_AGEMA_signal_4034), .B0_t (LED_128_Instance_SBox_Instance_15_L8), .B0_f (new_AGEMA_signal_4617), .B1_t (new_AGEMA_signal_4618), .B1_f (new_AGEMA_signal_4619), .Z0_t (LED_128_Instance_subcells_out[62]), .Z0_f (new_AGEMA_signal_4746), .Z1_t (new_AGEMA_signal_4747), .Z1_f (new_AGEMA_signal_4748) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_15_XOR14_U1 ( .A0_t (LED_128_Instance_SBox_Instance_15_L4), .A0_f (new_AGEMA_signal_4038), .A1_t (new_AGEMA_signal_4039), .A1_f (new_AGEMA_signal_4040), .B0_t (LED_128_Instance_SBox_Instance_15_T3), .B0_f (new_AGEMA_signal_4614), .B1_t (new_AGEMA_signal_4615), .B1_f (new_AGEMA_signal_4616), .Z0_t (LED_128_Instance_subcells_out[61]), .Z0_f (new_AGEMA_signal_4749), .Z1_t (new_AGEMA_signal_4750), .Z1_f (new_AGEMA_signal_4751) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_SBox_Instance_15_XOR15_U1 ( .A0_t (LED_128_Instance_SBox_Instance_15_L3), .A0_f (new_AGEMA_signal_4035), .A1_t (new_AGEMA_signal_4036), .A1_f (new_AGEMA_signal_4037), .B0_t (LED_128_Instance_SBox_Instance_15_T2), .B0_f (new_AGEMA_signal_4041), .B1_t (new_AGEMA_signal_4042), .B1_f (new_AGEMA_signal_4043), .Z0_t (LED_128_Instance_subcells_out[60]), .Z0_f (new_AGEMA_signal_4281), .Z1_t (new_AGEMA_signal_4282), .Z1_f (new_AGEMA_signal_4283) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U58 ( .A0_t (LED_128_Instance_subcells_out[2]), .A0_f (new_AGEMA_signal_4623), .A1_t (new_AGEMA_signal_4624), .A1_f (new_AGEMA_signal_4625), .B0_t (LED_128_Instance_MCS_Instance_0_n42), .B0_f (new_AGEMA_signal_5139), .B1_t (new_AGEMA_signal_5140), .B1_f (new_AGEMA_signal_5141), .Z0_t (LED_128_Instance_mixcolumns_out[1]), .Z0_f (new_AGEMA_signal_5319), .Z1_t (new_AGEMA_signal_5320), .Z1_f (new_AGEMA_signal_5321) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U57 ( .A0_t (LED_128_Instance_MCS_Instance_0_n41), .A0_f (new_AGEMA_signal_5334), .A1_t (new_AGEMA_signal_5335), .A1_f (new_AGEMA_signal_5336), .B0_t (LED_128_Instance_subcells_out[62]), .B0_f (new_AGEMA_signal_4746), .B1_t (new_AGEMA_signal_4747), .B1_f (new_AGEMA_signal_4748), .Z0_t (LED_128_Instance_mixcolumns_out[19]), .Z0_f (new_AGEMA_signal_5556), .Z1_t (new_AGEMA_signal_5557), .Z1_f (new_AGEMA_signal_5558) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U56 ( .A0_t (LED_128_Instance_subcells_out[61]), .A0_f (new_AGEMA_signal_4749), .A1_t (new_AGEMA_signal_4750), .A1_f (new_AGEMA_signal_4751), .B0_t (LED_128_Instance_MCS_Instance_0_n40), .B0_f (new_AGEMA_signal_5322), .B1_t (new_AGEMA_signal_5323), .B1_f (new_AGEMA_signal_5324), .Z0_t (LED_128_Instance_mixcolumns_out[18]), .Z0_f (new_AGEMA_signal_5559), .Z1_t (new_AGEMA_signal_5560), .Z1_f (new_AGEMA_signal_5561) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U55 ( .A0_t (LED_128_Instance_MCS_Instance_0_n39), .A0_f (new_AGEMA_signal_5142), .A1_t (new_AGEMA_signal_5143), .A1_f (new_AGEMA_signal_5144), .B0_t (LED_128_Instance_MCS_Instance_0_n42), .B0_f (new_AGEMA_signal_5139), .B1_t (new_AGEMA_signal_5140), .B1_f (new_AGEMA_signal_5141), .Z0_t (LED_128_Instance_MCS_Instance_0_n40), .Z0_f (new_AGEMA_signal_5322), .Z1_t (new_AGEMA_signal_5323), .Z1_f (new_AGEMA_signal_5324) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U54 ( .A0_t (LED_128_Instance_MCS_Instance_0_n38), .A0_f (new_AGEMA_signal_5004), .A1_t (new_AGEMA_signal_5005), .A1_f (new_AGEMA_signal_5006), .B0_t (LED_128_Instance_MCS_Instance_0_n37), .B0_f (new_AGEMA_signal_4905), .B1_t (new_AGEMA_signal_4906), .B1_f (new_AGEMA_signal_4907), .Z0_t (LED_128_Instance_MCS_Instance_0_n42), .Z0_f (new_AGEMA_signal_5139), .Z1_t (new_AGEMA_signal_5140), .Z1_f (new_AGEMA_signal_5141) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U53 ( .A0_t (LED_128_Instance_MCS_Instance_0_n36), .A0_f (new_AGEMA_signal_5016), .A1_t (new_AGEMA_signal_5017), .A1_f (new_AGEMA_signal_5018), .B0_t (LED_128_Instance_MCS_Instance_0_n35), .B0_f (new_AGEMA_signal_4839), .B1_t (new_AGEMA_signal_4840), .B1_f (new_AGEMA_signal_4841), .Z0_t (LED_128_Instance_MCS_Instance_0_n39), .Z0_f (new_AGEMA_signal_5142), .Z1_t (new_AGEMA_signal_5143), .Z1_f (new_AGEMA_signal_5144) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U52 ( .A0_t (LED_128_Instance_MCS_Instance_0_n34), .A0_f (new_AGEMA_signal_5145), .A1_t (new_AGEMA_signal_5146), .A1_f (new_AGEMA_signal_5147), .B0_t (LED_128_Instance_MCS_Instance_0_n36), .B0_f (new_AGEMA_signal_5016), .B1_t (new_AGEMA_signal_5017), .B1_f (new_AGEMA_signal_5018), .Z0_t (LED_128_Instance_mixcolumns_out[35]), .Z0_f (new_AGEMA_signal_5325), .Z1_t (new_AGEMA_signal_5326), .Z1_f (new_AGEMA_signal_5327) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U51 ( .A0_t (LED_128_Instance_MCS_Instance_0_n33), .A0_f (new_AGEMA_signal_4995), .A1_t (new_AGEMA_signal_4996), .A1_f (new_AGEMA_signal_4997), .B0_t (LED_128_Instance_MCS_Instance_0_n32), .B0_f (new_AGEMA_signal_4992), .B1_t (new_AGEMA_signal_4993), .B1_f (new_AGEMA_signal_4994), .Z0_t (LED_128_Instance_MCS_Instance_0_n34), .Z0_f (new_AGEMA_signal_5145), .Z1_t (new_AGEMA_signal_5146), .Z1_f (new_AGEMA_signal_5147) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U50 ( .A0_t (LED_128_Instance_MCS_Instance_0_n31), .A0_f (new_AGEMA_signal_4902), .A1_t (new_AGEMA_signal_4903), .A1_f (new_AGEMA_signal_4904), .B0_t (LED_128_Instance_subcells_out[22]), .B0_f (new_AGEMA_signal_4776), .B1_t (new_AGEMA_signal_4777), .B1_f (new_AGEMA_signal_4778), .Z0_t (LED_128_Instance_MCS_Instance_0_n32), .Z0_f (new_AGEMA_signal_4992), .Z1_t (new_AGEMA_signal_4993), .Z1_f (new_AGEMA_signal_4994) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U49 ( .A0_t (LED_128_Instance_MCS_Instance_0_n30), .A0_f (new_AGEMA_signal_4416), .A1_t (new_AGEMA_signal_4417), .A1_f (new_AGEMA_signal_4418), .B0_t (LED_128_Instance_MCS_Instance_0_n29), .B0_f (new_AGEMA_signal_4899), .B1_t (new_AGEMA_signal_4900), .B1_f (new_AGEMA_signal_4901), .Z0_t (LED_128_Instance_MCS_Instance_0_n33), .Z0_f (new_AGEMA_signal_4995), .Z1_t (new_AGEMA_signal_4996), .Z1_f (new_AGEMA_signal_4997) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U48 ( .A0_t (LED_128_Instance_MCS_Instance_0_n28), .A0_f (new_AGEMA_signal_4998), .A1_t (new_AGEMA_signal_4999), .A1_f (new_AGEMA_signal_5000), .B0_t (LED_128_Instance_MCS_Instance_0_n27), .B0_f (new_AGEMA_signal_5151), .B1_t (new_AGEMA_signal_5152), .B1_f (new_AGEMA_signal_5153), .Z0_t (LED_128_Instance_mixcolumns_out[34]), .Z0_f (new_AGEMA_signal_5328), .Z1_t (new_AGEMA_signal_5329), .Z1_f (new_AGEMA_signal_5330) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U47 ( .A0_t (LED_128_Instance_MCS_Instance_0_n26), .A0_f (new_AGEMA_signal_4917), .A1_t (new_AGEMA_signal_4918), .A1_f (new_AGEMA_signal_4919), .B0_t (LED_128_Instance_MCS_Instance_0_n25), .B0_f (new_AGEMA_signal_4824), .B1_t (new_AGEMA_signal_4825), .B1_f (new_AGEMA_signal_4826), .Z0_t (LED_128_Instance_MCS_Instance_0_n28), .Z0_f (new_AGEMA_signal_4998), .Z1_t (new_AGEMA_signal_4999), .Z1_f (new_AGEMA_signal_5000) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U46 ( .A0_t (LED_128_Instance_subcells_out[42]), .A0_f (new_AGEMA_signal_4704), .A1_t (new_AGEMA_signal_4705), .A1_f (new_AGEMA_signal_4706), .B0_t (LED_128_Instance_subcells_out[20]), .B0_f (new_AGEMA_signal_4335), .B1_t (new_AGEMA_signal_4336), .B1_f (new_AGEMA_signal_4337), .Z0_t (LED_128_Instance_MCS_Instance_0_n25), .Z0_f (new_AGEMA_signal_4824), .Z1_t (new_AGEMA_signal_4825), .Z1_f (new_AGEMA_signal_4826) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U45 ( .A0_t (LED_128_Instance_MCS_Instance_0_n24), .A0_f (new_AGEMA_signal_5331), .A1_t (new_AGEMA_signal_5332), .A1_f (new_AGEMA_signal_5333), .B0_t (LED_128_Instance_MCS_Instance_0_n23), .B0_f (new_AGEMA_signal_4833), .B1_t (new_AGEMA_signal_4834), .B1_f (new_AGEMA_signal_4835), .Z0_t (LED_128_Instance_mixcolumns_out[33]), .Z0_f (new_AGEMA_signal_5562), .Z1_t (new_AGEMA_signal_5563), .Z1_f (new_AGEMA_signal_5564) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U44 ( .A0_t (LED_128_Instance_MCS_Instance_0_n22), .A0_f (new_AGEMA_signal_5001), .A1_t (new_AGEMA_signal_5002), .A1_f (new_AGEMA_signal_5003), .B0_t (LED_128_Instance_MCS_Instance_0_n21), .B0_f (new_AGEMA_signal_5148), .B1_t (new_AGEMA_signal_5149), .B1_f (new_AGEMA_signal_5150), .Z0_t (LED_128_Instance_MCS_Instance_0_n24), .Z0_f (new_AGEMA_signal_5331), .Z1_t (new_AGEMA_signal_5332), .Z1_f (new_AGEMA_signal_5333) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U43 ( .A0_t (LED_128_Instance_MCS_Instance_0_n38), .A0_f (new_AGEMA_signal_5004), .A1_t (new_AGEMA_signal_5005), .A1_f (new_AGEMA_signal_5006), .B0_t (LED_128_Instance_subcells_out[41]), .B0_f (new_AGEMA_signal_4707), .B1_t (new_AGEMA_signal_4708), .B1_f (new_AGEMA_signal_4709), .Z0_t (LED_128_Instance_MCS_Instance_0_n21), .Z0_f (new_AGEMA_signal_5148), .Z1_t (new_AGEMA_signal_5149), .Z1_f (new_AGEMA_signal_5150) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U42 ( .A0_t (LED_128_Instance_MCS_Instance_0_n29), .A0_f (new_AGEMA_signal_4899), .A1_t (new_AGEMA_signal_4900), .A1_f (new_AGEMA_signal_4901), .B0_t (LED_128_Instance_subcells_out[40]), .B0_f (new_AGEMA_signal_4206), .B1_t (new_AGEMA_signal_4207), .B1_f (new_AGEMA_signal_4208), .Z0_t (LED_128_Instance_MCS_Instance_0_n22), .Z0_f (new_AGEMA_signal_5001), .Z1_t (new_AGEMA_signal_5002), .Z1_f (new_AGEMA_signal_5003) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U41 ( .A0_t (LED_128_Instance_subcells_out[0]), .A0_f (new_AGEMA_signal_4056), .A1_t (new_AGEMA_signal_4057), .A1_f (new_AGEMA_signal_4058), .B0_t (LED_128_Instance_MCS_Instance_0_n35), .B0_f (new_AGEMA_signal_4839), .B1_t (new_AGEMA_signal_4840), .B1_f (new_AGEMA_signal_4841), .Z0_t (LED_128_Instance_MCS_Instance_0_n29), .Z0_f (new_AGEMA_signal_4899), .Z1_t (new_AGEMA_signal_4900), .Z1_f (new_AGEMA_signal_4901) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U40 ( .A0_t (LED_128_Instance_MCS_Instance_0_n20), .A0_f (new_AGEMA_signal_5565), .A1_t (new_AGEMA_signal_5566), .A1_f (new_AGEMA_signal_5567), .B0_t (LED_128_Instance_MCS_Instance_0_n19), .B0_f (new_AGEMA_signal_4836), .B1_t (new_AGEMA_signal_4837), .B1_f (new_AGEMA_signal_4838), .Z0_t (LED_128_Instance_mixcolumns_out[32]), .Z0_f (new_AGEMA_signal_5820), .Z1_t (new_AGEMA_signal_5821), .Z1_f (new_AGEMA_signal_5822) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U39 ( .A0_t (LED_128_Instance_MCS_Instance_0_n41), .A0_f (new_AGEMA_signal_5334), .A1_t (new_AGEMA_signal_5335), .A1_f (new_AGEMA_signal_5336), .B0_t (LED_128_Instance_subcells_out[23]), .B0_f (new_AGEMA_signal_4890), .B1_t (new_AGEMA_signal_4891), .B1_f (new_AGEMA_signal_4892), .Z0_t (LED_128_Instance_MCS_Instance_0_n20), .Z0_f (new_AGEMA_signal_5565), .Z1_t (new_AGEMA_signal_5566), .Z1_f (new_AGEMA_signal_5567) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U38 ( .A0_t (LED_128_Instance_MCS_Instance_0_n18), .A0_f (new_AGEMA_signal_4830), .A1_t (new_AGEMA_signal_4831), .A1_f (new_AGEMA_signal_4832), .B0_t (LED_128_Instance_MCS_Instance_0_n27), .B0_f (new_AGEMA_signal_5151), .B1_t (new_AGEMA_signal_5152), .B1_f (new_AGEMA_signal_5153), .Z0_t (LED_128_Instance_MCS_Instance_0_n41), .Z0_f (new_AGEMA_signal_5334), .Z1_t (new_AGEMA_signal_5335), .Z1_f (new_AGEMA_signal_5336) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U37 ( .A0_t (LED_128_Instance_MCS_Instance_0_n38), .A0_f (new_AGEMA_signal_5004), .A1_t (new_AGEMA_signal_5005), .A1_f (new_AGEMA_signal_5006), .B0_t (LED_128_Instance_MCS_Instance_0_n17), .B0_f (new_AGEMA_signal_4911), .B1_t (new_AGEMA_signal_4912), .B1_f (new_AGEMA_signal_4913), .Z0_t (LED_128_Instance_MCS_Instance_0_n27), .Z0_f (new_AGEMA_signal_5151), .Z1_t (new_AGEMA_signal_5152), .Z1_f (new_AGEMA_signal_5153) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U36 ( .A0_t (LED_128_Instance_subcells_out[3]), .A0_f (new_AGEMA_signal_4752), .A1_t (new_AGEMA_signal_4753), .A1_f (new_AGEMA_signal_4754), .B0_t (LED_128_Instance_MCS_Instance_0_n31), .B0_f (new_AGEMA_signal_4902), .B1_t (new_AGEMA_signal_4903), .B1_f (new_AGEMA_signal_4904), .Z0_t (LED_128_Instance_MCS_Instance_0_n38), .Z0_f (new_AGEMA_signal_5004), .Z1_t (new_AGEMA_signal_5005), .Z1_f (new_AGEMA_signal_5006) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U35 ( .A0_t (LED_128_Instance_subcells_out[43]), .A0_f (new_AGEMA_signal_4800), .A1_t (new_AGEMA_signal_4801), .A1_f (new_AGEMA_signal_4802), .B0_t (LED_128_Instance_subcells_out[21]), .B0_f (new_AGEMA_signal_4779), .B1_t (new_AGEMA_signal_4780), .B1_f (new_AGEMA_signal_4781), .Z0_t (LED_128_Instance_MCS_Instance_0_n31), .Z0_f (new_AGEMA_signal_4902), .Z1_t (new_AGEMA_signal_4903), .Z1_f (new_AGEMA_signal_4904) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U34 ( .A0_t (LED_128_Instance_MCS_Instance_0_n16), .A0_f (new_AGEMA_signal_5154), .A1_t (new_AGEMA_signal_5155), .A1_f (new_AGEMA_signal_5156), .B0_t (LED_128_Instance_MCS_Instance_0_n30), .B0_f (new_AGEMA_signal_4416), .B1_t (new_AGEMA_signal_4417), .B1_f (new_AGEMA_signal_4418), .Z0_t (LED_128_Instance_mixcolumns_out[51]), .Z0_f (new_AGEMA_signal_5337), .Z1_t (new_AGEMA_signal_5338), .Z1_f (new_AGEMA_signal_5339) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U33 ( .A0_t (LED_128_Instance_MCS_Instance_0_n15), .A0_f (new_AGEMA_signal_5013), .A1_t (new_AGEMA_signal_5014), .A1_f (new_AGEMA_signal_5015), .B0_t (LED_128_Instance_subcells_out[2]), .B0_f (new_AGEMA_signal_4623), .B1_t (new_AGEMA_signal_4624), .B1_f (new_AGEMA_signal_4625), .Z0_t (LED_128_Instance_MCS_Instance_0_n16), .Z0_f (new_AGEMA_signal_5154), .Z1_t (new_AGEMA_signal_5155), .Z1_f (new_AGEMA_signal_5156) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U32 ( .A0_t (LED_128_Instance_subcells_out[23]), .A0_f (new_AGEMA_signal_4890), .A1_t (new_AGEMA_signal_4891), .A1_f (new_AGEMA_signal_4892), .B0_t (LED_128_Instance_MCS_Instance_0_n14), .B0_f (new_AGEMA_signal_5340), .B1_t (new_AGEMA_signal_5341), .B1_f (new_AGEMA_signal_5342), .Z0_t (LED_128_Instance_mixcolumns_out[49]), .Z0_f (new_AGEMA_signal_5568), .Z1_t (new_AGEMA_signal_5569), .Z1_f (new_AGEMA_signal_5570) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U31 ( .A0_t (LED_128_Instance_MCS_Instance_0_n13), .A0_f (new_AGEMA_signal_5157), .A1_t (new_AGEMA_signal_5158), .A1_f (new_AGEMA_signal_5159), .B0_t (LED_128_Instance_MCS_Instance_0_n12), .B0_f (new_AGEMA_signal_4827), .B1_t (new_AGEMA_signal_4828), .B1_f (new_AGEMA_signal_4829), .Z0_t (LED_128_Instance_MCS_Instance_0_n14), .Z0_f (new_AGEMA_signal_5340), .Z1_t (new_AGEMA_signal_5341), .Z1_f (new_AGEMA_signal_5342) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U30 ( .A0_t (LED_128_Instance_subcells_out[0]), .A0_f (new_AGEMA_signal_4056), .A1_t (new_AGEMA_signal_4057), .A1_f (new_AGEMA_signal_4058), .B0_t (LED_128_Instance_subcells_out[62]), .B0_f (new_AGEMA_signal_4746), .B1_t (new_AGEMA_signal_4747), .B1_f (new_AGEMA_signal_4748), .Z0_t (LED_128_Instance_MCS_Instance_0_n12), .Z0_f (new_AGEMA_signal_4827), .Z1_t (new_AGEMA_signal_4828), .Z1_f (new_AGEMA_signal_4829) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U29 ( .A0_t (LED_128_Instance_MCS_Instance_0_n11), .A0_f (new_AGEMA_signal_5007), .A1_t (new_AGEMA_signal_5008), .A1_f (new_AGEMA_signal_5009), .B0_t (LED_128_Instance_subcells_out[20]), .B0_f (new_AGEMA_signal_4335), .B1_t (new_AGEMA_signal_4336), .B1_f (new_AGEMA_signal_4337), .Z0_t (LED_128_Instance_MCS_Instance_0_n13), .Z0_f (new_AGEMA_signal_5157), .Z1_t (new_AGEMA_signal_5158), .Z1_f (new_AGEMA_signal_5159) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U28 ( .A0_t (LED_128_Instance_subcells_out[43]), .A0_f (new_AGEMA_signal_4800), .A1_t (new_AGEMA_signal_4801), .A1_f (new_AGEMA_signal_4802), .B0_t (LED_128_Instance_MCS_Instance_0_n10), .B0_f (new_AGEMA_signal_5343), .B1_t (new_AGEMA_signal_5344), .B1_f (new_AGEMA_signal_5345), .Z0_t (LED_128_Instance_mixcolumns_out[48]), .Z0_f (new_AGEMA_signal_5571), .Z1_t (new_AGEMA_signal_5572), .Z1_f (new_AGEMA_signal_5573) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U27 ( .A0_t (LED_128_Instance_MCS_Instance_0_n9), .A0_f (new_AGEMA_signal_5160), .A1_t (new_AGEMA_signal_5161), .A1_f (new_AGEMA_signal_5162), .B0_t (LED_128_Instance_MCS_Instance_0_n36), .B0_f (new_AGEMA_signal_5016), .B1_t (new_AGEMA_signal_5017), .B1_f (new_AGEMA_signal_5018), .Z0_t (LED_128_Instance_MCS_Instance_0_n10), .Z0_f (new_AGEMA_signal_5343), .Z1_t (new_AGEMA_signal_5344), .Z1_f (new_AGEMA_signal_5345) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U26 ( .A0_t (LED_128_Instance_MCS_Instance_0_n11), .A0_f (new_AGEMA_signal_5007), .A1_t (new_AGEMA_signal_5008), .A1_f (new_AGEMA_signal_5009), .B0_t (LED_128_Instance_MCS_Instance_0_n8), .B0_f (new_AGEMA_signal_4842), .B1_t (new_AGEMA_signal_4843), .B1_f (new_AGEMA_signal_4844), .Z0_t (LED_128_Instance_MCS_Instance_0_n9), .Z0_f (new_AGEMA_signal_5160), .Z1_t (new_AGEMA_signal_5161), .Z1_f (new_AGEMA_signal_5162) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U25 ( .A0_t (LED_128_Instance_subcells_out[3]), .A0_f (new_AGEMA_signal_4752), .A1_t (new_AGEMA_signal_4753), .A1_f (new_AGEMA_signal_4754), .B0_t (LED_128_Instance_MCS_Instance_0_n37), .B0_f (new_AGEMA_signal_4905), .B1_t (new_AGEMA_signal_4906), .B1_f (new_AGEMA_signal_4907), .Z0_t (LED_128_Instance_MCS_Instance_0_n11), .Z0_f (new_AGEMA_signal_5007), .Z1_t (new_AGEMA_signal_5008), .Z1_f (new_AGEMA_signal_5009) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U24 ( .A0_t (LED_128_Instance_subcells_out[63]), .A0_f (new_AGEMA_signal_4821), .A1_t (new_AGEMA_signal_4822), .A1_f (new_AGEMA_signal_4823), .B0_t (LED_128_Instance_MCS_Instance_0_n30), .B0_f (new_AGEMA_signal_4416), .B1_t (new_AGEMA_signal_4417), .B1_f (new_AGEMA_signal_4418), .Z0_t (LED_128_Instance_MCS_Instance_0_n37), .Z0_f (new_AGEMA_signal_4905), .Z1_t (new_AGEMA_signal_4906), .Z1_f (new_AGEMA_signal_4907) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U23 ( .A0_t (LED_128_Instance_subcells_out[60]), .A0_f (new_AGEMA_signal_4281), .A1_t (new_AGEMA_signal_4282), .A1_f (new_AGEMA_signal_4283), .B0_t (LED_128_Instance_subcells_out[40]), .B0_f (new_AGEMA_signal_4206), .B1_t (new_AGEMA_signal_4207), .B1_f (new_AGEMA_signal_4208), .Z0_t (LED_128_Instance_MCS_Instance_0_n30), .Z0_f (new_AGEMA_signal_4416), .Z1_t (new_AGEMA_signal_4417), .Z1_f (new_AGEMA_signal_4418) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U22 ( .A0_t (LED_128_Instance_MCS_Instance_0_n7), .A0_f (new_AGEMA_signal_4908), .A1_t (new_AGEMA_signal_4909), .A1_f (new_AGEMA_signal_4910), .B0_t (LED_128_Instance_MCS_Instance_0_n17), .B0_f (new_AGEMA_signal_4911), .B1_t (new_AGEMA_signal_4912), .B1_f (new_AGEMA_signal_4913), .Z0_t (LED_128_Instance_mixcolumns_out[2]), .Z0_f (new_AGEMA_signal_5010), .Z1_t (new_AGEMA_signal_5011), .Z1_f (new_AGEMA_signal_5012) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U21 ( .A0_t (LED_128_Instance_MCS_Instance_0_n18), .A0_f (new_AGEMA_signal_4830), .A1_t (new_AGEMA_signal_4831), .A1_f (new_AGEMA_signal_4832), .B0_t (LED_128_Instance_subcells_out[3]), .B0_f (new_AGEMA_signal_4752), .B1_t (new_AGEMA_signal_4753), .B1_f (new_AGEMA_signal_4754), .Z0_t (LED_128_Instance_MCS_Instance_0_n7), .Z0_f (new_AGEMA_signal_4908), .Z1_t (new_AGEMA_signal_4909), .Z1_f (new_AGEMA_signal_4910) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U20 ( .A0_t (LED_128_Instance_subcells_out[0]), .A0_f (new_AGEMA_signal_4056), .A1_t (new_AGEMA_signal_4057), .A1_f (new_AGEMA_signal_4058), .B0_t (LED_128_Instance_subcells_out[61]), .B0_f (new_AGEMA_signal_4749), .B1_t (new_AGEMA_signal_4750), .B1_f (new_AGEMA_signal_4751), .Z0_t (LED_128_Instance_MCS_Instance_0_n18), .Z0_f (new_AGEMA_signal_4830), .Z1_t (new_AGEMA_signal_4831), .Z1_f (new_AGEMA_signal_4832) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U19 ( .A0_t (LED_128_Instance_MCS_Instance_0_n6), .A0_f (new_AGEMA_signal_5163), .A1_t (new_AGEMA_signal_5164), .A1_f (new_AGEMA_signal_5165), .B0_t (LED_128_Instance_MCS_Instance_0_n5), .B0_f (new_AGEMA_signal_4914), .B1_t (new_AGEMA_signal_4915), .B1_f (new_AGEMA_signal_4916), .Z0_t (LED_128_Instance_mixcolumns_out[17]), .Z0_f (new_AGEMA_signal_5346), .Z1_t (new_AGEMA_signal_5347), .Z1_f (new_AGEMA_signal_5348) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U18 ( .A0_t (LED_128_Instance_MCS_Instance_0_n19), .A0_f (new_AGEMA_signal_4836), .A1_t (new_AGEMA_signal_4837), .A1_f (new_AGEMA_signal_4838), .B0_t (LED_128_Instance_MCS_Instance_0_n15), .B0_f (new_AGEMA_signal_5013), .B1_t (new_AGEMA_signal_5014), .B1_f (new_AGEMA_signal_5015), .Z0_t (LED_128_Instance_MCS_Instance_0_n6), .Z0_f (new_AGEMA_signal_5163), .Z1_t (new_AGEMA_signal_5164), .Z1_f (new_AGEMA_signal_5165) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U17 ( .A0_t (LED_128_Instance_MCS_Instance_0_n17), .A0_f (new_AGEMA_signal_4911), .A1_t (new_AGEMA_signal_4912), .A1_f (new_AGEMA_signal_4913), .B0_t (LED_128_Instance_MCS_Instance_0_n23), .B0_f (new_AGEMA_signal_4833), .B1_t (new_AGEMA_signal_4834), .B1_f (new_AGEMA_signal_4835), .Z0_t (LED_128_Instance_MCS_Instance_0_n15), .Z0_f (new_AGEMA_signal_5013), .Z1_t (new_AGEMA_signal_5014), .Z1_f (new_AGEMA_signal_5015) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U16 ( .A0_t (LED_128_Instance_subcells_out[62]), .A0_f (new_AGEMA_signal_4746), .A1_t (new_AGEMA_signal_4747), .A1_f (new_AGEMA_signal_4748), .B0_t (LED_128_Instance_subcells_out[42]), .B0_f (new_AGEMA_signal_4704), .B1_t (new_AGEMA_signal_4705), .B1_f (new_AGEMA_signal_4706), .Z0_t (LED_128_Instance_MCS_Instance_0_n23), .Z0_f (new_AGEMA_signal_4833), .Z1_t (new_AGEMA_signal_4834), .Z1_f (new_AGEMA_signal_4835) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U15 ( .A0_t (LED_128_Instance_subcells_out[41]), .A0_f (new_AGEMA_signal_4707), .A1_t (new_AGEMA_signal_4708), .A1_f (new_AGEMA_signal_4709), .B0_t (LED_128_Instance_subcells_out[22]), .B0_f (new_AGEMA_signal_4776), .B1_t (new_AGEMA_signal_4777), .B1_f (new_AGEMA_signal_4778), .Z0_t (LED_128_Instance_MCS_Instance_0_n17), .Z0_f (new_AGEMA_signal_4911), .Z1_t (new_AGEMA_signal_4912), .Z1_f (new_AGEMA_signal_4913) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U14 ( .A0_t (LED_128_Instance_subcells_out[60]), .A0_f (new_AGEMA_signal_4281), .A1_t (new_AGEMA_signal_4282), .A1_f (new_AGEMA_signal_4283), .B0_t (LED_128_Instance_subcells_out[1]), .B0_f (new_AGEMA_signal_4626), .B1_t (new_AGEMA_signal_4627), .B1_f (new_AGEMA_signal_4628), .Z0_t (LED_128_Instance_MCS_Instance_0_n19), .Z0_f (new_AGEMA_signal_4836), .Z1_t (new_AGEMA_signal_4837), .Z1_f (new_AGEMA_signal_4838) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U13 ( .A0_t (LED_128_Instance_subcells_out[1]), .A0_f (new_AGEMA_signal_4626), .A1_t (new_AGEMA_signal_4627), .A1_f (new_AGEMA_signal_4628), .B0_t (LED_128_Instance_MCS_Instance_0_n4), .B0_f (new_AGEMA_signal_5166), .B1_t (new_AGEMA_signal_5167), .B1_f (new_AGEMA_signal_5168), .Z0_t (LED_128_Instance_mixcolumns_out[3]), .Z0_f (new_AGEMA_signal_5349), .Z1_t (new_AGEMA_signal_5350), .Z1_f (new_AGEMA_signal_5351) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U12 ( .A0_t (LED_128_Instance_MCS_Instance_0_n3), .A0_f (new_AGEMA_signal_5352), .A1_t (new_AGEMA_signal_5353), .A1_f (new_AGEMA_signal_5354), .B0_t (LED_128_Instance_MCS_Instance_0_n2), .B0_f (new_AGEMA_signal_5022), .B1_t (new_AGEMA_signal_5023), .B1_f (new_AGEMA_signal_5024), .Z0_t (LED_128_Instance_mixcolumns_out[16]), .Z0_f (new_AGEMA_signal_5574), .Z1_t (new_AGEMA_signal_5575), .Z1_f (new_AGEMA_signal_5576) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U11 ( .A0_t (LED_128_Instance_subcells_out[22]), .A0_f (new_AGEMA_signal_4776), .A1_t (new_AGEMA_signal_4777), .A1_f (new_AGEMA_signal_4778), .B0_t (LED_128_Instance_MCS_Instance_0_n4), .B0_f (new_AGEMA_signal_5166), .B1_t (new_AGEMA_signal_5167), .B1_f (new_AGEMA_signal_5168), .Z0_t (LED_128_Instance_MCS_Instance_0_n3), .Z0_f (new_AGEMA_signal_5352), .Z1_t (new_AGEMA_signal_5353), .Z1_f (new_AGEMA_signal_5354) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U10 ( .A0_t (LED_128_Instance_subcells_out[62]), .A0_f (new_AGEMA_signal_4746), .A1_t (new_AGEMA_signal_4747), .A1_f (new_AGEMA_signal_4748), .B0_t (LED_128_Instance_MCS_Instance_0_n36), .B0_f (new_AGEMA_signal_5016), .B1_t (new_AGEMA_signal_5017), .B1_f (new_AGEMA_signal_5018), .Z0_t (LED_128_Instance_MCS_Instance_0_n4), .Z0_f (new_AGEMA_signal_5166), .Z1_t (new_AGEMA_signal_5167), .Z1_f (new_AGEMA_signal_5168) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U9 ( .A0_t (LED_128_Instance_subcells_out[23]), .A0_f (new_AGEMA_signal_4890), .A1_t (new_AGEMA_signal_4891), .A1_f (new_AGEMA_signal_4892), .B0_t (LED_128_Instance_subcells_out[42]), .B0_f (new_AGEMA_signal_4704), .B1_t (new_AGEMA_signal_4705), .B1_f (new_AGEMA_signal_4706), .Z0_t (LED_128_Instance_MCS_Instance_0_n36), .Z0_f (new_AGEMA_signal_5016), .Z1_t (new_AGEMA_signal_5017), .Z1_f (new_AGEMA_signal_5018) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U8 ( .A0_t (LED_128_Instance_subcells_out[63]), .A0_f (new_AGEMA_signal_4821), .A1_t (new_AGEMA_signal_4822), .A1_f (new_AGEMA_signal_4823), .B0_t (LED_128_Instance_MCS_Instance_0_n5), .B0_f (new_AGEMA_signal_4914), .B1_t (new_AGEMA_signal_4915), .B1_f (new_AGEMA_signal_4916), .Z0_t (LED_128_Instance_mixcolumns_out[0]), .Z0_f (new_AGEMA_signal_5019), .Z1_t (new_AGEMA_signal_5020), .Z1_f (new_AGEMA_signal_5021) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U7 ( .A0_t (LED_128_Instance_subcells_out[43]), .A0_f (new_AGEMA_signal_4800), .A1_t (new_AGEMA_signal_4801), .A1_f (new_AGEMA_signal_4802), .B0_t (LED_128_Instance_MCS_Instance_0_n35), .B0_f (new_AGEMA_signal_4839), .B1_t (new_AGEMA_signal_4840), .B1_f (new_AGEMA_signal_4841), .Z0_t (LED_128_Instance_MCS_Instance_0_n5), .Z0_f (new_AGEMA_signal_4914), .Z1_t (new_AGEMA_signal_4915), .Z1_f (new_AGEMA_signal_4916) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U6 ( .A0_t (LED_128_Instance_subcells_out[2]), .A0_f (new_AGEMA_signal_4623), .A1_t (new_AGEMA_signal_4624), .A1_f (new_AGEMA_signal_4625), .B0_t (LED_128_Instance_subcells_out[20]), .B0_f (new_AGEMA_signal_4335), .B1_t (new_AGEMA_signal_4336), .B1_f (new_AGEMA_signal_4337), .Z0_t (LED_128_Instance_MCS_Instance_0_n35), .Z0_f (new_AGEMA_signal_4839), .Z1_t (new_AGEMA_signal_4840), .Z1_f (new_AGEMA_signal_4841) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U5 ( .A0_t (LED_128_Instance_MCS_Instance_0_n1), .A0_f (new_AGEMA_signal_5169), .A1_t (new_AGEMA_signal_5170), .A1_f (new_AGEMA_signal_5171), .B0_t (LED_128_Instance_MCS_Instance_0_n8), .B0_f (new_AGEMA_signal_4842), .B1_t (new_AGEMA_signal_4843), .B1_f (new_AGEMA_signal_4844), .Z0_t (LED_128_Instance_mixcolumns_out[50]), .Z0_f (new_AGEMA_signal_5355), .Z1_t (new_AGEMA_signal_5356), .Z1_f (new_AGEMA_signal_5357) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U4 ( .A0_t (LED_128_Instance_subcells_out[61]), .A0_f (new_AGEMA_signal_4749), .A1_t (new_AGEMA_signal_4750), .A1_f (new_AGEMA_signal_4751), .B0_t (LED_128_Instance_subcells_out[41]), .B0_f (new_AGEMA_signal_4707), .B1_t (new_AGEMA_signal_4708), .B1_f (new_AGEMA_signal_4709), .Z0_t (LED_128_Instance_MCS_Instance_0_n8), .Z0_f (new_AGEMA_signal_4842), .Z1_t (new_AGEMA_signal_4843), .Z1_f (new_AGEMA_signal_4844) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U3 ( .A0_t (LED_128_Instance_subcells_out[21]), .A0_f (new_AGEMA_signal_4779), .A1_t (new_AGEMA_signal_4780), .A1_f (new_AGEMA_signal_4781), .B0_t (LED_128_Instance_MCS_Instance_0_n2), .B0_f (new_AGEMA_signal_5022), .B1_t (new_AGEMA_signal_5023), .B1_f (new_AGEMA_signal_5024), .Z0_t (LED_128_Instance_MCS_Instance_0_n1), .Z0_f (new_AGEMA_signal_5169), .Z1_t (new_AGEMA_signal_5170), .Z1_f (new_AGEMA_signal_5171) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U2 ( .A0_t (LED_128_Instance_subcells_out[40]), .A0_f (new_AGEMA_signal_4206), .A1_t (new_AGEMA_signal_4207), .A1_f (new_AGEMA_signal_4208), .B0_t (LED_128_Instance_MCS_Instance_0_n26), .B0_f (new_AGEMA_signal_4917), .B1_t (new_AGEMA_signal_4918), .B1_f (new_AGEMA_signal_4919), .Z0_t (LED_128_Instance_MCS_Instance_0_n2), .Z0_f (new_AGEMA_signal_5022), .Z1_t (new_AGEMA_signal_5023), .Z1_f (new_AGEMA_signal_5024) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_0_U1 ( .A0_t (LED_128_Instance_subcells_out[1]), .A0_f (new_AGEMA_signal_4626), .A1_t (new_AGEMA_signal_4627), .A1_f (new_AGEMA_signal_4628), .B0_t (LED_128_Instance_subcells_out[63]), .B0_f (new_AGEMA_signal_4821), .B1_t (new_AGEMA_signal_4822), .B1_f (new_AGEMA_signal_4823), .Z0_t (LED_128_Instance_MCS_Instance_0_n26), .Z0_f (new_AGEMA_signal_4917), .Z1_t (new_AGEMA_signal_4918), .Z1_f (new_AGEMA_signal_4919) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U58 ( .A0_t (LED_128_Instance_subcells_out[6]), .A0_f (new_AGEMA_signal_4758), .A1_t (new_AGEMA_signal_4759), .A1_f (new_AGEMA_signal_4760), .B0_t (LED_128_Instance_MCS_Instance_1_n42), .B0_f (new_AGEMA_signal_5172), .B1_t (new_AGEMA_signal_5173), .B1_f (new_AGEMA_signal_5174), .Z0_t (LED_128_Instance_mixcolumns_out[5]), .Z0_f (new_AGEMA_signal_5358), .Z1_t (new_AGEMA_signal_5359), .Z1_f (new_AGEMA_signal_5360) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U57 ( .A0_t (LED_128_Instance_MCS_Instance_1_n41), .A0_f (new_AGEMA_signal_5373), .A1_t (new_AGEMA_signal_5374), .A1_f (new_AGEMA_signal_5375), .B0_t (LED_128_Instance_subcells_out[50]), .B0_f (new_AGEMA_signal_4722), .B1_t (new_AGEMA_signal_4723), .B1_f (new_AGEMA_signal_4724), .Z0_t (LED_128_Instance_mixcolumns_out[23]), .Z0_f (new_AGEMA_signal_5577), .Z1_t (new_AGEMA_signal_5578), .Z1_f (new_AGEMA_signal_5579) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U56 ( .A0_t (LED_128_Instance_subcells_out[49]), .A0_f (new_AGEMA_signal_4725), .A1_t (new_AGEMA_signal_4726), .A1_f (new_AGEMA_signal_4727), .B0_t (LED_128_Instance_MCS_Instance_1_n40), .B0_f (new_AGEMA_signal_5361), .B1_t (new_AGEMA_signal_5362), .B1_f (new_AGEMA_signal_5363), .Z0_t (LED_128_Instance_mixcolumns_out[22]), .Z0_f (new_AGEMA_signal_5580), .Z1_t (new_AGEMA_signal_5581), .Z1_f (new_AGEMA_signal_5582) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U55 ( .A0_t (LED_128_Instance_MCS_Instance_1_n39), .A0_f (new_AGEMA_signal_5025), .A1_t (new_AGEMA_signal_5026), .A1_f (new_AGEMA_signal_5027), .B0_t (LED_128_Instance_MCS_Instance_1_n42), .B0_f (new_AGEMA_signal_5172), .B1_t (new_AGEMA_signal_5173), .B1_f (new_AGEMA_signal_5174), .Z0_t (LED_128_Instance_MCS_Instance_1_n40), .Z0_f (new_AGEMA_signal_5361), .Z1_t (new_AGEMA_signal_5362), .Z1_f (new_AGEMA_signal_5363) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U54 ( .A0_t (LED_128_Instance_MCS_Instance_1_n38), .A0_f (new_AGEMA_signal_5037), .A1_t (new_AGEMA_signal_5038), .A1_f (new_AGEMA_signal_5039), .B0_t (LED_128_Instance_MCS_Instance_1_n37), .B0_f (new_AGEMA_signal_4923), .B1_t (new_AGEMA_signal_4924), .B1_f (new_AGEMA_signal_4925), .Z0_t (LED_128_Instance_MCS_Instance_1_n42), .Z0_f (new_AGEMA_signal_5172), .Z1_t (new_AGEMA_signal_5173), .Z1_f (new_AGEMA_signal_5174) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U53 ( .A0_t (LED_128_Instance_MCS_Instance_1_n36), .A0_f (new_AGEMA_signal_4932), .A1_t (new_AGEMA_signal_4933), .A1_f (new_AGEMA_signal_4934), .B0_t (LED_128_Instance_MCS_Instance_1_n35), .B0_f (new_AGEMA_signal_4935), .B1_t (new_AGEMA_signal_4936), .B1_f (new_AGEMA_signal_4937), .Z0_t (LED_128_Instance_MCS_Instance_1_n39), .Z0_f (new_AGEMA_signal_5025), .Z1_t (new_AGEMA_signal_5026), .Z1_f (new_AGEMA_signal_5027) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U52 ( .A0_t (LED_128_Instance_MCS_Instance_1_n34), .A0_f (new_AGEMA_signal_5364), .A1_t (new_AGEMA_signal_5365), .A1_f (new_AGEMA_signal_5366), .B0_t (LED_128_Instance_MCS_Instance_1_n36), .B0_f (new_AGEMA_signal_4932), .B1_t (new_AGEMA_signal_4933), .B1_f (new_AGEMA_signal_4934), .Z0_t (LED_128_Instance_mixcolumns_out[39]), .Z0_f (new_AGEMA_signal_5583), .Z1_t (new_AGEMA_signal_5584), .Z1_f (new_AGEMA_signal_5585) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U51 ( .A0_t (LED_128_Instance_MCS_Instance_1_n33), .A0_f (new_AGEMA_signal_5175), .A1_t (new_AGEMA_signal_5176), .A1_f (new_AGEMA_signal_5177), .B0_t (LED_128_Instance_MCS_Instance_1_n32), .B0_f (new_AGEMA_signal_5028), .B1_t (new_AGEMA_signal_5029), .B1_f (new_AGEMA_signal_5030), .Z0_t (LED_128_Instance_MCS_Instance_1_n34), .Z0_f (new_AGEMA_signal_5364), .Z1_t (new_AGEMA_signal_5365), .Z1_f (new_AGEMA_signal_5366) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U50 ( .A0_t (LED_128_Instance_MCS_Instance_1_n31), .A0_f (new_AGEMA_signal_4920), .A1_t (new_AGEMA_signal_4921), .A1_f (new_AGEMA_signal_4922), .B0_t (LED_128_Instance_subcells_out[26]), .B0_f (new_AGEMA_signal_4671), .B1_t (new_AGEMA_signal_4672), .B1_f (new_AGEMA_signal_4673), .Z0_t (LED_128_Instance_MCS_Instance_1_n32), .Z0_f (new_AGEMA_signal_5028), .Z1_t (new_AGEMA_signal_5029), .Z1_f (new_AGEMA_signal_5030) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U49 ( .A0_t (LED_128_Instance_MCS_Instance_1_n30), .A0_f (new_AGEMA_signal_4419), .A1_t (new_AGEMA_signal_4420), .A1_f (new_AGEMA_signal_4421), .B0_t (LED_128_Instance_MCS_Instance_1_n29), .B0_f (new_AGEMA_signal_5034), .B1_t (new_AGEMA_signal_5035), .B1_f (new_AGEMA_signal_5036), .Z0_t (LED_128_Instance_MCS_Instance_1_n33), .Z0_f (new_AGEMA_signal_5175), .Z1_t (new_AGEMA_signal_5176), .Z1_f (new_AGEMA_signal_5177) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U48 ( .A0_t (LED_128_Instance_MCS_Instance_1_n28), .A0_f (new_AGEMA_signal_5031), .A1_t (new_AGEMA_signal_5032), .A1_f (new_AGEMA_signal_5033), .B0_t (LED_128_Instance_MCS_Instance_1_n27), .B0_f (new_AGEMA_signal_5184), .B1_t (new_AGEMA_signal_5185), .B1_f (new_AGEMA_signal_5186), .Z0_t (LED_128_Instance_mixcolumns_out[38]), .Z0_f (new_AGEMA_signal_5367), .Z1_t (new_AGEMA_signal_5368), .Z1_f (new_AGEMA_signal_5369) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U47 ( .A0_t (LED_128_Instance_MCS_Instance_1_n26), .A0_f (new_AGEMA_signal_4938), .A1_t (new_AGEMA_signal_4939), .A1_f (new_AGEMA_signal_4940), .B0_t (LED_128_Instance_MCS_Instance_1_n25), .B0_f (new_AGEMA_signal_4845), .B1_t (new_AGEMA_signal_4846), .B1_f (new_AGEMA_signal_4847), .Z0_t (LED_128_Instance_MCS_Instance_1_n28), .Z0_f (new_AGEMA_signal_5031), .Z1_t (new_AGEMA_signal_5032), .Z1_f (new_AGEMA_signal_5033) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U46 ( .A0_t (LED_128_Instance_subcells_out[46]), .A0_f (new_AGEMA_signal_4713), .A1_t (new_AGEMA_signal_4714), .A1_f (new_AGEMA_signal_4715), .B0_t (LED_128_Instance_subcells_out[24]), .B0_f (new_AGEMA_signal_4146), .B1_t (new_AGEMA_signal_4147), .B1_f (new_AGEMA_signal_4148), .Z0_t (LED_128_Instance_MCS_Instance_1_n25), .Z0_f (new_AGEMA_signal_4845), .Z1_t (new_AGEMA_signal_4846), .Z1_f (new_AGEMA_signal_4847) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U45 ( .A0_t (LED_128_Instance_MCS_Instance_1_n24), .A0_f (new_AGEMA_signal_5370), .A1_t (new_AGEMA_signal_5371), .A1_f (new_AGEMA_signal_5372), .B0_t (LED_128_Instance_MCS_Instance_1_n23), .B0_f (new_AGEMA_signal_4854), .B1_t (new_AGEMA_signal_4855), .B1_f (new_AGEMA_signal_4856), .Z0_t (LED_128_Instance_mixcolumns_out[37]), .Z0_f (new_AGEMA_signal_5586), .Z1_t (new_AGEMA_signal_5587), .Z1_f (new_AGEMA_signal_5588) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U44 ( .A0_t (LED_128_Instance_MCS_Instance_1_n22), .A0_f (new_AGEMA_signal_5181), .A1_t (new_AGEMA_signal_5182), .A1_f (new_AGEMA_signal_5183), .B0_t (LED_128_Instance_MCS_Instance_1_n21), .B0_f (new_AGEMA_signal_5178), .B1_t (new_AGEMA_signal_5179), .B1_f (new_AGEMA_signal_5180), .Z0_t (LED_128_Instance_MCS_Instance_1_n24), .Z0_f (new_AGEMA_signal_5370), .Z1_t (new_AGEMA_signal_5371), .Z1_f (new_AGEMA_signal_5372) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U43 ( .A0_t (LED_128_Instance_MCS_Instance_1_n38), .A0_f (new_AGEMA_signal_5037), .A1_t (new_AGEMA_signal_5038), .A1_f (new_AGEMA_signal_5039), .B0_t (LED_128_Instance_subcells_out[45]), .B0_f (new_AGEMA_signal_4716), .B1_t (new_AGEMA_signal_4717), .B1_f (new_AGEMA_signal_4718), .Z0_t (LED_128_Instance_MCS_Instance_1_n21), .Z0_f (new_AGEMA_signal_5178), .Z1_t (new_AGEMA_signal_5179), .Z1_f (new_AGEMA_signal_5180) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U42 ( .A0_t (LED_128_Instance_MCS_Instance_1_n29), .A0_f (new_AGEMA_signal_5034), .A1_t (new_AGEMA_signal_5035), .A1_f (new_AGEMA_signal_5036), .B0_t (LED_128_Instance_subcells_out[44]), .B0_f (new_AGEMA_signal_4221), .B1_t (new_AGEMA_signal_4222), .B1_f (new_AGEMA_signal_4223), .Z0_t (LED_128_Instance_MCS_Instance_1_n22), .Z0_f (new_AGEMA_signal_5181), .Z1_t (new_AGEMA_signal_5182), .Z1_f (new_AGEMA_signal_5183) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U41 ( .A0_t (LED_128_Instance_subcells_out[4]), .A0_f (new_AGEMA_signal_4302), .A1_t (new_AGEMA_signal_4303), .A1_f (new_AGEMA_signal_4304), .B0_t (LED_128_Instance_MCS_Instance_1_n35), .B0_f (new_AGEMA_signal_4935), .B1_t (new_AGEMA_signal_4936), .B1_f (new_AGEMA_signal_4937), .Z0_t (LED_128_Instance_MCS_Instance_1_n29), .Z0_f (new_AGEMA_signal_5034), .Z1_t (new_AGEMA_signal_5035), .Z1_f (new_AGEMA_signal_5036) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U40 ( .A0_t (LED_128_Instance_MCS_Instance_1_n20), .A0_f (new_AGEMA_signal_5589), .A1_t (new_AGEMA_signal_5590), .A1_f (new_AGEMA_signal_5591), .B0_t (LED_128_Instance_MCS_Instance_1_n19), .B0_f (new_AGEMA_signal_4929), .B1_t (new_AGEMA_signal_4930), .B1_f (new_AGEMA_signal_4931), .Z0_t (LED_128_Instance_mixcolumns_out[36]), .Z0_f (new_AGEMA_signal_5823), .Z1_t (new_AGEMA_signal_5824), .Z1_f (new_AGEMA_signal_5825) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U39 ( .A0_t (LED_128_Instance_MCS_Instance_1_n41), .A0_f (new_AGEMA_signal_5373), .A1_t (new_AGEMA_signal_5374), .A1_f (new_AGEMA_signal_5375), .B0_t (LED_128_Instance_subcells_out[27]), .B0_f (new_AGEMA_signal_4782), .B1_t (new_AGEMA_signal_4783), .B1_f (new_AGEMA_signal_4784), .Z0_t (LED_128_Instance_MCS_Instance_1_n20), .Z0_f (new_AGEMA_signal_5589), .Z1_t (new_AGEMA_signal_5590), .Z1_f (new_AGEMA_signal_5591) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U38 ( .A0_t (LED_128_Instance_MCS_Instance_1_n18), .A0_f (new_AGEMA_signal_4851), .A1_t (new_AGEMA_signal_4852), .A1_f (new_AGEMA_signal_4853), .B0_t (LED_128_Instance_MCS_Instance_1_n27), .B0_f (new_AGEMA_signal_5184), .B1_t (new_AGEMA_signal_5185), .B1_f (new_AGEMA_signal_5186), .Z0_t (LED_128_Instance_MCS_Instance_1_n41), .Z0_f (new_AGEMA_signal_5373), .Z1_t (new_AGEMA_signal_5374), .Z1_f (new_AGEMA_signal_5375) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U37 ( .A0_t (LED_128_Instance_MCS_Instance_1_n38), .A0_f (new_AGEMA_signal_5037), .A1_t (new_AGEMA_signal_5038), .A1_f (new_AGEMA_signal_5039), .B0_t (LED_128_Instance_MCS_Instance_1_n17), .B0_f (new_AGEMA_signal_4857), .B1_t (new_AGEMA_signal_4858), .B1_f (new_AGEMA_signal_4859), .Z0_t (LED_128_Instance_MCS_Instance_1_n27), .Z0_f (new_AGEMA_signal_5184), .Z1_t (new_AGEMA_signal_5185), .Z1_f (new_AGEMA_signal_5186) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U36 ( .A0_t (LED_128_Instance_subcells_out[7]), .A0_f (new_AGEMA_signal_4887), .A1_t (new_AGEMA_signal_4888), .A1_f (new_AGEMA_signal_4889), .B0_t (LED_128_Instance_MCS_Instance_1_n31), .B0_f (new_AGEMA_signal_4920), .B1_t (new_AGEMA_signal_4921), .B1_f (new_AGEMA_signal_4922), .Z0_t (LED_128_Instance_MCS_Instance_1_n38), .Z0_f (new_AGEMA_signal_5037), .Z1_t (new_AGEMA_signal_5038), .Z1_f (new_AGEMA_signal_5039) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U35 ( .A0_t (LED_128_Instance_subcells_out[47]), .A0_f (new_AGEMA_signal_4803), .A1_t (new_AGEMA_signal_4804), .A1_f (new_AGEMA_signal_4805), .B0_t (LED_128_Instance_subcells_out[25]), .B0_f (new_AGEMA_signal_4674), .B1_t (new_AGEMA_signal_4675), .B1_f (new_AGEMA_signal_4676), .Z0_t (LED_128_Instance_MCS_Instance_1_n31), .Z0_f (new_AGEMA_signal_4920), .Z1_t (new_AGEMA_signal_4921), .Z1_f (new_AGEMA_signal_4922) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U34 ( .A0_t (LED_128_Instance_MCS_Instance_1_n16), .A0_f (new_AGEMA_signal_5040), .A1_t (new_AGEMA_signal_5041), .A1_f (new_AGEMA_signal_5042), .B0_t (LED_128_Instance_MCS_Instance_1_n30), .B0_f (new_AGEMA_signal_4419), .B1_t (new_AGEMA_signal_4420), .B1_f (new_AGEMA_signal_4421), .Z0_t (LED_128_Instance_mixcolumns_out[55]), .Z0_f (new_AGEMA_signal_5187), .Z1_t (new_AGEMA_signal_5188), .Z1_f (new_AGEMA_signal_5189) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U33 ( .A0_t (LED_128_Instance_MCS_Instance_1_n15), .A0_f (new_AGEMA_signal_4926), .A1_t (new_AGEMA_signal_4927), .A1_f (new_AGEMA_signal_4928), .B0_t (LED_128_Instance_subcells_out[6]), .B0_f (new_AGEMA_signal_4758), .B1_t (new_AGEMA_signal_4759), .B1_f (new_AGEMA_signal_4760), .Z0_t (LED_128_Instance_MCS_Instance_1_n16), .Z0_f (new_AGEMA_signal_5040), .Z1_t (new_AGEMA_signal_5041), .Z1_f (new_AGEMA_signal_5042) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U32 ( .A0_t (LED_128_Instance_subcells_out[27]), .A0_f (new_AGEMA_signal_4782), .A1_t (new_AGEMA_signal_4783), .A1_f (new_AGEMA_signal_4784), .B0_t (LED_128_Instance_MCS_Instance_1_n14), .B0_f (new_AGEMA_signal_5376), .B1_t (new_AGEMA_signal_5377), .B1_f (new_AGEMA_signal_5378), .Z0_t (LED_128_Instance_mixcolumns_out[53]), .Z0_f (new_AGEMA_signal_5592), .Z1_t (new_AGEMA_signal_5593), .Z1_f (new_AGEMA_signal_5594) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U31 ( .A0_t (LED_128_Instance_MCS_Instance_1_n13), .A0_f (new_AGEMA_signal_5190), .A1_t (new_AGEMA_signal_5191), .A1_f (new_AGEMA_signal_5192), .B0_t (LED_128_Instance_MCS_Instance_1_n12), .B0_f (new_AGEMA_signal_4848), .B1_t (new_AGEMA_signal_4849), .B1_f (new_AGEMA_signal_4850), .Z0_t (LED_128_Instance_MCS_Instance_1_n14), .Z0_f (new_AGEMA_signal_5376), .Z1_t (new_AGEMA_signal_5377), .Z1_f (new_AGEMA_signal_5378) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U30 ( .A0_t (LED_128_Instance_subcells_out[4]), .A0_f (new_AGEMA_signal_4302), .A1_t (new_AGEMA_signal_4303), .A1_f (new_AGEMA_signal_4304), .B0_t (LED_128_Instance_subcells_out[50]), .B0_f (new_AGEMA_signal_4722), .B1_t (new_AGEMA_signal_4723), .B1_f (new_AGEMA_signal_4724), .Z0_t (LED_128_Instance_MCS_Instance_1_n12), .Z0_f (new_AGEMA_signal_4848), .Z1_t (new_AGEMA_signal_4849), .Z1_f (new_AGEMA_signal_4850) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U29 ( .A0_t (LED_128_Instance_MCS_Instance_1_n11), .A0_f (new_AGEMA_signal_5043), .A1_t (new_AGEMA_signal_5044), .A1_f (new_AGEMA_signal_5045), .B0_t (LED_128_Instance_subcells_out[24]), .B0_f (new_AGEMA_signal_4146), .B1_t (new_AGEMA_signal_4147), .B1_f (new_AGEMA_signal_4148), .Z0_t (LED_128_Instance_MCS_Instance_1_n13), .Z0_f (new_AGEMA_signal_5190), .Z1_t (new_AGEMA_signal_5191), .Z1_f (new_AGEMA_signal_5192) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U28 ( .A0_t (LED_128_Instance_subcells_out[47]), .A0_f (new_AGEMA_signal_4803), .A1_t (new_AGEMA_signal_4804), .A1_f (new_AGEMA_signal_4805), .B0_t (LED_128_Instance_MCS_Instance_1_n10), .B0_f (new_AGEMA_signal_5379), .B1_t (new_AGEMA_signal_5380), .B1_f (new_AGEMA_signal_5381), .Z0_t (LED_128_Instance_mixcolumns_out[52]), .Z0_f (new_AGEMA_signal_5595), .Z1_t (new_AGEMA_signal_5596), .Z1_f (new_AGEMA_signal_5597) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U27 ( .A0_t (LED_128_Instance_MCS_Instance_1_n9), .A0_f (new_AGEMA_signal_5193), .A1_t (new_AGEMA_signal_5194), .A1_f (new_AGEMA_signal_5195), .B0_t (LED_128_Instance_MCS_Instance_1_n36), .B0_f (new_AGEMA_signal_4932), .B1_t (new_AGEMA_signal_4933), .B1_f (new_AGEMA_signal_4934), .Z0_t (LED_128_Instance_MCS_Instance_1_n10), .Z0_f (new_AGEMA_signal_5379), .Z1_t (new_AGEMA_signal_5380), .Z1_f (new_AGEMA_signal_5381) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U26 ( .A0_t (LED_128_Instance_MCS_Instance_1_n11), .A0_f (new_AGEMA_signal_5043), .A1_t (new_AGEMA_signal_5044), .A1_f (new_AGEMA_signal_5045), .B0_t (LED_128_Instance_MCS_Instance_1_n8), .B0_f (new_AGEMA_signal_4860), .B1_t (new_AGEMA_signal_4861), .B1_f (new_AGEMA_signal_4862), .Z0_t (LED_128_Instance_MCS_Instance_1_n9), .Z0_f (new_AGEMA_signal_5193), .Z1_t (new_AGEMA_signal_5194), .Z1_f (new_AGEMA_signal_5195) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U25 ( .A0_t (LED_128_Instance_subcells_out[7]), .A0_f (new_AGEMA_signal_4887), .A1_t (new_AGEMA_signal_4888), .A1_f (new_AGEMA_signal_4889), .B0_t (LED_128_Instance_MCS_Instance_1_n37), .B0_f (new_AGEMA_signal_4923), .B1_t (new_AGEMA_signal_4924), .B1_f (new_AGEMA_signal_4925), .Z0_t (LED_128_Instance_MCS_Instance_1_n11), .Z0_f (new_AGEMA_signal_5043), .Z1_t (new_AGEMA_signal_5044), .Z1_f (new_AGEMA_signal_5045) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U24 ( .A0_t (LED_128_Instance_subcells_out[51]), .A0_f (new_AGEMA_signal_4806), .A1_t (new_AGEMA_signal_4807), .A1_f (new_AGEMA_signal_4808), .B0_t (LED_128_Instance_MCS_Instance_1_n30), .B0_f (new_AGEMA_signal_4419), .B1_t (new_AGEMA_signal_4420), .B1_f (new_AGEMA_signal_4421), .Z0_t (LED_128_Instance_MCS_Instance_1_n37), .Z0_f (new_AGEMA_signal_4923), .Z1_t (new_AGEMA_signal_4924), .Z1_f (new_AGEMA_signal_4925) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U23 ( .A0_t (LED_128_Instance_subcells_out[48]), .A0_f (new_AGEMA_signal_4236), .A1_t (new_AGEMA_signal_4237), .A1_f (new_AGEMA_signal_4238), .B0_t (LED_128_Instance_subcells_out[44]), .B0_f (new_AGEMA_signal_4221), .B1_t (new_AGEMA_signal_4222), .B1_f (new_AGEMA_signal_4223), .Z0_t (LED_128_Instance_MCS_Instance_1_n30), .Z0_f (new_AGEMA_signal_4419), .Z1_t (new_AGEMA_signal_4420), .Z1_f (new_AGEMA_signal_4421) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U22 ( .A0_t (LED_128_Instance_MCS_Instance_1_n7), .A0_f (new_AGEMA_signal_5046), .A1_t (new_AGEMA_signal_5047), .A1_f (new_AGEMA_signal_5048), .B0_t (LED_128_Instance_MCS_Instance_1_n17), .B0_f (new_AGEMA_signal_4857), .B1_t (new_AGEMA_signal_4858), .B1_f (new_AGEMA_signal_4859), .Z0_t (LED_128_Instance_mixcolumns_out[6]), .Z0_f (new_AGEMA_signal_5196), .Z1_t (new_AGEMA_signal_5197), .Z1_f (new_AGEMA_signal_5198) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U21 ( .A0_t (LED_128_Instance_MCS_Instance_1_n18), .A0_f (new_AGEMA_signal_4851), .A1_t (new_AGEMA_signal_4852), .A1_f (new_AGEMA_signal_4853), .B0_t (LED_128_Instance_subcells_out[7]), .B0_f (new_AGEMA_signal_4887), .B1_t (new_AGEMA_signal_4888), .B1_f (new_AGEMA_signal_4889), .Z0_t (LED_128_Instance_MCS_Instance_1_n7), .Z0_f (new_AGEMA_signal_5046), .Z1_t (new_AGEMA_signal_5047), .Z1_f (new_AGEMA_signal_5048) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U20 ( .A0_t (LED_128_Instance_subcells_out[4]), .A0_f (new_AGEMA_signal_4302), .A1_t (new_AGEMA_signal_4303), .A1_f (new_AGEMA_signal_4304), .B0_t (LED_128_Instance_subcells_out[49]), .B0_f (new_AGEMA_signal_4725), .B1_t (new_AGEMA_signal_4726), .B1_f (new_AGEMA_signal_4727), .Z0_t (LED_128_Instance_MCS_Instance_1_n18), .Z0_f (new_AGEMA_signal_4851), .Z1_t (new_AGEMA_signal_4852), .Z1_f (new_AGEMA_signal_4853) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U19 ( .A0_t (LED_128_Instance_MCS_Instance_1_n6), .A0_f (new_AGEMA_signal_5049), .A1_t (new_AGEMA_signal_5050), .A1_f (new_AGEMA_signal_5051), .B0_t (LED_128_Instance_MCS_Instance_1_n5), .B0_f (new_AGEMA_signal_5055), .B1_t (new_AGEMA_signal_5056), .B1_f (new_AGEMA_signal_5057), .Z0_t (LED_128_Instance_mixcolumns_out[21]), .Z0_f (new_AGEMA_signal_5199), .Z1_t (new_AGEMA_signal_5200), .Z1_f (new_AGEMA_signal_5201) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U18 ( .A0_t (LED_128_Instance_MCS_Instance_1_n19), .A0_f (new_AGEMA_signal_4929), .A1_t (new_AGEMA_signal_4930), .A1_f (new_AGEMA_signal_4931), .B0_t (LED_128_Instance_MCS_Instance_1_n15), .B0_f (new_AGEMA_signal_4926), .B1_t (new_AGEMA_signal_4927), .B1_f (new_AGEMA_signal_4928), .Z0_t (LED_128_Instance_MCS_Instance_1_n6), .Z0_f (new_AGEMA_signal_5049), .Z1_t (new_AGEMA_signal_5050), .Z1_f (new_AGEMA_signal_5051) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U17 ( .A0_t (LED_128_Instance_MCS_Instance_1_n17), .A0_f (new_AGEMA_signal_4857), .A1_t (new_AGEMA_signal_4858), .A1_f (new_AGEMA_signal_4859), .B0_t (LED_128_Instance_MCS_Instance_1_n23), .B0_f (new_AGEMA_signal_4854), .B1_t (new_AGEMA_signal_4855), .B1_f (new_AGEMA_signal_4856), .Z0_t (LED_128_Instance_MCS_Instance_1_n15), .Z0_f (new_AGEMA_signal_4926), .Z1_t (new_AGEMA_signal_4927), .Z1_f (new_AGEMA_signal_4928) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U16 ( .A0_t (LED_128_Instance_subcells_out[50]), .A0_f (new_AGEMA_signal_4722), .A1_t (new_AGEMA_signal_4723), .A1_f (new_AGEMA_signal_4724), .B0_t (LED_128_Instance_subcells_out[46]), .B0_f (new_AGEMA_signal_4713), .B1_t (new_AGEMA_signal_4714), .B1_f (new_AGEMA_signal_4715), .Z0_t (LED_128_Instance_MCS_Instance_1_n23), .Z0_f (new_AGEMA_signal_4854), .Z1_t (new_AGEMA_signal_4855), .Z1_f (new_AGEMA_signal_4856) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U15 ( .A0_t (LED_128_Instance_subcells_out[45]), .A0_f (new_AGEMA_signal_4716), .A1_t (new_AGEMA_signal_4717), .A1_f (new_AGEMA_signal_4718), .B0_t (LED_128_Instance_subcells_out[26]), .B0_f (new_AGEMA_signal_4671), .B1_t (new_AGEMA_signal_4672), .B1_f (new_AGEMA_signal_4673), .Z0_t (LED_128_Instance_MCS_Instance_1_n17), .Z0_f (new_AGEMA_signal_4857), .Z1_t (new_AGEMA_signal_4858), .Z1_f (new_AGEMA_signal_4859) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U14 ( .A0_t (LED_128_Instance_subcells_out[48]), .A0_f (new_AGEMA_signal_4236), .A1_t (new_AGEMA_signal_4237), .A1_f (new_AGEMA_signal_4238), .B0_t (LED_128_Instance_subcells_out[5]), .B0_f (new_AGEMA_signal_4761), .B1_t (new_AGEMA_signal_4762), .B1_f (new_AGEMA_signal_4763), .Z0_t (LED_128_Instance_MCS_Instance_1_n19), .Z0_f (new_AGEMA_signal_4929), .Z1_t (new_AGEMA_signal_4930), .Z1_f (new_AGEMA_signal_4931) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U13 ( .A0_t (LED_128_Instance_subcells_out[5]), .A0_f (new_AGEMA_signal_4761), .A1_t (new_AGEMA_signal_4762), .A1_f (new_AGEMA_signal_4763), .B0_t (LED_128_Instance_MCS_Instance_1_n4), .B0_f (new_AGEMA_signal_5052), .B1_t (new_AGEMA_signal_5053), .B1_f (new_AGEMA_signal_5054), .Z0_t (LED_128_Instance_mixcolumns_out[7]), .Z0_f (new_AGEMA_signal_5202), .Z1_t (new_AGEMA_signal_5203), .Z1_f (new_AGEMA_signal_5204) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U12 ( .A0_t (LED_128_Instance_MCS_Instance_1_n3), .A0_f (new_AGEMA_signal_5205), .A1_t (new_AGEMA_signal_5206), .A1_f (new_AGEMA_signal_5207), .B0_t (LED_128_Instance_MCS_Instance_1_n2), .B0_f (new_AGEMA_signal_5058), .B1_t (new_AGEMA_signal_5059), .B1_f (new_AGEMA_signal_5060), .Z0_t (LED_128_Instance_mixcolumns_out[20]), .Z0_f (new_AGEMA_signal_5382), .Z1_t (new_AGEMA_signal_5383), .Z1_f (new_AGEMA_signal_5384) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U11 ( .A0_t (LED_128_Instance_subcells_out[26]), .A0_f (new_AGEMA_signal_4671), .A1_t (new_AGEMA_signal_4672), .A1_f (new_AGEMA_signal_4673), .B0_t (LED_128_Instance_MCS_Instance_1_n4), .B0_f (new_AGEMA_signal_5052), .B1_t (new_AGEMA_signal_5053), .B1_f (new_AGEMA_signal_5054), .Z0_t (LED_128_Instance_MCS_Instance_1_n3), .Z0_f (new_AGEMA_signal_5205), .Z1_t (new_AGEMA_signal_5206), .Z1_f (new_AGEMA_signal_5207) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U10 ( .A0_t (LED_128_Instance_subcells_out[50]), .A0_f (new_AGEMA_signal_4722), .A1_t (new_AGEMA_signal_4723), .A1_f (new_AGEMA_signal_4724), .B0_t (LED_128_Instance_MCS_Instance_1_n36), .B0_f (new_AGEMA_signal_4932), .B1_t (new_AGEMA_signal_4933), .B1_f (new_AGEMA_signal_4934), .Z0_t (LED_128_Instance_MCS_Instance_1_n4), .Z0_f (new_AGEMA_signal_5052), .Z1_t (new_AGEMA_signal_5053), .Z1_f (new_AGEMA_signal_5054) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U9 ( .A0_t (LED_128_Instance_subcells_out[27]), .A0_f (new_AGEMA_signal_4782), .A1_t (new_AGEMA_signal_4783), .A1_f (new_AGEMA_signal_4784), .B0_t (LED_128_Instance_subcells_out[46]), .B0_f (new_AGEMA_signal_4713), .B1_t (new_AGEMA_signal_4714), .B1_f (new_AGEMA_signal_4715), .Z0_t (LED_128_Instance_MCS_Instance_1_n36), .Z0_f (new_AGEMA_signal_4932), .Z1_t (new_AGEMA_signal_4933), .Z1_f (new_AGEMA_signal_4934) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U8 ( .A0_t (LED_128_Instance_subcells_out[51]), .A0_f (new_AGEMA_signal_4806), .A1_t (new_AGEMA_signal_4807), .A1_f (new_AGEMA_signal_4808), .B0_t (LED_128_Instance_MCS_Instance_1_n5), .B0_f (new_AGEMA_signal_5055), .B1_t (new_AGEMA_signal_5056), .B1_f (new_AGEMA_signal_5057), .Z0_t (LED_128_Instance_mixcolumns_out[4]), .Z0_f (new_AGEMA_signal_5208), .Z1_t (new_AGEMA_signal_5209), .Z1_f (new_AGEMA_signal_5210) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U7 ( .A0_t (LED_128_Instance_subcells_out[47]), .A0_f (new_AGEMA_signal_4803), .A1_t (new_AGEMA_signal_4804), .A1_f (new_AGEMA_signal_4805), .B0_t (LED_128_Instance_MCS_Instance_1_n35), .B0_f (new_AGEMA_signal_4935), .B1_t (new_AGEMA_signal_4936), .B1_f (new_AGEMA_signal_4937), .Z0_t (LED_128_Instance_MCS_Instance_1_n5), .Z0_f (new_AGEMA_signal_5055), .Z1_t (new_AGEMA_signal_5056), .Z1_f (new_AGEMA_signal_5057) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U6 ( .A0_t (LED_128_Instance_subcells_out[6]), .A0_f (new_AGEMA_signal_4758), .A1_t (new_AGEMA_signal_4759), .A1_f (new_AGEMA_signal_4760), .B0_t (LED_128_Instance_subcells_out[24]), .B0_f (new_AGEMA_signal_4146), .B1_t (new_AGEMA_signal_4147), .B1_f (new_AGEMA_signal_4148), .Z0_t (LED_128_Instance_MCS_Instance_1_n35), .Z0_f (new_AGEMA_signal_4935), .Z1_t (new_AGEMA_signal_4936), .Z1_f (new_AGEMA_signal_4937) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U5 ( .A0_t (LED_128_Instance_MCS_Instance_1_n1), .A0_f (new_AGEMA_signal_5211), .A1_t (new_AGEMA_signal_5212), .A1_f (new_AGEMA_signal_5213), .B0_t (LED_128_Instance_MCS_Instance_1_n8), .B0_f (new_AGEMA_signal_4860), .B1_t (new_AGEMA_signal_4861), .B1_f (new_AGEMA_signal_4862), .Z0_t (LED_128_Instance_mixcolumns_out[54]), .Z0_f (new_AGEMA_signal_5385), .Z1_t (new_AGEMA_signal_5386), .Z1_f (new_AGEMA_signal_5387) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U4 ( .A0_t (LED_128_Instance_subcells_out[49]), .A0_f (new_AGEMA_signal_4725), .A1_t (new_AGEMA_signal_4726), .A1_f (new_AGEMA_signal_4727), .B0_t (LED_128_Instance_subcells_out[45]), .B0_f (new_AGEMA_signal_4716), .B1_t (new_AGEMA_signal_4717), .B1_f (new_AGEMA_signal_4718), .Z0_t (LED_128_Instance_MCS_Instance_1_n8), .Z0_f (new_AGEMA_signal_4860), .Z1_t (new_AGEMA_signal_4861), .Z1_f (new_AGEMA_signal_4862) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U3 ( .A0_t (LED_128_Instance_subcells_out[25]), .A0_f (new_AGEMA_signal_4674), .A1_t (new_AGEMA_signal_4675), .A1_f (new_AGEMA_signal_4676), .B0_t (LED_128_Instance_MCS_Instance_1_n2), .B0_f (new_AGEMA_signal_5058), .B1_t (new_AGEMA_signal_5059), .B1_f (new_AGEMA_signal_5060), .Z0_t (LED_128_Instance_MCS_Instance_1_n1), .Z0_f (new_AGEMA_signal_5211), .Z1_t (new_AGEMA_signal_5212), .Z1_f (new_AGEMA_signal_5213) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U2 ( .A0_t (LED_128_Instance_subcells_out[44]), .A0_f (new_AGEMA_signal_4221), .A1_t (new_AGEMA_signal_4222), .A1_f (new_AGEMA_signal_4223), .B0_t (LED_128_Instance_MCS_Instance_1_n26), .B0_f (new_AGEMA_signal_4938), .B1_t (new_AGEMA_signal_4939), .B1_f (new_AGEMA_signal_4940), .Z0_t (LED_128_Instance_MCS_Instance_1_n2), .Z0_f (new_AGEMA_signal_5058), .Z1_t (new_AGEMA_signal_5059), .Z1_f (new_AGEMA_signal_5060) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_1_U1 ( .A0_t (LED_128_Instance_subcells_out[5]), .A0_f (new_AGEMA_signal_4761), .A1_t (new_AGEMA_signal_4762), .A1_f (new_AGEMA_signal_4763), .B0_t (LED_128_Instance_subcells_out[51]), .B0_f (new_AGEMA_signal_4806), .B1_t (new_AGEMA_signal_4807), .B1_f (new_AGEMA_signal_4808), .Z0_t (LED_128_Instance_MCS_Instance_1_n26), .Z0_f (new_AGEMA_signal_4938), .Z1_t (new_AGEMA_signal_4939), .Z1_f (new_AGEMA_signal_4940) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U58 ( .A0_t (LED_128_Instance_subcells_out[10]), .A0_f (new_AGEMA_signal_4638), .A1_t (new_AGEMA_signal_4639), .A1_f (new_AGEMA_signal_4640), .B0_t (LED_128_Instance_MCS_Instance_2_n42), .B0_f (new_AGEMA_signal_5214), .B1_t (new_AGEMA_signal_5215), .B1_f (new_AGEMA_signal_5216), .Z0_t (LED_128_Instance_mixcolumns_out[9]), .Z0_f (new_AGEMA_signal_5388), .Z1_t (new_AGEMA_signal_5389), .Z1_f (new_AGEMA_signal_5390) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U57 ( .A0_t (LED_128_Instance_MCS_Instance_2_n41), .A0_f (new_AGEMA_signal_5403), .A1_t (new_AGEMA_signal_5404), .A1_f (new_AGEMA_signal_5405), .B0_t (LED_128_Instance_subcells_out[54]), .B0_f (new_AGEMA_signal_4812), .B1_t (new_AGEMA_signal_4813), .B1_f (new_AGEMA_signal_4814), .Z0_t (LED_128_Instance_mixcolumns_out[27]), .Z0_f (new_AGEMA_signal_5598), .Z1_t (new_AGEMA_signal_5599), .Z1_f (new_AGEMA_signal_5600) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U56 ( .A0_t (LED_128_Instance_subcells_out[53]), .A0_f (new_AGEMA_signal_4815), .A1_t (new_AGEMA_signal_4816), .A1_f (new_AGEMA_signal_4817), .B0_t (LED_128_Instance_MCS_Instance_2_n40), .B0_f (new_AGEMA_signal_5391), .B1_t (new_AGEMA_signal_5392), .B1_f (new_AGEMA_signal_5393), .Z0_t (LED_128_Instance_mixcolumns_out[26]), .Z0_f (new_AGEMA_signal_5601), .Z1_t (new_AGEMA_signal_5602), .Z1_f (new_AGEMA_signal_5603) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U55 ( .A0_t (LED_128_Instance_MCS_Instance_2_n39), .A0_f (new_AGEMA_signal_5061), .A1_t (new_AGEMA_signal_5062), .A1_f (new_AGEMA_signal_5063), .B0_t (LED_128_Instance_MCS_Instance_2_n42), .B0_f (new_AGEMA_signal_5214), .B1_t (new_AGEMA_signal_5215), .B1_f (new_AGEMA_signal_5216), .Z0_t (LED_128_Instance_MCS_Instance_2_n40), .Z0_f (new_AGEMA_signal_5391), .Z1_t (new_AGEMA_signal_5392), .Z1_f (new_AGEMA_signal_5393) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U54 ( .A0_t (LED_128_Instance_MCS_Instance_2_n38), .A0_f (new_AGEMA_signal_5073), .A1_t (new_AGEMA_signal_5074), .A1_f (new_AGEMA_signal_5075), .B0_t (LED_128_Instance_MCS_Instance_2_n37), .B0_f (new_AGEMA_signal_5076), .B1_t (new_AGEMA_signal_5077), .B1_f (new_AGEMA_signal_5078), .Z0_t (LED_128_Instance_MCS_Instance_2_n42), .Z0_f (new_AGEMA_signal_5214), .Z1_t (new_AGEMA_signal_5215), .Z1_f (new_AGEMA_signal_5216) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U53 ( .A0_t (LED_128_Instance_MCS_Instance_2_n36), .A0_f (new_AGEMA_signal_4956), .A1_t (new_AGEMA_signal_4957), .A1_f (new_AGEMA_signal_4958), .B0_t (LED_128_Instance_MCS_Instance_2_n35), .B0_f (new_AGEMA_signal_4872), .B1_t (new_AGEMA_signal_4873), .B1_f (new_AGEMA_signal_4874), .Z0_t (LED_128_Instance_MCS_Instance_2_n39), .Z0_f (new_AGEMA_signal_5061), .Z1_t (new_AGEMA_signal_5062), .Z1_f (new_AGEMA_signal_5063) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U52 ( .A0_t (LED_128_Instance_MCS_Instance_2_n34), .A0_f (new_AGEMA_signal_5217), .A1_t (new_AGEMA_signal_5218), .A1_f (new_AGEMA_signal_5219), .B0_t (LED_128_Instance_MCS_Instance_2_n36), .B0_f (new_AGEMA_signal_4956), .B1_t (new_AGEMA_signal_4957), .B1_f (new_AGEMA_signal_4958), .Z0_t (LED_128_Instance_mixcolumns_out[43]), .Z0_f (new_AGEMA_signal_5394), .Z1_t (new_AGEMA_signal_5395), .Z1_f (new_AGEMA_signal_5396) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U51 ( .A0_t (LED_128_Instance_MCS_Instance_2_n33), .A0_f (new_AGEMA_signal_5067), .A1_t (new_AGEMA_signal_5068), .A1_f (new_AGEMA_signal_5069), .B0_t (LED_128_Instance_MCS_Instance_2_n32), .B0_f (new_AGEMA_signal_5064), .B1_t (new_AGEMA_signal_5065), .B1_f (new_AGEMA_signal_5066), .Z0_t (LED_128_Instance_MCS_Instance_2_n34), .Z0_f (new_AGEMA_signal_5217), .Z1_t (new_AGEMA_signal_5218), .Z1_f (new_AGEMA_signal_5219) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U50 ( .A0_t (LED_128_Instance_MCS_Instance_2_n31), .A0_f (new_AGEMA_signal_4944), .A1_t (new_AGEMA_signal_4945), .A1_f (new_AGEMA_signal_4946), .B0_t (LED_128_Instance_subcells_out[30]), .B0_f (new_AGEMA_signal_4680), .B1_t (new_AGEMA_signal_4681), .B1_f (new_AGEMA_signal_4682), .Z0_t (LED_128_Instance_MCS_Instance_2_n32), .Z0_f (new_AGEMA_signal_5064), .Z1_t (new_AGEMA_signal_5065), .Z1_f (new_AGEMA_signal_5066) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U49 ( .A0_t (LED_128_Instance_MCS_Instance_2_n30), .A0_f (new_AGEMA_signal_4518), .A1_t (new_AGEMA_signal_4519), .A1_f (new_AGEMA_signal_4520), .B0_t (LED_128_Instance_MCS_Instance_2_n29), .B0_f (new_AGEMA_signal_4941), .B1_t (new_AGEMA_signal_4942), .B1_f (new_AGEMA_signal_4943), .Z0_t (LED_128_Instance_MCS_Instance_2_n33), .Z0_f (new_AGEMA_signal_5067), .Z1_t (new_AGEMA_signal_5068), .Z1_f (new_AGEMA_signal_5069) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U48 ( .A0_t (LED_128_Instance_MCS_Instance_2_n28), .A0_f (new_AGEMA_signal_5220), .A1_t (new_AGEMA_signal_5221), .A1_f (new_AGEMA_signal_5222), .B0_t (LED_128_Instance_MCS_Instance_2_n27), .B0_f (new_AGEMA_signal_5226), .B1_t (new_AGEMA_signal_5227), .B1_f (new_AGEMA_signal_5228), .Z0_t (LED_128_Instance_mixcolumns_out[42]), .Z0_f (new_AGEMA_signal_5397), .Z1_t (new_AGEMA_signal_5398), .Z1_f (new_AGEMA_signal_5399) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U47 ( .A0_t (LED_128_Instance_MCS_Instance_2_n26), .A0_f (new_AGEMA_signal_5091), .A1_t (new_AGEMA_signal_5092), .A1_f (new_AGEMA_signal_5093), .B0_t (LED_128_Instance_MCS_Instance_2_n25), .B0_f (new_AGEMA_signal_4863), .B1_t (new_AGEMA_signal_4864), .B1_f (new_AGEMA_signal_4865), .Z0_t (LED_128_Instance_MCS_Instance_2_n28), .Z0_f (new_AGEMA_signal_5220), .Z1_t (new_AGEMA_signal_5221), .Z1_f (new_AGEMA_signal_5222) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U46 ( .A0_t (LED_128_Instance_subcells_out[34]), .A0_f (new_AGEMA_signal_4689), .A1_t (new_AGEMA_signal_4690), .A1_f (new_AGEMA_signal_4691), .B0_t (LED_128_Instance_subcells_out[28]), .B0_f (new_AGEMA_signal_4161), .B1_t (new_AGEMA_signal_4162), .B1_f (new_AGEMA_signal_4163), .Z0_t (LED_128_Instance_MCS_Instance_2_n25), .Z0_f (new_AGEMA_signal_4863), .Z1_t (new_AGEMA_signal_4864), .Z1_f (new_AGEMA_signal_4865) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U45 ( .A0_t (LED_128_Instance_MCS_Instance_2_n24), .A0_f (new_AGEMA_signal_5400), .A1_t (new_AGEMA_signal_5401), .A1_f (new_AGEMA_signal_5402), .B0_t (LED_128_Instance_MCS_Instance_2_n23), .B0_f (new_AGEMA_signal_4953), .B1_t (new_AGEMA_signal_4954), .B1_f (new_AGEMA_signal_4955), .Z0_t (LED_128_Instance_mixcolumns_out[41]), .Z0_f (new_AGEMA_signal_5604), .Z1_t (new_AGEMA_signal_5605), .Z1_f (new_AGEMA_signal_5606) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U44 ( .A0_t (LED_128_Instance_MCS_Instance_2_n22), .A0_f (new_AGEMA_signal_5070), .A1_t (new_AGEMA_signal_5071), .A1_f (new_AGEMA_signal_5072), .B0_t (LED_128_Instance_MCS_Instance_2_n21), .B0_f (new_AGEMA_signal_5223), .B1_t (new_AGEMA_signal_5224), .B1_f (new_AGEMA_signal_5225), .Z0_t (LED_128_Instance_MCS_Instance_2_n24), .Z0_f (new_AGEMA_signal_5400), .Z1_t (new_AGEMA_signal_5401), .Z1_f (new_AGEMA_signal_5402) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U43 ( .A0_t (LED_128_Instance_MCS_Instance_2_n38), .A0_f (new_AGEMA_signal_5073), .A1_t (new_AGEMA_signal_5074), .A1_f (new_AGEMA_signal_5075), .B0_t (LED_128_Instance_subcells_out[33]), .B0_f (new_AGEMA_signal_4692), .B1_t (new_AGEMA_signal_4693), .B1_f (new_AGEMA_signal_4694), .Z0_t (LED_128_Instance_MCS_Instance_2_n21), .Z0_f (new_AGEMA_signal_5223), .Z1_t (new_AGEMA_signal_5224), .Z1_f (new_AGEMA_signal_5225) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U42 ( .A0_t (LED_128_Instance_MCS_Instance_2_n29), .A0_f (new_AGEMA_signal_4941), .A1_t (new_AGEMA_signal_4942), .A1_f (new_AGEMA_signal_4943), .B0_t (LED_128_Instance_subcells_out[32]), .B0_f (new_AGEMA_signal_4176), .B1_t (new_AGEMA_signal_4177), .B1_f (new_AGEMA_signal_4178), .Z0_t (LED_128_Instance_MCS_Instance_2_n22), .Z0_f (new_AGEMA_signal_5070), .Z1_t (new_AGEMA_signal_5071), .Z1_f (new_AGEMA_signal_5072) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U41 ( .A0_t (LED_128_Instance_subcells_out[8]), .A0_f (new_AGEMA_signal_4086), .A1_t (new_AGEMA_signal_4087), .A1_f (new_AGEMA_signal_4088), .B0_t (LED_128_Instance_MCS_Instance_2_n35), .B0_f (new_AGEMA_signal_4872), .B1_t (new_AGEMA_signal_4873), .B1_f (new_AGEMA_signal_4874), .Z0_t (LED_128_Instance_MCS_Instance_2_n29), .Z0_f (new_AGEMA_signal_4941), .Z1_t (new_AGEMA_signal_4942), .Z1_f (new_AGEMA_signal_4943) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U40 ( .A0_t (LED_128_Instance_MCS_Instance_2_n20), .A0_f (new_AGEMA_signal_5607), .A1_t (new_AGEMA_signal_5608), .A1_f (new_AGEMA_signal_5609), .B0_t (LED_128_Instance_MCS_Instance_2_n19), .B0_f (new_AGEMA_signal_4869), .B1_t (new_AGEMA_signal_4870), .B1_f (new_AGEMA_signal_4871), .Z0_t (LED_128_Instance_mixcolumns_out[40]), .Z0_f (new_AGEMA_signal_5826), .Z1_t (new_AGEMA_signal_5827), .Z1_f (new_AGEMA_signal_5828) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U39 ( .A0_t (LED_128_Instance_MCS_Instance_2_n41), .A0_f (new_AGEMA_signal_5403), .A1_t (new_AGEMA_signal_5404), .A1_f (new_AGEMA_signal_5405), .B0_t (LED_128_Instance_subcells_out[31]), .B0_f (new_AGEMA_signal_4785), .B1_t (new_AGEMA_signal_4786), .B1_f (new_AGEMA_signal_4787), .Z0_t (LED_128_Instance_MCS_Instance_2_n20), .Z0_f (new_AGEMA_signal_5607), .Z1_t (new_AGEMA_signal_5608), .Z1_f (new_AGEMA_signal_5609) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U38 ( .A0_t (LED_128_Instance_MCS_Instance_2_n18), .A0_f (new_AGEMA_signal_4950), .A1_t (new_AGEMA_signal_4951), .A1_f (new_AGEMA_signal_4952), .B0_t (LED_128_Instance_MCS_Instance_2_n27), .B0_f (new_AGEMA_signal_5226), .B1_t (new_AGEMA_signal_5227), .B1_f (new_AGEMA_signal_5228), .Z0_t (LED_128_Instance_MCS_Instance_2_n41), .Z0_f (new_AGEMA_signal_5403), .Z1_t (new_AGEMA_signal_5404), .Z1_f (new_AGEMA_signal_5405) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U37 ( .A0_t (LED_128_Instance_MCS_Instance_2_n38), .A0_f (new_AGEMA_signal_5073), .A1_t (new_AGEMA_signal_5074), .A1_f (new_AGEMA_signal_5075), .B0_t (LED_128_Instance_MCS_Instance_2_n17), .B0_f (new_AGEMA_signal_4866), .B1_t (new_AGEMA_signal_4867), .B1_f (new_AGEMA_signal_4868), .Z0_t (LED_128_Instance_MCS_Instance_2_n27), .Z0_f (new_AGEMA_signal_5226), .Z1_t (new_AGEMA_signal_5227), .Z1_f (new_AGEMA_signal_5228) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U36 ( .A0_t (LED_128_Instance_subcells_out[11]), .A0_f (new_AGEMA_signal_4764), .A1_t (new_AGEMA_signal_4765), .A1_f (new_AGEMA_signal_4766), .B0_t (LED_128_Instance_MCS_Instance_2_n31), .B0_f (new_AGEMA_signal_4944), .B1_t (new_AGEMA_signal_4945), .B1_f (new_AGEMA_signal_4946), .Z0_t (LED_128_Instance_MCS_Instance_2_n38), .Z0_f (new_AGEMA_signal_5073), .Z1_t (new_AGEMA_signal_5074), .Z1_f (new_AGEMA_signal_5075) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U35 ( .A0_t (LED_128_Instance_subcells_out[35]), .A0_f (new_AGEMA_signal_4788), .A1_t (new_AGEMA_signal_4789), .A1_f (new_AGEMA_signal_4790), .B0_t (LED_128_Instance_subcells_out[29]), .B0_f (new_AGEMA_signal_4683), .B1_t (new_AGEMA_signal_4684), .B1_f (new_AGEMA_signal_4685), .Z0_t (LED_128_Instance_MCS_Instance_2_n31), .Z0_f (new_AGEMA_signal_4944), .Z1_t (new_AGEMA_signal_4945), .Z1_f (new_AGEMA_signal_4946) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U34 ( .A0_t (LED_128_Instance_MCS_Instance_2_n16), .A0_f (new_AGEMA_signal_5229), .A1_t (new_AGEMA_signal_5230), .A1_f (new_AGEMA_signal_5231), .B0_t (LED_128_Instance_MCS_Instance_2_n30), .B0_f (new_AGEMA_signal_4518), .B1_t (new_AGEMA_signal_4519), .B1_f (new_AGEMA_signal_4520), .Z0_t (LED_128_Instance_mixcolumns_out[59]), .Z0_f (new_AGEMA_signal_5406), .Z1_t (new_AGEMA_signal_5407), .Z1_f (new_AGEMA_signal_5408) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U33 ( .A0_t (LED_128_Instance_MCS_Instance_2_n15), .A0_f (new_AGEMA_signal_5082), .A1_t (new_AGEMA_signal_5083), .A1_f (new_AGEMA_signal_5084), .B0_t (LED_128_Instance_subcells_out[10]), .B0_f (new_AGEMA_signal_4638), .B1_t (new_AGEMA_signal_4639), .B1_f (new_AGEMA_signal_4640), .Z0_t (LED_128_Instance_MCS_Instance_2_n16), .Z0_f (new_AGEMA_signal_5229), .Z1_t (new_AGEMA_signal_5230), .Z1_f (new_AGEMA_signal_5231) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U32 ( .A0_t (LED_128_Instance_subcells_out[31]), .A0_f (new_AGEMA_signal_4785), .A1_t (new_AGEMA_signal_4786), .A1_f (new_AGEMA_signal_4787), .B0_t (LED_128_Instance_MCS_Instance_2_n14), .B0_f (new_AGEMA_signal_5610), .B1_t (new_AGEMA_signal_5611), .B1_f (new_AGEMA_signal_5612), .Z0_t (LED_128_Instance_mixcolumns_out[57]), .Z0_f (new_AGEMA_signal_5829), .Z1_t (new_AGEMA_signal_5830), .Z1_f (new_AGEMA_signal_5831) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U31 ( .A0_t (LED_128_Instance_MCS_Instance_2_n13), .A0_f (new_AGEMA_signal_5409), .A1_t (new_AGEMA_signal_5410), .A1_f (new_AGEMA_signal_5411), .B0_t (LED_128_Instance_MCS_Instance_2_n12), .B0_f (new_AGEMA_signal_4947), .B1_t (new_AGEMA_signal_4948), .B1_f (new_AGEMA_signal_4949), .Z0_t (LED_128_Instance_MCS_Instance_2_n14), .Z0_f (new_AGEMA_signal_5610), .Z1_t (new_AGEMA_signal_5611), .Z1_f (new_AGEMA_signal_5612) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U30 ( .A0_t (LED_128_Instance_subcells_out[8]), .A0_f (new_AGEMA_signal_4086), .A1_t (new_AGEMA_signal_4087), .A1_f (new_AGEMA_signal_4088), .B0_t (LED_128_Instance_subcells_out[54]), .B0_f (new_AGEMA_signal_4812), .B1_t (new_AGEMA_signal_4813), .B1_f (new_AGEMA_signal_4814), .Z0_t (LED_128_Instance_MCS_Instance_2_n12), .Z0_f (new_AGEMA_signal_4947), .Z1_t (new_AGEMA_signal_4948), .Z1_f (new_AGEMA_signal_4949) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U29 ( .A0_t (LED_128_Instance_MCS_Instance_2_n11), .A0_f (new_AGEMA_signal_5232), .A1_t (new_AGEMA_signal_5233), .A1_f (new_AGEMA_signal_5234), .B0_t (LED_128_Instance_subcells_out[28]), .B0_f (new_AGEMA_signal_4161), .B1_t (new_AGEMA_signal_4162), .B1_f (new_AGEMA_signal_4163), .Z0_t (LED_128_Instance_MCS_Instance_2_n13), .Z0_f (new_AGEMA_signal_5409), .Z1_t (new_AGEMA_signal_5410), .Z1_f (new_AGEMA_signal_5411) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U28 ( .A0_t (LED_128_Instance_subcells_out[35]), .A0_f (new_AGEMA_signal_4788), .A1_t (new_AGEMA_signal_4789), .A1_f (new_AGEMA_signal_4790), .B0_t (LED_128_Instance_MCS_Instance_2_n10), .B0_f (new_AGEMA_signal_5613), .B1_t (new_AGEMA_signal_5614), .B1_f (new_AGEMA_signal_5615), .Z0_t (LED_128_Instance_mixcolumns_out[56]), .Z0_f (new_AGEMA_signal_5832), .Z1_t (new_AGEMA_signal_5833), .Z1_f (new_AGEMA_signal_5834) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U27 ( .A0_t (LED_128_Instance_MCS_Instance_2_n9), .A0_f (new_AGEMA_signal_5412), .A1_t (new_AGEMA_signal_5413), .A1_f (new_AGEMA_signal_5414), .B0_t (LED_128_Instance_MCS_Instance_2_n36), .B0_f (new_AGEMA_signal_4956), .B1_t (new_AGEMA_signal_4957), .B1_f (new_AGEMA_signal_4958), .Z0_t (LED_128_Instance_MCS_Instance_2_n10), .Z0_f (new_AGEMA_signal_5613), .Z1_t (new_AGEMA_signal_5614), .Z1_f (new_AGEMA_signal_5615) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U26 ( .A0_t (LED_128_Instance_MCS_Instance_2_n11), .A0_f (new_AGEMA_signal_5232), .A1_t (new_AGEMA_signal_5233), .A1_f (new_AGEMA_signal_5234), .B0_t (LED_128_Instance_MCS_Instance_2_n8), .B0_f (new_AGEMA_signal_4962), .B1_t (new_AGEMA_signal_4963), .B1_f (new_AGEMA_signal_4964), .Z0_t (LED_128_Instance_MCS_Instance_2_n9), .Z0_f (new_AGEMA_signal_5412), .Z1_t (new_AGEMA_signal_5413), .Z1_f (new_AGEMA_signal_5414) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U25 ( .A0_t (LED_128_Instance_subcells_out[11]), .A0_f (new_AGEMA_signal_4764), .A1_t (new_AGEMA_signal_4765), .A1_f (new_AGEMA_signal_4766), .B0_t (LED_128_Instance_MCS_Instance_2_n37), .B0_f (new_AGEMA_signal_5076), .B1_t (new_AGEMA_signal_5077), .B1_f (new_AGEMA_signal_5078), .Z0_t (LED_128_Instance_MCS_Instance_2_n11), .Z0_f (new_AGEMA_signal_5232), .Z1_t (new_AGEMA_signal_5233), .Z1_f (new_AGEMA_signal_5234) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U24 ( .A0_t (LED_128_Instance_subcells_out[55]), .A0_f (new_AGEMA_signal_4896), .A1_t (new_AGEMA_signal_4897), .A1_f (new_AGEMA_signal_4898), .B0_t (LED_128_Instance_MCS_Instance_2_n30), .B0_f (new_AGEMA_signal_4518), .B1_t (new_AGEMA_signal_4519), .B1_f (new_AGEMA_signal_4520), .Z0_t (LED_128_Instance_MCS_Instance_2_n37), .Z0_f (new_AGEMA_signal_5076), .Z1_t (new_AGEMA_signal_5077), .Z1_f (new_AGEMA_signal_5078) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U23 ( .A0_t (LED_128_Instance_subcells_out[52]), .A0_f (new_AGEMA_signal_4401), .A1_t (new_AGEMA_signal_4402), .A1_f (new_AGEMA_signal_4403), .B0_t (LED_128_Instance_subcells_out[32]), .B0_f (new_AGEMA_signal_4176), .B1_t (new_AGEMA_signal_4177), .B1_f (new_AGEMA_signal_4178), .Z0_t (LED_128_Instance_MCS_Instance_2_n30), .Z0_f (new_AGEMA_signal_4518), .Z1_t (new_AGEMA_signal_4519), .Z1_f (new_AGEMA_signal_4520) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U22 ( .A0_t (LED_128_Instance_MCS_Instance_2_n7), .A0_f (new_AGEMA_signal_5079), .A1_t (new_AGEMA_signal_5080), .A1_f (new_AGEMA_signal_5081), .B0_t (LED_128_Instance_MCS_Instance_2_n17), .B0_f (new_AGEMA_signal_4866), .B1_t (new_AGEMA_signal_4867), .B1_f (new_AGEMA_signal_4868), .Z0_t (LED_128_Instance_mixcolumns_out[10]), .Z0_f (new_AGEMA_signal_5235), .Z1_t (new_AGEMA_signal_5236), .Z1_f (new_AGEMA_signal_5237) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U21 ( .A0_t (LED_128_Instance_MCS_Instance_2_n18), .A0_f (new_AGEMA_signal_4950), .A1_t (new_AGEMA_signal_4951), .A1_f (new_AGEMA_signal_4952), .B0_t (LED_128_Instance_subcells_out[11]), .B0_f (new_AGEMA_signal_4764), .B1_t (new_AGEMA_signal_4765), .B1_f (new_AGEMA_signal_4766), .Z0_t (LED_128_Instance_MCS_Instance_2_n7), .Z0_f (new_AGEMA_signal_5079), .Z1_t (new_AGEMA_signal_5080), .Z1_f (new_AGEMA_signal_5081) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U20 ( .A0_t (LED_128_Instance_subcells_out[8]), .A0_f (new_AGEMA_signal_4086), .A1_t (new_AGEMA_signal_4087), .A1_f (new_AGEMA_signal_4088), .B0_t (LED_128_Instance_subcells_out[53]), .B0_f (new_AGEMA_signal_4815), .B1_t (new_AGEMA_signal_4816), .B1_f (new_AGEMA_signal_4817), .Z0_t (LED_128_Instance_MCS_Instance_2_n18), .Z0_f (new_AGEMA_signal_4950), .Z1_t (new_AGEMA_signal_4951), .Z1_f (new_AGEMA_signal_4952) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U19 ( .A0_t (LED_128_Instance_MCS_Instance_2_n6), .A0_f (new_AGEMA_signal_5238), .A1_t (new_AGEMA_signal_5239), .A1_f (new_AGEMA_signal_5240), .B0_t (LED_128_Instance_MCS_Instance_2_n5), .B0_f (new_AGEMA_signal_4959), .B1_t (new_AGEMA_signal_4960), .B1_f (new_AGEMA_signal_4961), .Z0_t (LED_128_Instance_mixcolumns_out[25]), .Z0_f (new_AGEMA_signal_5415), .Z1_t (new_AGEMA_signal_5416), .Z1_f (new_AGEMA_signal_5417) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U18 ( .A0_t (LED_128_Instance_MCS_Instance_2_n19), .A0_f (new_AGEMA_signal_4869), .A1_t (new_AGEMA_signal_4870), .A1_f (new_AGEMA_signal_4871), .B0_t (LED_128_Instance_MCS_Instance_2_n15), .B0_f (new_AGEMA_signal_5082), .B1_t (new_AGEMA_signal_5083), .B1_f (new_AGEMA_signal_5084), .Z0_t (LED_128_Instance_MCS_Instance_2_n6), .Z0_f (new_AGEMA_signal_5238), .Z1_t (new_AGEMA_signal_5239), .Z1_f (new_AGEMA_signal_5240) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U17 ( .A0_t (LED_128_Instance_MCS_Instance_2_n17), .A0_f (new_AGEMA_signal_4866), .A1_t (new_AGEMA_signal_4867), .A1_f (new_AGEMA_signal_4868), .B0_t (LED_128_Instance_MCS_Instance_2_n23), .B0_f (new_AGEMA_signal_4953), .B1_t (new_AGEMA_signal_4954), .B1_f (new_AGEMA_signal_4955), .Z0_t (LED_128_Instance_MCS_Instance_2_n15), .Z0_f (new_AGEMA_signal_5082), .Z1_t (new_AGEMA_signal_5083), .Z1_f (new_AGEMA_signal_5084) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U16 ( .A0_t (LED_128_Instance_subcells_out[54]), .A0_f (new_AGEMA_signal_4812), .A1_t (new_AGEMA_signal_4813), .A1_f (new_AGEMA_signal_4814), .B0_t (LED_128_Instance_subcells_out[34]), .B0_f (new_AGEMA_signal_4689), .B1_t (new_AGEMA_signal_4690), .B1_f (new_AGEMA_signal_4691), .Z0_t (LED_128_Instance_MCS_Instance_2_n23), .Z0_f (new_AGEMA_signal_4953), .Z1_t (new_AGEMA_signal_4954), .Z1_f (new_AGEMA_signal_4955) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U15 ( .A0_t (LED_128_Instance_subcells_out[33]), .A0_f (new_AGEMA_signal_4692), .A1_t (new_AGEMA_signal_4693), .A1_f (new_AGEMA_signal_4694), .B0_t (LED_128_Instance_subcells_out[30]), .B0_f (new_AGEMA_signal_4680), .B1_t (new_AGEMA_signal_4681), .B1_f (new_AGEMA_signal_4682), .Z0_t (LED_128_Instance_MCS_Instance_2_n17), .Z0_f (new_AGEMA_signal_4866), .Z1_t (new_AGEMA_signal_4867), .Z1_f (new_AGEMA_signal_4868) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U14 ( .A0_t (LED_128_Instance_subcells_out[52]), .A0_f (new_AGEMA_signal_4401), .A1_t (new_AGEMA_signal_4402), .A1_f (new_AGEMA_signal_4403), .B0_t (LED_128_Instance_subcells_out[9]), .B0_f (new_AGEMA_signal_4641), .B1_t (new_AGEMA_signal_4642), .B1_f (new_AGEMA_signal_4643), .Z0_t (LED_128_Instance_MCS_Instance_2_n19), .Z0_f (new_AGEMA_signal_4869), .Z1_t (new_AGEMA_signal_4870), .Z1_f (new_AGEMA_signal_4871) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U13 ( .A0_t (LED_128_Instance_subcells_out[9]), .A0_f (new_AGEMA_signal_4641), .A1_t (new_AGEMA_signal_4642), .A1_f (new_AGEMA_signal_4643), .B0_t (LED_128_Instance_MCS_Instance_2_n4), .B0_f (new_AGEMA_signal_5085), .B1_t (new_AGEMA_signal_5086), .B1_f (new_AGEMA_signal_5087), .Z0_t (LED_128_Instance_mixcolumns_out[11]), .Z0_f (new_AGEMA_signal_5241), .Z1_t (new_AGEMA_signal_5242), .Z1_f (new_AGEMA_signal_5243) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U12 ( .A0_t (LED_128_Instance_MCS_Instance_2_n3), .A0_f (new_AGEMA_signal_5244), .A1_t (new_AGEMA_signal_5245), .A1_f (new_AGEMA_signal_5246), .B0_t (LED_128_Instance_MCS_Instance_2_n2), .B0_f (new_AGEMA_signal_5247), .B1_t (new_AGEMA_signal_5248), .B1_f (new_AGEMA_signal_5249), .Z0_t (LED_128_Instance_mixcolumns_out[24]), .Z0_f (new_AGEMA_signal_5418), .Z1_t (new_AGEMA_signal_5419), .Z1_f (new_AGEMA_signal_5420) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U11 ( .A0_t (LED_128_Instance_subcells_out[30]), .A0_f (new_AGEMA_signal_4680), .A1_t (new_AGEMA_signal_4681), .A1_f (new_AGEMA_signal_4682), .B0_t (LED_128_Instance_MCS_Instance_2_n4), .B0_f (new_AGEMA_signal_5085), .B1_t (new_AGEMA_signal_5086), .B1_f (new_AGEMA_signal_5087), .Z0_t (LED_128_Instance_MCS_Instance_2_n3), .Z0_f (new_AGEMA_signal_5244), .Z1_t (new_AGEMA_signal_5245), .Z1_f (new_AGEMA_signal_5246) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U10 ( .A0_t (LED_128_Instance_subcells_out[54]), .A0_f (new_AGEMA_signal_4812), .A1_t (new_AGEMA_signal_4813), .A1_f (new_AGEMA_signal_4814), .B0_t (LED_128_Instance_MCS_Instance_2_n36), .B0_f (new_AGEMA_signal_4956), .B1_t (new_AGEMA_signal_4957), .B1_f (new_AGEMA_signal_4958), .Z0_t (LED_128_Instance_MCS_Instance_2_n4), .Z0_f (new_AGEMA_signal_5085), .Z1_t (new_AGEMA_signal_5086), .Z1_f (new_AGEMA_signal_5087) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U9 ( .A0_t (LED_128_Instance_subcells_out[31]), .A0_f (new_AGEMA_signal_4785), .A1_t (new_AGEMA_signal_4786), .A1_f (new_AGEMA_signal_4787), .B0_t (LED_128_Instance_subcells_out[34]), .B0_f (new_AGEMA_signal_4689), .B1_t (new_AGEMA_signal_4690), .B1_f (new_AGEMA_signal_4691), .Z0_t (LED_128_Instance_MCS_Instance_2_n36), .Z0_f (new_AGEMA_signal_4956), .Z1_t (new_AGEMA_signal_4957), .Z1_f (new_AGEMA_signal_4958) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U8 ( .A0_t (LED_128_Instance_subcells_out[55]), .A0_f (new_AGEMA_signal_4896), .A1_t (new_AGEMA_signal_4897), .A1_f (new_AGEMA_signal_4898), .B0_t (LED_128_Instance_MCS_Instance_2_n5), .B0_f (new_AGEMA_signal_4959), .B1_t (new_AGEMA_signal_4960), .B1_f (new_AGEMA_signal_4961), .Z0_t (LED_128_Instance_mixcolumns_out[8]), .Z0_f (new_AGEMA_signal_5088), .Z1_t (new_AGEMA_signal_5089), .Z1_f (new_AGEMA_signal_5090) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U7 ( .A0_t (LED_128_Instance_subcells_out[35]), .A0_f (new_AGEMA_signal_4788), .A1_t (new_AGEMA_signal_4789), .A1_f (new_AGEMA_signal_4790), .B0_t (LED_128_Instance_MCS_Instance_2_n35), .B0_f (new_AGEMA_signal_4872), .B1_t (new_AGEMA_signal_4873), .B1_f (new_AGEMA_signal_4874), .Z0_t (LED_128_Instance_MCS_Instance_2_n5), .Z0_f (new_AGEMA_signal_4959), .Z1_t (new_AGEMA_signal_4960), .Z1_f (new_AGEMA_signal_4961) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U6 ( .A0_t (LED_128_Instance_subcells_out[10]), .A0_f (new_AGEMA_signal_4638), .A1_t (new_AGEMA_signal_4639), .A1_f (new_AGEMA_signal_4640), .B0_t (LED_128_Instance_subcells_out[28]), .B0_f (new_AGEMA_signal_4161), .B1_t (new_AGEMA_signal_4162), .B1_f (new_AGEMA_signal_4163), .Z0_t (LED_128_Instance_MCS_Instance_2_n35), .Z0_f (new_AGEMA_signal_4872), .Z1_t (new_AGEMA_signal_4873), .Z1_f (new_AGEMA_signal_4874) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U5 ( .A0_t (LED_128_Instance_MCS_Instance_2_n1), .A0_f (new_AGEMA_signal_5421), .A1_t (new_AGEMA_signal_5422), .A1_f (new_AGEMA_signal_5423), .B0_t (LED_128_Instance_MCS_Instance_2_n8), .B0_f (new_AGEMA_signal_4962), .B1_t (new_AGEMA_signal_4963), .B1_f (new_AGEMA_signal_4964), .Z0_t (LED_128_Instance_mixcolumns_out[58]), .Z0_f (new_AGEMA_signal_5616), .Z1_t (new_AGEMA_signal_5617), .Z1_f (new_AGEMA_signal_5618) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U4 ( .A0_t (LED_128_Instance_subcells_out[53]), .A0_f (new_AGEMA_signal_4815), .A1_t (new_AGEMA_signal_4816), .A1_f (new_AGEMA_signal_4817), .B0_t (LED_128_Instance_subcells_out[33]), .B0_f (new_AGEMA_signal_4692), .B1_t (new_AGEMA_signal_4693), .B1_f (new_AGEMA_signal_4694), .Z0_t (LED_128_Instance_MCS_Instance_2_n8), .Z0_f (new_AGEMA_signal_4962), .Z1_t (new_AGEMA_signal_4963), .Z1_f (new_AGEMA_signal_4964) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U3 ( .A0_t (LED_128_Instance_subcells_out[29]), .A0_f (new_AGEMA_signal_4683), .A1_t (new_AGEMA_signal_4684), .A1_f (new_AGEMA_signal_4685), .B0_t (LED_128_Instance_MCS_Instance_2_n2), .B0_f (new_AGEMA_signal_5247), .B1_t (new_AGEMA_signal_5248), .B1_f (new_AGEMA_signal_5249), .Z0_t (LED_128_Instance_MCS_Instance_2_n1), .Z0_f (new_AGEMA_signal_5421), .Z1_t (new_AGEMA_signal_5422), .Z1_f (new_AGEMA_signal_5423) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U2 ( .A0_t (LED_128_Instance_subcells_out[32]), .A0_f (new_AGEMA_signal_4176), .A1_t (new_AGEMA_signal_4177), .A1_f (new_AGEMA_signal_4178), .B0_t (LED_128_Instance_MCS_Instance_2_n26), .B0_f (new_AGEMA_signal_5091), .B1_t (new_AGEMA_signal_5092), .B1_f (new_AGEMA_signal_5093), .Z0_t (LED_128_Instance_MCS_Instance_2_n2), .Z0_f (new_AGEMA_signal_5247), .Z1_t (new_AGEMA_signal_5248), .Z1_f (new_AGEMA_signal_5249) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_2_U1 ( .A0_t (LED_128_Instance_subcells_out[9]), .A0_f (new_AGEMA_signal_4641), .A1_t (new_AGEMA_signal_4642), .A1_f (new_AGEMA_signal_4643), .B0_t (LED_128_Instance_subcells_out[55]), .B0_f (new_AGEMA_signal_4896), .B1_t (new_AGEMA_signal_4897), .B1_f (new_AGEMA_signal_4898), .Z0_t (LED_128_Instance_MCS_Instance_2_n26), .Z0_f (new_AGEMA_signal_5091), .Z1_t (new_AGEMA_signal_5092), .Z1_f (new_AGEMA_signal_5093) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U58 ( .A0_t (LED_128_Instance_subcells_out[14]), .A0_f (new_AGEMA_signal_4647), .A1_t (new_AGEMA_signal_4648), .A1_f (new_AGEMA_signal_4649), .B0_t (LED_128_Instance_MCS_Instance_3_n42), .B0_f (new_AGEMA_signal_5424), .B1_t (new_AGEMA_signal_5425), .B1_f (new_AGEMA_signal_5426), .Z0_t (LED_128_Instance_mixcolumns_out[13]), .Z0_f (new_AGEMA_signal_5619), .Z1_t (new_AGEMA_signal_5620), .Z1_f (new_AGEMA_signal_5621) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U57 ( .A0_t (LED_128_Instance_MCS_Instance_3_n41), .A0_f (new_AGEMA_signal_5634), .A1_t (new_AGEMA_signal_5635), .A1_f (new_AGEMA_signal_5636), .B0_t (LED_128_Instance_subcells_out[58]), .B0_f (new_AGEMA_signal_4737), .B1_t (new_AGEMA_signal_4738), .B1_f (new_AGEMA_signal_4739), .Z0_t (LED_128_Instance_mixcolumns_out[31]), .Z0_f (new_AGEMA_signal_5835), .Z1_t (new_AGEMA_signal_5836), .Z1_f (new_AGEMA_signal_5837) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U56 ( .A0_t (LED_128_Instance_subcells_out[57]), .A0_f (new_AGEMA_signal_4740), .A1_t (new_AGEMA_signal_4741), .A1_f (new_AGEMA_signal_4742), .B0_t (LED_128_Instance_MCS_Instance_3_n40), .B0_f (new_AGEMA_signal_5622), .B1_t (new_AGEMA_signal_5623), .B1_f (new_AGEMA_signal_5624), .Z0_t (LED_128_Instance_mixcolumns_out[30]), .Z0_f (new_AGEMA_signal_5838), .Z1_t (new_AGEMA_signal_5839), .Z1_f (new_AGEMA_signal_5840) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U55 ( .A0_t (LED_128_Instance_MCS_Instance_3_n39), .A0_f (new_AGEMA_signal_5094), .A1_t (new_AGEMA_signal_5095), .A1_f (new_AGEMA_signal_5096), .B0_t (LED_128_Instance_MCS_Instance_3_n42), .B0_f (new_AGEMA_signal_5424), .B1_t (new_AGEMA_signal_5425), .B1_f (new_AGEMA_signal_5426), .Z0_t (LED_128_Instance_MCS_Instance_3_n40), .Z0_f (new_AGEMA_signal_5622), .Z1_t (new_AGEMA_signal_5623), .Z1_f (new_AGEMA_signal_5624) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U54 ( .A0_t (LED_128_Instance_MCS_Instance_3_n38), .A0_f (new_AGEMA_signal_5253), .A1_t (new_AGEMA_signal_5254), .A1_f (new_AGEMA_signal_5255), .B0_t (LED_128_Instance_MCS_Instance_3_n37), .B0_f (new_AGEMA_signal_4971), .B1_t (new_AGEMA_signal_4972), .B1_f (new_AGEMA_signal_4973), .Z0_t (LED_128_Instance_MCS_Instance_3_n42), .Z0_f (new_AGEMA_signal_5424), .Z1_t (new_AGEMA_signal_5425), .Z1_f (new_AGEMA_signal_5426) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U53 ( .A0_t (LED_128_Instance_MCS_Instance_3_n36), .A0_f (new_AGEMA_signal_4983), .A1_t (new_AGEMA_signal_4984), .A1_f (new_AGEMA_signal_4985), .B0_t (LED_128_Instance_MCS_Instance_3_n35), .B0_f (new_AGEMA_signal_4884), .B1_t (new_AGEMA_signal_4885), .B1_f (new_AGEMA_signal_4886), .Z0_t (LED_128_Instance_MCS_Instance_3_n39), .Z0_f (new_AGEMA_signal_5094), .Z1_t (new_AGEMA_signal_5095), .Z1_f (new_AGEMA_signal_5096) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U52 ( .A0_t (LED_128_Instance_MCS_Instance_3_n34), .A0_f (new_AGEMA_signal_5427), .A1_t (new_AGEMA_signal_5428), .A1_f (new_AGEMA_signal_5429), .B0_t (LED_128_Instance_MCS_Instance_3_n36), .B0_f (new_AGEMA_signal_4983), .B1_t (new_AGEMA_signal_4984), .B1_f (new_AGEMA_signal_4985), .Z0_t (LED_128_Instance_mixcolumns_out[47]), .Z0_f (new_AGEMA_signal_5625), .Z1_t (new_AGEMA_signal_5626), .Z1_f (new_AGEMA_signal_5627) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U51 ( .A0_t (LED_128_Instance_MCS_Instance_3_n33), .A0_f (new_AGEMA_signal_5097), .A1_t (new_AGEMA_signal_5098), .A1_f (new_AGEMA_signal_5099), .B0_t (LED_128_Instance_MCS_Instance_3_n32), .B0_f (new_AGEMA_signal_5250), .B1_t (new_AGEMA_signal_5251), .B1_f (new_AGEMA_signal_5252), .Z0_t (LED_128_Instance_MCS_Instance_3_n34), .Z0_f (new_AGEMA_signal_5427), .Z1_t (new_AGEMA_signal_5428), .Z1_f (new_AGEMA_signal_5429) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U50 ( .A0_t (LED_128_Instance_MCS_Instance_3_n31), .A0_f (new_AGEMA_signal_5106), .A1_t (new_AGEMA_signal_5107), .A1_f (new_AGEMA_signal_5108), .B0_t (LED_128_Instance_subcells_out[18]), .B0_f (new_AGEMA_signal_4656), .B1_t (new_AGEMA_signal_4657), .B1_f (new_AGEMA_signal_4658), .Z0_t (LED_128_Instance_MCS_Instance_3_n32), .Z0_f (new_AGEMA_signal_5250), .Z1_t (new_AGEMA_signal_5251), .Z1_f (new_AGEMA_signal_5252) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U49 ( .A0_t (LED_128_Instance_MCS_Instance_3_n30), .A0_f (new_AGEMA_signal_4521), .A1_t (new_AGEMA_signal_4522), .A1_f (new_AGEMA_signal_4523), .B0_t (LED_128_Instance_MCS_Instance_3_n29), .B0_f (new_AGEMA_signal_4968), .B1_t (new_AGEMA_signal_4969), .B1_f (new_AGEMA_signal_4970), .Z0_t (LED_128_Instance_MCS_Instance_3_n33), .Z0_f (new_AGEMA_signal_5097), .Z1_t (new_AGEMA_signal_5098), .Z1_f (new_AGEMA_signal_5099) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U48 ( .A0_t (LED_128_Instance_MCS_Instance_3_n28), .A0_f (new_AGEMA_signal_5100), .A1_t (new_AGEMA_signal_5101), .A1_f (new_AGEMA_signal_5102), .B0_t (LED_128_Instance_MCS_Instance_3_n27), .B0_f (new_AGEMA_signal_5433), .B1_t (new_AGEMA_signal_5434), .B1_f (new_AGEMA_signal_5435), .Z0_t (LED_128_Instance_mixcolumns_out[46]), .Z0_f (new_AGEMA_signal_5628), .Z1_t (new_AGEMA_signal_5629), .Z1_f (new_AGEMA_signal_5630) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U47 ( .A0_t (LED_128_Instance_MCS_Instance_3_n26), .A0_f (new_AGEMA_signal_4989), .A1_t (new_AGEMA_signal_4990), .A1_f (new_AGEMA_signal_4991), .B0_t (LED_128_Instance_MCS_Instance_3_n25), .B0_f (new_AGEMA_signal_4965), .B1_t (new_AGEMA_signal_4966), .B1_f (new_AGEMA_signal_4967), .Z0_t (LED_128_Instance_MCS_Instance_3_n28), .Z0_f (new_AGEMA_signal_5100), .Z1_t (new_AGEMA_signal_5101), .Z1_f (new_AGEMA_signal_5102) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U46 ( .A0_t (LED_128_Instance_subcells_out[38]), .A0_f (new_AGEMA_signal_4794), .A1_t (new_AGEMA_signal_4795), .A1_f (new_AGEMA_signal_4796), .B0_t (LED_128_Instance_subcells_out[16]), .B0_f (new_AGEMA_signal_4116), .B1_t (new_AGEMA_signal_4117), .B1_f (new_AGEMA_signal_4118), .Z0_t (LED_128_Instance_MCS_Instance_3_n25), .Z0_f (new_AGEMA_signal_4965), .Z1_t (new_AGEMA_signal_4966), .Z1_f (new_AGEMA_signal_4967) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U45 ( .A0_t (LED_128_Instance_MCS_Instance_3_n24), .A0_f (new_AGEMA_signal_5631), .A1_t (new_AGEMA_signal_5632), .A1_f (new_AGEMA_signal_5633), .B0_t (LED_128_Instance_MCS_Instance_3_n23), .B0_f (new_AGEMA_signal_4977), .B1_t (new_AGEMA_signal_4978), .B1_f (new_AGEMA_signal_4979), .Z0_t (LED_128_Instance_mixcolumns_out[45]), .Z0_f (new_AGEMA_signal_5841), .Z1_t (new_AGEMA_signal_5842), .Z1_f (new_AGEMA_signal_5843) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U44 ( .A0_t (LED_128_Instance_MCS_Instance_3_n22), .A0_f (new_AGEMA_signal_5103), .A1_t (new_AGEMA_signal_5104), .A1_f (new_AGEMA_signal_5105), .B0_t (LED_128_Instance_MCS_Instance_3_n21), .B0_f (new_AGEMA_signal_5430), .B1_t (new_AGEMA_signal_5431), .B1_f (new_AGEMA_signal_5432), .Z0_t (LED_128_Instance_MCS_Instance_3_n24), .Z0_f (new_AGEMA_signal_5631), .Z1_t (new_AGEMA_signal_5632), .Z1_f (new_AGEMA_signal_5633) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U43 ( .A0_t (LED_128_Instance_MCS_Instance_3_n38), .A0_f (new_AGEMA_signal_5253), .A1_t (new_AGEMA_signal_5254), .A1_f (new_AGEMA_signal_5255), .B0_t (LED_128_Instance_subcells_out[37]), .B0_f (new_AGEMA_signal_4797), .B1_t (new_AGEMA_signal_4798), .B1_f (new_AGEMA_signal_4799), .Z0_t (LED_128_Instance_MCS_Instance_3_n21), .Z0_f (new_AGEMA_signal_5430), .Z1_t (new_AGEMA_signal_5431), .Z1_f (new_AGEMA_signal_5432) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U42 ( .A0_t (LED_128_Instance_MCS_Instance_3_n29), .A0_f (new_AGEMA_signal_4968), .A1_t (new_AGEMA_signal_4969), .A1_f (new_AGEMA_signal_4970), .B0_t (LED_128_Instance_subcells_out[36]), .B0_f (new_AGEMA_signal_4368), .B1_t (new_AGEMA_signal_4369), .B1_f (new_AGEMA_signal_4370), .Z0_t (LED_128_Instance_MCS_Instance_3_n22), .Z0_f (new_AGEMA_signal_5103), .Z1_t (new_AGEMA_signal_5104), .Z1_f (new_AGEMA_signal_5105) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U41 ( .A0_t (LED_128_Instance_subcells_out[12]), .A0_f (new_AGEMA_signal_4101), .A1_t (new_AGEMA_signal_4102), .A1_f (new_AGEMA_signal_4103), .B0_t (LED_128_Instance_MCS_Instance_3_n35), .B0_f (new_AGEMA_signal_4884), .B1_t (new_AGEMA_signal_4885), .B1_f (new_AGEMA_signal_4886), .Z0_t (LED_128_Instance_MCS_Instance_3_n29), .Z0_f (new_AGEMA_signal_4968), .Z1_t (new_AGEMA_signal_4969), .Z1_f (new_AGEMA_signal_4970) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U40 ( .A0_t (LED_128_Instance_MCS_Instance_3_n20), .A0_f (new_AGEMA_signal_5844), .A1_t (new_AGEMA_signal_5845), .A1_f (new_AGEMA_signal_5846), .B0_t (LED_128_Instance_MCS_Instance_3_n19), .B0_f (new_AGEMA_signal_4881), .B1_t (new_AGEMA_signal_4882), .B1_f (new_AGEMA_signal_4883), .Z0_t (LED_128_Instance_mixcolumns_out[44]), .Z0_f (new_AGEMA_signal_6063), .Z1_t (new_AGEMA_signal_6064), .Z1_f (new_AGEMA_signal_6065) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U39 ( .A0_t (LED_128_Instance_MCS_Instance_3_n41), .A0_f (new_AGEMA_signal_5634), .A1_t (new_AGEMA_signal_5635), .A1_f (new_AGEMA_signal_5636), .B0_t (LED_128_Instance_subcells_out[19]), .B0_f (new_AGEMA_signal_4770), .B1_t (new_AGEMA_signal_4771), .B1_f (new_AGEMA_signal_4772), .Z0_t (LED_128_Instance_MCS_Instance_3_n20), .Z0_f (new_AGEMA_signal_5844), .Z1_t (new_AGEMA_signal_5845), .Z1_f (new_AGEMA_signal_5846) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U38 ( .A0_t (LED_128_Instance_MCS_Instance_3_n18), .A0_f (new_AGEMA_signal_4878), .A1_t (new_AGEMA_signal_4879), .A1_f (new_AGEMA_signal_4880), .B0_t (LED_128_Instance_MCS_Instance_3_n27), .B0_f (new_AGEMA_signal_5433), .B1_t (new_AGEMA_signal_5434), .B1_f (new_AGEMA_signal_5435), .Z0_t (LED_128_Instance_MCS_Instance_3_n41), .Z0_f (new_AGEMA_signal_5634), .Z1_t (new_AGEMA_signal_5635), .Z1_f (new_AGEMA_signal_5636) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U37 ( .A0_t (LED_128_Instance_MCS_Instance_3_n38), .A0_f (new_AGEMA_signal_5253), .A1_t (new_AGEMA_signal_5254), .A1_f (new_AGEMA_signal_5255), .B0_t (LED_128_Instance_MCS_Instance_3_n17), .B0_f (new_AGEMA_signal_4980), .B1_t (new_AGEMA_signal_4981), .B1_f (new_AGEMA_signal_4982), .Z0_t (LED_128_Instance_MCS_Instance_3_n27), .Z0_f (new_AGEMA_signal_5433), .Z1_t (new_AGEMA_signal_5434), .Z1_f (new_AGEMA_signal_5435) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U36 ( .A0_t (LED_128_Instance_subcells_out[15]), .A0_f (new_AGEMA_signal_4767), .A1_t (new_AGEMA_signal_4768), .A1_f (new_AGEMA_signal_4769), .B0_t (LED_128_Instance_MCS_Instance_3_n31), .B0_f (new_AGEMA_signal_5106), .B1_t (new_AGEMA_signal_5107), .B1_f (new_AGEMA_signal_5108), .Z0_t (LED_128_Instance_MCS_Instance_3_n38), .Z0_f (new_AGEMA_signal_5253), .Z1_t (new_AGEMA_signal_5254), .Z1_f (new_AGEMA_signal_5255) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U35 ( .A0_t (LED_128_Instance_subcells_out[39]), .A0_f (new_AGEMA_signal_4893), .A1_t (new_AGEMA_signal_4894), .A1_f (new_AGEMA_signal_4895), .B0_t (LED_128_Instance_subcells_out[17]), .B0_f (new_AGEMA_signal_4659), .B1_t (new_AGEMA_signal_4660), .B1_f (new_AGEMA_signal_4661), .Z0_t (LED_128_Instance_MCS_Instance_3_n31), .Z0_f (new_AGEMA_signal_5106), .Z1_t (new_AGEMA_signal_5107), .Z1_f (new_AGEMA_signal_5108) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U34 ( .A0_t (LED_128_Instance_MCS_Instance_3_n16), .A0_f (new_AGEMA_signal_5256), .A1_t (new_AGEMA_signal_5257), .A1_f (new_AGEMA_signal_5258), .B0_t (LED_128_Instance_MCS_Instance_3_n30), .B0_f (new_AGEMA_signal_4521), .B1_t (new_AGEMA_signal_4522), .B1_f (new_AGEMA_signal_4523), .Z0_t (LED_128_Instance_mixcolumns_out[63]), .Z0_f (new_AGEMA_signal_5436), .Z1_t (new_AGEMA_signal_5437), .Z1_f (new_AGEMA_signal_5438) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U33 ( .A0_t (LED_128_Instance_MCS_Instance_3_n15), .A0_f (new_AGEMA_signal_5115), .A1_t (new_AGEMA_signal_5116), .A1_f (new_AGEMA_signal_5117), .B0_t (LED_128_Instance_subcells_out[14]), .B0_f (new_AGEMA_signal_4647), .B1_t (new_AGEMA_signal_4648), .B1_f (new_AGEMA_signal_4649), .Z0_t (LED_128_Instance_MCS_Instance_3_n16), .Z0_f (new_AGEMA_signal_5256), .Z1_t (new_AGEMA_signal_5257), .Z1_f (new_AGEMA_signal_5258) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U32 ( .A0_t (LED_128_Instance_subcells_out[19]), .A0_f (new_AGEMA_signal_4770), .A1_t (new_AGEMA_signal_4771), .A1_f (new_AGEMA_signal_4772), .B0_t (LED_128_Instance_MCS_Instance_3_n14), .B0_f (new_AGEMA_signal_5439), .B1_t (new_AGEMA_signal_5440), .B1_f (new_AGEMA_signal_5441), .Z0_t (LED_128_Instance_mixcolumns_out[61]), .Z0_f (new_AGEMA_signal_5637), .Z1_t (new_AGEMA_signal_5638), .Z1_f (new_AGEMA_signal_5639) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U31 ( .A0_t (LED_128_Instance_MCS_Instance_3_n13), .A0_f (new_AGEMA_signal_5259), .A1_t (new_AGEMA_signal_5260), .A1_f (new_AGEMA_signal_5261), .B0_t (LED_128_Instance_MCS_Instance_3_n12), .B0_f (new_AGEMA_signal_4875), .B1_t (new_AGEMA_signal_4876), .B1_f (new_AGEMA_signal_4877), .Z0_t (LED_128_Instance_MCS_Instance_3_n14), .Z0_f (new_AGEMA_signal_5439), .Z1_t (new_AGEMA_signal_5440), .Z1_f (new_AGEMA_signal_5441) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U30 ( .A0_t (LED_128_Instance_subcells_out[12]), .A0_f (new_AGEMA_signal_4101), .A1_t (new_AGEMA_signal_4102), .A1_f (new_AGEMA_signal_4103), .B0_t (LED_128_Instance_subcells_out[58]), .B0_f (new_AGEMA_signal_4737), .B1_t (new_AGEMA_signal_4738), .B1_f (new_AGEMA_signal_4739), .Z0_t (LED_128_Instance_MCS_Instance_3_n12), .Z0_f (new_AGEMA_signal_4875), .Z1_t (new_AGEMA_signal_4876), .Z1_f (new_AGEMA_signal_4877) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U29 ( .A0_t (LED_128_Instance_MCS_Instance_3_n11), .A0_f (new_AGEMA_signal_5109), .A1_t (new_AGEMA_signal_5110), .A1_f (new_AGEMA_signal_5111), .B0_t (LED_128_Instance_subcells_out[16]), .B0_f (new_AGEMA_signal_4116), .B1_t (new_AGEMA_signal_4117), .B1_f (new_AGEMA_signal_4118), .Z0_t (LED_128_Instance_MCS_Instance_3_n13), .Z0_f (new_AGEMA_signal_5259), .Z1_t (new_AGEMA_signal_5260), .Z1_f (new_AGEMA_signal_5261) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U28 ( .A0_t (LED_128_Instance_subcells_out[39]), .A0_f (new_AGEMA_signal_4893), .A1_t (new_AGEMA_signal_4894), .A1_f (new_AGEMA_signal_4895), .B0_t (LED_128_Instance_MCS_Instance_3_n10), .B0_f (new_AGEMA_signal_5442), .B1_t (new_AGEMA_signal_5443), .B1_f (new_AGEMA_signal_5444), .Z0_t (LED_128_Instance_mixcolumns_out[60]), .Z0_f (new_AGEMA_signal_5640), .Z1_t (new_AGEMA_signal_5641), .Z1_f (new_AGEMA_signal_5642) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U27 ( .A0_t (LED_128_Instance_MCS_Instance_3_n9), .A0_f (new_AGEMA_signal_5262), .A1_t (new_AGEMA_signal_5263), .A1_f (new_AGEMA_signal_5264), .B0_t (LED_128_Instance_MCS_Instance_3_n36), .B0_f (new_AGEMA_signal_4983), .B1_t (new_AGEMA_signal_4984), .B1_f (new_AGEMA_signal_4985), .Z0_t (LED_128_Instance_MCS_Instance_3_n10), .Z0_f (new_AGEMA_signal_5442), .Z1_t (new_AGEMA_signal_5443), .Z1_f (new_AGEMA_signal_5444) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U26 ( .A0_t (LED_128_Instance_MCS_Instance_3_n11), .A0_f (new_AGEMA_signal_5109), .A1_t (new_AGEMA_signal_5110), .A1_f (new_AGEMA_signal_5111), .B0_t (LED_128_Instance_MCS_Instance_3_n8), .B0_f (new_AGEMA_signal_4986), .B1_t (new_AGEMA_signal_4987), .B1_f (new_AGEMA_signal_4988), .Z0_t (LED_128_Instance_MCS_Instance_3_n9), .Z0_f (new_AGEMA_signal_5262), .Z1_t (new_AGEMA_signal_5263), .Z1_f (new_AGEMA_signal_5264) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U25 ( .A0_t (LED_128_Instance_subcells_out[15]), .A0_f (new_AGEMA_signal_4767), .A1_t (new_AGEMA_signal_4768), .A1_f (new_AGEMA_signal_4769), .B0_t (LED_128_Instance_MCS_Instance_3_n37), .B0_f (new_AGEMA_signal_4971), .B1_t (new_AGEMA_signal_4972), .B1_f (new_AGEMA_signal_4973), .Z0_t (LED_128_Instance_MCS_Instance_3_n11), .Z0_f (new_AGEMA_signal_5109), .Z1_t (new_AGEMA_signal_5110), .Z1_f (new_AGEMA_signal_5111) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U24 ( .A0_t (LED_128_Instance_subcells_out[59]), .A0_f (new_AGEMA_signal_4818), .A1_t (new_AGEMA_signal_4819), .A1_f (new_AGEMA_signal_4820), .B0_t (LED_128_Instance_MCS_Instance_3_n30), .B0_f (new_AGEMA_signal_4521), .B1_t (new_AGEMA_signal_4522), .B1_f (new_AGEMA_signal_4523), .Z0_t (LED_128_Instance_MCS_Instance_3_n37), .Z0_f (new_AGEMA_signal_4971), .Z1_t (new_AGEMA_signal_4972), .Z1_f (new_AGEMA_signal_4973) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U23 ( .A0_t (LED_128_Instance_subcells_out[56]), .A0_f (new_AGEMA_signal_4266), .A1_t (new_AGEMA_signal_4267), .A1_f (new_AGEMA_signal_4268), .B0_t (LED_128_Instance_subcells_out[36]), .B0_f (new_AGEMA_signal_4368), .B1_t (new_AGEMA_signal_4369), .B1_f (new_AGEMA_signal_4370), .Z0_t (LED_128_Instance_MCS_Instance_3_n30), .Z0_f (new_AGEMA_signal_4521), .Z1_t (new_AGEMA_signal_4522), .Z1_f (new_AGEMA_signal_4523) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U22 ( .A0_t (LED_128_Instance_MCS_Instance_3_n7), .A0_f (new_AGEMA_signal_4974), .A1_t (new_AGEMA_signal_4975), .A1_f (new_AGEMA_signal_4976), .B0_t (LED_128_Instance_MCS_Instance_3_n17), .B0_f (new_AGEMA_signal_4980), .B1_t (new_AGEMA_signal_4981), .B1_f (new_AGEMA_signal_4982), .Z0_t (LED_128_Instance_mixcolumns_out[14]), .Z0_f (new_AGEMA_signal_5112), .Z1_t (new_AGEMA_signal_5113), .Z1_f (new_AGEMA_signal_5114) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U21 ( .A0_t (LED_128_Instance_MCS_Instance_3_n18), .A0_f (new_AGEMA_signal_4878), .A1_t (new_AGEMA_signal_4879), .A1_f (new_AGEMA_signal_4880), .B0_t (LED_128_Instance_subcells_out[15]), .B0_f (new_AGEMA_signal_4767), .B1_t (new_AGEMA_signal_4768), .B1_f (new_AGEMA_signal_4769), .Z0_t (LED_128_Instance_MCS_Instance_3_n7), .Z0_f (new_AGEMA_signal_4974), .Z1_t (new_AGEMA_signal_4975), .Z1_f (new_AGEMA_signal_4976) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U20 ( .A0_t (LED_128_Instance_subcells_out[12]), .A0_f (new_AGEMA_signal_4101), .A1_t (new_AGEMA_signal_4102), .A1_f (new_AGEMA_signal_4103), .B0_t (LED_128_Instance_subcells_out[57]), .B0_f (new_AGEMA_signal_4740), .B1_t (new_AGEMA_signal_4741), .B1_f (new_AGEMA_signal_4742), .Z0_t (LED_128_Instance_MCS_Instance_3_n18), .Z0_f (new_AGEMA_signal_4878), .Z1_t (new_AGEMA_signal_4879), .Z1_f (new_AGEMA_signal_4880) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U19 ( .A0_t (LED_128_Instance_MCS_Instance_3_n6), .A0_f (new_AGEMA_signal_5265), .A1_t (new_AGEMA_signal_5266), .A1_f (new_AGEMA_signal_5267), .B0_t (LED_128_Instance_MCS_Instance_3_n5), .B0_f (new_AGEMA_signal_5121), .B1_t (new_AGEMA_signal_5122), .B1_f (new_AGEMA_signal_5123), .Z0_t (LED_128_Instance_mixcolumns_out[29]), .Z0_f (new_AGEMA_signal_5445), .Z1_t (new_AGEMA_signal_5446), .Z1_f (new_AGEMA_signal_5447) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U18 ( .A0_t (LED_128_Instance_MCS_Instance_3_n19), .A0_f (new_AGEMA_signal_4881), .A1_t (new_AGEMA_signal_4882), .A1_f (new_AGEMA_signal_4883), .B0_t (LED_128_Instance_MCS_Instance_3_n15), .B0_f (new_AGEMA_signal_5115), .B1_t (new_AGEMA_signal_5116), .B1_f (new_AGEMA_signal_5117), .Z0_t (LED_128_Instance_MCS_Instance_3_n6), .Z0_f (new_AGEMA_signal_5265), .Z1_t (new_AGEMA_signal_5266), .Z1_f (new_AGEMA_signal_5267) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U17 ( .A0_t (LED_128_Instance_MCS_Instance_3_n17), .A0_f (new_AGEMA_signal_4980), .A1_t (new_AGEMA_signal_4981), .A1_f (new_AGEMA_signal_4982), .B0_t (LED_128_Instance_MCS_Instance_3_n23), .B0_f (new_AGEMA_signal_4977), .B1_t (new_AGEMA_signal_4978), .B1_f (new_AGEMA_signal_4979), .Z0_t (LED_128_Instance_MCS_Instance_3_n15), .Z0_f (new_AGEMA_signal_5115), .Z1_t (new_AGEMA_signal_5116), .Z1_f (new_AGEMA_signal_5117) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U16 ( .A0_t (LED_128_Instance_subcells_out[58]), .A0_f (new_AGEMA_signal_4737), .A1_t (new_AGEMA_signal_4738), .A1_f (new_AGEMA_signal_4739), .B0_t (LED_128_Instance_subcells_out[38]), .B0_f (new_AGEMA_signal_4794), .B1_t (new_AGEMA_signal_4795), .B1_f (new_AGEMA_signal_4796), .Z0_t (LED_128_Instance_MCS_Instance_3_n23), .Z0_f (new_AGEMA_signal_4977), .Z1_t (new_AGEMA_signal_4978), .Z1_f (new_AGEMA_signal_4979) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U15 ( .A0_t (LED_128_Instance_subcells_out[37]), .A0_f (new_AGEMA_signal_4797), .A1_t (new_AGEMA_signal_4798), .A1_f (new_AGEMA_signal_4799), .B0_t (LED_128_Instance_subcells_out[18]), .B0_f (new_AGEMA_signal_4656), .B1_t (new_AGEMA_signal_4657), .B1_f (new_AGEMA_signal_4658), .Z0_t (LED_128_Instance_MCS_Instance_3_n17), .Z0_f (new_AGEMA_signal_4980), .Z1_t (new_AGEMA_signal_4981), .Z1_f (new_AGEMA_signal_4982) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U14 ( .A0_t (LED_128_Instance_subcells_out[56]), .A0_f (new_AGEMA_signal_4266), .A1_t (new_AGEMA_signal_4267), .A1_f (new_AGEMA_signal_4268), .B0_t (LED_128_Instance_subcells_out[13]), .B0_f (new_AGEMA_signal_4650), .B1_t (new_AGEMA_signal_4651), .B1_f (new_AGEMA_signal_4652), .Z0_t (LED_128_Instance_MCS_Instance_3_n19), .Z0_f (new_AGEMA_signal_4881), .Z1_t (new_AGEMA_signal_4882), .Z1_f (new_AGEMA_signal_4883) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U13 ( .A0_t (LED_128_Instance_subcells_out[13]), .A0_f (new_AGEMA_signal_4650), .A1_t (new_AGEMA_signal_4651), .A1_f (new_AGEMA_signal_4652), .B0_t (LED_128_Instance_MCS_Instance_3_n4), .B0_f (new_AGEMA_signal_5118), .B1_t (new_AGEMA_signal_5119), .B1_f (new_AGEMA_signal_5120), .Z0_t (LED_128_Instance_mixcolumns_out[15]), .Z0_f (new_AGEMA_signal_5268), .Z1_t (new_AGEMA_signal_5269), .Z1_f (new_AGEMA_signal_5270) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U12 ( .A0_t (LED_128_Instance_MCS_Instance_3_n3), .A0_f (new_AGEMA_signal_5271), .A1_t (new_AGEMA_signal_5272), .A1_f (new_AGEMA_signal_5273), .B0_t (LED_128_Instance_MCS_Instance_3_n2), .B0_f (new_AGEMA_signal_5124), .B1_t (new_AGEMA_signal_5125), .B1_f (new_AGEMA_signal_5126), .Z0_t (LED_128_Instance_mixcolumns_out[28]), .Z0_f (new_AGEMA_signal_5448), .Z1_t (new_AGEMA_signal_5449), .Z1_f (new_AGEMA_signal_5450) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U11 ( .A0_t (LED_128_Instance_subcells_out[18]), .A0_f (new_AGEMA_signal_4656), .A1_t (new_AGEMA_signal_4657), .A1_f (new_AGEMA_signal_4658), .B0_t (LED_128_Instance_MCS_Instance_3_n4), .B0_f (new_AGEMA_signal_5118), .B1_t (new_AGEMA_signal_5119), .B1_f (new_AGEMA_signal_5120), .Z0_t (LED_128_Instance_MCS_Instance_3_n3), .Z0_f (new_AGEMA_signal_5271), .Z1_t (new_AGEMA_signal_5272), .Z1_f (new_AGEMA_signal_5273) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U10 ( .A0_t (LED_128_Instance_subcells_out[58]), .A0_f (new_AGEMA_signal_4737), .A1_t (new_AGEMA_signal_4738), .A1_f (new_AGEMA_signal_4739), .B0_t (LED_128_Instance_MCS_Instance_3_n36), .B0_f (new_AGEMA_signal_4983), .B1_t (new_AGEMA_signal_4984), .B1_f (new_AGEMA_signal_4985), .Z0_t (LED_128_Instance_MCS_Instance_3_n4), .Z0_f (new_AGEMA_signal_5118), .Z1_t (new_AGEMA_signal_5119), .Z1_f (new_AGEMA_signal_5120) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U9 ( .A0_t (LED_128_Instance_subcells_out[19]), .A0_f (new_AGEMA_signal_4770), .A1_t (new_AGEMA_signal_4771), .A1_f (new_AGEMA_signal_4772), .B0_t (LED_128_Instance_subcells_out[38]), .B0_f (new_AGEMA_signal_4794), .B1_t (new_AGEMA_signal_4795), .B1_f (new_AGEMA_signal_4796), .Z0_t (LED_128_Instance_MCS_Instance_3_n36), .Z0_f (new_AGEMA_signal_4983), .Z1_t (new_AGEMA_signal_4984), .Z1_f (new_AGEMA_signal_4985) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U8 ( .A0_t (LED_128_Instance_subcells_out[59]), .A0_f (new_AGEMA_signal_4818), .A1_t (new_AGEMA_signal_4819), .A1_f (new_AGEMA_signal_4820), .B0_t (LED_128_Instance_MCS_Instance_3_n5), .B0_f (new_AGEMA_signal_5121), .B1_t (new_AGEMA_signal_5122), .B1_f (new_AGEMA_signal_5123), .Z0_t (LED_128_Instance_mixcolumns_out[12]), .Z0_f (new_AGEMA_signal_5274), .Z1_t (new_AGEMA_signal_5275), .Z1_f (new_AGEMA_signal_5276) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U7 ( .A0_t (LED_128_Instance_subcells_out[39]), .A0_f (new_AGEMA_signal_4893), .A1_t (new_AGEMA_signal_4894), .A1_f (new_AGEMA_signal_4895), .B0_t (LED_128_Instance_MCS_Instance_3_n35), .B0_f (new_AGEMA_signal_4884), .B1_t (new_AGEMA_signal_4885), .B1_f (new_AGEMA_signal_4886), .Z0_t (LED_128_Instance_MCS_Instance_3_n5), .Z0_f (new_AGEMA_signal_5121), .Z1_t (new_AGEMA_signal_5122), .Z1_f (new_AGEMA_signal_5123) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U6 ( .A0_t (LED_128_Instance_subcells_out[14]), .A0_f (new_AGEMA_signal_4647), .A1_t (new_AGEMA_signal_4648), .A1_f (new_AGEMA_signal_4649), .B0_t (LED_128_Instance_subcells_out[16]), .B0_f (new_AGEMA_signal_4116), .B1_t (new_AGEMA_signal_4117), .B1_f (new_AGEMA_signal_4118), .Z0_t (LED_128_Instance_MCS_Instance_3_n35), .Z0_f (new_AGEMA_signal_4884), .Z1_t (new_AGEMA_signal_4885), .Z1_f (new_AGEMA_signal_4886) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U5 ( .A0_t (LED_128_Instance_MCS_Instance_3_n1), .A0_f (new_AGEMA_signal_5277), .A1_t (new_AGEMA_signal_5278), .A1_f (new_AGEMA_signal_5279), .B0_t (LED_128_Instance_MCS_Instance_3_n8), .B0_f (new_AGEMA_signal_4986), .B1_t (new_AGEMA_signal_4987), .B1_f (new_AGEMA_signal_4988), .Z0_t (LED_128_Instance_mixcolumns_out[62]), .Z0_f (new_AGEMA_signal_5451), .Z1_t (new_AGEMA_signal_5452), .Z1_f (new_AGEMA_signal_5453) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U4 ( .A0_t (LED_128_Instance_subcells_out[57]), .A0_f (new_AGEMA_signal_4740), .A1_t (new_AGEMA_signal_4741), .A1_f (new_AGEMA_signal_4742), .B0_t (LED_128_Instance_subcells_out[37]), .B0_f (new_AGEMA_signal_4797), .B1_t (new_AGEMA_signal_4798), .B1_f (new_AGEMA_signal_4799), .Z0_t (LED_128_Instance_MCS_Instance_3_n8), .Z0_f (new_AGEMA_signal_4986), .Z1_t (new_AGEMA_signal_4987), .Z1_f (new_AGEMA_signal_4988) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U3 ( .A0_t (LED_128_Instance_subcells_out[17]), .A0_f (new_AGEMA_signal_4659), .A1_t (new_AGEMA_signal_4660), .A1_f (new_AGEMA_signal_4661), .B0_t (LED_128_Instance_MCS_Instance_3_n2), .B0_f (new_AGEMA_signal_5124), .B1_t (new_AGEMA_signal_5125), .B1_f (new_AGEMA_signal_5126), .Z0_t (LED_128_Instance_MCS_Instance_3_n1), .Z0_f (new_AGEMA_signal_5277), .Z1_t (new_AGEMA_signal_5278), .Z1_f (new_AGEMA_signal_5279) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U2 ( .A0_t (LED_128_Instance_subcells_out[36]), .A0_f (new_AGEMA_signal_4368), .A1_t (new_AGEMA_signal_4369), .A1_f (new_AGEMA_signal_4370), .B0_t (LED_128_Instance_MCS_Instance_3_n26), .B0_f (new_AGEMA_signal_4989), .B1_t (new_AGEMA_signal_4990), .B1_f (new_AGEMA_signal_4991), .Z0_t (LED_128_Instance_MCS_Instance_3_n2), .Z0_f (new_AGEMA_signal_5124), .Z1_t (new_AGEMA_signal_5125), .Z1_f (new_AGEMA_signal_5126) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) LED_128_Instance_MCS_Instance_3_U1 ( .A0_t (LED_128_Instance_subcells_out[13]), .A0_f (new_AGEMA_signal_4650), .A1_t (new_AGEMA_signal_4651), .A1_f (new_AGEMA_signal_4652), .B0_t (LED_128_Instance_subcells_out[59]), .B0_f (new_AGEMA_signal_4818), .B1_t (new_AGEMA_signal_4819), .B1_f (new_AGEMA_signal_4820), .Z0_t (LED_128_Instance_MCS_Instance_3_n26), .Z0_f (new_AGEMA_signal_4989), .Z1_t (new_AGEMA_signal_4990), .Z1_f (new_AGEMA_signal_4991) ) ;

    /* register cells */
endmodule
