/* modified netlist. Source: module present in file /mnt/c/Users/amirm/Desktop/Papers_in_progress/SAUBER/Design for our FPGA/11-PRESENT80_nibble_serial_encryption_PortParallel/4-AGEMA/present.v */
/* 0 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 1 register stage(s) in total */

module present_SAUBER_Pipeline_d1 (data_in, key, reset, data_out, done);
    input [63:0] data_in ;
    input [79:0] key ;
    input reset ;
    output [63:0] data_out ;
    output done ;
    wire selSbox ;
    wire intDone ;
    wire fsm_n14 ;
    wire fsm_n13 ;
    wire fsm_n12 ;
    wire fsm_n11 ;
    wire fsm_n10 ;
    wire fsm_n9 ;
    wire fsm_n8 ;
    wire fsm_n7 ;
    wire fsm_n6 ;
    wire fsm_n5 ;
    wire fsm_n4 ;
    wire fsm_rst_countSerial ;
    wire fsm_en_countRound ;
    wire fsm_n16 ;
    wire fsm_ps_state_0_ ;
    wire fsm_cnt_rnd_n12 ;
    wire fsm_cnt_rnd_n10 ;
    wire fsm_cnt_rnd_n9 ;
    wire fsm_cnt_rnd_n8 ;
    wire fsm_cnt_rnd_n7 ;
    wire fsm_cnt_rnd_n6 ;
    wire fsm_cnt_rnd_n5 ;
    wire fsm_cnt_rnd_n4 ;
    wire fsm_cnt_rnd_n3 ;
    wire fsm_cnt_ser_n9 ;
    wire fsm_cnt_ser_n7 ;
    wire fsm_cnt_ser_n6 ;
    wire fsm_cnt_ser_n5 ;
    wire fsm_cnt_ser_n4 ;
    wire fsm_cnt_ser_n3 ;
    wire fsm_cnt_ser_n2 ;
    wire stateFF_state_gff_1_MUX_inst1_mux_inst_0_U1_Y ;
    wire stateFF_state_gff_1_MUX_inst1_mux_inst_0_U1_X ;
    wire stateFF_state_gff_1_MUX_inst1_mux_inst_1_U1_Y ;
    wire stateFF_state_gff_1_MUX_inst1_mux_inst_1_U1_X ;
    wire stateFF_state_gff_1_MUX_inst1_mux_inst_2_U1_Y ;
    wire stateFF_state_gff_1_MUX_inst1_mux_inst_2_U1_X ;
    wire stateFF_state_gff_1_MUX_inst1_mux_inst_3_U1_Y ;
    wire stateFF_state_gff_1_MUX_inst1_mux_inst_3_U1_X ;
    wire stateFF_state_gff_2_MUX_inst1_mux_inst_0_U1_Y ;
    wire stateFF_state_gff_2_MUX_inst1_mux_inst_0_U1_X ;
    wire stateFF_state_gff_2_MUX_inst1_mux_inst_1_U1_Y ;
    wire stateFF_state_gff_2_MUX_inst1_mux_inst_1_U1_X ;
    wire stateFF_state_gff_2_MUX_inst1_mux_inst_2_U1_Y ;
    wire stateFF_state_gff_2_MUX_inst1_mux_inst_2_U1_X ;
    wire stateFF_state_gff_2_MUX_inst1_mux_inst_3_U1_Y ;
    wire stateFF_state_gff_2_MUX_inst1_mux_inst_3_U1_X ;
    wire stateFF_state_gff_3_MUX_inst1_mux_inst_0_U1_Y ;
    wire stateFF_state_gff_3_MUX_inst1_mux_inst_0_U1_X ;
    wire stateFF_state_gff_3_MUX_inst1_mux_inst_1_U1_Y ;
    wire stateFF_state_gff_3_MUX_inst1_mux_inst_1_U1_X ;
    wire stateFF_state_gff_3_MUX_inst1_mux_inst_2_U1_Y ;
    wire stateFF_state_gff_3_MUX_inst1_mux_inst_2_U1_X ;
    wire stateFF_state_gff_3_MUX_inst1_mux_inst_3_U1_Y ;
    wire stateFF_state_gff_3_MUX_inst1_mux_inst_3_U1_X ;
    wire stateFF_state_gff_4_MUX_inst1_mux_inst_0_U1_Y ;
    wire stateFF_state_gff_4_MUX_inst1_mux_inst_0_U1_X ;
    wire stateFF_state_gff_4_MUX_inst1_mux_inst_1_U1_Y ;
    wire stateFF_state_gff_4_MUX_inst1_mux_inst_1_U1_X ;
    wire stateFF_state_gff_4_MUX_inst1_mux_inst_2_U1_Y ;
    wire stateFF_state_gff_4_MUX_inst1_mux_inst_2_U1_X ;
    wire stateFF_state_gff_4_MUX_inst1_mux_inst_3_U1_Y ;
    wire stateFF_state_gff_4_MUX_inst1_mux_inst_3_U1_X ;
    wire stateFF_state_gff_5_MUX_inst1_mux_inst_0_U1_Y ;
    wire stateFF_state_gff_5_MUX_inst1_mux_inst_0_U1_X ;
    wire stateFF_state_gff_5_MUX_inst1_mux_inst_1_U1_Y ;
    wire stateFF_state_gff_5_MUX_inst1_mux_inst_1_U1_X ;
    wire stateFF_state_gff_5_MUX_inst1_mux_inst_2_U1_Y ;
    wire stateFF_state_gff_5_MUX_inst1_mux_inst_2_U1_X ;
    wire stateFF_state_gff_5_MUX_inst1_mux_inst_3_U1_Y ;
    wire stateFF_state_gff_5_MUX_inst1_mux_inst_3_U1_X ;
    wire stateFF_state_gff_6_MUX_inst1_mux_inst_0_U1_Y ;
    wire stateFF_state_gff_6_MUX_inst1_mux_inst_0_U1_X ;
    wire stateFF_state_gff_6_MUX_inst1_mux_inst_1_U1_Y ;
    wire stateFF_state_gff_6_MUX_inst1_mux_inst_1_U1_X ;
    wire stateFF_state_gff_6_MUX_inst1_mux_inst_2_U1_Y ;
    wire stateFF_state_gff_6_MUX_inst1_mux_inst_2_U1_X ;
    wire stateFF_state_gff_6_MUX_inst1_mux_inst_3_U1_Y ;
    wire stateFF_state_gff_6_MUX_inst1_mux_inst_3_U1_X ;
    wire stateFF_state_gff_7_MUX_inst1_mux_inst_0_U1_Y ;
    wire stateFF_state_gff_7_MUX_inst1_mux_inst_0_U1_X ;
    wire stateFF_state_gff_7_MUX_inst1_mux_inst_1_U1_Y ;
    wire stateFF_state_gff_7_MUX_inst1_mux_inst_1_U1_X ;
    wire stateFF_state_gff_7_MUX_inst1_mux_inst_2_U1_Y ;
    wire stateFF_state_gff_7_MUX_inst1_mux_inst_2_U1_X ;
    wire stateFF_state_gff_7_MUX_inst1_mux_inst_3_U1_Y ;
    wire stateFF_state_gff_7_MUX_inst1_mux_inst_3_U1_X ;
    wire stateFF_state_gff_8_MUX_inst1_mux_inst_0_U1_Y ;
    wire stateFF_state_gff_8_MUX_inst1_mux_inst_0_U1_X ;
    wire stateFF_state_gff_8_MUX_inst1_mux_inst_1_U1_Y ;
    wire stateFF_state_gff_8_MUX_inst1_mux_inst_1_U1_X ;
    wire stateFF_state_gff_8_MUX_inst1_mux_inst_2_U1_Y ;
    wire stateFF_state_gff_8_MUX_inst1_mux_inst_2_U1_X ;
    wire stateFF_state_gff_8_MUX_inst1_mux_inst_3_U1_Y ;
    wire stateFF_state_gff_8_MUX_inst1_mux_inst_3_U1_X ;
    wire stateFF_state_gff_9_MUX_inst1_mux_inst_0_U1_Y ;
    wire stateFF_state_gff_9_MUX_inst1_mux_inst_0_U1_X ;
    wire stateFF_state_gff_9_MUX_inst1_mux_inst_1_U1_Y ;
    wire stateFF_state_gff_9_MUX_inst1_mux_inst_1_U1_X ;
    wire stateFF_state_gff_9_MUX_inst1_mux_inst_2_U1_Y ;
    wire stateFF_state_gff_9_MUX_inst1_mux_inst_2_U1_X ;
    wire stateFF_state_gff_9_MUX_inst1_mux_inst_3_U1_Y ;
    wire stateFF_state_gff_9_MUX_inst1_mux_inst_3_U1_X ;
    wire stateFF_state_gff_10_MUX_inst1_mux_inst_0_U1_Y ;
    wire stateFF_state_gff_10_MUX_inst1_mux_inst_0_U1_X ;
    wire stateFF_state_gff_10_MUX_inst1_mux_inst_1_U1_Y ;
    wire stateFF_state_gff_10_MUX_inst1_mux_inst_1_U1_X ;
    wire stateFF_state_gff_10_MUX_inst1_mux_inst_2_U1_Y ;
    wire stateFF_state_gff_10_MUX_inst1_mux_inst_2_U1_X ;
    wire stateFF_state_gff_10_MUX_inst1_mux_inst_3_U1_Y ;
    wire stateFF_state_gff_10_MUX_inst1_mux_inst_3_U1_X ;
    wire stateFF_state_gff_11_MUX_inst1_mux_inst_0_U1_Y ;
    wire stateFF_state_gff_11_MUX_inst1_mux_inst_0_U1_X ;
    wire stateFF_state_gff_11_MUX_inst1_mux_inst_1_U1_Y ;
    wire stateFF_state_gff_11_MUX_inst1_mux_inst_1_U1_X ;
    wire stateFF_state_gff_11_MUX_inst1_mux_inst_2_U1_Y ;
    wire stateFF_state_gff_11_MUX_inst1_mux_inst_2_U1_X ;
    wire stateFF_state_gff_11_MUX_inst1_mux_inst_3_U1_Y ;
    wire stateFF_state_gff_11_MUX_inst1_mux_inst_3_U1_X ;
    wire stateFF_state_gff_12_MUX_inst1_mux_inst_0_U1_Y ;
    wire stateFF_state_gff_12_MUX_inst1_mux_inst_0_U1_X ;
    wire stateFF_state_gff_12_MUX_inst1_mux_inst_1_U1_Y ;
    wire stateFF_state_gff_12_MUX_inst1_mux_inst_1_U1_X ;
    wire stateFF_state_gff_12_MUX_inst1_mux_inst_2_U1_Y ;
    wire stateFF_state_gff_12_MUX_inst1_mux_inst_2_U1_X ;
    wire stateFF_state_gff_12_MUX_inst1_mux_inst_3_U1_Y ;
    wire stateFF_state_gff_12_MUX_inst1_mux_inst_3_U1_X ;
    wire stateFF_state_gff_13_MUX_inst1_mux_inst_0_U1_Y ;
    wire stateFF_state_gff_13_MUX_inst1_mux_inst_0_U1_X ;
    wire stateFF_state_gff_13_MUX_inst1_mux_inst_1_U1_Y ;
    wire stateFF_state_gff_13_MUX_inst1_mux_inst_1_U1_X ;
    wire stateFF_state_gff_13_MUX_inst1_mux_inst_2_U1_Y ;
    wire stateFF_state_gff_13_MUX_inst1_mux_inst_2_U1_X ;
    wire stateFF_state_gff_13_MUX_inst1_mux_inst_3_U1_Y ;
    wire stateFF_state_gff_13_MUX_inst1_mux_inst_3_U1_X ;
    wire stateFF_state_gff_14_MUX_inst1_mux_inst_0_U1_Y ;
    wire stateFF_state_gff_14_MUX_inst1_mux_inst_0_U1_X ;
    wire stateFF_state_gff_14_MUX_inst1_mux_inst_1_U1_Y ;
    wire stateFF_state_gff_14_MUX_inst1_mux_inst_1_U1_X ;
    wire stateFF_state_gff_14_MUX_inst1_mux_inst_2_U1_Y ;
    wire stateFF_state_gff_14_MUX_inst1_mux_inst_2_U1_X ;
    wire stateFF_state_gff_14_MUX_inst1_mux_inst_3_U1_Y ;
    wire stateFF_state_gff_14_MUX_inst1_mux_inst_3_U1_X ;
    wire stateFF_state_gff_15_MUX_inst1_mux_inst_0_U1_Y ;
    wire stateFF_state_gff_15_MUX_inst1_mux_inst_0_U1_X ;
    wire stateFF_state_gff_15_MUX_inst1_mux_inst_1_U1_Y ;
    wire stateFF_state_gff_15_MUX_inst1_mux_inst_1_U1_X ;
    wire stateFF_state_gff_15_MUX_inst1_mux_inst_2_U1_Y ;
    wire stateFF_state_gff_15_MUX_inst1_mux_inst_2_U1_X ;
    wire stateFF_state_gff_15_MUX_inst1_mux_inst_3_U1_Y ;
    wire stateFF_state_gff_15_MUX_inst1_mux_inst_3_U1_X ;
    wire stateFF_state_gff_16_MUX_inst1_mux_inst_0_U1_Y ;
    wire stateFF_state_gff_16_MUX_inst1_mux_inst_0_U1_X ;
    wire stateFF_state_gff_16_MUX_inst1_mux_inst_1_U1_Y ;
    wire stateFF_state_gff_16_MUX_inst1_mux_inst_1_U1_X ;
    wire stateFF_state_gff_16_MUX_inst1_mux_inst_2_U1_Y ;
    wire stateFF_state_gff_16_MUX_inst1_mux_inst_2_U1_X ;
    wire stateFF_state_gff_16_MUX_inst1_mux_inst_3_U1_Y ;
    wire stateFF_state_gff_16_MUX_inst1_mux_inst_3_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_0_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_0_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_1_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_1_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_2_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_2_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_3_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_3_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_4_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_4_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_5_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_5_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_6_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_6_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_7_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_7_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_8_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_8_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_9_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_9_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_10_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_10_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_11_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_11_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_12_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_12_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_13_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_13_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_14_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_14_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_15_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_15_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_16_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_16_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_17_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_17_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_18_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_18_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_19_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_19_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_20_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_20_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_21_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_21_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_22_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_22_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_23_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_23_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_24_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_24_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_25_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_25_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_26_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_26_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_27_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_27_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_28_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_28_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_29_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_29_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_30_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_30_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_31_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_31_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_32_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_32_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_33_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_33_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_34_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_34_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_35_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_35_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_36_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_36_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_37_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_37_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_38_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_38_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_39_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_39_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_40_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_40_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_41_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_41_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_42_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_42_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_43_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_43_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_44_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_44_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_45_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_45_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_46_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_46_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_47_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_47_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_48_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_48_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_49_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_49_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_50_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_50_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_51_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_51_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_52_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_52_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_53_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_53_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_54_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_54_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_55_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_55_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_56_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_56_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_57_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_57_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_58_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_58_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_59_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_59_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_60_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_60_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_61_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_61_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_62_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_62_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_63_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_63_U1_X ;
    wire keyFF_keystate_gff_1_MUX_inst1_mux_inst_0_U1_Y ;
    wire keyFF_keystate_gff_1_MUX_inst1_mux_inst_0_U1_X ;
    wire keyFF_keystate_gff_1_MUX_inst1_mux_inst_1_U1_Y ;
    wire keyFF_keystate_gff_1_MUX_inst1_mux_inst_1_U1_X ;
    wire keyFF_keystate_gff_1_MUX_inst1_mux_inst_2_U1_Y ;
    wire keyFF_keystate_gff_1_MUX_inst1_mux_inst_2_U1_X ;
    wire keyFF_keystate_gff_1_MUX_inst1_mux_inst_3_U1_Y ;
    wire keyFF_keystate_gff_1_MUX_inst1_mux_inst_3_U1_X ;
    wire keyFF_keystate_gff_2_MUX_inst1_mux_inst_0_U1_Y ;
    wire keyFF_keystate_gff_2_MUX_inst1_mux_inst_0_U1_X ;
    wire keyFF_keystate_gff_2_MUX_inst1_mux_inst_1_U1_Y ;
    wire keyFF_keystate_gff_2_MUX_inst1_mux_inst_1_U1_X ;
    wire keyFF_keystate_gff_2_MUX_inst1_mux_inst_2_U1_Y ;
    wire keyFF_keystate_gff_2_MUX_inst1_mux_inst_2_U1_X ;
    wire keyFF_keystate_gff_2_MUX_inst1_mux_inst_3_U1_Y ;
    wire keyFF_keystate_gff_2_MUX_inst1_mux_inst_3_U1_X ;
    wire keyFF_keystate_gff_3_MUX_inst1_mux_inst_0_U1_Y ;
    wire keyFF_keystate_gff_3_MUX_inst1_mux_inst_0_U1_X ;
    wire keyFF_keystate_gff_3_MUX_inst1_mux_inst_1_U1_Y ;
    wire keyFF_keystate_gff_3_MUX_inst1_mux_inst_1_U1_X ;
    wire keyFF_keystate_gff_3_MUX_inst1_mux_inst_2_U1_Y ;
    wire keyFF_keystate_gff_3_MUX_inst1_mux_inst_2_U1_X ;
    wire keyFF_keystate_gff_3_MUX_inst1_mux_inst_3_U1_Y ;
    wire keyFF_keystate_gff_3_MUX_inst1_mux_inst_3_U1_X ;
    wire keyFF_keystate_gff_4_MUX_inst1_mux_inst_0_U1_Y ;
    wire keyFF_keystate_gff_4_MUX_inst1_mux_inst_0_U1_X ;
    wire keyFF_keystate_gff_4_MUX_inst1_mux_inst_1_U1_Y ;
    wire keyFF_keystate_gff_4_MUX_inst1_mux_inst_1_U1_X ;
    wire keyFF_keystate_gff_4_MUX_inst1_mux_inst_2_U1_Y ;
    wire keyFF_keystate_gff_4_MUX_inst1_mux_inst_2_U1_X ;
    wire keyFF_keystate_gff_4_MUX_inst1_mux_inst_3_U1_Y ;
    wire keyFF_keystate_gff_4_MUX_inst1_mux_inst_3_U1_X ;
    wire keyFF_keystate_gff_5_MUX_inst1_mux_inst_0_U1_Y ;
    wire keyFF_keystate_gff_5_MUX_inst1_mux_inst_0_U1_X ;
    wire keyFF_keystate_gff_5_MUX_inst1_mux_inst_1_U1_Y ;
    wire keyFF_keystate_gff_5_MUX_inst1_mux_inst_1_U1_X ;
    wire keyFF_keystate_gff_5_MUX_inst1_mux_inst_2_U1_Y ;
    wire keyFF_keystate_gff_5_MUX_inst1_mux_inst_2_U1_X ;
    wire keyFF_keystate_gff_5_MUX_inst1_mux_inst_3_U1_Y ;
    wire keyFF_keystate_gff_5_MUX_inst1_mux_inst_3_U1_X ;
    wire keyFF_keystate_gff_6_MUX_inst1_mux_inst_0_U1_Y ;
    wire keyFF_keystate_gff_6_MUX_inst1_mux_inst_0_U1_X ;
    wire keyFF_keystate_gff_6_MUX_inst1_mux_inst_1_U1_Y ;
    wire keyFF_keystate_gff_6_MUX_inst1_mux_inst_1_U1_X ;
    wire keyFF_keystate_gff_6_MUX_inst1_mux_inst_2_U1_Y ;
    wire keyFF_keystate_gff_6_MUX_inst1_mux_inst_2_U1_X ;
    wire keyFF_keystate_gff_6_MUX_inst1_mux_inst_3_U1_Y ;
    wire keyFF_keystate_gff_6_MUX_inst1_mux_inst_3_U1_X ;
    wire keyFF_keystate_gff_7_MUX_inst1_mux_inst_0_U1_Y ;
    wire keyFF_keystate_gff_7_MUX_inst1_mux_inst_0_U1_X ;
    wire keyFF_keystate_gff_7_MUX_inst1_mux_inst_1_U1_Y ;
    wire keyFF_keystate_gff_7_MUX_inst1_mux_inst_1_U1_X ;
    wire keyFF_keystate_gff_7_MUX_inst1_mux_inst_2_U1_Y ;
    wire keyFF_keystate_gff_7_MUX_inst1_mux_inst_2_U1_X ;
    wire keyFF_keystate_gff_7_MUX_inst1_mux_inst_3_U1_Y ;
    wire keyFF_keystate_gff_7_MUX_inst1_mux_inst_3_U1_X ;
    wire keyFF_keystate_gff_8_MUX_inst1_mux_inst_0_U1_Y ;
    wire keyFF_keystate_gff_8_MUX_inst1_mux_inst_0_U1_X ;
    wire keyFF_keystate_gff_8_MUX_inst1_mux_inst_1_U1_Y ;
    wire keyFF_keystate_gff_8_MUX_inst1_mux_inst_1_U1_X ;
    wire keyFF_keystate_gff_8_MUX_inst1_mux_inst_2_U1_Y ;
    wire keyFF_keystate_gff_8_MUX_inst1_mux_inst_2_U1_X ;
    wire keyFF_keystate_gff_8_MUX_inst1_mux_inst_3_U1_Y ;
    wire keyFF_keystate_gff_8_MUX_inst1_mux_inst_3_U1_X ;
    wire keyFF_keystate_gff_9_MUX_inst1_mux_inst_0_U1_Y ;
    wire keyFF_keystate_gff_9_MUX_inst1_mux_inst_0_U1_X ;
    wire keyFF_keystate_gff_9_MUX_inst1_mux_inst_1_U1_Y ;
    wire keyFF_keystate_gff_9_MUX_inst1_mux_inst_1_U1_X ;
    wire keyFF_keystate_gff_9_MUX_inst1_mux_inst_2_U1_Y ;
    wire keyFF_keystate_gff_9_MUX_inst1_mux_inst_2_U1_X ;
    wire keyFF_keystate_gff_9_MUX_inst1_mux_inst_3_U1_Y ;
    wire keyFF_keystate_gff_9_MUX_inst1_mux_inst_3_U1_X ;
    wire keyFF_keystate_gff_10_MUX_inst1_mux_inst_0_U1_Y ;
    wire keyFF_keystate_gff_10_MUX_inst1_mux_inst_0_U1_X ;
    wire keyFF_keystate_gff_10_MUX_inst1_mux_inst_1_U1_Y ;
    wire keyFF_keystate_gff_10_MUX_inst1_mux_inst_1_U1_X ;
    wire keyFF_keystate_gff_10_MUX_inst1_mux_inst_2_U1_Y ;
    wire keyFF_keystate_gff_10_MUX_inst1_mux_inst_2_U1_X ;
    wire keyFF_keystate_gff_10_MUX_inst1_mux_inst_3_U1_Y ;
    wire keyFF_keystate_gff_10_MUX_inst1_mux_inst_3_U1_X ;
    wire keyFF_keystate_gff_11_MUX_inst1_mux_inst_0_U1_Y ;
    wire keyFF_keystate_gff_11_MUX_inst1_mux_inst_0_U1_X ;
    wire keyFF_keystate_gff_11_MUX_inst1_mux_inst_1_U1_Y ;
    wire keyFF_keystate_gff_11_MUX_inst1_mux_inst_1_U1_X ;
    wire keyFF_keystate_gff_11_MUX_inst1_mux_inst_2_U1_Y ;
    wire keyFF_keystate_gff_11_MUX_inst1_mux_inst_2_U1_X ;
    wire keyFF_keystate_gff_11_MUX_inst1_mux_inst_3_U1_Y ;
    wire keyFF_keystate_gff_11_MUX_inst1_mux_inst_3_U1_X ;
    wire keyFF_keystate_gff_12_MUX_inst1_mux_inst_0_U1_Y ;
    wire keyFF_keystate_gff_12_MUX_inst1_mux_inst_0_U1_X ;
    wire keyFF_keystate_gff_12_MUX_inst1_mux_inst_1_U1_Y ;
    wire keyFF_keystate_gff_12_MUX_inst1_mux_inst_1_U1_X ;
    wire keyFF_keystate_gff_12_MUX_inst1_mux_inst_2_U1_Y ;
    wire keyFF_keystate_gff_12_MUX_inst1_mux_inst_2_U1_X ;
    wire keyFF_keystate_gff_12_MUX_inst1_mux_inst_3_U1_Y ;
    wire keyFF_keystate_gff_12_MUX_inst1_mux_inst_3_U1_X ;
    wire keyFF_keystate_gff_13_MUX_inst1_mux_inst_0_U1_Y ;
    wire keyFF_keystate_gff_13_MUX_inst1_mux_inst_0_U1_X ;
    wire keyFF_keystate_gff_13_MUX_inst1_mux_inst_1_U1_Y ;
    wire keyFF_keystate_gff_13_MUX_inst1_mux_inst_1_U1_X ;
    wire keyFF_keystate_gff_13_MUX_inst1_mux_inst_2_U1_Y ;
    wire keyFF_keystate_gff_13_MUX_inst1_mux_inst_2_U1_X ;
    wire keyFF_keystate_gff_13_MUX_inst1_mux_inst_3_U1_Y ;
    wire keyFF_keystate_gff_13_MUX_inst1_mux_inst_3_U1_X ;
    wire keyFF_keystate_gff_14_MUX_inst1_mux_inst_0_U1_Y ;
    wire keyFF_keystate_gff_14_MUX_inst1_mux_inst_0_U1_X ;
    wire keyFF_keystate_gff_14_MUX_inst1_mux_inst_1_U1_Y ;
    wire keyFF_keystate_gff_14_MUX_inst1_mux_inst_1_U1_X ;
    wire keyFF_keystate_gff_14_MUX_inst1_mux_inst_2_U1_Y ;
    wire keyFF_keystate_gff_14_MUX_inst1_mux_inst_2_U1_X ;
    wire keyFF_keystate_gff_14_MUX_inst1_mux_inst_3_U1_Y ;
    wire keyFF_keystate_gff_14_MUX_inst1_mux_inst_3_U1_X ;
    wire keyFF_keystate_gff_15_MUX_inst1_mux_inst_0_U1_Y ;
    wire keyFF_keystate_gff_15_MUX_inst1_mux_inst_0_U1_X ;
    wire keyFF_keystate_gff_15_MUX_inst1_mux_inst_1_U1_Y ;
    wire keyFF_keystate_gff_15_MUX_inst1_mux_inst_1_U1_X ;
    wire keyFF_keystate_gff_15_MUX_inst1_mux_inst_2_U1_Y ;
    wire keyFF_keystate_gff_15_MUX_inst1_mux_inst_2_U1_X ;
    wire keyFF_keystate_gff_15_MUX_inst1_mux_inst_3_U1_Y ;
    wire keyFF_keystate_gff_15_MUX_inst1_mux_inst_3_U1_X ;
    wire keyFF_keystate_gff_16_MUX_inst1_mux_inst_0_U1_Y ;
    wire keyFF_keystate_gff_16_MUX_inst1_mux_inst_0_U1_X ;
    wire keyFF_keystate_gff_16_MUX_inst1_mux_inst_1_U1_Y ;
    wire keyFF_keystate_gff_16_MUX_inst1_mux_inst_1_U1_X ;
    wire keyFF_keystate_gff_16_MUX_inst1_mux_inst_2_U1_Y ;
    wire keyFF_keystate_gff_16_MUX_inst1_mux_inst_2_U1_X ;
    wire keyFF_keystate_gff_16_MUX_inst1_mux_inst_3_U1_Y ;
    wire keyFF_keystate_gff_16_MUX_inst1_mux_inst_3_U1_X ;
    wire keyFF_keystate_gff_17_MUX_inst1_mux_inst_0_U1_Y ;
    wire keyFF_keystate_gff_17_MUX_inst1_mux_inst_0_U1_X ;
    wire keyFF_keystate_gff_17_MUX_inst1_mux_inst_1_U1_Y ;
    wire keyFF_keystate_gff_17_MUX_inst1_mux_inst_1_U1_X ;
    wire keyFF_keystate_gff_17_MUX_inst1_mux_inst_2_U1_Y ;
    wire keyFF_keystate_gff_17_MUX_inst1_mux_inst_2_U1_X ;
    wire keyFF_keystate_gff_17_MUX_inst1_mux_inst_3_U1_Y ;
    wire keyFF_keystate_gff_17_MUX_inst1_mux_inst_3_U1_X ;
    wire keyFF_keystate_gff_18_MUX_inst1_mux_inst_0_U1_Y ;
    wire keyFF_keystate_gff_18_MUX_inst1_mux_inst_0_U1_X ;
    wire keyFF_keystate_gff_18_MUX_inst1_mux_inst_1_U1_Y ;
    wire keyFF_keystate_gff_18_MUX_inst1_mux_inst_1_U1_X ;
    wire keyFF_keystate_gff_18_MUX_inst1_mux_inst_2_U1_Y ;
    wire keyFF_keystate_gff_18_MUX_inst1_mux_inst_2_U1_X ;
    wire keyFF_keystate_gff_18_MUX_inst1_mux_inst_3_U1_Y ;
    wire keyFF_keystate_gff_18_MUX_inst1_mux_inst_3_U1_X ;
    wire keyFF_keystate_gff_19_MUX_inst1_mux_inst_0_U1_Y ;
    wire keyFF_keystate_gff_19_MUX_inst1_mux_inst_0_U1_X ;
    wire keyFF_keystate_gff_19_MUX_inst1_mux_inst_1_U1_Y ;
    wire keyFF_keystate_gff_19_MUX_inst1_mux_inst_1_U1_X ;
    wire keyFF_keystate_gff_19_MUX_inst1_mux_inst_2_U1_Y ;
    wire keyFF_keystate_gff_19_MUX_inst1_mux_inst_2_U1_X ;
    wire keyFF_keystate_gff_19_MUX_inst1_mux_inst_3_U1_Y ;
    wire keyFF_keystate_gff_19_MUX_inst1_mux_inst_3_U1_X ;
    wire keyFF_keystate_gff_20_MUX_inst1_mux_inst_0_U1_Y ;
    wire keyFF_keystate_gff_20_MUX_inst1_mux_inst_0_U1_X ;
    wire keyFF_keystate_gff_20_MUX_inst1_mux_inst_1_U1_Y ;
    wire keyFF_keystate_gff_20_MUX_inst1_mux_inst_1_U1_X ;
    wire keyFF_keystate_gff_20_MUX_inst1_mux_inst_2_U1_Y ;
    wire keyFF_keystate_gff_20_MUX_inst1_mux_inst_2_U1_X ;
    wire keyFF_keystate_gff_20_MUX_inst1_mux_inst_3_U1_Y ;
    wire keyFF_keystate_gff_20_MUX_inst1_mux_inst_3_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_0_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_0_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_1_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_1_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_2_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_2_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_3_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_3_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_4_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_4_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_5_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_5_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_6_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_6_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_7_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_7_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_8_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_8_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_9_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_9_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_10_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_10_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_11_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_11_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_12_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_12_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_13_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_13_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_14_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_14_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_15_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_15_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_16_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_16_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_17_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_17_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_18_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_18_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_19_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_19_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_20_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_20_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_21_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_21_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_22_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_22_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_23_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_23_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_24_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_24_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_25_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_25_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_26_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_26_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_27_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_27_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_28_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_28_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_29_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_29_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_30_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_30_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_31_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_31_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_32_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_32_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_33_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_33_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_34_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_34_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_35_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_35_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_36_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_36_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_37_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_37_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_38_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_38_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_39_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_39_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_40_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_40_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_41_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_41_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_42_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_42_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_43_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_43_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_44_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_44_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_45_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_45_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_46_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_46_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_47_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_47_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_48_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_48_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_49_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_49_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_50_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_50_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_51_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_51_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_52_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_52_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_53_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_53_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_54_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_54_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_55_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_55_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_56_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_56_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_57_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_57_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_58_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_58_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_59_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_59_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_60_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_60_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_61_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_61_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_62_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_62_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_63_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_63_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_64_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_64_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_65_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_65_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_66_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_66_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_67_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_67_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_68_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_68_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_69_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_69_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_70_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_70_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_71_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_71_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_72_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_72_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_73_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_73_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_74_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_74_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_75_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_75_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_76_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_76_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_77_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_77_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_78_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_78_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_79_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_79_U1_X ;
    wire sboxInst_L8 ;
    wire sboxInst_L7 ;
    wire sboxInst_T3 ;
    wire sboxInst_T1 ;
    wire sboxInst_Q7 ;
    wire sboxInst_Q6 ;
    wire sboxInst_L5 ;
    wire sboxInst_T2 ;
    wire sboxInst_L4 ;
    wire sboxInst_Q3 ;
    wire sboxInst_L3 ;
    wire sboxInst_Q2 ;
    wire sboxInst_T0 ;
    wire sboxInst_L2 ;
    wire sboxInst_L1 ;
    wire sboxInst_L0 ;
    wire MUX_sboxin_mux_inst_0_U1_Y ;
    wire MUX_sboxin_mux_inst_0_U1_X ;
    wire MUX_sboxin_mux_inst_1_U1_Y ;
    wire MUX_sboxin_mux_inst_1_U1_X ;
    wire MUX_sboxin_mux_inst_2_U1_Y ;
    wire MUX_sboxin_mux_inst_2_U1_X ;
    wire MUX_sboxin_mux_inst_3_U1_Y ;
    wire MUX_sboxin_mux_inst_3_U1_X ;
    wire MUX_serialIn_mux_inst_0_U1_Y ;
    wire MUX_serialIn_mux_inst_0_U1_X ;
    wire MUX_serialIn_mux_inst_1_U1_Y ;
    wire MUX_serialIn_mux_inst_1_U1_X ;
    wire MUX_serialIn_mux_inst_2_U1_Y ;
    wire MUX_serialIn_mux_inst_2_U1_X ;
    wire MUX_serialIn_mux_inst_3_U1_Y ;
    wire MUX_serialIn_mux_inst_3_U1_X ;
    wire [4:0] counter ;
    wire [3:0] serialIn ;
    wire [3:0] sboxOut ;
    wire [3:0] roundkey ;
    wire [3:1] keyRegKS ;
    wire [3:0] sboxIn ;
    wire [3:0] stateXORroundkey ;
    wire [3:0] fsm_countSerial ;
    wire [63:0] stateFF_inputPar ;
    wire [4:0] keyFF_counterAdd ;
    wire [75:3] keyFF_outputPar ;
    wire [79:0] keyFF_inputPar ;

    /* cells in depth 0 */
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U9 ( .A0_t (roundkey[1]), .B0_t (data_out[61]), .Z0_t (stateXORroundkey[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U10 ( .A0_t (roundkey[2]), .B0_t (data_out[62]), .Z0_t (stateXORroundkey[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U11 ( .A0_t (roundkey[0]), .B0_t (data_out[60]), .Z0_t (stateXORroundkey[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U12 ( .A0_t (roundkey[3]), .B0_t (data_out[63]), .Z0_t (stateXORroundkey[3]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) fsm_U19 ( .A0_t (reset), .B0_t (fsm_n14), .Z0_t (fsm_n16) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) fsm_U18 ( .A0_t (fsm_n16), .B0_t (fsm_n13), .Z0_t (fsm_n14) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) fsm_U17 ( .A0_t (fsm_n12), .B0_t (fsm_n11), .Z0_t (fsm_n13) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) fsm_U16 ( .A0_t (counter[3]), .B0_t (fsm_ps_state_0_), .Z0_t (fsm_n11) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) fsm_U15 ( .A0_t (fsm_n10), .B0_t (fsm_n9), .Z0_t (fsm_n12) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) fsm_U14 ( .A0_t (counter[4]), .B0_t (counter[0]), .Z0_t (fsm_n9) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) fsm_U13 ( .A0_t (counter[1]), .B0_t (counter[2]), .Z0_t (fsm_n10) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) fsm_U12 ( .A0_t (fsm_n16), .B0_t (fsm_ps_state_0_), .Z0_t (intDone) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) fsm_U11 ( .A0_t (fsm_n8), .B0_t (fsm_n16), .Z0_t (fsm_en_countRound) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) fsm_U10 ( .A0_t (reset), .B0_t (fsm_n7), .Z0_t (fsm_ps_state_0_) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) fsm_U9 ( .A0_t (fsm_n8), .B0_t (done), .Z0_t (fsm_n7) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) fsm_U8 ( .A0_t (fsm_countSerial[1]), .B0_t (fsm_n6), .Z0_t (fsm_n8) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) fsm_U7 ( .A0_t (fsm_n5), .B0_t (fsm_n4), .Z0_t (fsm_n6) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) fsm_U6 ( .A0_t (fsm_countSerial[3]), .B0_t (fsm_countSerial[2]), .Z0_t (fsm_n4) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) fsm_U5 ( .A0_t (fsm_ps_state_0_), .B0_t (fsm_countSerial[0]), .Z0_t (fsm_n5) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) fsm_U4 ( .A0_t (fsm_ps_state_0_), .B0_t (fsm_n16), .Z0_t (done) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) fsm_U2 ( .A0_t (reset), .B0_t (selSbox), .Z0_t (fsm_rst_countSerial) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) fsm_U1 ( .A0_t (fsm_ps_state_0_), .B0_t (fsm_n16), .Z0_t (selSbox) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) fsm_cnt_rnd_U15 ( .A0_t (fsm_cnt_rnd_n12), .B0_t (reset), .Z0_t (counter[2]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b0)) fsm_cnt_rnd_U14 ( .A0_t (fsm_cnt_rnd_n10), .B0_t (counter[2]), .Z0_t (fsm_cnt_rnd_n12) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) fsm_cnt_rnd_U13 ( .A0_t (fsm_cnt_rnd_n9), .B0_t (reset), .Z0_t (counter[0]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b0)) fsm_cnt_rnd_U12 ( .A0_t (counter[0]), .B0_t (fsm_en_countRound), .Z0_t (fsm_cnt_rnd_n9) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) fsm_cnt_rnd_U11 ( .A0_t (fsm_cnt_rnd_n8), .B0_t (reset), .Z0_t (counter[4]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b0)) fsm_cnt_rnd_U10 ( .A0_t (counter[4]), .B0_t (fsm_cnt_rnd_n7), .Z0_t (fsm_cnt_rnd_n8) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) fsm_cnt_rnd_U9 ( .A0_t (counter[3]), .B0_t (fsm_cnt_rnd_n6), .Z0_t (fsm_cnt_rnd_n7) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) fsm_cnt_rnd_U8 ( .A0_t (reset), .B0_t (fsm_cnt_rnd_n5), .Z0_t (counter[1]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) fsm_cnt_rnd_U7 ( .A0_t (counter[1]), .B0_t (fsm_cnt_rnd_n4), .Z0_t (fsm_cnt_rnd_n5) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) fsm_cnt_rnd_U6 ( .A0_t (fsm_cnt_rnd_n3), .B0_t (reset), .Z0_t (counter[3]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b0)) fsm_cnt_rnd_U4 ( .A0_t (fsm_cnt_rnd_n6), .B0_t (counter[3]), .Z0_t (fsm_cnt_rnd_n3) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) fsm_cnt_rnd_U3 ( .A0_t (fsm_cnt_rnd_n10), .B0_t (counter[2]), .Z0_t (fsm_cnt_rnd_n6) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) fsm_cnt_rnd_U2 ( .A0_t (counter[1]), .B0_t (fsm_cnt_rnd_n4), .Z0_t (fsm_cnt_rnd_n10) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) fsm_cnt_rnd_U1 ( .A0_t (counter[0]), .B0_t (fsm_en_countRound), .Z0_t (fsm_cnt_rnd_n4) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) fsm_cnt_ser_U12 ( .A0_t (fsm_cnt_ser_n9), .B0_t (fsm_rst_countSerial), .Z0_t (fsm_countSerial[0]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b0)) fsm_cnt_ser_U11 ( .A0_t (fsm_ps_state_0_), .B0_t (fsm_countSerial[0]), .Z0_t (fsm_cnt_ser_n9) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) fsm_cnt_ser_U10 ( .A0_t (fsm_cnt_ser_n7), .B0_t (fsm_rst_countSerial), .Z0_t (fsm_countSerial[1]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b0)) fsm_cnt_ser_U9 ( .A0_t (fsm_cnt_ser_n6), .B0_t (fsm_countSerial[1]), .Z0_t (fsm_cnt_ser_n7) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) fsm_cnt_ser_U8 ( .A0_t (fsm_cnt_ser_n5), .B0_t (fsm_rst_countSerial), .Z0_t (fsm_countSerial[3]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b0)) fsm_cnt_ser_U7 ( .A0_t (fsm_countSerial[3]), .B0_t (fsm_cnt_ser_n4), .Z0_t (fsm_cnt_ser_n5) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) fsm_cnt_ser_U6 ( .A0_t (fsm_countSerial[2]), .B0_t (fsm_cnt_ser_n3), .Z0_t (fsm_cnt_ser_n4) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) fsm_cnt_ser_U5 ( .A0_t (fsm_cnt_ser_n2), .B0_t (fsm_rst_countSerial), .Z0_t (fsm_countSerial[2]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b0)) fsm_cnt_ser_U3 ( .A0_t (fsm_cnt_ser_n3), .B0_t (fsm_countSerial[2]), .Z0_t (fsm_cnt_ser_n2) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) fsm_cnt_ser_U2 ( .A0_t (fsm_cnt_ser_n6), .B0_t (fsm_countSerial[1]), .Z0_t (fsm_cnt_ser_n3) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) fsm_cnt_ser_U1 ( .A0_t (fsm_ps_state_0_), .B0_t (fsm_countSerial[0]), .Z0_t (fsm_cnt_ser_n6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_1_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (serialIn[0]), .B0_t (stateFF_inputPar[0]), .Z0_t (stateFF_state_gff_1_MUX_inst1_mux_inst_0_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_1_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (stateFF_state_gff_1_MUX_inst1_mux_inst_0_U1_X), .Z0_t (stateFF_state_gff_1_MUX_inst1_mux_inst_0_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_1_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_1_MUX_inst1_mux_inst_0_U1_Y), .B0_t (serialIn[0]), .Z0_t (data_out[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_1_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (serialIn[1]), .B0_t (stateFF_inputPar[1]), .Z0_t (stateFF_state_gff_1_MUX_inst1_mux_inst_1_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_1_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (stateFF_state_gff_1_MUX_inst1_mux_inst_1_U1_X), .Z0_t (stateFF_state_gff_1_MUX_inst1_mux_inst_1_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_1_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_1_MUX_inst1_mux_inst_1_U1_Y), .B0_t (serialIn[1]), .Z0_t (data_out[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_1_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (serialIn[2]), .B0_t (stateFF_inputPar[2]), .Z0_t (stateFF_state_gff_1_MUX_inst1_mux_inst_2_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_1_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (stateFF_state_gff_1_MUX_inst1_mux_inst_2_U1_X), .Z0_t (stateFF_state_gff_1_MUX_inst1_mux_inst_2_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_1_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_1_MUX_inst1_mux_inst_2_U1_Y), .B0_t (serialIn[2]), .Z0_t (data_out[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_1_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (serialIn[3]), .B0_t (stateFF_inputPar[3]), .Z0_t (stateFF_state_gff_1_MUX_inst1_mux_inst_3_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_1_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (stateFF_state_gff_1_MUX_inst1_mux_inst_3_U1_X), .Z0_t (stateFF_state_gff_1_MUX_inst1_mux_inst_3_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_1_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_1_MUX_inst1_mux_inst_3_U1_Y), .B0_t (serialIn[3]), .Z0_t (data_out[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_2_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (data_out[0]), .B0_t (stateFF_inputPar[4]), .Z0_t (stateFF_state_gff_2_MUX_inst1_mux_inst_0_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_2_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (stateFF_state_gff_2_MUX_inst1_mux_inst_0_U1_X), .Z0_t (stateFF_state_gff_2_MUX_inst1_mux_inst_0_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_2_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_2_MUX_inst1_mux_inst_0_U1_Y), .B0_t (data_out[0]), .Z0_t (data_out[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_2_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (data_out[1]), .B0_t (stateFF_inputPar[5]), .Z0_t (stateFF_state_gff_2_MUX_inst1_mux_inst_1_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_2_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (stateFF_state_gff_2_MUX_inst1_mux_inst_1_U1_X), .Z0_t (stateFF_state_gff_2_MUX_inst1_mux_inst_1_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_2_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_2_MUX_inst1_mux_inst_1_U1_Y), .B0_t (data_out[1]), .Z0_t (data_out[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_2_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (data_out[2]), .B0_t (stateFF_inputPar[6]), .Z0_t (stateFF_state_gff_2_MUX_inst1_mux_inst_2_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_2_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (stateFF_state_gff_2_MUX_inst1_mux_inst_2_U1_X), .Z0_t (stateFF_state_gff_2_MUX_inst1_mux_inst_2_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_2_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_2_MUX_inst1_mux_inst_2_U1_Y), .B0_t (data_out[2]), .Z0_t (data_out[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_2_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (data_out[3]), .B0_t (stateFF_inputPar[7]), .Z0_t (stateFF_state_gff_2_MUX_inst1_mux_inst_3_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_2_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (stateFF_state_gff_2_MUX_inst1_mux_inst_3_U1_X), .Z0_t (stateFF_state_gff_2_MUX_inst1_mux_inst_3_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_2_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_2_MUX_inst1_mux_inst_3_U1_Y), .B0_t (data_out[3]), .Z0_t (data_out[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_3_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (data_out[4]), .B0_t (stateFF_inputPar[8]), .Z0_t (stateFF_state_gff_3_MUX_inst1_mux_inst_0_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_3_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (stateFF_state_gff_3_MUX_inst1_mux_inst_0_U1_X), .Z0_t (stateFF_state_gff_3_MUX_inst1_mux_inst_0_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_3_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_3_MUX_inst1_mux_inst_0_U1_Y), .B0_t (data_out[4]), .Z0_t (data_out[8]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_3_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (data_out[5]), .B0_t (stateFF_inputPar[9]), .Z0_t (stateFF_state_gff_3_MUX_inst1_mux_inst_1_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_3_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (stateFF_state_gff_3_MUX_inst1_mux_inst_1_U1_X), .Z0_t (stateFF_state_gff_3_MUX_inst1_mux_inst_1_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_3_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_3_MUX_inst1_mux_inst_1_U1_Y), .B0_t (data_out[5]), .Z0_t (data_out[9]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_3_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (data_out[6]), .B0_t (stateFF_inputPar[10]), .Z0_t (stateFF_state_gff_3_MUX_inst1_mux_inst_2_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_3_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (stateFF_state_gff_3_MUX_inst1_mux_inst_2_U1_X), .Z0_t (stateFF_state_gff_3_MUX_inst1_mux_inst_2_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_3_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_3_MUX_inst1_mux_inst_2_U1_Y), .B0_t (data_out[6]), .Z0_t (data_out[10]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_3_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (data_out[7]), .B0_t (stateFF_inputPar[11]), .Z0_t (stateFF_state_gff_3_MUX_inst1_mux_inst_3_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_3_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (stateFF_state_gff_3_MUX_inst1_mux_inst_3_U1_X), .Z0_t (stateFF_state_gff_3_MUX_inst1_mux_inst_3_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_3_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_3_MUX_inst1_mux_inst_3_U1_Y), .B0_t (data_out[7]), .Z0_t (data_out[11]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_4_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (data_out[8]), .B0_t (stateFF_inputPar[12]), .Z0_t (stateFF_state_gff_4_MUX_inst1_mux_inst_0_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_4_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (stateFF_state_gff_4_MUX_inst1_mux_inst_0_U1_X), .Z0_t (stateFF_state_gff_4_MUX_inst1_mux_inst_0_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_4_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_4_MUX_inst1_mux_inst_0_U1_Y), .B0_t (data_out[8]), .Z0_t (data_out[12]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_4_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (data_out[9]), .B0_t (stateFF_inputPar[13]), .Z0_t (stateFF_state_gff_4_MUX_inst1_mux_inst_1_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_4_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (stateFF_state_gff_4_MUX_inst1_mux_inst_1_U1_X), .Z0_t (stateFF_state_gff_4_MUX_inst1_mux_inst_1_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_4_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_4_MUX_inst1_mux_inst_1_U1_Y), .B0_t (data_out[9]), .Z0_t (data_out[13]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_4_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (data_out[10]), .B0_t (stateFF_inputPar[14]), .Z0_t (stateFF_state_gff_4_MUX_inst1_mux_inst_2_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_4_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (stateFF_state_gff_4_MUX_inst1_mux_inst_2_U1_X), .Z0_t (stateFF_state_gff_4_MUX_inst1_mux_inst_2_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_4_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_4_MUX_inst1_mux_inst_2_U1_Y), .B0_t (data_out[10]), .Z0_t (data_out[14]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_4_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (data_out[11]), .B0_t (stateFF_inputPar[15]), .Z0_t (stateFF_state_gff_4_MUX_inst1_mux_inst_3_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_4_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (stateFF_state_gff_4_MUX_inst1_mux_inst_3_U1_X), .Z0_t (stateFF_state_gff_4_MUX_inst1_mux_inst_3_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_4_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_4_MUX_inst1_mux_inst_3_U1_Y), .B0_t (data_out[11]), .Z0_t (data_out[15]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_5_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (data_out[12]), .B0_t (stateFF_inputPar[16]), .Z0_t (stateFF_state_gff_5_MUX_inst1_mux_inst_0_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_5_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (stateFF_state_gff_5_MUX_inst1_mux_inst_0_U1_X), .Z0_t (stateFF_state_gff_5_MUX_inst1_mux_inst_0_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_5_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_5_MUX_inst1_mux_inst_0_U1_Y), .B0_t (data_out[12]), .Z0_t (data_out[16]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_5_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (data_out[13]), .B0_t (stateFF_inputPar[17]), .Z0_t (stateFF_state_gff_5_MUX_inst1_mux_inst_1_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_5_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (stateFF_state_gff_5_MUX_inst1_mux_inst_1_U1_X), .Z0_t (stateFF_state_gff_5_MUX_inst1_mux_inst_1_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_5_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_5_MUX_inst1_mux_inst_1_U1_Y), .B0_t (data_out[13]), .Z0_t (data_out[17]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_5_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (data_out[14]), .B0_t (stateFF_inputPar[18]), .Z0_t (stateFF_state_gff_5_MUX_inst1_mux_inst_2_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_5_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (stateFF_state_gff_5_MUX_inst1_mux_inst_2_U1_X), .Z0_t (stateFF_state_gff_5_MUX_inst1_mux_inst_2_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_5_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_5_MUX_inst1_mux_inst_2_U1_Y), .B0_t (data_out[14]), .Z0_t (data_out[18]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_5_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (data_out[15]), .B0_t (stateFF_inputPar[19]), .Z0_t (stateFF_state_gff_5_MUX_inst1_mux_inst_3_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_5_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (stateFF_state_gff_5_MUX_inst1_mux_inst_3_U1_X), .Z0_t (stateFF_state_gff_5_MUX_inst1_mux_inst_3_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_5_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_5_MUX_inst1_mux_inst_3_U1_Y), .B0_t (data_out[15]), .Z0_t (data_out[19]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_6_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (data_out[16]), .B0_t (stateFF_inputPar[20]), .Z0_t (stateFF_state_gff_6_MUX_inst1_mux_inst_0_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_6_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (stateFF_state_gff_6_MUX_inst1_mux_inst_0_U1_X), .Z0_t (stateFF_state_gff_6_MUX_inst1_mux_inst_0_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_6_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_6_MUX_inst1_mux_inst_0_U1_Y), .B0_t (data_out[16]), .Z0_t (data_out[20]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_6_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (data_out[17]), .B0_t (stateFF_inputPar[21]), .Z0_t (stateFF_state_gff_6_MUX_inst1_mux_inst_1_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_6_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (stateFF_state_gff_6_MUX_inst1_mux_inst_1_U1_X), .Z0_t (stateFF_state_gff_6_MUX_inst1_mux_inst_1_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_6_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_6_MUX_inst1_mux_inst_1_U1_Y), .B0_t (data_out[17]), .Z0_t (data_out[21]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_6_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (data_out[18]), .B0_t (stateFF_inputPar[22]), .Z0_t (stateFF_state_gff_6_MUX_inst1_mux_inst_2_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_6_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (stateFF_state_gff_6_MUX_inst1_mux_inst_2_U1_X), .Z0_t (stateFF_state_gff_6_MUX_inst1_mux_inst_2_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_6_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_6_MUX_inst1_mux_inst_2_U1_Y), .B0_t (data_out[18]), .Z0_t (data_out[22]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_6_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (data_out[19]), .B0_t (stateFF_inputPar[23]), .Z0_t (stateFF_state_gff_6_MUX_inst1_mux_inst_3_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_6_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (stateFF_state_gff_6_MUX_inst1_mux_inst_3_U1_X), .Z0_t (stateFF_state_gff_6_MUX_inst1_mux_inst_3_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_6_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_6_MUX_inst1_mux_inst_3_U1_Y), .B0_t (data_out[19]), .Z0_t (data_out[23]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_7_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (data_out[20]), .B0_t (stateFF_inputPar[24]), .Z0_t (stateFF_state_gff_7_MUX_inst1_mux_inst_0_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_7_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (stateFF_state_gff_7_MUX_inst1_mux_inst_0_U1_X), .Z0_t (stateFF_state_gff_7_MUX_inst1_mux_inst_0_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_7_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_7_MUX_inst1_mux_inst_0_U1_Y), .B0_t (data_out[20]), .Z0_t (data_out[24]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_7_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (data_out[21]), .B0_t (stateFF_inputPar[25]), .Z0_t (stateFF_state_gff_7_MUX_inst1_mux_inst_1_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_7_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (stateFF_state_gff_7_MUX_inst1_mux_inst_1_U1_X), .Z0_t (stateFF_state_gff_7_MUX_inst1_mux_inst_1_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_7_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_7_MUX_inst1_mux_inst_1_U1_Y), .B0_t (data_out[21]), .Z0_t (data_out[25]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_7_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (data_out[22]), .B0_t (stateFF_inputPar[26]), .Z0_t (stateFF_state_gff_7_MUX_inst1_mux_inst_2_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_7_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (stateFF_state_gff_7_MUX_inst1_mux_inst_2_U1_X), .Z0_t (stateFF_state_gff_7_MUX_inst1_mux_inst_2_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_7_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_7_MUX_inst1_mux_inst_2_U1_Y), .B0_t (data_out[22]), .Z0_t (data_out[26]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_7_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (data_out[23]), .B0_t (stateFF_inputPar[27]), .Z0_t (stateFF_state_gff_7_MUX_inst1_mux_inst_3_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_7_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (stateFF_state_gff_7_MUX_inst1_mux_inst_3_U1_X), .Z0_t (stateFF_state_gff_7_MUX_inst1_mux_inst_3_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_7_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_7_MUX_inst1_mux_inst_3_U1_Y), .B0_t (data_out[23]), .Z0_t (data_out[27]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_8_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (data_out[24]), .B0_t (stateFF_inputPar[28]), .Z0_t (stateFF_state_gff_8_MUX_inst1_mux_inst_0_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_8_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (stateFF_state_gff_8_MUX_inst1_mux_inst_0_U1_X), .Z0_t (stateFF_state_gff_8_MUX_inst1_mux_inst_0_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_8_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_8_MUX_inst1_mux_inst_0_U1_Y), .B0_t (data_out[24]), .Z0_t (data_out[28]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_8_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (data_out[25]), .B0_t (stateFF_inputPar[29]), .Z0_t (stateFF_state_gff_8_MUX_inst1_mux_inst_1_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_8_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (stateFF_state_gff_8_MUX_inst1_mux_inst_1_U1_X), .Z0_t (stateFF_state_gff_8_MUX_inst1_mux_inst_1_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_8_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_8_MUX_inst1_mux_inst_1_U1_Y), .B0_t (data_out[25]), .Z0_t (data_out[29]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_8_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (data_out[26]), .B0_t (stateFF_inputPar[30]), .Z0_t (stateFF_state_gff_8_MUX_inst1_mux_inst_2_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_8_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (stateFF_state_gff_8_MUX_inst1_mux_inst_2_U1_X), .Z0_t (stateFF_state_gff_8_MUX_inst1_mux_inst_2_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_8_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_8_MUX_inst1_mux_inst_2_U1_Y), .B0_t (data_out[26]), .Z0_t (data_out[30]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_8_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (data_out[27]), .B0_t (stateFF_inputPar[31]), .Z0_t (stateFF_state_gff_8_MUX_inst1_mux_inst_3_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_8_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (stateFF_state_gff_8_MUX_inst1_mux_inst_3_U1_X), .Z0_t (stateFF_state_gff_8_MUX_inst1_mux_inst_3_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_8_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_8_MUX_inst1_mux_inst_3_U1_Y), .B0_t (data_out[27]), .Z0_t (data_out[31]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_9_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (data_out[28]), .B0_t (stateFF_inputPar[32]), .Z0_t (stateFF_state_gff_9_MUX_inst1_mux_inst_0_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_9_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (stateFF_state_gff_9_MUX_inst1_mux_inst_0_U1_X), .Z0_t (stateFF_state_gff_9_MUX_inst1_mux_inst_0_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_9_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_9_MUX_inst1_mux_inst_0_U1_Y), .B0_t (data_out[28]), .Z0_t (data_out[32]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_9_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (data_out[29]), .B0_t (stateFF_inputPar[33]), .Z0_t (stateFF_state_gff_9_MUX_inst1_mux_inst_1_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_9_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (stateFF_state_gff_9_MUX_inst1_mux_inst_1_U1_X), .Z0_t (stateFF_state_gff_9_MUX_inst1_mux_inst_1_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_9_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_9_MUX_inst1_mux_inst_1_U1_Y), .B0_t (data_out[29]), .Z0_t (data_out[33]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_9_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (data_out[30]), .B0_t (stateFF_inputPar[34]), .Z0_t (stateFF_state_gff_9_MUX_inst1_mux_inst_2_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_9_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (stateFF_state_gff_9_MUX_inst1_mux_inst_2_U1_X), .Z0_t (stateFF_state_gff_9_MUX_inst1_mux_inst_2_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_9_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_9_MUX_inst1_mux_inst_2_U1_Y), .B0_t (data_out[30]), .Z0_t (data_out[34]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_9_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (data_out[31]), .B0_t (stateFF_inputPar[35]), .Z0_t (stateFF_state_gff_9_MUX_inst1_mux_inst_3_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_9_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (stateFF_state_gff_9_MUX_inst1_mux_inst_3_U1_X), .Z0_t (stateFF_state_gff_9_MUX_inst1_mux_inst_3_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_9_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_9_MUX_inst1_mux_inst_3_U1_Y), .B0_t (data_out[31]), .Z0_t (data_out[35]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_10_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (data_out[32]), .B0_t (stateFF_inputPar[36]), .Z0_t (stateFF_state_gff_10_MUX_inst1_mux_inst_0_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_10_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (stateFF_state_gff_10_MUX_inst1_mux_inst_0_U1_X), .Z0_t (stateFF_state_gff_10_MUX_inst1_mux_inst_0_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_10_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_10_MUX_inst1_mux_inst_0_U1_Y), .B0_t (data_out[32]), .Z0_t (data_out[36]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_10_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (data_out[33]), .B0_t (stateFF_inputPar[37]), .Z0_t (stateFF_state_gff_10_MUX_inst1_mux_inst_1_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_10_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (stateFF_state_gff_10_MUX_inst1_mux_inst_1_U1_X), .Z0_t (stateFF_state_gff_10_MUX_inst1_mux_inst_1_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_10_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_10_MUX_inst1_mux_inst_1_U1_Y), .B0_t (data_out[33]), .Z0_t (data_out[37]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_10_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (data_out[34]), .B0_t (stateFF_inputPar[38]), .Z0_t (stateFF_state_gff_10_MUX_inst1_mux_inst_2_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_10_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (stateFF_state_gff_10_MUX_inst1_mux_inst_2_U1_X), .Z0_t (stateFF_state_gff_10_MUX_inst1_mux_inst_2_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_10_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_10_MUX_inst1_mux_inst_2_U1_Y), .B0_t (data_out[34]), .Z0_t (data_out[38]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_10_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (data_out[35]), .B0_t (stateFF_inputPar[39]), .Z0_t (stateFF_state_gff_10_MUX_inst1_mux_inst_3_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_10_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (stateFF_state_gff_10_MUX_inst1_mux_inst_3_U1_X), .Z0_t (stateFF_state_gff_10_MUX_inst1_mux_inst_3_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_10_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_10_MUX_inst1_mux_inst_3_U1_Y), .B0_t (data_out[35]), .Z0_t (data_out[39]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_11_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (data_out[36]), .B0_t (stateFF_inputPar[40]), .Z0_t (stateFF_state_gff_11_MUX_inst1_mux_inst_0_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_11_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (stateFF_state_gff_11_MUX_inst1_mux_inst_0_U1_X), .Z0_t (stateFF_state_gff_11_MUX_inst1_mux_inst_0_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_11_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_11_MUX_inst1_mux_inst_0_U1_Y), .B0_t (data_out[36]), .Z0_t (data_out[40]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_11_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (data_out[37]), .B0_t (stateFF_inputPar[41]), .Z0_t (stateFF_state_gff_11_MUX_inst1_mux_inst_1_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_11_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (stateFF_state_gff_11_MUX_inst1_mux_inst_1_U1_X), .Z0_t (stateFF_state_gff_11_MUX_inst1_mux_inst_1_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_11_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_11_MUX_inst1_mux_inst_1_U1_Y), .B0_t (data_out[37]), .Z0_t (data_out[41]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_11_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (data_out[38]), .B0_t (stateFF_inputPar[42]), .Z0_t (stateFF_state_gff_11_MUX_inst1_mux_inst_2_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_11_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (stateFF_state_gff_11_MUX_inst1_mux_inst_2_U1_X), .Z0_t (stateFF_state_gff_11_MUX_inst1_mux_inst_2_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_11_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_11_MUX_inst1_mux_inst_2_U1_Y), .B0_t (data_out[38]), .Z0_t (data_out[42]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_11_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (data_out[39]), .B0_t (stateFF_inputPar[43]), .Z0_t (stateFF_state_gff_11_MUX_inst1_mux_inst_3_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_11_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (stateFF_state_gff_11_MUX_inst1_mux_inst_3_U1_X), .Z0_t (stateFF_state_gff_11_MUX_inst1_mux_inst_3_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_11_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_11_MUX_inst1_mux_inst_3_U1_Y), .B0_t (data_out[39]), .Z0_t (data_out[43]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_12_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (data_out[40]), .B0_t (stateFF_inputPar[44]), .Z0_t (stateFF_state_gff_12_MUX_inst1_mux_inst_0_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_12_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (stateFF_state_gff_12_MUX_inst1_mux_inst_0_U1_X), .Z0_t (stateFF_state_gff_12_MUX_inst1_mux_inst_0_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_12_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_12_MUX_inst1_mux_inst_0_U1_Y), .B0_t (data_out[40]), .Z0_t (data_out[44]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_12_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (data_out[41]), .B0_t (stateFF_inputPar[45]), .Z0_t (stateFF_state_gff_12_MUX_inst1_mux_inst_1_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_12_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (stateFF_state_gff_12_MUX_inst1_mux_inst_1_U1_X), .Z0_t (stateFF_state_gff_12_MUX_inst1_mux_inst_1_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_12_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_12_MUX_inst1_mux_inst_1_U1_Y), .B0_t (data_out[41]), .Z0_t (data_out[45]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_12_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (data_out[42]), .B0_t (stateFF_inputPar[46]), .Z0_t (stateFF_state_gff_12_MUX_inst1_mux_inst_2_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_12_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (stateFF_state_gff_12_MUX_inst1_mux_inst_2_U1_X), .Z0_t (stateFF_state_gff_12_MUX_inst1_mux_inst_2_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_12_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_12_MUX_inst1_mux_inst_2_U1_Y), .B0_t (data_out[42]), .Z0_t (data_out[46]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_12_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (data_out[43]), .B0_t (stateFF_inputPar[47]), .Z0_t (stateFF_state_gff_12_MUX_inst1_mux_inst_3_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_12_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (stateFF_state_gff_12_MUX_inst1_mux_inst_3_U1_X), .Z0_t (stateFF_state_gff_12_MUX_inst1_mux_inst_3_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_12_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_12_MUX_inst1_mux_inst_3_U1_Y), .B0_t (data_out[43]), .Z0_t (data_out[47]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_13_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (data_out[44]), .B0_t (stateFF_inputPar[48]), .Z0_t (stateFF_state_gff_13_MUX_inst1_mux_inst_0_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_13_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (stateFF_state_gff_13_MUX_inst1_mux_inst_0_U1_X), .Z0_t (stateFF_state_gff_13_MUX_inst1_mux_inst_0_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_13_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_13_MUX_inst1_mux_inst_0_U1_Y), .B0_t (data_out[44]), .Z0_t (data_out[48]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_13_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (data_out[45]), .B0_t (stateFF_inputPar[49]), .Z0_t (stateFF_state_gff_13_MUX_inst1_mux_inst_1_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_13_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (stateFF_state_gff_13_MUX_inst1_mux_inst_1_U1_X), .Z0_t (stateFF_state_gff_13_MUX_inst1_mux_inst_1_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_13_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_13_MUX_inst1_mux_inst_1_U1_Y), .B0_t (data_out[45]), .Z0_t (data_out[49]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_13_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (data_out[46]), .B0_t (stateFF_inputPar[50]), .Z0_t (stateFF_state_gff_13_MUX_inst1_mux_inst_2_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_13_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (stateFF_state_gff_13_MUX_inst1_mux_inst_2_U1_X), .Z0_t (stateFF_state_gff_13_MUX_inst1_mux_inst_2_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_13_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_13_MUX_inst1_mux_inst_2_U1_Y), .B0_t (data_out[46]), .Z0_t (data_out[50]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_13_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (data_out[47]), .B0_t (stateFF_inputPar[51]), .Z0_t (stateFF_state_gff_13_MUX_inst1_mux_inst_3_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_13_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (stateFF_state_gff_13_MUX_inst1_mux_inst_3_U1_X), .Z0_t (stateFF_state_gff_13_MUX_inst1_mux_inst_3_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_13_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_13_MUX_inst1_mux_inst_3_U1_Y), .B0_t (data_out[47]), .Z0_t (data_out[51]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_14_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (data_out[48]), .B0_t (stateFF_inputPar[52]), .Z0_t (stateFF_state_gff_14_MUX_inst1_mux_inst_0_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_14_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (stateFF_state_gff_14_MUX_inst1_mux_inst_0_U1_X), .Z0_t (stateFF_state_gff_14_MUX_inst1_mux_inst_0_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_14_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_14_MUX_inst1_mux_inst_0_U1_Y), .B0_t (data_out[48]), .Z0_t (data_out[52]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_14_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (data_out[49]), .B0_t (stateFF_inputPar[53]), .Z0_t (stateFF_state_gff_14_MUX_inst1_mux_inst_1_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_14_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (stateFF_state_gff_14_MUX_inst1_mux_inst_1_U1_X), .Z0_t (stateFF_state_gff_14_MUX_inst1_mux_inst_1_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_14_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_14_MUX_inst1_mux_inst_1_U1_Y), .B0_t (data_out[49]), .Z0_t (data_out[53]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_14_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (data_out[50]), .B0_t (stateFF_inputPar[54]), .Z0_t (stateFF_state_gff_14_MUX_inst1_mux_inst_2_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_14_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (stateFF_state_gff_14_MUX_inst1_mux_inst_2_U1_X), .Z0_t (stateFF_state_gff_14_MUX_inst1_mux_inst_2_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_14_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_14_MUX_inst1_mux_inst_2_U1_Y), .B0_t (data_out[50]), .Z0_t (data_out[54]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_14_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (data_out[51]), .B0_t (stateFF_inputPar[55]), .Z0_t (stateFF_state_gff_14_MUX_inst1_mux_inst_3_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_14_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (stateFF_state_gff_14_MUX_inst1_mux_inst_3_U1_X), .Z0_t (stateFF_state_gff_14_MUX_inst1_mux_inst_3_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_14_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_14_MUX_inst1_mux_inst_3_U1_Y), .B0_t (data_out[51]), .Z0_t (data_out[55]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_15_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (data_out[52]), .B0_t (stateFF_inputPar[56]), .Z0_t (stateFF_state_gff_15_MUX_inst1_mux_inst_0_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_15_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (stateFF_state_gff_15_MUX_inst1_mux_inst_0_U1_X), .Z0_t (stateFF_state_gff_15_MUX_inst1_mux_inst_0_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_15_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_15_MUX_inst1_mux_inst_0_U1_Y), .B0_t (data_out[52]), .Z0_t (data_out[56]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_15_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (data_out[53]), .B0_t (stateFF_inputPar[57]), .Z0_t (stateFF_state_gff_15_MUX_inst1_mux_inst_1_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_15_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (stateFF_state_gff_15_MUX_inst1_mux_inst_1_U1_X), .Z0_t (stateFF_state_gff_15_MUX_inst1_mux_inst_1_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_15_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_15_MUX_inst1_mux_inst_1_U1_Y), .B0_t (data_out[53]), .Z0_t (data_out[57]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_15_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (data_out[54]), .B0_t (stateFF_inputPar[58]), .Z0_t (stateFF_state_gff_15_MUX_inst1_mux_inst_2_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_15_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (stateFF_state_gff_15_MUX_inst1_mux_inst_2_U1_X), .Z0_t (stateFF_state_gff_15_MUX_inst1_mux_inst_2_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_15_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_15_MUX_inst1_mux_inst_2_U1_Y), .B0_t (data_out[54]), .Z0_t (data_out[58]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_15_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (data_out[55]), .B0_t (stateFF_inputPar[59]), .Z0_t (stateFF_state_gff_15_MUX_inst1_mux_inst_3_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_15_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (stateFF_state_gff_15_MUX_inst1_mux_inst_3_U1_X), .Z0_t (stateFF_state_gff_15_MUX_inst1_mux_inst_3_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_15_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_15_MUX_inst1_mux_inst_3_U1_Y), .B0_t (data_out[55]), .Z0_t (data_out[59]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_16_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (data_out[56]), .B0_t (stateFF_inputPar[60]), .Z0_t (stateFF_state_gff_16_MUX_inst1_mux_inst_0_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_16_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (stateFF_state_gff_16_MUX_inst1_mux_inst_0_U1_X), .Z0_t (stateFF_state_gff_16_MUX_inst1_mux_inst_0_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_16_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_16_MUX_inst1_mux_inst_0_U1_Y), .B0_t (data_out[56]), .Z0_t (data_out[60]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_16_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (data_out[57]), .B0_t (stateFF_inputPar[61]), .Z0_t (stateFF_state_gff_16_MUX_inst1_mux_inst_1_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_16_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (stateFF_state_gff_16_MUX_inst1_mux_inst_1_U1_X), .Z0_t (stateFF_state_gff_16_MUX_inst1_mux_inst_1_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_16_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_16_MUX_inst1_mux_inst_1_U1_Y), .B0_t (data_out[57]), .Z0_t (data_out[61]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_16_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (data_out[58]), .B0_t (stateFF_inputPar[62]), .Z0_t (stateFF_state_gff_16_MUX_inst1_mux_inst_2_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_16_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (stateFF_state_gff_16_MUX_inst1_mux_inst_2_U1_X), .Z0_t (stateFF_state_gff_16_MUX_inst1_mux_inst_2_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_16_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_16_MUX_inst1_mux_inst_2_U1_Y), .B0_t (data_out[58]), .Z0_t (data_out[62]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_16_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (data_out[59]), .B0_t (stateFF_inputPar[63]), .Z0_t (stateFF_state_gff_16_MUX_inst1_mux_inst_3_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_16_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (stateFF_state_gff_16_MUX_inst1_mux_inst_3_U1_X), .Z0_t (stateFF_state_gff_16_MUX_inst1_mux_inst_3_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_16_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_16_MUX_inst1_mux_inst_3_U1_Y), .B0_t (data_out[59]), .Z0_t (data_out[63]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_0_U1_XOR1_U1 ( .A0_t (data_out[0]), .B0_t (data_in[0]), .Z0_t (stateFF_MUX_inputPar_mux_inst_0_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_0_U1_AND1_U1 ( .A0_t (reset), .B0_t (stateFF_MUX_inputPar_mux_inst_0_U1_X), .Z0_t (stateFF_MUX_inputPar_mux_inst_0_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_0_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_0_U1_Y), .B0_t (data_out[0]), .Z0_t (stateFF_inputPar[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_1_U1_XOR1_U1 ( .A0_t (data_out[4]), .B0_t (data_in[1]), .Z0_t (stateFF_MUX_inputPar_mux_inst_1_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_1_U1_AND1_U1 ( .A0_t (reset), .B0_t (stateFF_MUX_inputPar_mux_inst_1_U1_X), .Z0_t (stateFF_MUX_inputPar_mux_inst_1_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_1_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_1_U1_Y), .B0_t (data_out[4]), .Z0_t (stateFF_inputPar[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_2_U1_XOR1_U1 ( .A0_t (data_out[8]), .B0_t (data_in[2]), .Z0_t (stateFF_MUX_inputPar_mux_inst_2_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_2_U1_AND1_U1 ( .A0_t (reset), .B0_t (stateFF_MUX_inputPar_mux_inst_2_U1_X), .Z0_t (stateFF_MUX_inputPar_mux_inst_2_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_2_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_2_U1_Y), .B0_t (data_out[8]), .Z0_t (stateFF_inputPar[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_3_U1_XOR1_U1 ( .A0_t (data_out[12]), .B0_t (data_in[3]), .Z0_t (stateFF_MUX_inputPar_mux_inst_3_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_3_U1_AND1_U1 ( .A0_t (reset), .B0_t (stateFF_MUX_inputPar_mux_inst_3_U1_X), .Z0_t (stateFF_MUX_inputPar_mux_inst_3_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_3_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_3_U1_Y), .B0_t (data_out[12]), .Z0_t (stateFF_inputPar[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_4_U1_XOR1_U1 ( .A0_t (data_out[16]), .B0_t (data_in[4]), .Z0_t (stateFF_MUX_inputPar_mux_inst_4_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_4_U1_AND1_U1 ( .A0_t (reset), .B0_t (stateFF_MUX_inputPar_mux_inst_4_U1_X), .Z0_t (stateFF_MUX_inputPar_mux_inst_4_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_4_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_4_U1_Y), .B0_t (data_out[16]), .Z0_t (stateFF_inputPar[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_5_U1_XOR1_U1 ( .A0_t (data_out[20]), .B0_t (data_in[5]), .Z0_t (stateFF_MUX_inputPar_mux_inst_5_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_5_U1_AND1_U1 ( .A0_t (reset), .B0_t (stateFF_MUX_inputPar_mux_inst_5_U1_X), .Z0_t (stateFF_MUX_inputPar_mux_inst_5_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_5_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_5_U1_Y), .B0_t (data_out[20]), .Z0_t (stateFF_inputPar[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_6_U1_XOR1_U1 ( .A0_t (data_out[24]), .B0_t (data_in[6]), .Z0_t (stateFF_MUX_inputPar_mux_inst_6_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_6_U1_AND1_U1 ( .A0_t (reset), .B0_t (stateFF_MUX_inputPar_mux_inst_6_U1_X), .Z0_t (stateFF_MUX_inputPar_mux_inst_6_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_6_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_6_U1_Y), .B0_t (data_out[24]), .Z0_t (stateFF_inputPar[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_7_U1_XOR1_U1 ( .A0_t (data_out[28]), .B0_t (data_in[7]), .Z0_t (stateFF_MUX_inputPar_mux_inst_7_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_7_U1_AND1_U1 ( .A0_t (reset), .B0_t (stateFF_MUX_inputPar_mux_inst_7_U1_X), .Z0_t (stateFF_MUX_inputPar_mux_inst_7_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_7_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_7_U1_Y), .B0_t (data_out[28]), .Z0_t (stateFF_inputPar[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_8_U1_XOR1_U1 ( .A0_t (data_out[32]), .B0_t (data_in[8]), .Z0_t (stateFF_MUX_inputPar_mux_inst_8_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_8_U1_AND1_U1 ( .A0_t (reset), .B0_t (stateFF_MUX_inputPar_mux_inst_8_U1_X), .Z0_t (stateFF_MUX_inputPar_mux_inst_8_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_8_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_8_U1_Y), .B0_t (data_out[32]), .Z0_t (stateFF_inputPar[8]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_9_U1_XOR1_U1 ( .A0_t (data_out[36]), .B0_t (data_in[9]), .Z0_t (stateFF_MUX_inputPar_mux_inst_9_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_9_U1_AND1_U1 ( .A0_t (reset), .B0_t (stateFF_MUX_inputPar_mux_inst_9_U1_X), .Z0_t (stateFF_MUX_inputPar_mux_inst_9_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_9_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_9_U1_Y), .B0_t (data_out[36]), .Z0_t (stateFF_inputPar[9]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_10_U1_XOR1_U1 ( .A0_t (data_out[40]), .B0_t (data_in[10]), .Z0_t (stateFF_MUX_inputPar_mux_inst_10_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_10_U1_AND1_U1 ( .A0_t (reset), .B0_t (stateFF_MUX_inputPar_mux_inst_10_U1_X), .Z0_t (stateFF_MUX_inputPar_mux_inst_10_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_10_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_10_U1_Y), .B0_t (data_out[40]), .Z0_t (stateFF_inputPar[10]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_11_U1_XOR1_U1 ( .A0_t (data_out[44]), .B0_t (data_in[11]), .Z0_t (stateFF_MUX_inputPar_mux_inst_11_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_11_U1_AND1_U1 ( .A0_t (reset), .B0_t (stateFF_MUX_inputPar_mux_inst_11_U1_X), .Z0_t (stateFF_MUX_inputPar_mux_inst_11_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_11_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_11_U1_Y), .B0_t (data_out[44]), .Z0_t (stateFF_inputPar[11]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_12_U1_XOR1_U1 ( .A0_t (data_out[48]), .B0_t (data_in[12]), .Z0_t (stateFF_MUX_inputPar_mux_inst_12_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_12_U1_AND1_U1 ( .A0_t (reset), .B0_t (stateFF_MUX_inputPar_mux_inst_12_U1_X), .Z0_t (stateFF_MUX_inputPar_mux_inst_12_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_12_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_12_U1_Y), .B0_t (data_out[48]), .Z0_t (stateFF_inputPar[12]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_13_U1_XOR1_U1 ( .A0_t (data_out[52]), .B0_t (data_in[13]), .Z0_t (stateFF_MUX_inputPar_mux_inst_13_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_13_U1_AND1_U1 ( .A0_t (reset), .B0_t (stateFF_MUX_inputPar_mux_inst_13_U1_X), .Z0_t (stateFF_MUX_inputPar_mux_inst_13_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_13_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_13_U1_Y), .B0_t (data_out[52]), .Z0_t (stateFF_inputPar[13]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_14_U1_XOR1_U1 ( .A0_t (data_out[56]), .B0_t (data_in[14]), .Z0_t (stateFF_MUX_inputPar_mux_inst_14_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_14_U1_AND1_U1 ( .A0_t (reset), .B0_t (stateFF_MUX_inputPar_mux_inst_14_U1_X), .Z0_t (stateFF_MUX_inputPar_mux_inst_14_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_14_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_14_U1_Y), .B0_t (data_out[56]), .Z0_t (stateFF_inputPar[14]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_15_U1_XOR1_U1 ( .A0_t (data_out[60]), .B0_t (data_in[15]), .Z0_t (stateFF_MUX_inputPar_mux_inst_15_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_15_U1_AND1_U1 ( .A0_t (reset), .B0_t (stateFF_MUX_inputPar_mux_inst_15_U1_X), .Z0_t (stateFF_MUX_inputPar_mux_inst_15_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_15_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_15_U1_Y), .B0_t (data_out[60]), .Z0_t (stateFF_inputPar[15]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_16_U1_XOR1_U1 ( .A0_t (data_out[1]), .B0_t (data_in[16]), .Z0_t (stateFF_MUX_inputPar_mux_inst_16_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_16_U1_AND1_U1 ( .A0_t (reset), .B0_t (stateFF_MUX_inputPar_mux_inst_16_U1_X), .Z0_t (stateFF_MUX_inputPar_mux_inst_16_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_16_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_16_U1_Y), .B0_t (data_out[1]), .Z0_t (stateFF_inputPar[16]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_17_U1_XOR1_U1 ( .A0_t (data_out[5]), .B0_t (data_in[17]), .Z0_t (stateFF_MUX_inputPar_mux_inst_17_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_17_U1_AND1_U1 ( .A0_t (reset), .B0_t (stateFF_MUX_inputPar_mux_inst_17_U1_X), .Z0_t (stateFF_MUX_inputPar_mux_inst_17_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_17_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_17_U1_Y), .B0_t (data_out[5]), .Z0_t (stateFF_inputPar[17]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_18_U1_XOR1_U1 ( .A0_t (data_out[9]), .B0_t (data_in[18]), .Z0_t (stateFF_MUX_inputPar_mux_inst_18_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_18_U1_AND1_U1 ( .A0_t (reset), .B0_t (stateFF_MUX_inputPar_mux_inst_18_U1_X), .Z0_t (stateFF_MUX_inputPar_mux_inst_18_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_18_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_18_U1_Y), .B0_t (data_out[9]), .Z0_t (stateFF_inputPar[18]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_19_U1_XOR1_U1 ( .A0_t (data_out[13]), .B0_t (data_in[19]), .Z0_t (stateFF_MUX_inputPar_mux_inst_19_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_19_U1_AND1_U1 ( .A0_t (reset), .B0_t (stateFF_MUX_inputPar_mux_inst_19_U1_X), .Z0_t (stateFF_MUX_inputPar_mux_inst_19_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_19_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_19_U1_Y), .B0_t (data_out[13]), .Z0_t (stateFF_inputPar[19]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_20_U1_XOR1_U1 ( .A0_t (data_out[17]), .B0_t (data_in[20]), .Z0_t (stateFF_MUX_inputPar_mux_inst_20_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_20_U1_AND1_U1 ( .A0_t (reset), .B0_t (stateFF_MUX_inputPar_mux_inst_20_U1_X), .Z0_t (stateFF_MUX_inputPar_mux_inst_20_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_20_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_20_U1_Y), .B0_t (data_out[17]), .Z0_t (stateFF_inputPar[20]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_21_U1_XOR1_U1 ( .A0_t (data_out[21]), .B0_t (data_in[21]), .Z0_t (stateFF_MUX_inputPar_mux_inst_21_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_21_U1_AND1_U1 ( .A0_t (reset), .B0_t (stateFF_MUX_inputPar_mux_inst_21_U1_X), .Z0_t (stateFF_MUX_inputPar_mux_inst_21_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_21_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_21_U1_Y), .B0_t (data_out[21]), .Z0_t (stateFF_inputPar[21]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_22_U1_XOR1_U1 ( .A0_t (data_out[25]), .B0_t (data_in[22]), .Z0_t (stateFF_MUX_inputPar_mux_inst_22_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_22_U1_AND1_U1 ( .A0_t (reset), .B0_t (stateFF_MUX_inputPar_mux_inst_22_U1_X), .Z0_t (stateFF_MUX_inputPar_mux_inst_22_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_22_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_22_U1_Y), .B0_t (data_out[25]), .Z0_t (stateFF_inputPar[22]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_23_U1_XOR1_U1 ( .A0_t (data_out[29]), .B0_t (data_in[23]), .Z0_t (stateFF_MUX_inputPar_mux_inst_23_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_23_U1_AND1_U1 ( .A0_t (reset), .B0_t (stateFF_MUX_inputPar_mux_inst_23_U1_X), .Z0_t (stateFF_MUX_inputPar_mux_inst_23_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_23_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_23_U1_Y), .B0_t (data_out[29]), .Z0_t (stateFF_inputPar[23]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_24_U1_XOR1_U1 ( .A0_t (data_out[33]), .B0_t (data_in[24]), .Z0_t (stateFF_MUX_inputPar_mux_inst_24_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_24_U1_AND1_U1 ( .A0_t (reset), .B0_t (stateFF_MUX_inputPar_mux_inst_24_U1_X), .Z0_t (stateFF_MUX_inputPar_mux_inst_24_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_24_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_24_U1_Y), .B0_t (data_out[33]), .Z0_t (stateFF_inputPar[24]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_25_U1_XOR1_U1 ( .A0_t (data_out[37]), .B0_t (data_in[25]), .Z0_t (stateFF_MUX_inputPar_mux_inst_25_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_25_U1_AND1_U1 ( .A0_t (reset), .B0_t (stateFF_MUX_inputPar_mux_inst_25_U1_X), .Z0_t (stateFF_MUX_inputPar_mux_inst_25_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_25_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_25_U1_Y), .B0_t (data_out[37]), .Z0_t (stateFF_inputPar[25]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_26_U1_XOR1_U1 ( .A0_t (data_out[41]), .B0_t (data_in[26]), .Z0_t (stateFF_MUX_inputPar_mux_inst_26_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_26_U1_AND1_U1 ( .A0_t (reset), .B0_t (stateFF_MUX_inputPar_mux_inst_26_U1_X), .Z0_t (stateFF_MUX_inputPar_mux_inst_26_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_26_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_26_U1_Y), .B0_t (data_out[41]), .Z0_t (stateFF_inputPar[26]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_27_U1_XOR1_U1 ( .A0_t (data_out[45]), .B0_t (data_in[27]), .Z0_t (stateFF_MUX_inputPar_mux_inst_27_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_27_U1_AND1_U1 ( .A0_t (reset), .B0_t (stateFF_MUX_inputPar_mux_inst_27_U1_X), .Z0_t (stateFF_MUX_inputPar_mux_inst_27_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_27_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_27_U1_Y), .B0_t (data_out[45]), .Z0_t (stateFF_inputPar[27]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_28_U1_XOR1_U1 ( .A0_t (data_out[49]), .B0_t (data_in[28]), .Z0_t (stateFF_MUX_inputPar_mux_inst_28_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_28_U1_AND1_U1 ( .A0_t (reset), .B0_t (stateFF_MUX_inputPar_mux_inst_28_U1_X), .Z0_t (stateFF_MUX_inputPar_mux_inst_28_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_28_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_28_U1_Y), .B0_t (data_out[49]), .Z0_t (stateFF_inputPar[28]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_29_U1_XOR1_U1 ( .A0_t (data_out[53]), .B0_t (data_in[29]), .Z0_t (stateFF_MUX_inputPar_mux_inst_29_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_29_U1_AND1_U1 ( .A0_t (reset), .B0_t (stateFF_MUX_inputPar_mux_inst_29_U1_X), .Z0_t (stateFF_MUX_inputPar_mux_inst_29_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_29_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_29_U1_Y), .B0_t (data_out[53]), .Z0_t (stateFF_inputPar[29]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_30_U1_XOR1_U1 ( .A0_t (data_out[57]), .B0_t (data_in[30]), .Z0_t (stateFF_MUX_inputPar_mux_inst_30_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_30_U1_AND1_U1 ( .A0_t (reset), .B0_t (stateFF_MUX_inputPar_mux_inst_30_U1_X), .Z0_t (stateFF_MUX_inputPar_mux_inst_30_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_30_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_30_U1_Y), .B0_t (data_out[57]), .Z0_t (stateFF_inputPar[30]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_31_U1_XOR1_U1 ( .A0_t (data_out[61]), .B0_t (data_in[31]), .Z0_t (stateFF_MUX_inputPar_mux_inst_31_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_31_U1_AND1_U1 ( .A0_t (reset), .B0_t (stateFF_MUX_inputPar_mux_inst_31_U1_X), .Z0_t (stateFF_MUX_inputPar_mux_inst_31_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_31_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_31_U1_Y), .B0_t (data_out[61]), .Z0_t (stateFF_inputPar[31]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_32_U1_XOR1_U1 ( .A0_t (data_out[2]), .B0_t (data_in[32]), .Z0_t (stateFF_MUX_inputPar_mux_inst_32_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_32_U1_AND1_U1 ( .A0_t (reset), .B0_t (stateFF_MUX_inputPar_mux_inst_32_U1_X), .Z0_t (stateFF_MUX_inputPar_mux_inst_32_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_32_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_32_U1_Y), .B0_t (data_out[2]), .Z0_t (stateFF_inputPar[32]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_33_U1_XOR1_U1 ( .A0_t (data_out[6]), .B0_t (data_in[33]), .Z0_t (stateFF_MUX_inputPar_mux_inst_33_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_33_U1_AND1_U1 ( .A0_t (reset), .B0_t (stateFF_MUX_inputPar_mux_inst_33_U1_X), .Z0_t (stateFF_MUX_inputPar_mux_inst_33_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_33_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_33_U1_Y), .B0_t (data_out[6]), .Z0_t (stateFF_inputPar[33]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_34_U1_XOR1_U1 ( .A0_t (data_out[10]), .B0_t (data_in[34]), .Z0_t (stateFF_MUX_inputPar_mux_inst_34_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_34_U1_AND1_U1 ( .A0_t (reset), .B0_t (stateFF_MUX_inputPar_mux_inst_34_U1_X), .Z0_t (stateFF_MUX_inputPar_mux_inst_34_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_34_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_34_U1_Y), .B0_t (data_out[10]), .Z0_t (stateFF_inputPar[34]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_35_U1_XOR1_U1 ( .A0_t (data_out[14]), .B0_t (data_in[35]), .Z0_t (stateFF_MUX_inputPar_mux_inst_35_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_35_U1_AND1_U1 ( .A0_t (reset), .B0_t (stateFF_MUX_inputPar_mux_inst_35_U1_X), .Z0_t (stateFF_MUX_inputPar_mux_inst_35_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_35_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_35_U1_Y), .B0_t (data_out[14]), .Z0_t (stateFF_inputPar[35]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_36_U1_XOR1_U1 ( .A0_t (data_out[18]), .B0_t (data_in[36]), .Z0_t (stateFF_MUX_inputPar_mux_inst_36_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_36_U1_AND1_U1 ( .A0_t (reset), .B0_t (stateFF_MUX_inputPar_mux_inst_36_U1_X), .Z0_t (stateFF_MUX_inputPar_mux_inst_36_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_36_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_36_U1_Y), .B0_t (data_out[18]), .Z0_t (stateFF_inputPar[36]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_37_U1_XOR1_U1 ( .A0_t (data_out[22]), .B0_t (data_in[37]), .Z0_t (stateFF_MUX_inputPar_mux_inst_37_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_37_U1_AND1_U1 ( .A0_t (reset), .B0_t (stateFF_MUX_inputPar_mux_inst_37_U1_X), .Z0_t (stateFF_MUX_inputPar_mux_inst_37_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_37_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_37_U1_Y), .B0_t (data_out[22]), .Z0_t (stateFF_inputPar[37]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_38_U1_XOR1_U1 ( .A0_t (data_out[26]), .B0_t (data_in[38]), .Z0_t (stateFF_MUX_inputPar_mux_inst_38_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_38_U1_AND1_U1 ( .A0_t (reset), .B0_t (stateFF_MUX_inputPar_mux_inst_38_U1_X), .Z0_t (stateFF_MUX_inputPar_mux_inst_38_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_38_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_38_U1_Y), .B0_t (data_out[26]), .Z0_t (stateFF_inputPar[38]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_39_U1_XOR1_U1 ( .A0_t (data_out[30]), .B0_t (data_in[39]), .Z0_t (stateFF_MUX_inputPar_mux_inst_39_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_39_U1_AND1_U1 ( .A0_t (reset), .B0_t (stateFF_MUX_inputPar_mux_inst_39_U1_X), .Z0_t (stateFF_MUX_inputPar_mux_inst_39_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_39_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_39_U1_Y), .B0_t (data_out[30]), .Z0_t (stateFF_inputPar[39]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_40_U1_XOR1_U1 ( .A0_t (data_out[34]), .B0_t (data_in[40]), .Z0_t (stateFF_MUX_inputPar_mux_inst_40_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_40_U1_AND1_U1 ( .A0_t (reset), .B0_t (stateFF_MUX_inputPar_mux_inst_40_U1_X), .Z0_t (stateFF_MUX_inputPar_mux_inst_40_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_40_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_40_U1_Y), .B0_t (data_out[34]), .Z0_t (stateFF_inputPar[40]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_41_U1_XOR1_U1 ( .A0_t (data_out[38]), .B0_t (data_in[41]), .Z0_t (stateFF_MUX_inputPar_mux_inst_41_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_41_U1_AND1_U1 ( .A0_t (reset), .B0_t (stateFF_MUX_inputPar_mux_inst_41_U1_X), .Z0_t (stateFF_MUX_inputPar_mux_inst_41_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_41_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_41_U1_Y), .B0_t (data_out[38]), .Z0_t (stateFF_inputPar[41]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_42_U1_XOR1_U1 ( .A0_t (data_out[42]), .B0_t (data_in[42]), .Z0_t (stateFF_MUX_inputPar_mux_inst_42_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_42_U1_AND1_U1 ( .A0_t (reset), .B0_t (stateFF_MUX_inputPar_mux_inst_42_U1_X), .Z0_t (stateFF_MUX_inputPar_mux_inst_42_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_42_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_42_U1_Y), .B0_t (data_out[42]), .Z0_t (stateFF_inputPar[42]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_43_U1_XOR1_U1 ( .A0_t (data_out[46]), .B0_t (data_in[43]), .Z0_t (stateFF_MUX_inputPar_mux_inst_43_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_43_U1_AND1_U1 ( .A0_t (reset), .B0_t (stateFF_MUX_inputPar_mux_inst_43_U1_X), .Z0_t (stateFF_MUX_inputPar_mux_inst_43_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_43_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_43_U1_Y), .B0_t (data_out[46]), .Z0_t (stateFF_inputPar[43]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_44_U1_XOR1_U1 ( .A0_t (data_out[50]), .B0_t (data_in[44]), .Z0_t (stateFF_MUX_inputPar_mux_inst_44_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_44_U1_AND1_U1 ( .A0_t (reset), .B0_t (stateFF_MUX_inputPar_mux_inst_44_U1_X), .Z0_t (stateFF_MUX_inputPar_mux_inst_44_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_44_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_44_U1_Y), .B0_t (data_out[50]), .Z0_t (stateFF_inputPar[44]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_45_U1_XOR1_U1 ( .A0_t (data_out[54]), .B0_t (data_in[45]), .Z0_t (stateFF_MUX_inputPar_mux_inst_45_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_45_U1_AND1_U1 ( .A0_t (reset), .B0_t (stateFF_MUX_inputPar_mux_inst_45_U1_X), .Z0_t (stateFF_MUX_inputPar_mux_inst_45_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_45_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_45_U1_Y), .B0_t (data_out[54]), .Z0_t (stateFF_inputPar[45]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_46_U1_XOR1_U1 ( .A0_t (data_out[58]), .B0_t (data_in[46]), .Z0_t (stateFF_MUX_inputPar_mux_inst_46_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_46_U1_AND1_U1 ( .A0_t (reset), .B0_t (stateFF_MUX_inputPar_mux_inst_46_U1_X), .Z0_t (stateFF_MUX_inputPar_mux_inst_46_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_46_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_46_U1_Y), .B0_t (data_out[58]), .Z0_t (stateFF_inputPar[46]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_47_U1_XOR1_U1 ( .A0_t (data_out[62]), .B0_t (data_in[47]), .Z0_t (stateFF_MUX_inputPar_mux_inst_47_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_47_U1_AND1_U1 ( .A0_t (reset), .B0_t (stateFF_MUX_inputPar_mux_inst_47_U1_X), .Z0_t (stateFF_MUX_inputPar_mux_inst_47_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_47_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_47_U1_Y), .B0_t (data_out[62]), .Z0_t (stateFF_inputPar[47]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_48_U1_XOR1_U1 ( .A0_t (data_out[3]), .B0_t (data_in[48]), .Z0_t (stateFF_MUX_inputPar_mux_inst_48_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_48_U1_AND1_U1 ( .A0_t (reset), .B0_t (stateFF_MUX_inputPar_mux_inst_48_U1_X), .Z0_t (stateFF_MUX_inputPar_mux_inst_48_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_48_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_48_U1_Y), .B0_t (data_out[3]), .Z0_t (stateFF_inputPar[48]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_49_U1_XOR1_U1 ( .A0_t (data_out[7]), .B0_t (data_in[49]), .Z0_t (stateFF_MUX_inputPar_mux_inst_49_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_49_U1_AND1_U1 ( .A0_t (reset), .B0_t (stateFF_MUX_inputPar_mux_inst_49_U1_X), .Z0_t (stateFF_MUX_inputPar_mux_inst_49_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_49_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_49_U1_Y), .B0_t (data_out[7]), .Z0_t (stateFF_inputPar[49]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_50_U1_XOR1_U1 ( .A0_t (data_out[11]), .B0_t (data_in[50]), .Z0_t (stateFF_MUX_inputPar_mux_inst_50_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_50_U1_AND1_U1 ( .A0_t (reset), .B0_t (stateFF_MUX_inputPar_mux_inst_50_U1_X), .Z0_t (stateFF_MUX_inputPar_mux_inst_50_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_50_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_50_U1_Y), .B0_t (data_out[11]), .Z0_t (stateFF_inputPar[50]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_51_U1_XOR1_U1 ( .A0_t (data_out[15]), .B0_t (data_in[51]), .Z0_t (stateFF_MUX_inputPar_mux_inst_51_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_51_U1_AND1_U1 ( .A0_t (reset), .B0_t (stateFF_MUX_inputPar_mux_inst_51_U1_X), .Z0_t (stateFF_MUX_inputPar_mux_inst_51_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_51_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_51_U1_Y), .B0_t (data_out[15]), .Z0_t (stateFF_inputPar[51]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_52_U1_XOR1_U1 ( .A0_t (data_out[19]), .B0_t (data_in[52]), .Z0_t (stateFF_MUX_inputPar_mux_inst_52_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_52_U1_AND1_U1 ( .A0_t (reset), .B0_t (stateFF_MUX_inputPar_mux_inst_52_U1_X), .Z0_t (stateFF_MUX_inputPar_mux_inst_52_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_52_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_52_U1_Y), .B0_t (data_out[19]), .Z0_t (stateFF_inputPar[52]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_53_U1_XOR1_U1 ( .A0_t (data_out[23]), .B0_t (data_in[53]), .Z0_t (stateFF_MUX_inputPar_mux_inst_53_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_53_U1_AND1_U1 ( .A0_t (reset), .B0_t (stateFF_MUX_inputPar_mux_inst_53_U1_X), .Z0_t (stateFF_MUX_inputPar_mux_inst_53_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_53_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_53_U1_Y), .B0_t (data_out[23]), .Z0_t (stateFF_inputPar[53]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_54_U1_XOR1_U1 ( .A0_t (data_out[27]), .B0_t (data_in[54]), .Z0_t (stateFF_MUX_inputPar_mux_inst_54_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_54_U1_AND1_U1 ( .A0_t (reset), .B0_t (stateFF_MUX_inputPar_mux_inst_54_U1_X), .Z0_t (stateFF_MUX_inputPar_mux_inst_54_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_54_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_54_U1_Y), .B0_t (data_out[27]), .Z0_t (stateFF_inputPar[54]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_55_U1_XOR1_U1 ( .A0_t (data_out[31]), .B0_t (data_in[55]), .Z0_t (stateFF_MUX_inputPar_mux_inst_55_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_55_U1_AND1_U1 ( .A0_t (reset), .B0_t (stateFF_MUX_inputPar_mux_inst_55_U1_X), .Z0_t (stateFF_MUX_inputPar_mux_inst_55_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_55_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_55_U1_Y), .B0_t (data_out[31]), .Z0_t (stateFF_inputPar[55]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_56_U1_XOR1_U1 ( .A0_t (data_out[35]), .B0_t (data_in[56]), .Z0_t (stateFF_MUX_inputPar_mux_inst_56_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_56_U1_AND1_U1 ( .A0_t (reset), .B0_t (stateFF_MUX_inputPar_mux_inst_56_U1_X), .Z0_t (stateFF_MUX_inputPar_mux_inst_56_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_56_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_56_U1_Y), .B0_t (data_out[35]), .Z0_t (stateFF_inputPar[56]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_57_U1_XOR1_U1 ( .A0_t (data_out[39]), .B0_t (data_in[57]), .Z0_t (stateFF_MUX_inputPar_mux_inst_57_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_57_U1_AND1_U1 ( .A0_t (reset), .B0_t (stateFF_MUX_inputPar_mux_inst_57_U1_X), .Z0_t (stateFF_MUX_inputPar_mux_inst_57_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_57_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_57_U1_Y), .B0_t (data_out[39]), .Z0_t (stateFF_inputPar[57]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_58_U1_XOR1_U1 ( .A0_t (data_out[43]), .B0_t (data_in[58]), .Z0_t (stateFF_MUX_inputPar_mux_inst_58_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_58_U1_AND1_U1 ( .A0_t (reset), .B0_t (stateFF_MUX_inputPar_mux_inst_58_U1_X), .Z0_t (stateFF_MUX_inputPar_mux_inst_58_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_58_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_58_U1_Y), .B0_t (data_out[43]), .Z0_t (stateFF_inputPar[58]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_59_U1_XOR1_U1 ( .A0_t (data_out[47]), .B0_t (data_in[59]), .Z0_t (stateFF_MUX_inputPar_mux_inst_59_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_59_U1_AND1_U1 ( .A0_t (reset), .B0_t (stateFF_MUX_inputPar_mux_inst_59_U1_X), .Z0_t (stateFF_MUX_inputPar_mux_inst_59_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_59_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_59_U1_Y), .B0_t (data_out[47]), .Z0_t (stateFF_inputPar[59]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_60_U1_XOR1_U1 ( .A0_t (data_out[51]), .B0_t (data_in[60]), .Z0_t (stateFF_MUX_inputPar_mux_inst_60_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_60_U1_AND1_U1 ( .A0_t (reset), .B0_t (stateFF_MUX_inputPar_mux_inst_60_U1_X), .Z0_t (stateFF_MUX_inputPar_mux_inst_60_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_60_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_60_U1_Y), .B0_t (data_out[51]), .Z0_t (stateFF_inputPar[60]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_61_U1_XOR1_U1 ( .A0_t (data_out[55]), .B0_t (data_in[61]), .Z0_t (stateFF_MUX_inputPar_mux_inst_61_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_61_U1_AND1_U1 ( .A0_t (reset), .B0_t (stateFF_MUX_inputPar_mux_inst_61_U1_X), .Z0_t (stateFF_MUX_inputPar_mux_inst_61_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_61_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_61_U1_Y), .B0_t (data_out[55]), .Z0_t (stateFF_inputPar[61]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_62_U1_XOR1_U1 ( .A0_t (data_out[59]), .B0_t (data_in[62]), .Z0_t (stateFF_MUX_inputPar_mux_inst_62_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_62_U1_AND1_U1 ( .A0_t (reset), .B0_t (stateFF_MUX_inputPar_mux_inst_62_U1_X), .Z0_t (stateFF_MUX_inputPar_mux_inst_62_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_62_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_62_U1_Y), .B0_t (data_out[59]), .Z0_t (stateFF_inputPar[62]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_63_U1_XOR1_U1 ( .A0_t (data_out[63]), .B0_t (data_in[63]), .Z0_t (stateFF_MUX_inputPar_mux_inst_63_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_63_U1_AND1_U1 ( .A0_t (reset), .B0_t (stateFF_MUX_inputPar_mux_inst_63_U1_X), .Z0_t (stateFF_MUX_inputPar_mux_inst_63_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_63_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_63_U1_Y), .B0_t (data_out[63]), .Z0_t (stateFF_inputPar[63]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_U5 ( .A0_t (counter[3]), .B0_t (keyFF_outputPar[21]), .Z0_t (keyFF_counterAdd[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_U4 ( .A0_t (counter[1]), .B0_t (keyFF_outputPar[19]), .Z0_t (keyFF_counterAdd[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_U3 ( .A0_t (counter[4]), .B0_t (keyFF_outputPar[22]), .Z0_t (keyFF_counterAdd[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_U2 ( .A0_t (counter[0]), .B0_t (keyFF_outputPar[18]), .Z0_t (keyFF_counterAdd[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_U1 ( .A0_t (counter[2]), .B0_t (keyFF_outputPar[20]), .Z0_t (keyFF_counterAdd[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_1_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (roundkey[0]), .B0_t (keyFF_inputPar[0]), .Z0_t (keyFF_keystate_gff_1_MUX_inst1_mux_inst_0_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_1_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_1_MUX_inst1_mux_inst_0_U1_X), .Z0_t (keyFF_keystate_gff_1_MUX_inst1_mux_inst_0_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_1_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_1_MUX_inst1_mux_inst_0_U1_Y), .B0_t (roundkey[0]), .Z0_t (keyRegKS[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_1_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (roundkey[1]), .B0_t (keyFF_inputPar[1]), .Z0_t (keyFF_keystate_gff_1_MUX_inst1_mux_inst_1_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_1_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_1_MUX_inst1_mux_inst_1_U1_X), .Z0_t (keyFF_keystate_gff_1_MUX_inst1_mux_inst_1_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_1_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_1_MUX_inst1_mux_inst_1_U1_Y), .B0_t (roundkey[1]), .Z0_t (keyRegKS[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_1_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (roundkey[2]), .B0_t (keyFF_inputPar[2]), .Z0_t (keyFF_keystate_gff_1_MUX_inst1_mux_inst_2_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_1_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_1_MUX_inst1_mux_inst_2_U1_X), .Z0_t (keyFF_keystate_gff_1_MUX_inst1_mux_inst_2_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_1_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_1_MUX_inst1_mux_inst_2_U1_Y), .B0_t (roundkey[2]), .Z0_t (keyRegKS[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_1_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (roundkey[3]), .B0_t (keyFF_inputPar[3]), .Z0_t (keyFF_keystate_gff_1_MUX_inst1_mux_inst_3_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_1_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_1_MUX_inst1_mux_inst_3_U1_X), .Z0_t (keyFF_keystate_gff_1_MUX_inst1_mux_inst_3_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_1_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_1_MUX_inst1_mux_inst_3_U1_Y), .B0_t (roundkey[3]), .Z0_t (keyFF_outputPar[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_2_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (keyRegKS[1]), .B0_t (keyFF_inputPar[4]), .Z0_t (keyFF_keystate_gff_2_MUX_inst1_mux_inst_0_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_2_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_2_MUX_inst1_mux_inst_0_U1_X), .Z0_t (keyFF_keystate_gff_2_MUX_inst1_mux_inst_0_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_2_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_2_MUX_inst1_mux_inst_0_U1_Y), .B0_t (keyRegKS[1]), .Z0_t (keyFF_outputPar[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_2_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (keyRegKS[2]), .B0_t (keyFF_inputPar[5]), .Z0_t (keyFF_keystate_gff_2_MUX_inst1_mux_inst_1_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_2_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_2_MUX_inst1_mux_inst_1_U1_X), .Z0_t (keyFF_keystate_gff_2_MUX_inst1_mux_inst_1_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_2_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_2_MUX_inst1_mux_inst_1_U1_Y), .B0_t (keyRegKS[2]), .Z0_t (keyFF_outputPar[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_2_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (keyRegKS[3]), .B0_t (keyFF_inputPar[6]), .Z0_t (keyFF_keystate_gff_2_MUX_inst1_mux_inst_2_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_2_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_2_MUX_inst1_mux_inst_2_U1_X), .Z0_t (keyFF_keystate_gff_2_MUX_inst1_mux_inst_2_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_2_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_2_MUX_inst1_mux_inst_2_U1_Y), .B0_t (keyRegKS[3]), .Z0_t (keyFF_outputPar[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_2_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[3]), .B0_t (keyFF_inputPar[7]), .Z0_t (keyFF_keystate_gff_2_MUX_inst1_mux_inst_3_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_2_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_2_MUX_inst1_mux_inst_3_U1_X), .Z0_t (keyFF_keystate_gff_2_MUX_inst1_mux_inst_3_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_2_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_2_MUX_inst1_mux_inst_3_U1_Y), .B0_t (keyFF_outputPar[3]), .Z0_t (keyFF_outputPar[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_3_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[4]), .B0_t (keyFF_inputPar[8]), .Z0_t (keyFF_keystate_gff_3_MUX_inst1_mux_inst_0_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_3_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_3_MUX_inst1_mux_inst_0_U1_X), .Z0_t (keyFF_keystate_gff_3_MUX_inst1_mux_inst_0_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_3_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_3_MUX_inst1_mux_inst_0_U1_Y), .B0_t (keyFF_outputPar[4]), .Z0_t (keyFF_outputPar[8]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_3_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[5]), .B0_t (keyFF_inputPar[9]), .Z0_t (keyFF_keystate_gff_3_MUX_inst1_mux_inst_1_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_3_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_3_MUX_inst1_mux_inst_1_U1_X), .Z0_t (keyFF_keystate_gff_3_MUX_inst1_mux_inst_1_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_3_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_3_MUX_inst1_mux_inst_1_U1_Y), .B0_t (keyFF_outputPar[5]), .Z0_t (keyFF_outputPar[9]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_3_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[6]), .B0_t (keyFF_inputPar[10]), .Z0_t (keyFF_keystate_gff_3_MUX_inst1_mux_inst_2_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_3_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_3_MUX_inst1_mux_inst_2_U1_X), .Z0_t (keyFF_keystate_gff_3_MUX_inst1_mux_inst_2_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_3_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_3_MUX_inst1_mux_inst_2_U1_Y), .B0_t (keyFF_outputPar[6]), .Z0_t (keyFF_outputPar[10]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_3_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[7]), .B0_t (keyFF_inputPar[11]), .Z0_t (keyFF_keystate_gff_3_MUX_inst1_mux_inst_3_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_3_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_3_MUX_inst1_mux_inst_3_U1_X), .Z0_t (keyFF_keystate_gff_3_MUX_inst1_mux_inst_3_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_3_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_3_MUX_inst1_mux_inst_3_U1_Y), .B0_t (keyFF_outputPar[7]), .Z0_t (keyFF_outputPar[11]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_4_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[8]), .B0_t (keyFF_inputPar[12]), .Z0_t (keyFF_keystate_gff_4_MUX_inst1_mux_inst_0_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_4_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_4_MUX_inst1_mux_inst_0_U1_X), .Z0_t (keyFF_keystate_gff_4_MUX_inst1_mux_inst_0_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_4_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_4_MUX_inst1_mux_inst_0_U1_Y), .B0_t (keyFF_outputPar[8]), .Z0_t (keyFF_outputPar[12]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_4_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[9]), .B0_t (keyFF_inputPar[13]), .Z0_t (keyFF_keystate_gff_4_MUX_inst1_mux_inst_1_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_4_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_4_MUX_inst1_mux_inst_1_U1_X), .Z0_t (keyFF_keystate_gff_4_MUX_inst1_mux_inst_1_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_4_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_4_MUX_inst1_mux_inst_1_U1_Y), .B0_t (keyFF_outputPar[9]), .Z0_t (keyFF_outputPar[13]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_4_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[10]), .B0_t (keyFF_inputPar[14]), .Z0_t (keyFF_keystate_gff_4_MUX_inst1_mux_inst_2_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_4_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_4_MUX_inst1_mux_inst_2_U1_X), .Z0_t (keyFF_keystate_gff_4_MUX_inst1_mux_inst_2_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_4_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_4_MUX_inst1_mux_inst_2_U1_Y), .B0_t (keyFF_outputPar[10]), .Z0_t (keyFF_outputPar[14]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_4_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[11]), .B0_t (keyFF_inputPar[15]), .Z0_t (keyFF_keystate_gff_4_MUX_inst1_mux_inst_3_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_4_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_4_MUX_inst1_mux_inst_3_U1_X), .Z0_t (keyFF_keystate_gff_4_MUX_inst1_mux_inst_3_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_4_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_4_MUX_inst1_mux_inst_3_U1_Y), .B0_t (keyFF_outputPar[11]), .Z0_t (keyFF_outputPar[15]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_5_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[12]), .B0_t (keyFF_inputPar[16]), .Z0_t (keyFF_keystate_gff_5_MUX_inst1_mux_inst_0_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_5_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_5_MUX_inst1_mux_inst_0_U1_X), .Z0_t (keyFF_keystate_gff_5_MUX_inst1_mux_inst_0_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_5_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_5_MUX_inst1_mux_inst_0_U1_Y), .B0_t (keyFF_outputPar[12]), .Z0_t (keyFF_outputPar[16]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_5_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[13]), .B0_t (keyFF_inputPar[17]), .Z0_t (keyFF_keystate_gff_5_MUX_inst1_mux_inst_1_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_5_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_5_MUX_inst1_mux_inst_1_U1_X), .Z0_t (keyFF_keystate_gff_5_MUX_inst1_mux_inst_1_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_5_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_5_MUX_inst1_mux_inst_1_U1_Y), .B0_t (keyFF_outputPar[13]), .Z0_t (keyFF_outputPar[17]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_5_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[14]), .B0_t (keyFF_inputPar[18]), .Z0_t (keyFF_keystate_gff_5_MUX_inst1_mux_inst_2_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_5_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_5_MUX_inst1_mux_inst_2_U1_X), .Z0_t (keyFF_keystate_gff_5_MUX_inst1_mux_inst_2_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_5_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_5_MUX_inst1_mux_inst_2_U1_Y), .B0_t (keyFF_outputPar[14]), .Z0_t (keyFF_outputPar[18]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_5_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[15]), .B0_t (keyFF_inputPar[19]), .Z0_t (keyFF_keystate_gff_5_MUX_inst1_mux_inst_3_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_5_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_5_MUX_inst1_mux_inst_3_U1_X), .Z0_t (keyFF_keystate_gff_5_MUX_inst1_mux_inst_3_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_5_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_5_MUX_inst1_mux_inst_3_U1_Y), .B0_t (keyFF_outputPar[15]), .Z0_t (keyFF_outputPar[19]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_6_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[16]), .B0_t (keyFF_inputPar[20]), .Z0_t (keyFF_keystate_gff_6_MUX_inst1_mux_inst_0_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_6_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_6_MUX_inst1_mux_inst_0_U1_X), .Z0_t (keyFF_keystate_gff_6_MUX_inst1_mux_inst_0_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_6_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_6_MUX_inst1_mux_inst_0_U1_Y), .B0_t (keyFF_outputPar[16]), .Z0_t (keyFF_outputPar[20]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_6_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[17]), .B0_t (keyFF_inputPar[21]), .Z0_t (keyFF_keystate_gff_6_MUX_inst1_mux_inst_1_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_6_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_6_MUX_inst1_mux_inst_1_U1_X), .Z0_t (keyFF_keystate_gff_6_MUX_inst1_mux_inst_1_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_6_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_6_MUX_inst1_mux_inst_1_U1_Y), .B0_t (keyFF_outputPar[17]), .Z0_t (keyFF_outputPar[21]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_6_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[18]), .B0_t (keyFF_inputPar[22]), .Z0_t (keyFF_keystate_gff_6_MUX_inst1_mux_inst_2_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_6_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_6_MUX_inst1_mux_inst_2_U1_X), .Z0_t (keyFF_keystate_gff_6_MUX_inst1_mux_inst_2_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_6_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_6_MUX_inst1_mux_inst_2_U1_Y), .B0_t (keyFF_outputPar[18]), .Z0_t (keyFF_outputPar[22]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_6_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[19]), .B0_t (keyFF_inputPar[23]), .Z0_t (keyFF_keystate_gff_6_MUX_inst1_mux_inst_3_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_6_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_6_MUX_inst1_mux_inst_3_U1_X), .Z0_t (keyFF_keystate_gff_6_MUX_inst1_mux_inst_3_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_6_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_6_MUX_inst1_mux_inst_3_U1_Y), .B0_t (keyFF_outputPar[19]), .Z0_t (keyFF_outputPar[23]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_7_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[20]), .B0_t (keyFF_inputPar[24]), .Z0_t (keyFF_keystate_gff_7_MUX_inst1_mux_inst_0_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_7_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_7_MUX_inst1_mux_inst_0_U1_X), .Z0_t (keyFF_keystate_gff_7_MUX_inst1_mux_inst_0_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_7_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_7_MUX_inst1_mux_inst_0_U1_Y), .B0_t (keyFF_outputPar[20]), .Z0_t (keyFF_outputPar[24]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_7_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[21]), .B0_t (keyFF_inputPar[25]), .Z0_t (keyFF_keystate_gff_7_MUX_inst1_mux_inst_1_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_7_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_7_MUX_inst1_mux_inst_1_U1_X), .Z0_t (keyFF_keystate_gff_7_MUX_inst1_mux_inst_1_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_7_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_7_MUX_inst1_mux_inst_1_U1_Y), .B0_t (keyFF_outputPar[21]), .Z0_t (keyFF_outputPar[25]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_7_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[22]), .B0_t (keyFF_inputPar[26]), .Z0_t (keyFF_keystate_gff_7_MUX_inst1_mux_inst_2_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_7_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_7_MUX_inst1_mux_inst_2_U1_X), .Z0_t (keyFF_keystate_gff_7_MUX_inst1_mux_inst_2_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_7_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_7_MUX_inst1_mux_inst_2_U1_Y), .B0_t (keyFF_outputPar[22]), .Z0_t (keyFF_outputPar[26]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_7_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[23]), .B0_t (keyFF_inputPar[27]), .Z0_t (keyFF_keystate_gff_7_MUX_inst1_mux_inst_3_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_7_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_7_MUX_inst1_mux_inst_3_U1_X), .Z0_t (keyFF_keystate_gff_7_MUX_inst1_mux_inst_3_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_7_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_7_MUX_inst1_mux_inst_3_U1_Y), .B0_t (keyFF_outputPar[23]), .Z0_t (keyFF_outputPar[27]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_8_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[24]), .B0_t (keyFF_inputPar[28]), .Z0_t (keyFF_keystate_gff_8_MUX_inst1_mux_inst_0_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_8_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_8_MUX_inst1_mux_inst_0_U1_X), .Z0_t (keyFF_keystate_gff_8_MUX_inst1_mux_inst_0_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_8_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_8_MUX_inst1_mux_inst_0_U1_Y), .B0_t (keyFF_outputPar[24]), .Z0_t (keyFF_outputPar[28]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_8_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[25]), .B0_t (keyFF_inputPar[29]), .Z0_t (keyFF_keystate_gff_8_MUX_inst1_mux_inst_1_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_8_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_8_MUX_inst1_mux_inst_1_U1_X), .Z0_t (keyFF_keystate_gff_8_MUX_inst1_mux_inst_1_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_8_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_8_MUX_inst1_mux_inst_1_U1_Y), .B0_t (keyFF_outputPar[25]), .Z0_t (keyFF_outputPar[29]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_8_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[26]), .B0_t (keyFF_inputPar[30]), .Z0_t (keyFF_keystate_gff_8_MUX_inst1_mux_inst_2_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_8_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_8_MUX_inst1_mux_inst_2_U1_X), .Z0_t (keyFF_keystate_gff_8_MUX_inst1_mux_inst_2_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_8_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_8_MUX_inst1_mux_inst_2_U1_Y), .B0_t (keyFF_outputPar[26]), .Z0_t (keyFF_outputPar[30]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_8_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[27]), .B0_t (keyFF_inputPar[31]), .Z0_t (keyFF_keystate_gff_8_MUX_inst1_mux_inst_3_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_8_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_8_MUX_inst1_mux_inst_3_U1_X), .Z0_t (keyFF_keystate_gff_8_MUX_inst1_mux_inst_3_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_8_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_8_MUX_inst1_mux_inst_3_U1_Y), .B0_t (keyFF_outputPar[27]), .Z0_t (keyFF_outputPar[31]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_9_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[28]), .B0_t (keyFF_inputPar[32]), .Z0_t (keyFF_keystate_gff_9_MUX_inst1_mux_inst_0_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_9_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_9_MUX_inst1_mux_inst_0_U1_X), .Z0_t (keyFF_keystate_gff_9_MUX_inst1_mux_inst_0_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_9_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_9_MUX_inst1_mux_inst_0_U1_Y), .B0_t (keyFF_outputPar[28]), .Z0_t (keyFF_outputPar[32]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_9_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[29]), .B0_t (keyFF_inputPar[33]), .Z0_t (keyFF_keystate_gff_9_MUX_inst1_mux_inst_1_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_9_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_9_MUX_inst1_mux_inst_1_U1_X), .Z0_t (keyFF_keystate_gff_9_MUX_inst1_mux_inst_1_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_9_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_9_MUX_inst1_mux_inst_1_U1_Y), .B0_t (keyFF_outputPar[29]), .Z0_t (keyFF_outputPar[33]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_9_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[30]), .B0_t (keyFF_inputPar[34]), .Z0_t (keyFF_keystate_gff_9_MUX_inst1_mux_inst_2_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_9_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_9_MUX_inst1_mux_inst_2_U1_X), .Z0_t (keyFF_keystate_gff_9_MUX_inst1_mux_inst_2_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_9_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_9_MUX_inst1_mux_inst_2_U1_Y), .B0_t (keyFF_outputPar[30]), .Z0_t (keyFF_outputPar[34]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_9_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[31]), .B0_t (keyFF_inputPar[35]), .Z0_t (keyFF_keystate_gff_9_MUX_inst1_mux_inst_3_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_9_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_9_MUX_inst1_mux_inst_3_U1_X), .Z0_t (keyFF_keystate_gff_9_MUX_inst1_mux_inst_3_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_9_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_9_MUX_inst1_mux_inst_3_U1_Y), .B0_t (keyFF_outputPar[31]), .Z0_t (keyFF_outputPar[35]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_10_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[32]), .B0_t (keyFF_inputPar[36]), .Z0_t (keyFF_keystate_gff_10_MUX_inst1_mux_inst_0_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_10_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_10_MUX_inst1_mux_inst_0_U1_X), .Z0_t (keyFF_keystate_gff_10_MUX_inst1_mux_inst_0_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_10_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_10_MUX_inst1_mux_inst_0_U1_Y), .B0_t (keyFF_outputPar[32]), .Z0_t (keyFF_outputPar[36]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_10_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[33]), .B0_t (keyFF_inputPar[37]), .Z0_t (keyFF_keystate_gff_10_MUX_inst1_mux_inst_1_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_10_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_10_MUX_inst1_mux_inst_1_U1_X), .Z0_t (keyFF_keystate_gff_10_MUX_inst1_mux_inst_1_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_10_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_10_MUX_inst1_mux_inst_1_U1_Y), .B0_t (keyFF_outputPar[33]), .Z0_t (keyFF_outputPar[37]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_10_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[34]), .B0_t (keyFF_inputPar[38]), .Z0_t (keyFF_keystate_gff_10_MUX_inst1_mux_inst_2_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_10_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_10_MUX_inst1_mux_inst_2_U1_X), .Z0_t (keyFF_keystate_gff_10_MUX_inst1_mux_inst_2_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_10_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_10_MUX_inst1_mux_inst_2_U1_Y), .B0_t (keyFF_outputPar[34]), .Z0_t (keyFF_outputPar[38]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_10_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[35]), .B0_t (keyFF_inputPar[39]), .Z0_t (keyFF_keystate_gff_10_MUX_inst1_mux_inst_3_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_10_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_10_MUX_inst1_mux_inst_3_U1_X), .Z0_t (keyFF_keystate_gff_10_MUX_inst1_mux_inst_3_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_10_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_10_MUX_inst1_mux_inst_3_U1_Y), .B0_t (keyFF_outputPar[35]), .Z0_t (keyFF_outputPar[39]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_11_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[36]), .B0_t (keyFF_inputPar[40]), .Z0_t (keyFF_keystate_gff_11_MUX_inst1_mux_inst_0_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_11_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_11_MUX_inst1_mux_inst_0_U1_X), .Z0_t (keyFF_keystate_gff_11_MUX_inst1_mux_inst_0_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_11_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_11_MUX_inst1_mux_inst_0_U1_Y), .B0_t (keyFF_outputPar[36]), .Z0_t (keyFF_outputPar[40]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_11_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[37]), .B0_t (keyFF_inputPar[41]), .Z0_t (keyFF_keystate_gff_11_MUX_inst1_mux_inst_1_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_11_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_11_MUX_inst1_mux_inst_1_U1_X), .Z0_t (keyFF_keystate_gff_11_MUX_inst1_mux_inst_1_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_11_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_11_MUX_inst1_mux_inst_1_U1_Y), .B0_t (keyFF_outputPar[37]), .Z0_t (keyFF_outputPar[41]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_11_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[38]), .B0_t (keyFF_inputPar[42]), .Z0_t (keyFF_keystate_gff_11_MUX_inst1_mux_inst_2_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_11_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_11_MUX_inst1_mux_inst_2_U1_X), .Z0_t (keyFF_keystate_gff_11_MUX_inst1_mux_inst_2_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_11_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_11_MUX_inst1_mux_inst_2_U1_Y), .B0_t (keyFF_outputPar[38]), .Z0_t (keyFF_outputPar[42]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_11_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[39]), .B0_t (keyFF_inputPar[43]), .Z0_t (keyFF_keystate_gff_11_MUX_inst1_mux_inst_3_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_11_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_11_MUX_inst1_mux_inst_3_U1_X), .Z0_t (keyFF_keystate_gff_11_MUX_inst1_mux_inst_3_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_11_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_11_MUX_inst1_mux_inst_3_U1_Y), .B0_t (keyFF_outputPar[39]), .Z0_t (keyFF_outputPar[43]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_12_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[40]), .B0_t (keyFF_inputPar[44]), .Z0_t (keyFF_keystate_gff_12_MUX_inst1_mux_inst_0_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_12_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_12_MUX_inst1_mux_inst_0_U1_X), .Z0_t (keyFF_keystate_gff_12_MUX_inst1_mux_inst_0_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_12_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_12_MUX_inst1_mux_inst_0_U1_Y), .B0_t (keyFF_outputPar[40]), .Z0_t (keyFF_outputPar[44]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_12_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[41]), .B0_t (keyFF_inputPar[45]), .Z0_t (keyFF_keystate_gff_12_MUX_inst1_mux_inst_1_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_12_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_12_MUX_inst1_mux_inst_1_U1_X), .Z0_t (keyFF_keystate_gff_12_MUX_inst1_mux_inst_1_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_12_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_12_MUX_inst1_mux_inst_1_U1_Y), .B0_t (keyFF_outputPar[41]), .Z0_t (keyFF_outputPar[45]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_12_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[42]), .B0_t (keyFF_inputPar[46]), .Z0_t (keyFF_keystate_gff_12_MUX_inst1_mux_inst_2_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_12_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_12_MUX_inst1_mux_inst_2_U1_X), .Z0_t (keyFF_keystate_gff_12_MUX_inst1_mux_inst_2_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_12_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_12_MUX_inst1_mux_inst_2_U1_Y), .B0_t (keyFF_outputPar[42]), .Z0_t (keyFF_outputPar[46]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_12_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[43]), .B0_t (keyFF_inputPar[47]), .Z0_t (keyFF_keystate_gff_12_MUX_inst1_mux_inst_3_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_12_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_12_MUX_inst1_mux_inst_3_U1_X), .Z0_t (keyFF_keystate_gff_12_MUX_inst1_mux_inst_3_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_12_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_12_MUX_inst1_mux_inst_3_U1_Y), .B0_t (keyFF_outputPar[43]), .Z0_t (keyFF_outputPar[47]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_13_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[44]), .B0_t (keyFF_inputPar[48]), .Z0_t (keyFF_keystate_gff_13_MUX_inst1_mux_inst_0_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_13_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_13_MUX_inst1_mux_inst_0_U1_X), .Z0_t (keyFF_keystate_gff_13_MUX_inst1_mux_inst_0_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_13_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_13_MUX_inst1_mux_inst_0_U1_Y), .B0_t (keyFF_outputPar[44]), .Z0_t (keyFF_outputPar[48]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_13_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[45]), .B0_t (keyFF_inputPar[49]), .Z0_t (keyFF_keystate_gff_13_MUX_inst1_mux_inst_1_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_13_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_13_MUX_inst1_mux_inst_1_U1_X), .Z0_t (keyFF_keystate_gff_13_MUX_inst1_mux_inst_1_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_13_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_13_MUX_inst1_mux_inst_1_U1_Y), .B0_t (keyFF_outputPar[45]), .Z0_t (keyFF_outputPar[49]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_13_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[46]), .B0_t (keyFF_inputPar[50]), .Z0_t (keyFF_keystate_gff_13_MUX_inst1_mux_inst_2_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_13_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_13_MUX_inst1_mux_inst_2_U1_X), .Z0_t (keyFF_keystate_gff_13_MUX_inst1_mux_inst_2_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_13_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_13_MUX_inst1_mux_inst_2_U1_Y), .B0_t (keyFF_outputPar[46]), .Z0_t (keyFF_outputPar[50]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_13_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[47]), .B0_t (keyFF_inputPar[51]), .Z0_t (keyFF_keystate_gff_13_MUX_inst1_mux_inst_3_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_13_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_13_MUX_inst1_mux_inst_3_U1_X), .Z0_t (keyFF_keystate_gff_13_MUX_inst1_mux_inst_3_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_13_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_13_MUX_inst1_mux_inst_3_U1_Y), .B0_t (keyFF_outputPar[47]), .Z0_t (keyFF_outputPar[51]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_14_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[48]), .B0_t (keyFF_inputPar[52]), .Z0_t (keyFF_keystate_gff_14_MUX_inst1_mux_inst_0_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_14_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_14_MUX_inst1_mux_inst_0_U1_X), .Z0_t (keyFF_keystate_gff_14_MUX_inst1_mux_inst_0_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_14_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_14_MUX_inst1_mux_inst_0_U1_Y), .B0_t (keyFF_outputPar[48]), .Z0_t (keyFF_outputPar[52]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_14_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[49]), .B0_t (keyFF_inputPar[53]), .Z0_t (keyFF_keystate_gff_14_MUX_inst1_mux_inst_1_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_14_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_14_MUX_inst1_mux_inst_1_U1_X), .Z0_t (keyFF_keystate_gff_14_MUX_inst1_mux_inst_1_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_14_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_14_MUX_inst1_mux_inst_1_U1_Y), .B0_t (keyFF_outputPar[49]), .Z0_t (keyFF_outputPar[53]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_14_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[50]), .B0_t (keyFF_inputPar[54]), .Z0_t (keyFF_keystate_gff_14_MUX_inst1_mux_inst_2_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_14_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_14_MUX_inst1_mux_inst_2_U1_X), .Z0_t (keyFF_keystate_gff_14_MUX_inst1_mux_inst_2_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_14_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_14_MUX_inst1_mux_inst_2_U1_Y), .B0_t (keyFF_outputPar[50]), .Z0_t (keyFF_outputPar[54]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_14_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[51]), .B0_t (keyFF_inputPar[55]), .Z0_t (keyFF_keystate_gff_14_MUX_inst1_mux_inst_3_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_14_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_14_MUX_inst1_mux_inst_3_U1_X), .Z0_t (keyFF_keystate_gff_14_MUX_inst1_mux_inst_3_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_14_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_14_MUX_inst1_mux_inst_3_U1_Y), .B0_t (keyFF_outputPar[51]), .Z0_t (keyFF_outputPar[55]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_15_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[52]), .B0_t (keyFF_inputPar[56]), .Z0_t (keyFF_keystate_gff_15_MUX_inst1_mux_inst_0_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_15_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_15_MUX_inst1_mux_inst_0_U1_X), .Z0_t (keyFF_keystate_gff_15_MUX_inst1_mux_inst_0_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_15_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_15_MUX_inst1_mux_inst_0_U1_Y), .B0_t (keyFF_outputPar[52]), .Z0_t (keyFF_outputPar[56]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_15_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[53]), .B0_t (keyFF_inputPar[57]), .Z0_t (keyFF_keystate_gff_15_MUX_inst1_mux_inst_1_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_15_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_15_MUX_inst1_mux_inst_1_U1_X), .Z0_t (keyFF_keystate_gff_15_MUX_inst1_mux_inst_1_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_15_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_15_MUX_inst1_mux_inst_1_U1_Y), .B0_t (keyFF_outputPar[53]), .Z0_t (keyFF_outputPar[57]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_15_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[54]), .B0_t (keyFF_inputPar[58]), .Z0_t (keyFF_keystate_gff_15_MUX_inst1_mux_inst_2_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_15_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_15_MUX_inst1_mux_inst_2_U1_X), .Z0_t (keyFF_keystate_gff_15_MUX_inst1_mux_inst_2_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_15_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_15_MUX_inst1_mux_inst_2_U1_Y), .B0_t (keyFF_outputPar[54]), .Z0_t (keyFF_outputPar[58]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_15_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[55]), .B0_t (keyFF_inputPar[59]), .Z0_t (keyFF_keystate_gff_15_MUX_inst1_mux_inst_3_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_15_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_15_MUX_inst1_mux_inst_3_U1_X), .Z0_t (keyFF_keystate_gff_15_MUX_inst1_mux_inst_3_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_15_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_15_MUX_inst1_mux_inst_3_U1_Y), .B0_t (keyFF_outputPar[55]), .Z0_t (keyFF_outputPar[59]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_16_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[56]), .B0_t (keyFF_inputPar[60]), .Z0_t (keyFF_keystate_gff_16_MUX_inst1_mux_inst_0_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_16_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_16_MUX_inst1_mux_inst_0_U1_X), .Z0_t (keyFF_keystate_gff_16_MUX_inst1_mux_inst_0_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_16_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_16_MUX_inst1_mux_inst_0_U1_Y), .B0_t (keyFF_outputPar[56]), .Z0_t (keyFF_outputPar[60]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_16_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[57]), .B0_t (keyFF_inputPar[61]), .Z0_t (keyFF_keystate_gff_16_MUX_inst1_mux_inst_1_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_16_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_16_MUX_inst1_mux_inst_1_U1_X), .Z0_t (keyFF_keystate_gff_16_MUX_inst1_mux_inst_1_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_16_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_16_MUX_inst1_mux_inst_1_U1_Y), .B0_t (keyFF_outputPar[57]), .Z0_t (keyFF_outputPar[61]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_16_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[58]), .B0_t (keyFF_inputPar[62]), .Z0_t (keyFF_keystate_gff_16_MUX_inst1_mux_inst_2_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_16_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_16_MUX_inst1_mux_inst_2_U1_X), .Z0_t (keyFF_keystate_gff_16_MUX_inst1_mux_inst_2_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_16_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_16_MUX_inst1_mux_inst_2_U1_Y), .B0_t (keyFF_outputPar[58]), .Z0_t (keyFF_outputPar[62]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_16_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[59]), .B0_t (keyFF_inputPar[63]), .Z0_t (keyFF_keystate_gff_16_MUX_inst1_mux_inst_3_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_16_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_16_MUX_inst1_mux_inst_3_U1_X), .Z0_t (keyFF_keystate_gff_16_MUX_inst1_mux_inst_3_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_16_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_16_MUX_inst1_mux_inst_3_U1_Y), .B0_t (keyFF_outputPar[59]), .Z0_t (keyFF_outputPar[63]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_17_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[60]), .B0_t (keyFF_inputPar[64]), .Z0_t (keyFF_keystate_gff_17_MUX_inst1_mux_inst_0_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_17_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_17_MUX_inst1_mux_inst_0_U1_X), .Z0_t (keyFF_keystate_gff_17_MUX_inst1_mux_inst_0_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_17_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_17_MUX_inst1_mux_inst_0_U1_Y), .B0_t (keyFF_outputPar[60]), .Z0_t (keyFF_outputPar[64]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_17_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[61]), .B0_t (keyFF_inputPar[65]), .Z0_t (keyFF_keystate_gff_17_MUX_inst1_mux_inst_1_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_17_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_17_MUX_inst1_mux_inst_1_U1_X), .Z0_t (keyFF_keystate_gff_17_MUX_inst1_mux_inst_1_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_17_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_17_MUX_inst1_mux_inst_1_U1_Y), .B0_t (keyFF_outputPar[61]), .Z0_t (keyFF_outputPar[65]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_17_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[62]), .B0_t (keyFF_inputPar[66]), .Z0_t (keyFF_keystate_gff_17_MUX_inst1_mux_inst_2_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_17_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_17_MUX_inst1_mux_inst_2_U1_X), .Z0_t (keyFF_keystate_gff_17_MUX_inst1_mux_inst_2_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_17_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_17_MUX_inst1_mux_inst_2_U1_Y), .B0_t (keyFF_outputPar[62]), .Z0_t (keyFF_outputPar[66]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_17_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[63]), .B0_t (keyFF_inputPar[67]), .Z0_t (keyFF_keystate_gff_17_MUX_inst1_mux_inst_3_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_17_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_17_MUX_inst1_mux_inst_3_U1_X), .Z0_t (keyFF_keystate_gff_17_MUX_inst1_mux_inst_3_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_17_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_17_MUX_inst1_mux_inst_3_U1_Y), .B0_t (keyFF_outputPar[63]), .Z0_t (keyFF_outputPar[67]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_18_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[64]), .B0_t (keyFF_inputPar[68]), .Z0_t (keyFF_keystate_gff_18_MUX_inst1_mux_inst_0_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_18_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_18_MUX_inst1_mux_inst_0_U1_X), .Z0_t (keyFF_keystate_gff_18_MUX_inst1_mux_inst_0_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_18_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_18_MUX_inst1_mux_inst_0_U1_Y), .B0_t (keyFF_outputPar[64]), .Z0_t (keyFF_outputPar[68]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_18_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[65]), .B0_t (keyFF_inputPar[69]), .Z0_t (keyFF_keystate_gff_18_MUX_inst1_mux_inst_1_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_18_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_18_MUX_inst1_mux_inst_1_U1_X), .Z0_t (keyFF_keystate_gff_18_MUX_inst1_mux_inst_1_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_18_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_18_MUX_inst1_mux_inst_1_U1_Y), .B0_t (keyFF_outputPar[65]), .Z0_t (keyFF_outputPar[69]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_18_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[66]), .B0_t (keyFF_inputPar[70]), .Z0_t (keyFF_keystate_gff_18_MUX_inst1_mux_inst_2_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_18_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_18_MUX_inst1_mux_inst_2_U1_X), .Z0_t (keyFF_keystate_gff_18_MUX_inst1_mux_inst_2_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_18_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_18_MUX_inst1_mux_inst_2_U1_Y), .B0_t (keyFF_outputPar[66]), .Z0_t (keyFF_outputPar[70]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_18_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[67]), .B0_t (keyFF_inputPar[71]), .Z0_t (keyFF_keystate_gff_18_MUX_inst1_mux_inst_3_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_18_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_18_MUX_inst1_mux_inst_3_U1_X), .Z0_t (keyFF_keystate_gff_18_MUX_inst1_mux_inst_3_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_18_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_18_MUX_inst1_mux_inst_3_U1_Y), .B0_t (keyFF_outputPar[67]), .Z0_t (keyFF_outputPar[71]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_19_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[68]), .B0_t (keyFF_inputPar[72]), .Z0_t (keyFF_keystate_gff_19_MUX_inst1_mux_inst_0_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_19_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_19_MUX_inst1_mux_inst_0_U1_X), .Z0_t (keyFF_keystate_gff_19_MUX_inst1_mux_inst_0_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_19_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_19_MUX_inst1_mux_inst_0_U1_Y), .B0_t (keyFF_outputPar[68]), .Z0_t (keyFF_outputPar[72]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_19_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[69]), .B0_t (keyFF_inputPar[73]), .Z0_t (keyFF_keystate_gff_19_MUX_inst1_mux_inst_1_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_19_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_19_MUX_inst1_mux_inst_1_U1_X), .Z0_t (keyFF_keystate_gff_19_MUX_inst1_mux_inst_1_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_19_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_19_MUX_inst1_mux_inst_1_U1_Y), .B0_t (keyFF_outputPar[69]), .Z0_t (keyFF_outputPar[73]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_19_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[70]), .B0_t (keyFF_inputPar[74]), .Z0_t (keyFF_keystate_gff_19_MUX_inst1_mux_inst_2_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_19_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_19_MUX_inst1_mux_inst_2_U1_X), .Z0_t (keyFF_keystate_gff_19_MUX_inst1_mux_inst_2_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_19_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_19_MUX_inst1_mux_inst_2_U1_Y), .B0_t (keyFF_outputPar[70]), .Z0_t (keyFF_outputPar[74]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_19_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[71]), .B0_t (keyFF_inputPar[75]), .Z0_t (keyFF_keystate_gff_19_MUX_inst1_mux_inst_3_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_19_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_19_MUX_inst1_mux_inst_3_U1_X), .Z0_t (keyFF_keystate_gff_19_MUX_inst1_mux_inst_3_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_19_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_19_MUX_inst1_mux_inst_3_U1_Y), .B0_t (keyFF_outputPar[71]), .Z0_t (keyFF_outputPar[75]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_20_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[72]), .B0_t (keyFF_inputPar[76]), .Z0_t (keyFF_keystate_gff_20_MUX_inst1_mux_inst_0_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_20_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_20_MUX_inst1_mux_inst_0_U1_X), .Z0_t (keyFF_keystate_gff_20_MUX_inst1_mux_inst_0_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_20_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_20_MUX_inst1_mux_inst_0_U1_Y), .B0_t (keyFF_outputPar[72]), .Z0_t (roundkey[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_20_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[73]), .B0_t (keyFF_inputPar[77]), .Z0_t (keyFF_keystate_gff_20_MUX_inst1_mux_inst_1_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_20_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_20_MUX_inst1_mux_inst_1_U1_X), .Z0_t (keyFF_keystate_gff_20_MUX_inst1_mux_inst_1_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_20_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_20_MUX_inst1_mux_inst_1_U1_Y), .B0_t (keyFF_outputPar[73]), .Z0_t (roundkey[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_20_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[74]), .B0_t (keyFF_inputPar[78]), .Z0_t (keyFF_keystate_gff_20_MUX_inst1_mux_inst_2_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_20_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_20_MUX_inst1_mux_inst_2_U1_X), .Z0_t (keyFF_keystate_gff_20_MUX_inst1_mux_inst_2_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_20_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_20_MUX_inst1_mux_inst_2_U1_Y), .B0_t (keyFF_outputPar[74]), .Z0_t (roundkey[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_20_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[75]), .B0_t (keyFF_inputPar[79]), .Z0_t (keyFF_keystate_gff_20_MUX_inst1_mux_inst_3_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_20_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (fsm_rst_countSerial), .B0_t (keyFF_keystate_gff_20_MUX_inst1_mux_inst_3_U1_X), .Z0_t (keyFF_keystate_gff_20_MUX_inst1_mux_inst_3_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_20_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_20_MUX_inst1_mux_inst_3_U1_Y), .B0_t (keyFF_outputPar[75]), .Z0_t (roundkey[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_0_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[3]), .B0_t (key[0]), .Z0_t (keyFF_MUX_inputPar_mux_inst_0_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_0_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_0_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_0_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_0_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_0_U1_Y), .B0_t (keyFF_outputPar[3]), .Z0_t (keyFF_inputPar[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_1_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[4]), .B0_t (key[1]), .Z0_t (keyFF_MUX_inputPar_mux_inst_1_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_1_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_1_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_1_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_1_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_1_U1_Y), .B0_t (keyFF_outputPar[4]), .Z0_t (keyFF_inputPar[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_2_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[5]), .B0_t (key[2]), .Z0_t (keyFF_MUX_inputPar_mux_inst_2_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_2_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_2_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_2_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_2_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_2_U1_Y), .B0_t (keyFF_outputPar[5]), .Z0_t (keyFF_inputPar[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_3_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[6]), .B0_t (key[3]), .Z0_t (keyFF_MUX_inputPar_mux_inst_3_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_3_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_3_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_3_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_3_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_3_U1_Y), .B0_t (keyFF_outputPar[6]), .Z0_t (keyFF_inputPar[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_4_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[7]), .B0_t (key[4]), .Z0_t (keyFF_MUX_inputPar_mux_inst_4_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_4_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_4_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_4_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_4_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_4_U1_Y), .B0_t (keyFF_outputPar[7]), .Z0_t (keyFF_inputPar[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_5_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[8]), .B0_t (key[5]), .Z0_t (keyFF_MUX_inputPar_mux_inst_5_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_5_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_5_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_5_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_5_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_5_U1_Y), .B0_t (keyFF_outputPar[8]), .Z0_t (keyFF_inputPar[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_6_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[9]), .B0_t (key[6]), .Z0_t (keyFF_MUX_inputPar_mux_inst_6_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_6_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_6_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_6_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_6_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_6_U1_Y), .B0_t (keyFF_outputPar[9]), .Z0_t (keyFF_inputPar[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_7_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[10]), .B0_t (key[7]), .Z0_t (keyFF_MUX_inputPar_mux_inst_7_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_7_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_7_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_7_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_7_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_7_U1_Y), .B0_t (keyFF_outputPar[10]), .Z0_t (keyFF_inputPar[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_8_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[11]), .B0_t (key[8]), .Z0_t (keyFF_MUX_inputPar_mux_inst_8_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_8_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_8_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_8_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_8_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_8_U1_Y), .B0_t (keyFF_outputPar[11]), .Z0_t (keyFF_inputPar[8]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_9_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[12]), .B0_t (key[9]), .Z0_t (keyFF_MUX_inputPar_mux_inst_9_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_9_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_9_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_9_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_9_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_9_U1_Y), .B0_t (keyFF_outputPar[12]), .Z0_t (keyFF_inputPar[9]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_10_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[13]), .B0_t (key[10]), .Z0_t (keyFF_MUX_inputPar_mux_inst_10_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_10_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_10_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_10_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_10_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_10_U1_Y), .B0_t (keyFF_outputPar[13]), .Z0_t (keyFF_inputPar[10]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_11_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[14]), .B0_t (key[11]), .Z0_t (keyFF_MUX_inputPar_mux_inst_11_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_11_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_11_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_11_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_11_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_11_U1_Y), .B0_t (keyFF_outputPar[14]), .Z0_t (keyFF_inputPar[11]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_12_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[15]), .B0_t (key[12]), .Z0_t (keyFF_MUX_inputPar_mux_inst_12_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_12_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_12_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_12_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_12_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_12_U1_Y), .B0_t (keyFF_outputPar[15]), .Z0_t (keyFF_inputPar[12]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_13_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[16]), .B0_t (key[13]), .Z0_t (keyFF_MUX_inputPar_mux_inst_13_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_13_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_13_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_13_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_13_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_13_U1_Y), .B0_t (keyFF_outputPar[16]), .Z0_t (keyFF_inputPar[13]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_14_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[17]), .B0_t (key[14]), .Z0_t (keyFF_MUX_inputPar_mux_inst_14_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_14_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_14_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_14_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_14_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_14_U1_Y), .B0_t (keyFF_outputPar[17]), .Z0_t (keyFF_inputPar[14]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_15_U1_XOR1_U1 ( .A0_t (keyFF_counterAdd[0]), .B0_t (key[15]), .Z0_t (keyFF_MUX_inputPar_mux_inst_15_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_15_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_15_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_15_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_15_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_15_U1_Y), .B0_t (keyFF_counterAdd[0]), .Z0_t (keyFF_inputPar[15]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_16_U1_XOR1_U1 ( .A0_t (keyFF_counterAdd[1]), .B0_t (key[16]), .Z0_t (keyFF_MUX_inputPar_mux_inst_16_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_16_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_16_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_16_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_16_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_16_U1_Y), .B0_t (keyFF_counterAdd[1]), .Z0_t (keyFF_inputPar[16]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_17_U1_XOR1_U1 ( .A0_t (keyFF_counterAdd[2]), .B0_t (key[17]), .Z0_t (keyFF_MUX_inputPar_mux_inst_17_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_17_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_17_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_17_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_17_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_17_U1_Y), .B0_t (keyFF_counterAdd[2]), .Z0_t (keyFF_inputPar[17]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_18_U1_XOR1_U1 ( .A0_t (keyFF_counterAdd[3]), .B0_t (key[18]), .Z0_t (keyFF_MUX_inputPar_mux_inst_18_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_18_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_18_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_18_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_18_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_18_U1_Y), .B0_t (keyFF_counterAdd[3]), .Z0_t (keyFF_inputPar[18]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_19_U1_XOR1_U1 ( .A0_t (keyFF_counterAdd[4]), .B0_t (key[19]), .Z0_t (keyFF_MUX_inputPar_mux_inst_19_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_19_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_19_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_19_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_19_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_19_U1_Y), .B0_t (keyFF_counterAdd[4]), .Z0_t (keyFF_inputPar[19]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_20_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[23]), .B0_t (key[20]), .Z0_t (keyFF_MUX_inputPar_mux_inst_20_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_20_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_20_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_20_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_20_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_20_U1_Y), .B0_t (keyFF_outputPar[23]), .Z0_t (keyFF_inputPar[20]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_21_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[24]), .B0_t (key[21]), .Z0_t (keyFF_MUX_inputPar_mux_inst_21_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_21_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_21_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_21_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_21_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_21_U1_Y), .B0_t (keyFF_outputPar[24]), .Z0_t (keyFF_inputPar[21]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_22_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[25]), .B0_t (key[22]), .Z0_t (keyFF_MUX_inputPar_mux_inst_22_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_22_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_22_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_22_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_22_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_22_U1_Y), .B0_t (keyFF_outputPar[25]), .Z0_t (keyFF_inputPar[22]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_23_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[26]), .B0_t (key[23]), .Z0_t (keyFF_MUX_inputPar_mux_inst_23_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_23_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_23_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_23_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_23_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_23_U1_Y), .B0_t (keyFF_outputPar[26]), .Z0_t (keyFF_inputPar[23]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_24_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[27]), .B0_t (key[24]), .Z0_t (keyFF_MUX_inputPar_mux_inst_24_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_24_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_24_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_24_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_24_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_24_U1_Y), .B0_t (keyFF_outputPar[27]), .Z0_t (keyFF_inputPar[24]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_25_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[28]), .B0_t (key[25]), .Z0_t (keyFF_MUX_inputPar_mux_inst_25_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_25_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_25_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_25_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_25_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_25_U1_Y), .B0_t (keyFF_outputPar[28]), .Z0_t (keyFF_inputPar[25]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_26_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[29]), .B0_t (key[26]), .Z0_t (keyFF_MUX_inputPar_mux_inst_26_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_26_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_26_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_26_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_26_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_26_U1_Y), .B0_t (keyFF_outputPar[29]), .Z0_t (keyFF_inputPar[26]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_27_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[30]), .B0_t (key[27]), .Z0_t (keyFF_MUX_inputPar_mux_inst_27_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_27_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_27_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_27_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_27_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_27_U1_Y), .B0_t (keyFF_outputPar[30]), .Z0_t (keyFF_inputPar[27]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_28_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[31]), .B0_t (key[28]), .Z0_t (keyFF_MUX_inputPar_mux_inst_28_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_28_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_28_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_28_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_28_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_28_U1_Y), .B0_t (keyFF_outputPar[31]), .Z0_t (keyFF_inputPar[28]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_29_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[32]), .B0_t (key[29]), .Z0_t (keyFF_MUX_inputPar_mux_inst_29_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_29_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_29_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_29_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_29_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_29_U1_Y), .B0_t (keyFF_outputPar[32]), .Z0_t (keyFF_inputPar[29]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_30_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[33]), .B0_t (key[30]), .Z0_t (keyFF_MUX_inputPar_mux_inst_30_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_30_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_30_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_30_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_30_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_30_U1_Y), .B0_t (keyFF_outputPar[33]), .Z0_t (keyFF_inputPar[30]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_31_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[34]), .B0_t (key[31]), .Z0_t (keyFF_MUX_inputPar_mux_inst_31_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_31_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_31_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_31_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_31_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_31_U1_Y), .B0_t (keyFF_outputPar[34]), .Z0_t (keyFF_inputPar[31]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_32_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[35]), .B0_t (key[32]), .Z0_t (keyFF_MUX_inputPar_mux_inst_32_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_32_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_32_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_32_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_32_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_32_U1_Y), .B0_t (keyFF_outputPar[35]), .Z0_t (keyFF_inputPar[32]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_33_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[36]), .B0_t (key[33]), .Z0_t (keyFF_MUX_inputPar_mux_inst_33_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_33_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_33_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_33_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_33_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_33_U1_Y), .B0_t (keyFF_outputPar[36]), .Z0_t (keyFF_inputPar[33]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_34_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[37]), .B0_t (key[34]), .Z0_t (keyFF_MUX_inputPar_mux_inst_34_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_34_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_34_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_34_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_34_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_34_U1_Y), .B0_t (keyFF_outputPar[37]), .Z0_t (keyFF_inputPar[34]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_35_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[38]), .B0_t (key[35]), .Z0_t (keyFF_MUX_inputPar_mux_inst_35_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_35_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_35_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_35_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_35_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_35_U1_Y), .B0_t (keyFF_outputPar[38]), .Z0_t (keyFF_inputPar[35]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_36_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[39]), .B0_t (key[36]), .Z0_t (keyFF_MUX_inputPar_mux_inst_36_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_36_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_36_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_36_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_36_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_36_U1_Y), .B0_t (keyFF_outputPar[39]), .Z0_t (keyFF_inputPar[36]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_37_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[40]), .B0_t (key[37]), .Z0_t (keyFF_MUX_inputPar_mux_inst_37_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_37_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_37_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_37_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_37_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_37_U1_Y), .B0_t (keyFF_outputPar[40]), .Z0_t (keyFF_inputPar[37]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_38_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[41]), .B0_t (key[38]), .Z0_t (keyFF_MUX_inputPar_mux_inst_38_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_38_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_38_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_38_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_38_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_38_U1_Y), .B0_t (keyFF_outputPar[41]), .Z0_t (keyFF_inputPar[38]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_39_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[42]), .B0_t (key[39]), .Z0_t (keyFF_MUX_inputPar_mux_inst_39_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_39_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_39_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_39_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_39_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_39_U1_Y), .B0_t (keyFF_outputPar[42]), .Z0_t (keyFF_inputPar[39]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_40_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[43]), .B0_t (key[40]), .Z0_t (keyFF_MUX_inputPar_mux_inst_40_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_40_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_40_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_40_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_40_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_40_U1_Y), .B0_t (keyFF_outputPar[43]), .Z0_t (keyFF_inputPar[40]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_41_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[44]), .B0_t (key[41]), .Z0_t (keyFF_MUX_inputPar_mux_inst_41_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_41_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_41_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_41_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_41_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_41_U1_Y), .B0_t (keyFF_outputPar[44]), .Z0_t (keyFF_inputPar[41]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_42_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[45]), .B0_t (key[42]), .Z0_t (keyFF_MUX_inputPar_mux_inst_42_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_42_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_42_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_42_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_42_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_42_U1_Y), .B0_t (keyFF_outputPar[45]), .Z0_t (keyFF_inputPar[42]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_43_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[46]), .B0_t (key[43]), .Z0_t (keyFF_MUX_inputPar_mux_inst_43_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_43_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_43_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_43_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_43_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_43_U1_Y), .B0_t (keyFF_outputPar[46]), .Z0_t (keyFF_inputPar[43]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_44_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[47]), .B0_t (key[44]), .Z0_t (keyFF_MUX_inputPar_mux_inst_44_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_44_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_44_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_44_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_44_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_44_U1_Y), .B0_t (keyFF_outputPar[47]), .Z0_t (keyFF_inputPar[44]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_45_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[48]), .B0_t (key[45]), .Z0_t (keyFF_MUX_inputPar_mux_inst_45_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_45_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_45_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_45_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_45_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_45_U1_Y), .B0_t (keyFF_outputPar[48]), .Z0_t (keyFF_inputPar[45]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_46_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[49]), .B0_t (key[46]), .Z0_t (keyFF_MUX_inputPar_mux_inst_46_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_46_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_46_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_46_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_46_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_46_U1_Y), .B0_t (keyFF_outputPar[49]), .Z0_t (keyFF_inputPar[46]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_47_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[50]), .B0_t (key[47]), .Z0_t (keyFF_MUX_inputPar_mux_inst_47_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_47_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_47_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_47_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_47_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_47_U1_Y), .B0_t (keyFF_outputPar[50]), .Z0_t (keyFF_inputPar[47]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_48_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[51]), .B0_t (key[48]), .Z0_t (keyFF_MUX_inputPar_mux_inst_48_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_48_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_48_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_48_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_48_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_48_U1_Y), .B0_t (keyFF_outputPar[51]), .Z0_t (keyFF_inputPar[48]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_49_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[52]), .B0_t (key[49]), .Z0_t (keyFF_MUX_inputPar_mux_inst_49_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_49_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_49_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_49_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_49_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_49_U1_Y), .B0_t (keyFF_outputPar[52]), .Z0_t (keyFF_inputPar[49]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_50_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[53]), .B0_t (key[50]), .Z0_t (keyFF_MUX_inputPar_mux_inst_50_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_50_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_50_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_50_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_50_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_50_U1_Y), .B0_t (keyFF_outputPar[53]), .Z0_t (keyFF_inputPar[50]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_51_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[54]), .B0_t (key[51]), .Z0_t (keyFF_MUX_inputPar_mux_inst_51_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_51_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_51_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_51_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_51_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_51_U1_Y), .B0_t (keyFF_outputPar[54]), .Z0_t (keyFF_inputPar[51]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_52_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[55]), .B0_t (key[52]), .Z0_t (keyFF_MUX_inputPar_mux_inst_52_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_52_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_52_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_52_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_52_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_52_U1_Y), .B0_t (keyFF_outputPar[55]), .Z0_t (keyFF_inputPar[52]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_53_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[56]), .B0_t (key[53]), .Z0_t (keyFF_MUX_inputPar_mux_inst_53_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_53_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_53_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_53_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_53_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_53_U1_Y), .B0_t (keyFF_outputPar[56]), .Z0_t (keyFF_inputPar[53]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_54_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[57]), .B0_t (key[54]), .Z0_t (keyFF_MUX_inputPar_mux_inst_54_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_54_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_54_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_54_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_54_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_54_U1_Y), .B0_t (keyFF_outputPar[57]), .Z0_t (keyFF_inputPar[54]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_55_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[58]), .B0_t (key[55]), .Z0_t (keyFF_MUX_inputPar_mux_inst_55_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_55_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_55_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_55_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_55_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_55_U1_Y), .B0_t (keyFF_outputPar[58]), .Z0_t (keyFF_inputPar[55]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_56_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[59]), .B0_t (key[56]), .Z0_t (keyFF_MUX_inputPar_mux_inst_56_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_56_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_56_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_56_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_56_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_56_U1_Y), .B0_t (keyFF_outputPar[59]), .Z0_t (keyFF_inputPar[56]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_57_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[60]), .B0_t (key[57]), .Z0_t (keyFF_MUX_inputPar_mux_inst_57_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_57_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_57_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_57_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_57_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_57_U1_Y), .B0_t (keyFF_outputPar[60]), .Z0_t (keyFF_inputPar[57]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_58_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[61]), .B0_t (key[58]), .Z0_t (keyFF_MUX_inputPar_mux_inst_58_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_58_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_58_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_58_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_58_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_58_U1_Y), .B0_t (keyFF_outputPar[61]), .Z0_t (keyFF_inputPar[58]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_59_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[62]), .B0_t (key[59]), .Z0_t (keyFF_MUX_inputPar_mux_inst_59_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_59_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_59_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_59_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_59_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_59_U1_Y), .B0_t (keyFF_outputPar[62]), .Z0_t (keyFF_inputPar[59]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_60_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[63]), .B0_t (key[60]), .Z0_t (keyFF_MUX_inputPar_mux_inst_60_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_60_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_60_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_60_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_60_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_60_U1_Y), .B0_t (keyFF_outputPar[63]), .Z0_t (keyFF_inputPar[60]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_61_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[64]), .B0_t (key[61]), .Z0_t (keyFF_MUX_inputPar_mux_inst_61_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_61_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_61_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_61_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_61_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_61_U1_Y), .B0_t (keyFF_outputPar[64]), .Z0_t (keyFF_inputPar[61]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_62_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[65]), .B0_t (key[62]), .Z0_t (keyFF_MUX_inputPar_mux_inst_62_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_62_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_62_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_62_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_62_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_62_U1_Y), .B0_t (keyFF_outputPar[65]), .Z0_t (keyFF_inputPar[62]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_63_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[66]), .B0_t (key[63]), .Z0_t (keyFF_MUX_inputPar_mux_inst_63_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_63_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_63_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_63_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_63_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_63_U1_Y), .B0_t (keyFF_outputPar[66]), .Z0_t (keyFF_inputPar[63]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_64_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[67]), .B0_t (key[64]), .Z0_t (keyFF_MUX_inputPar_mux_inst_64_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_64_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_64_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_64_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_64_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_64_U1_Y), .B0_t (keyFF_outputPar[67]), .Z0_t (keyFF_inputPar[64]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_65_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[68]), .B0_t (key[65]), .Z0_t (keyFF_MUX_inputPar_mux_inst_65_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_65_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_65_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_65_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_65_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_65_U1_Y), .B0_t (keyFF_outputPar[68]), .Z0_t (keyFF_inputPar[65]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_66_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[69]), .B0_t (key[66]), .Z0_t (keyFF_MUX_inputPar_mux_inst_66_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_66_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_66_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_66_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_66_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_66_U1_Y), .B0_t (keyFF_outputPar[69]), .Z0_t (keyFF_inputPar[66]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_67_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[70]), .B0_t (key[67]), .Z0_t (keyFF_MUX_inputPar_mux_inst_67_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_67_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_67_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_67_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_67_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_67_U1_Y), .B0_t (keyFF_outputPar[70]), .Z0_t (keyFF_inputPar[67]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_68_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[71]), .B0_t (key[68]), .Z0_t (keyFF_MUX_inputPar_mux_inst_68_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_68_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_68_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_68_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_68_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_68_U1_Y), .B0_t (keyFF_outputPar[71]), .Z0_t (keyFF_inputPar[68]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_69_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[72]), .B0_t (key[69]), .Z0_t (keyFF_MUX_inputPar_mux_inst_69_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_69_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_69_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_69_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_69_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_69_U1_Y), .B0_t (keyFF_outputPar[72]), .Z0_t (keyFF_inputPar[69]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_70_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[73]), .B0_t (key[70]), .Z0_t (keyFF_MUX_inputPar_mux_inst_70_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_70_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_70_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_70_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_70_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_70_U1_Y), .B0_t (keyFF_outputPar[73]), .Z0_t (keyFF_inputPar[70]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_71_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[74]), .B0_t (key[71]), .Z0_t (keyFF_MUX_inputPar_mux_inst_71_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_71_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_71_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_71_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_71_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_71_U1_Y), .B0_t (keyFF_outputPar[74]), .Z0_t (keyFF_inputPar[71]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_72_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[75]), .B0_t (key[72]), .Z0_t (keyFF_MUX_inputPar_mux_inst_72_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_72_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_72_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_72_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_72_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_72_U1_Y), .B0_t (keyFF_outputPar[75]), .Z0_t (keyFF_inputPar[72]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_73_U1_XOR1_U1 ( .A0_t (roundkey[0]), .B0_t (key[73]), .Z0_t (keyFF_MUX_inputPar_mux_inst_73_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_73_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_73_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_73_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_73_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_73_U1_Y), .B0_t (roundkey[0]), .Z0_t (keyFF_inputPar[73]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_74_U1_XOR1_U1 ( .A0_t (roundkey[1]), .B0_t (key[74]), .Z0_t (keyFF_MUX_inputPar_mux_inst_74_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_74_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_74_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_74_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_74_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_74_U1_Y), .B0_t (roundkey[1]), .Z0_t (keyFF_inputPar[74]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_75_U1_XOR1_U1 ( .A0_t (roundkey[2]), .B0_t (key[75]), .Z0_t (keyFF_MUX_inputPar_mux_inst_75_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_75_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_75_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_75_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_75_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_75_U1_Y), .B0_t (roundkey[2]), .Z0_t (keyFF_inputPar[75]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_76_U1_XOR1_U1 ( .A0_t (sboxOut[0]), .B0_t (key[76]), .Z0_t (keyFF_MUX_inputPar_mux_inst_76_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_76_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_76_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_76_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_76_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_76_U1_Y), .B0_t (sboxOut[0]), .Z0_t (keyFF_inputPar[76]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_77_U1_XOR1_U1 ( .A0_t (sboxOut[1]), .B0_t (key[77]), .Z0_t (keyFF_MUX_inputPar_mux_inst_77_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_77_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_77_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_77_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_77_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_77_U1_Y), .B0_t (sboxOut[1]), .Z0_t (keyFF_inputPar[77]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_78_U1_XOR1_U1 ( .A0_t (sboxOut[2]), .B0_t (key[78]), .Z0_t (keyFF_MUX_inputPar_mux_inst_78_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_78_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_78_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_78_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_78_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_78_U1_Y), .B0_t (sboxOut[2]), .Z0_t (keyFF_inputPar[78]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_79_U1_XOR1_U1 ( .A0_t (sboxOut[3]), .B0_t (key[79]), .Z0_t (keyFF_MUX_inputPar_mux_inst_79_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_79_U1_AND1_U1 ( .A0_t (reset), .B0_t (keyFF_MUX_inputPar_mux_inst_79_U1_X), .Z0_t (keyFF_MUX_inputPar_mux_inst_79_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_79_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_79_U1_Y), .B0_t (sboxOut[3]), .Z0_t (keyFF_inputPar[79]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) sboxInst_XOR1_U1 ( .A0_t (sboxIn[2]), .B0_t (sboxIn[1]), .Z0_t (sboxInst_L0) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) sboxInst_XOR2_U1 ( .A0_t (sboxIn[1]), .B0_t (sboxIn[0]), .Z0_t (sboxInst_L1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) sboxInst_XOR3_U1 ( .A0_t (sboxInst_L1), .B0_t (sboxIn[3]), .Z0_t (sboxInst_L2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) sboxInst_XOR16_U1 ( .A0_t (sboxInst_T0), .B0_t (sboxInst_L2), .Z0_t (sboxInst_Q2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) sboxInst_XOR4_U1 ( .A0_t (sboxIn[3]), .B0_t (sboxIn[0]), .Z0_t (sboxInst_L3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) sboxInst_XOR5_U1 ( .A0_t (sboxInst_L3), .B0_t (sboxInst_L0), .Z0_t (sboxInst_Q3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) sboxInst_XOR6_U1 ( .A0_t (sboxIn[3]), .B0_t (sboxIn[1]), .Z0_t (sboxInst_L4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) sboxInst_XOR7_U1 ( .A0_t (sboxInst_T0), .B0_t (sboxInst_T2), .Z0_t (sboxInst_L5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) sboxInst_XOR8_U1 ( .A0_t (sboxInst_L4), .B0_t (sboxInst_L5), .Z0_t (sboxInst_Q6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) sboxInst_XOR9_U1 ( .A0_t (sboxInst_L1), .B0_t (sboxIn[2]), .Z0_t (sboxInst_Q7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) sboxInst_AND1_U1 ( .A0_t (sboxInst_L0), .B0_t (sboxIn[3]), .Z0_t (sboxInst_T0) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) sboxInst_AND2_U1 ( .A0_t (sboxInst_Q2), .B0_t (sboxInst_Q3), .Z0_t (sboxInst_T1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) sboxInst_AND3_U1 ( .A0_t (sboxIn[1]), .B0_t (sboxIn[2]), .Z0_t (sboxInst_T2) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) sboxInst_AND4_U1 ( .A0_t (sboxInst_Q6), .B0_t (sboxInst_Q7), .Z0_t (sboxInst_T3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) sboxInst_XOR10_U1 ( .A0_t (sboxInst_L5), .B0_t (sboxInst_T3), .Z0_t (sboxInst_L7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) sboxInst_XOR11_U1 ( .A0_t (sboxIn[0]), .B0_t (sboxInst_L7), .Z0_t (sboxOut[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) sboxInst_XOR12_U1 ( .A0_t (sboxInst_L5), .B0_t (sboxInst_T1), .Z0_t (sboxInst_L8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) sboxInst_XOR13_U1 ( .A0_t (sboxInst_L1), .B0_t (sboxInst_L8), .Z0_t (sboxOut[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) sboxInst_XOR14_U1 ( .A0_t (sboxInst_L4), .B0_t (sboxInst_T3), .Z0_t (sboxOut[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) sboxInst_XOR15_U1 ( .A0_t (sboxInst_L3), .B0_t (sboxInst_T2), .Z0_t (sboxOut[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_sboxin_mux_inst_0_U1_XOR1_U1 ( .A0_t (stateXORroundkey[0]), .B0_t (roundkey[3]), .Z0_t (MUX_sboxin_mux_inst_0_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_sboxin_mux_inst_0_U1_AND1_U1 ( .A0_t (selSbox), .B0_t (MUX_sboxin_mux_inst_0_U1_X), .Z0_t (MUX_sboxin_mux_inst_0_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_sboxin_mux_inst_0_U1_XOR2_U1 ( .A0_t (MUX_sboxin_mux_inst_0_U1_Y), .B0_t (stateXORroundkey[0]), .Z0_t (sboxIn[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_sboxin_mux_inst_1_U1_XOR1_U1 ( .A0_t (stateXORroundkey[1]), .B0_t (keyRegKS[1]), .Z0_t (MUX_sboxin_mux_inst_1_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_sboxin_mux_inst_1_U1_AND1_U1 ( .A0_t (selSbox), .B0_t (MUX_sboxin_mux_inst_1_U1_X), .Z0_t (MUX_sboxin_mux_inst_1_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_sboxin_mux_inst_1_U1_XOR2_U1 ( .A0_t (MUX_sboxin_mux_inst_1_U1_Y), .B0_t (stateXORroundkey[1]), .Z0_t (sboxIn[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_sboxin_mux_inst_2_U1_XOR1_U1 ( .A0_t (stateXORroundkey[2]), .B0_t (keyRegKS[2]), .Z0_t (MUX_sboxin_mux_inst_2_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_sboxin_mux_inst_2_U1_AND1_U1 ( .A0_t (selSbox), .B0_t (MUX_sboxin_mux_inst_2_U1_X), .Z0_t (MUX_sboxin_mux_inst_2_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_sboxin_mux_inst_2_U1_XOR2_U1 ( .A0_t (MUX_sboxin_mux_inst_2_U1_Y), .B0_t (stateXORroundkey[2]), .Z0_t (sboxIn[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_sboxin_mux_inst_3_U1_XOR1_U1 ( .A0_t (stateXORroundkey[3]), .B0_t (keyRegKS[3]), .Z0_t (MUX_sboxin_mux_inst_3_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_sboxin_mux_inst_3_U1_AND1_U1 ( .A0_t (selSbox), .B0_t (MUX_sboxin_mux_inst_3_U1_X), .Z0_t (MUX_sboxin_mux_inst_3_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_sboxin_mux_inst_3_U1_XOR2_U1 ( .A0_t (MUX_sboxin_mux_inst_3_U1_Y), .B0_t (stateXORroundkey[3]), .Z0_t (sboxIn[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_serialIn_mux_inst_0_U1_XOR1_U1 ( .A0_t (sboxOut[0]), .B0_t (stateXORroundkey[0]), .Z0_t (MUX_serialIn_mux_inst_0_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_serialIn_mux_inst_0_U1_AND1_U1 ( .A0_t (intDone), .B0_t (MUX_serialIn_mux_inst_0_U1_X), .Z0_t (MUX_serialIn_mux_inst_0_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_serialIn_mux_inst_0_U1_XOR2_U1 ( .A0_t (MUX_serialIn_mux_inst_0_U1_Y), .B0_t (sboxOut[0]), .Z0_t (serialIn[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_serialIn_mux_inst_1_U1_XOR1_U1 ( .A0_t (sboxOut[1]), .B0_t (stateXORroundkey[1]), .Z0_t (MUX_serialIn_mux_inst_1_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_serialIn_mux_inst_1_U1_AND1_U1 ( .A0_t (intDone), .B0_t (MUX_serialIn_mux_inst_1_U1_X), .Z0_t (MUX_serialIn_mux_inst_1_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_serialIn_mux_inst_1_U1_XOR2_U1 ( .A0_t (MUX_serialIn_mux_inst_1_U1_Y), .B0_t (sboxOut[1]), .Z0_t (serialIn[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_serialIn_mux_inst_2_U1_XOR1_U1 ( .A0_t (sboxOut[2]), .B0_t (stateXORroundkey[2]), .Z0_t (MUX_serialIn_mux_inst_2_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_serialIn_mux_inst_2_U1_AND1_U1 ( .A0_t (intDone), .B0_t (MUX_serialIn_mux_inst_2_U1_X), .Z0_t (MUX_serialIn_mux_inst_2_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_serialIn_mux_inst_2_U1_XOR2_U1 ( .A0_t (MUX_serialIn_mux_inst_2_U1_Y), .B0_t (sboxOut[2]), .Z0_t (serialIn[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_serialIn_mux_inst_3_U1_XOR1_U1 ( .A0_t (sboxOut[3]), .B0_t (stateXORroundkey[3]), .Z0_t (MUX_serialIn_mux_inst_3_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_serialIn_mux_inst_3_U1_AND1_U1 ( .A0_t (intDone), .B0_t (MUX_serialIn_mux_inst_3_U1_X), .Z0_t (MUX_serialIn_mux_inst_3_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_serialIn_mux_inst_3_U1_XOR2_U1 ( .A0_t (MUX_serialIn_mux_inst_3_U1_Y), .B0_t (sboxOut[3]), .Z0_t (serialIn[3]) ) ;

    /* register cells */
endmodule
