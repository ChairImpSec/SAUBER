/* modified netlist. Source: module Keccak in file /mnt/c/Users/amirm/Desktop/Papers_in_progress/SAUBER/Design for our FPGA/8-Keccak-200_RoundBased_PortSerial/4-AGEMA/Keccak.v */
/* 0 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 1 register stage(s) in total */

module Keccak_SAUBER_Pipeline_d1 (InData, Reset, OutData, Ready);
    input [7:0] InData ;
    input Reset ;
    output [7:0] OutData ;
    output Ready ;
    wire IotaRC_7 ;
    wire IotaRC_3 ;
    wire n9 ;
    wire THETA_n200 ;
    wire THETA_n199 ;
    wire THETA_n198 ;
    wire THETA_n197 ;
    wire THETA_n196 ;
    wire THETA_n195 ;
    wire THETA_n194 ;
    wire THETA_n193 ;
    wire THETA_n192 ;
    wire THETA_n191 ;
    wire THETA_n190 ;
    wire THETA_n189 ;
    wire THETA_n188 ;
    wire THETA_n187 ;
    wire THETA_n186 ;
    wire THETA_n185 ;
    wire THETA_n184 ;
    wire THETA_n183 ;
    wire THETA_n182 ;
    wire THETA_n181 ;
    wire THETA_n180 ;
    wire THETA_n179 ;
    wire THETA_n178 ;
    wire THETA_n177 ;
    wire THETA_n176 ;
    wire THETA_n175 ;
    wire THETA_n174 ;
    wire THETA_n173 ;
    wire THETA_n172 ;
    wire THETA_n171 ;
    wire THETA_n170 ;
    wire THETA_n169 ;
    wire THETA_n168 ;
    wire THETA_n167 ;
    wire THETA_n166 ;
    wire THETA_n165 ;
    wire THETA_n164 ;
    wire THETA_n163 ;
    wire THETA_n162 ;
    wire THETA_n161 ;
    wire THETA_n160 ;
    wire THETA_n159 ;
    wire THETA_n158 ;
    wire THETA_n157 ;
    wire THETA_n156 ;
    wire THETA_n155 ;
    wire THETA_n154 ;
    wire THETA_n153 ;
    wire THETA_n152 ;
    wire THETA_n151 ;
    wire THETA_n150 ;
    wire THETA_n149 ;
    wire THETA_n148 ;
    wire THETA_n147 ;
    wire THETA_n146 ;
    wire THETA_n145 ;
    wire THETA_n144 ;
    wire THETA_n143 ;
    wire THETA_n142 ;
    wire THETA_n141 ;
    wire THETA_n140 ;
    wire THETA_n139 ;
    wire THETA_n138 ;
    wire THETA_n137 ;
    wire THETA_n136 ;
    wire THETA_n135 ;
    wire THETA_n134 ;
    wire THETA_n133 ;
    wire THETA_n132 ;
    wire THETA_n131 ;
    wire THETA_n130 ;
    wire THETA_n129 ;
    wire THETA_n128 ;
    wire THETA_n127 ;
    wire THETA_n126 ;
    wire THETA_n125 ;
    wire THETA_n124 ;
    wire THETA_n123 ;
    wire THETA_n122 ;
    wire THETA_n121 ;
    wire THETA_n120 ;
    wire THETA_n119 ;
    wire THETA_n118 ;
    wire THETA_n117 ;
    wire THETA_n116 ;
    wire THETA_n115 ;
    wire THETA_n114 ;
    wire THETA_n113 ;
    wire THETA_n112 ;
    wire THETA_n111 ;
    wire THETA_n110 ;
    wire THETA_n109 ;
    wire THETA_n108 ;
    wire THETA_n107 ;
    wire THETA_n106 ;
    wire THETA_n105 ;
    wire THETA_n104 ;
    wire THETA_n103 ;
    wire THETA_n102 ;
    wire THETA_n101 ;
    wire THETA_n100 ;
    wire THETA_n99 ;
    wire THETA_n98 ;
    wire THETA_n97 ;
    wire THETA_n96 ;
    wire THETA_n95 ;
    wire THETA_n94 ;
    wire THETA_n93 ;
    wire THETA_n92 ;
    wire THETA_n91 ;
    wire THETA_n90 ;
    wire THETA_n89 ;
    wire THETA_n88 ;
    wire THETA_n87 ;
    wire THETA_n86 ;
    wire THETA_n85 ;
    wire THETA_n84 ;
    wire THETA_n83 ;
    wire THETA_n82 ;
    wire THETA_n81 ;
    wire THETA_n80 ;
    wire THETA_n79 ;
    wire THETA_n78 ;
    wire THETA_n77 ;
    wire THETA_n76 ;
    wire THETA_n75 ;
    wire THETA_n74 ;
    wire THETA_n73 ;
    wire THETA_n72 ;
    wire THETA_n71 ;
    wire THETA_n70 ;
    wire THETA_n69 ;
    wire THETA_n68 ;
    wire THETA_n67 ;
    wire THETA_n66 ;
    wire THETA_n65 ;
    wire THETA_n64 ;
    wire THETA_n63 ;
    wire THETA_n62 ;
    wire THETA_n61 ;
    wire THETA_n60 ;
    wire THETA_n59 ;
    wire THETA_n58 ;
    wire THETA_n57 ;
    wire THETA_n56 ;
    wire THETA_n55 ;
    wire THETA_n54 ;
    wire THETA_n53 ;
    wire THETA_n52 ;
    wire THETA_n51 ;
    wire THETA_n50 ;
    wire THETA_n49 ;
    wire THETA_n48 ;
    wire THETA_n47 ;
    wire THETA_n46 ;
    wire THETA_n45 ;
    wire THETA_n44 ;
    wire THETA_n43 ;
    wire THETA_n42 ;
    wire THETA_n41 ;
    wire THETA_n40 ;
    wire THETA_n39 ;
    wire THETA_n38 ;
    wire THETA_n37 ;
    wire THETA_n36 ;
    wire THETA_n35 ;
    wire THETA_n34 ;
    wire THETA_n33 ;
    wire THETA_n32 ;
    wire THETA_n31 ;
    wire THETA_n30 ;
    wire THETA_n29 ;
    wire THETA_n28 ;
    wire THETA_n27 ;
    wire THETA_n26 ;
    wire THETA_n25 ;
    wire THETA_n24 ;
    wire THETA_n23 ;
    wire THETA_n22 ;
    wire THETA_n21 ;
    wire THETA_n20 ;
    wire THETA_n19 ;
    wire THETA_n18 ;
    wire THETA_n17 ;
    wire THETA_n16 ;
    wire THETA_n15 ;
    wire THETA_n14 ;
    wire THETA_n13 ;
    wire THETA_n12 ;
    wire THETA_n11 ;
    wire THETA_n10 ;
    wire THETA_n9 ;
    wire THETA_n8 ;
    wire THETA_n7 ;
    wire THETA_n6 ;
    wire THETA_n5 ;
    wire THETA_n4 ;
    wire THETA_n3 ;
    wire THETA_n2 ;
    wire THETA_n1 ;
    wire CHI_ChiOut_3 ;
    wire CHI_ChiOut_7 ;
    wire CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_1__GEN_ROWS_0__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_1__GEN_ROWS_0__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_1__GEN_ROWS_0__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_1__GEN_ROWS_0__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_1__GEN_ROWS_0__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_1__GEN_ROWS_1__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_1__GEN_ROWS_1__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_1__GEN_ROWS_1__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_1__GEN_ROWS_1__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_1__GEN_ROWS_1__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_1__GEN_ROWS_2__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_1__GEN_ROWS_2__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_1__GEN_ROWS_2__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_1__GEN_ROWS_2__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_1__GEN_ROWS_2__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_1__GEN_ROWS_3__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_1__GEN_ROWS_3__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_1__GEN_ROWS_3__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_1__GEN_ROWS_3__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_1__GEN_ROWS_3__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_1__GEN_ROWS_4__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_1__GEN_ROWS_4__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_1__GEN_ROWS_4__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_1__GEN_ROWS_4__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_1__GEN_ROWS_4__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_2__GEN_ROWS_0__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_2__GEN_ROWS_0__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_2__GEN_ROWS_0__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_2__GEN_ROWS_0__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_2__GEN_ROWS_0__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_2__GEN_ROWS_1__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_2__GEN_ROWS_1__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_2__GEN_ROWS_1__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_2__GEN_ROWS_1__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_2__GEN_ROWS_1__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_2__GEN_ROWS_2__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_2__GEN_ROWS_2__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_2__GEN_ROWS_2__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_2__GEN_ROWS_2__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_2__GEN_ROWS_2__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_2__GEN_ROWS_3__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_2__GEN_ROWS_3__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_2__GEN_ROWS_3__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_2__GEN_ROWS_3__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_2__GEN_ROWS_3__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_2__GEN_ROWS_4__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_2__GEN_ROWS_4__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_2__GEN_ROWS_4__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_2__GEN_ROWS_4__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_2__GEN_ROWS_4__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_3__GEN_ROWS_0__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_3__GEN_ROWS_0__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_3__GEN_ROWS_0__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_3__GEN_ROWS_0__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_3__GEN_ROWS_0__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_3__GEN_ROWS_1__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_3__GEN_ROWS_1__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_3__GEN_ROWS_1__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_3__GEN_ROWS_1__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_3__GEN_ROWS_1__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_3__GEN_ROWS_2__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_3__GEN_ROWS_2__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_3__GEN_ROWS_2__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_3__GEN_ROWS_2__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_3__GEN_ROWS_2__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_3__GEN_ROWS_3__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_3__GEN_ROWS_3__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_3__GEN_ROWS_3__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_3__GEN_ROWS_3__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_3__GEN_ROWS_3__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_3__GEN_ROWS_4__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_3__GEN_ROWS_4__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_3__GEN_ROWS_4__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_3__GEN_ROWS_4__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_3__GEN_ROWS_4__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_4__GEN_ROWS_0__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_4__GEN_ROWS_0__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_4__GEN_ROWS_0__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_4__GEN_ROWS_0__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_4__GEN_ROWS_0__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_4__GEN_ROWS_1__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_4__GEN_ROWS_1__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_4__GEN_ROWS_1__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_4__GEN_ROWS_1__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_4__GEN_ROWS_1__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_4__GEN_ROWS_2__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_4__GEN_ROWS_2__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_4__GEN_ROWS_2__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_4__GEN_ROWS_2__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_4__GEN_ROWS_2__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_4__GEN_ROWS_3__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_4__GEN_ROWS_3__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_4__GEN_ROWS_3__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_4__GEN_ROWS_3__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_4__GEN_ROWS_3__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_4__GEN_ROWS_4__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_4__GEN_ROWS_4__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_4__GEN_ROWS_4__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_4__GEN_ROWS_4__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_4__GEN_ROWS_4__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_5__GEN_ROWS_0__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_5__GEN_ROWS_0__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_5__GEN_ROWS_0__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_5__GEN_ROWS_0__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_5__GEN_ROWS_0__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_5__GEN_ROWS_1__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_5__GEN_ROWS_1__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_5__GEN_ROWS_1__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_5__GEN_ROWS_1__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_5__GEN_ROWS_1__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_5__GEN_ROWS_2__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_5__GEN_ROWS_2__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_5__GEN_ROWS_2__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_5__GEN_ROWS_2__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_5__GEN_ROWS_2__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_5__GEN_ROWS_3__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_5__GEN_ROWS_3__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_5__GEN_ROWS_3__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_5__GEN_ROWS_3__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_5__GEN_ROWS_3__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_5__GEN_ROWS_4__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_5__GEN_ROWS_4__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_5__GEN_ROWS_4__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_5__GEN_ROWS_4__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_5__GEN_ROWS_4__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_6__GEN_ROWS_0__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_6__GEN_ROWS_0__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_6__GEN_ROWS_0__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_6__GEN_ROWS_0__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_6__GEN_ROWS_0__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_6__GEN_ROWS_1__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_6__GEN_ROWS_1__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_6__GEN_ROWS_1__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_6__GEN_ROWS_1__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_6__GEN_ROWS_1__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_6__GEN_ROWS_2__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_6__GEN_ROWS_2__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_6__GEN_ROWS_2__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_6__GEN_ROWS_2__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_6__GEN_ROWS_2__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_6__GEN_ROWS_3__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_6__GEN_ROWS_3__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_6__GEN_ROWS_3__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_6__GEN_ROWS_3__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_6__GEN_ROWS_3__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_6__GEN_ROWS_4__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_6__GEN_ROWS_4__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_6__GEN_ROWS_4__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_6__GEN_ROWS_4__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_6__GEN_ROWS_4__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_7__GEN_ROWS_0__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_7__GEN_ROWS_0__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_7__GEN_ROWS_0__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_7__GEN_ROWS_0__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_7__GEN_ROWS_0__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_7__GEN_ROWS_1__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_7__GEN_ROWS_1__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_7__GEN_ROWS_1__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_7__GEN_ROWS_1__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_7__GEN_ROWS_1__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_7__GEN_ROWS_2__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_7__GEN_ROWS_2__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_7__GEN_ROWS_2__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_7__GEN_ROWS_2__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_7__GEN_ROWS_2__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_7__GEN_ROWS_3__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_7__GEN_ROWS_3__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_7__GEN_ROWS_3__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_7__GEN_ROWS_3__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_7__GEN_ROWS_3__sbox_and_xor_inst_e_nxy ;
    wire CHI_GEN_SLICES_7__GEN_ROWS_4__sbox_and_xor_inst_a_nxy ;
    wire CHI_GEN_SLICES_7__GEN_ROWS_4__sbox_and_xor_inst_b_nxy ;
    wire CHI_GEN_SLICES_7__GEN_ROWS_4__sbox_and_xor_inst_c_nxy ;
    wire CHI_GEN_SLICES_7__GEN_ROWS_4__sbox_and_xor_inst_d_nxy ;
    wire CHI_GEN_SLICES_7__GEN_ROWS_4__sbox_and_xor_inst_e_nxy ;
    wire KECCAK_CONTROL_n47 ;
    wire KECCAK_CONTROL_n45 ;
    wire KECCAK_CONTROL_n44 ;
    wire KECCAK_CONTROL_n43 ;
    wire KECCAK_CONTROL_n34 ;
    wire KECCAK_CONTROL_n33 ;
    wire KECCAK_CONTROL_n32 ;
    wire KECCAK_CONTROL_n30 ;
    wire KECCAK_CONTROL_n29 ;
    wire KECCAK_CONTROL_n28 ;
    wire KECCAK_CONTROL_n27 ;
    wire KECCAK_CONTROL_n25 ;
    wire KECCAK_CONTROL_n23 ;
    wire KECCAK_CONTROL_n22 ;
    wire KECCAK_CONTROL_n21 ;
    wire KECCAK_CONTROL_n20 ;
    wire KECCAK_CONTROL_n19 ;
    wire KECCAK_CONTROL_n18 ;
    wire KECCAK_CONTROL_n17 ;
    wire KECCAK_CONTROL_n16 ;
    wire KECCAK_CONTROL_n15 ;
    wire KECCAK_CONTROL_n14 ;
    wire KECCAK_CONTROL_n13 ;
    wire KECCAK_CONTROL_n11 ;
    wire KECCAK_CONTROL_n10 ;
    wire KECCAK_CONTROL_n8 ;
    wire KECCAK_CONTROL_CtrlStatexDP_reg_1__Q ;
    wire KECCAK_CONTROL_RoundCountLastxDP_reg_Q ;
    wire KECCAK_CONTROL_RC_GEN_n28 ;
    wire KECCAK_CONTROL_RC_GEN_n27 ;
    wire KECCAK_CONTROL_RC_GEN_n26 ;
    wire KECCAK_CONTROL_RC_GEN_n25 ;
    wire KECCAK_CONTROL_RC_GEN_n22 ;
    wire KECCAK_CONTROL_RC_GEN_n19 ;
    wire KECCAK_CONTROL_RC_GEN_n18 ;
    wire KECCAK_CONTROL_RC_GEN_n17 ;
    wire KECCAK_CONTROL_RC_GEN_n15 ;
    wire KECCAK_CONTROL_RC_GEN_n14 ;
    wire KECCAK_CONTROL_RC_GEN_n13 ;
    wire KECCAK_CONTROL_RC_GEN_n12 ;
    wire KECCAK_CONTROL_RC_GEN_n11 ;
    wire KECCAK_CONTROL_RC_GEN_n9 ;
    wire KECCAK_CONTROL_RC_GEN_n8 ;
    wire KECCAK_CONTROL_RC_GEN_n6 ;
    wire KECCAK_CONTROL_RC_GEN_n5 ;
    wire KECCAK_CONTROL_RC_GEN_n4 ;
    wire KECCAK_CONTROL_RC_GEN_n3 ;
    wire KECCAK_CONTROL_RC_GEN_n2 ;
    wire KECCAK_CONTROL_RC_GEN_n30 ;
    wire KECCAK_CONTROL_RC_GEN_n31 ;
    wire KECCAK_CONTROL_RC_GEN_n23 ;
    wire KECCAK_CONTROL_RC_GEN_n24 ;
    wire KECCAK_CONTROL_RC_GEN_n20 ;
    wire KECCAK_CONTROL_RC_GEN_n21 ;
    wire KECCAK_CONTROL_RC_GEN_U25_Y ;
    wire KECCAK_CONTROL_RC_GEN_U25_X ;
    wire KECCAK_CONTROL_RC_GEN_U28_Y ;
    wire KECCAK_CONTROL_RC_GEN_U28_X ;
    wire KECCAK_CONTROL_RC_GEN_U32_Y ;
    wire KECCAK_CONTROL_RC_GEN_U32_X ;
    wire U810_Y ;
    wire U810_X ;
    wire U812_Y ;
    wire U812_X ;
    wire U814_Y ;
    wire U814_X ;
    wire U816_Y ;
    wire U816_X ;
    wire U817_Y ;
    wire U817_X ;
    wire U818_Y ;
    wire U818_X ;
    wire U820_Y ;
    wire U820_X ;
    wire U821_Y ;
    wire U821_X ;
    wire U822_Y ;
    wire U822_X ;
    wire U823_Y ;
    wire U823_X ;
    wire U824_Y ;
    wire U824_X ;
    wire U825_Y ;
    wire U825_X ;
    wire U827_Y ;
    wire U827_X ;
    wire U828_Y ;
    wire U828_X ;
    wire U830_Y ;
    wire U830_X ;
    wire U831_Y ;
    wire U831_X ;
    wire U832_Y ;
    wire U832_X ;
    wire U833_Y ;
    wire U833_X ;
    wire U834_Y ;
    wire U834_X ;
    wire U835_Y ;
    wire U835_X ;
    wire U836_Y ;
    wire U836_X ;
    wire U837_Y ;
    wire U837_X ;
    wire U838_Y ;
    wire U838_X ;
    wire U839_Y ;
    wire U839_X ;
    wire U841_Y ;
    wire U841_X ;
    wire U842_Y ;
    wire U842_X ;
    wire U843_Y ;
    wire U843_X ;
    wire U844_Y ;
    wire U844_X ;
    wire U845_Y ;
    wire U845_X ;
    wire U846_Y ;
    wire U846_X ;
    wire U847_Y ;
    wire U847_X ;
    wire U848_Y ;
    wire U848_X ;
    wire U849_Y ;
    wire U849_X ;
    wire U850_Y ;
    wire U850_X ;
    wire U851_Y ;
    wire U851_X ;
    wire U852_Y ;
    wire U852_X ;
    wire U853_Y ;
    wire U853_X ;
    wire U854_Y ;
    wire U854_X ;
    wire U855_Y ;
    wire U855_X ;
    wire U856_Y ;
    wire U856_X ;
    wire U857_Y ;
    wire U857_X ;
    wire U858_Y ;
    wire U858_X ;
    wire U859_Y ;
    wire U859_X ;
    wire U860_Y ;
    wire U860_X ;
    wire U861_Y ;
    wire U861_X ;
    wire U862_Y ;
    wire U862_X ;
    wire U863_Y ;
    wire U863_X ;
    wire U864_Y ;
    wire U864_X ;
    wire U865_Y ;
    wire U865_X ;
    wire U866_Y ;
    wire U866_X ;
    wire U867_Y ;
    wire U867_X ;
    wire U868_Y ;
    wire U868_X ;
    wire U869_Y ;
    wire U869_X ;
    wire U870_Y ;
    wire U870_X ;
    wire U871_Y ;
    wire U871_X ;
    wire U872_Y ;
    wire U872_X ;
    wire U873_Y ;
    wire U873_X ;
    wire U874_Y ;
    wire U874_X ;
    wire U875_Y ;
    wire U875_X ;
    wire U876_Y ;
    wire U876_X ;
    wire U877_Y ;
    wire U877_X ;
    wire U878_Y ;
    wire U878_X ;
    wire U879_Y ;
    wire U879_X ;
    wire U880_Y ;
    wire U880_X ;
    wire U881_Y ;
    wire U881_X ;
    wire U882_Y ;
    wire U882_X ;
    wire U883_Y ;
    wire U883_X ;
    wire U884_Y ;
    wire U884_X ;
    wire U885_Y ;
    wire U885_X ;
    wire U886_Y ;
    wire U886_X ;
    wire U887_Y ;
    wire U887_X ;
    wire U888_Y ;
    wire U888_X ;
    wire U889_Y ;
    wire U889_X ;
    wire U890_Y ;
    wire U890_X ;
    wire U891_Y ;
    wire U891_X ;
    wire U892_Y ;
    wire U892_X ;
    wire U893_Y ;
    wire U893_X ;
    wire U894_Y ;
    wire U894_X ;
    wire U895_Y ;
    wire U895_X ;
    wire U896_Y ;
    wire U896_X ;
    wire U897_Y ;
    wire U897_X ;
    wire U898_Y ;
    wire U898_X ;
    wire U899_Y ;
    wire U899_X ;
    wire U900_Y ;
    wire U900_X ;
    wire U901_Y ;
    wire U901_X ;
    wire U902_Y ;
    wire U902_X ;
    wire U903_Y ;
    wire U903_X ;
    wire U904_Y ;
    wire U904_X ;
    wire U905_Y ;
    wire U905_X ;
    wire U906_Y ;
    wire U906_X ;
    wire U907_Y ;
    wire U907_X ;
    wire U908_Y ;
    wire U908_X ;
    wire U909_Y ;
    wire U909_X ;
    wire U910_Y ;
    wire U910_X ;
    wire U911_Y ;
    wire U911_X ;
    wire U912_Y ;
    wire U912_X ;
    wire U913_Y ;
    wire U913_X ;
    wire U914_Y ;
    wire U914_X ;
    wire U915_Y ;
    wire U915_X ;
    wire U916_Y ;
    wire U916_X ;
    wire U917_Y ;
    wire U917_X ;
    wire U918_Y ;
    wire U918_X ;
    wire U919_Y ;
    wire U919_X ;
    wire U920_Y ;
    wire U920_X ;
    wire U921_Y ;
    wire U921_X ;
    wire U922_Y ;
    wire U922_X ;
    wire U923_Y ;
    wire U923_X ;
    wire U924_Y ;
    wire U924_X ;
    wire U925_Y ;
    wire U925_X ;
    wire U926_Y ;
    wire U926_X ;
    wire U927_Y ;
    wire U927_X ;
    wire U928_Y ;
    wire U928_X ;
    wire U929_Y ;
    wire U929_X ;
    wire U930_Y ;
    wire U930_X ;
    wire U931_Y ;
    wire U931_X ;
    wire U932_Y ;
    wire U932_X ;
    wire U933_Y ;
    wire U933_X ;
    wire U934_Y ;
    wire U934_X ;
    wire U935_Y ;
    wire U935_X ;
    wire U936_Y ;
    wire U936_X ;
    wire U937_Y ;
    wire U937_X ;
    wire U938_Y ;
    wire U938_X ;
    wire U939_Y ;
    wire U939_X ;
    wire U940_Y ;
    wire U940_X ;
    wire U941_Y ;
    wire U941_X ;
    wire U942_Y ;
    wire U942_X ;
    wire U943_Y ;
    wire U943_X ;
    wire U944_Y ;
    wire U944_X ;
    wire U945_Y ;
    wire U945_X ;
    wire U946_Y ;
    wire U946_X ;
    wire U947_Y ;
    wire U947_X ;
    wire U948_Y ;
    wire U948_X ;
    wire U949_Y ;
    wire U949_X ;
    wire U950_Y ;
    wire U950_X ;
    wire U951_Y ;
    wire U951_X ;
    wire U952_Y ;
    wire U952_X ;
    wire U953_Y ;
    wire U953_X ;
    wire U954_Y ;
    wire U954_X ;
    wire U955_Y ;
    wire U955_X ;
    wire U956_Y ;
    wire U956_X ;
    wire U957_Y ;
    wire U957_X ;
    wire U958_Y ;
    wire U958_X ;
    wire U959_Y ;
    wire U959_X ;
    wire U960_Y ;
    wire U960_X ;
    wire U961_Y ;
    wire U961_X ;
    wire U962_Y ;
    wire U962_X ;
    wire U963_Y ;
    wire U963_X ;
    wire U964_Y ;
    wire U964_X ;
    wire U965_Y ;
    wire U965_X ;
    wire U966_Y ;
    wire U966_X ;
    wire U967_Y ;
    wire U967_X ;
    wire U968_Y ;
    wire U968_X ;
    wire U969_Y ;
    wire U969_X ;
    wire U970_Y ;
    wire U970_X ;
    wire U971_Y ;
    wire U971_X ;
    wire U972_Y ;
    wire U972_X ;
    wire U973_Y ;
    wire U973_X ;
    wire U974_Y ;
    wire U974_X ;
    wire U975_Y ;
    wire U975_X ;
    wire U976_Y ;
    wire U976_X ;
    wire U977_Y ;
    wire U977_X ;
    wire U978_Y ;
    wire U978_X ;
    wire U979_Y ;
    wire U979_X ;
    wire U980_Y ;
    wire U980_X ;
    wire U981_Y ;
    wire U981_X ;
    wire U982_Y ;
    wire U982_X ;
    wire U983_Y ;
    wire U983_X ;
    wire U984_Y ;
    wire U984_X ;
    wire U985_Y ;
    wire U985_X ;
    wire U986_Y ;
    wire U986_X ;
    wire U987_Y ;
    wire U987_X ;
    wire U988_Y ;
    wire U988_X ;
    wire U989_Y ;
    wire U989_X ;
    wire U990_Y ;
    wire U990_X ;
    wire U991_Y ;
    wire U991_X ;
    wire U992_Y ;
    wire U992_X ;
    wire U993_Y ;
    wire U993_X ;
    wire U994_Y ;
    wire U994_X ;
    wire U995_Y ;
    wire U995_X ;
    wire U996_Y ;
    wire U996_X ;
    wire U997_Y ;
    wire U997_X ;
    wire U998_Y ;
    wire U998_X ;
    wire U999_Y ;
    wire U999_X ;
    wire U1000_Y ;
    wire U1000_X ;
    wire U1001_Y ;
    wire U1001_X ;
    wire U1002_Y ;
    wire U1002_X ;
    wire U1003_Y ;
    wire U1003_X ;
    wire U1004_Y ;
    wire U1004_X ;
    wire U1005_Y ;
    wire U1005_X ;
    wire U1006_Y ;
    wire U1006_X ;
    wire U1007_Y ;
    wire U1007_X ;
    wire U1008_Y ;
    wire U1008_X ;
    wire U1009_Y ;
    wire U1009_X ;
    wire U1010_Y ;
    wire U1010_X ;
    wire U1011_Y ;
    wire U1011_X ;
    wire U1012_Y ;
    wire U1012_X ;
    wire U1013_Y ;
    wire U1013_X ;
    wire U1014_Y ;
    wire U1014_X ;
    wire U1015_Y ;
    wire U1015_X ;
    wire U1016_Y ;
    wire U1016_X ;
    wire [199:8] StateOut ;
    wire [199:0] StateFromRhoPi ;
    wire [199:0] StateFromChi ;
    wire [1:0] IotaRC ;
    wire [1:0] CHI_ChiOut ;
    wire [4:0] KECCAK_CONTROL_RoundCountxDP ;
    wire [2:0] KECCAK_CONTROL_CtrlStatexDP ;

    /* cells in depth 0 */
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) U5 ( .A0_t (Reset), .B0_t (Ready), .Z0_t (n9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U400 ( .A0_t (StateOut[199]), .B0_t (THETA_n200), .Z0_t (StateFromRhoPi[165]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U399 ( .A0_t (StateOut[191]), .B0_t (THETA_n200), .Z0_t (StateFromRhoPi[143]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U398 ( .A0_t (StateOut[183]), .B0_t (THETA_n200), .Z0_t (StateFromRhoPi[118]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U397 ( .A0_t (StateOut[175]), .B0_t (THETA_n200), .Z0_t (StateFromRhoPi[51]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U396 ( .A0_t (StateOut[167]), .B0_t (THETA_n200), .Z0_t (StateFromRhoPi[26]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U395 ( .A0_t (THETA_n199), .B0_t (THETA_n198), .Z0_t (THETA_n200) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U394 ( .A0_t (StateOut[78]), .B0_t (THETA_n197), .Z0_t (StateFromRhoPi[192]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U393 ( .A0_t (StateOut[70]), .B0_t (THETA_n197), .Z0_t (StateFromRhoPi[131]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U392 ( .A0_t (StateOut[62]), .B0_t (THETA_n197), .Z0_t (StateFromRhoPi[104]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U391 ( .A0_t (StateOut[54]), .B0_t (THETA_n197), .Z0_t (StateFromRhoPi[42]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U390 ( .A0_t (StateOut[46]), .B0_t (THETA_n197), .Z0_t (StateFromRhoPi[23]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U389 ( .A0_t (THETA_n196), .B0_t (THETA_n198), .Z0_t (THETA_n197) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U388 ( .A0_t (OutData[6]), .B0_t (THETA_n195), .Z0_t (THETA_n198) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U387 ( .A0_t (THETA_n194), .B0_t (THETA_n193), .Z0_t (THETA_n195) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U386 ( .A0_t (StateOut[14]), .B0_t (StateOut[22]), .Z0_t (THETA_n193) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U385 ( .A0_t (StateOut[38]), .B0_t (StateOut[30]), .Z0_t (THETA_n194) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U384 ( .A0_t (StateOut[112]), .B0_t (THETA_n192), .Z0_t (StateFromRhoPi[173]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U383 ( .A0_t (StateOut[104]), .B0_t (THETA_n192), .Z0_t (StateFromRhoPi[151]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U382 ( .A0_t (StateOut[96]), .B0_t (THETA_n192), .Z0_t (StateFromRhoPi[83]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U381 ( .A0_t (StateOut[88]), .B0_t (THETA_n192), .Z0_t (StateFromRhoPi[62]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U380 ( .A0_t (StateOut[80]), .B0_t (THETA_n192), .Z0_t (StateFromRhoPi[38]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U379 ( .A0_t (THETA_n191), .B0_t (THETA_n199), .Z0_t (THETA_n192) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U378 ( .A0_t (StateOut[127]), .B0_t (THETA_n190), .Z0_t (THETA_n199) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U377 ( .A0_t (THETA_n189), .B0_t (THETA_n188), .Z0_t (THETA_n190) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U376 ( .A0_t (StateOut[135]), .B0_t (StateOut[143]), .Z0_t (THETA_n188) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U375 ( .A0_t (StateOut[159]), .B0_t (StateOut[151]), .Z0_t (THETA_n189) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U374 ( .A0_t (StateOut[198]), .B0_t (THETA_n187), .Z0_t (StateFromRhoPi[164]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U373 ( .A0_t (StateOut[190]), .B0_t (THETA_n187), .Z0_t (StateFromRhoPi[142]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U372 ( .A0_t (StateOut[182]), .B0_t (THETA_n187), .Z0_t (StateFromRhoPi[117]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U371 ( .A0_t (StateOut[174]), .B0_t (THETA_n187), .Z0_t (StateFromRhoPi[50]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U370 ( .A0_t (StateOut[166]), .B0_t (THETA_n187), .Z0_t (StateFromRhoPi[25]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U369 ( .A0_t (THETA_n186), .B0_t (THETA_n185), .Z0_t (THETA_n187) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U368 ( .A0_t (StateOut[119]), .B0_t (THETA_n184), .Z0_t (StateFromRhoPi[172]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U367 ( .A0_t (StateOut[111]), .B0_t (THETA_n184), .Z0_t (StateFromRhoPi[150]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U366 ( .A0_t (StateOut[103]), .B0_t (THETA_n184), .Z0_t (StateFromRhoPi[82]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U365 ( .A0_t (StateOut[95]), .B0_t (THETA_n184), .Z0_t (StateFromRhoPi[61]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U364 ( .A0_t (StateOut[87]), .B0_t (THETA_n184), .Z0_t (StateFromRhoPi[37]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U363 ( .A0_t (THETA_n183), .B0_t (THETA_n185), .Z0_t (THETA_n184) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U362 ( .A0_t (StateOut[126]), .B0_t (THETA_n182), .Z0_t (THETA_n185) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U361 ( .A0_t (THETA_n181), .B0_t (THETA_n180), .Z0_t (THETA_n182) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U360 ( .A0_t (StateOut[134]), .B0_t (StateOut[142]), .Z0_t (THETA_n180) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U359 ( .A0_t (StateOut[158]), .B0_t (StateOut[150]), .Z0_t (THETA_n181) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U358 ( .A0_t (StateOut[196]), .B0_t (THETA_n179), .Z0_t (StateFromRhoPi[162]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U357 ( .A0_t (StateOut[188]), .B0_t (THETA_n179), .Z0_t (StateFromRhoPi[140]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U356 ( .A0_t (StateOut[180]), .B0_t (THETA_n179), .Z0_t (StateFromRhoPi[115]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U355 ( .A0_t (StateOut[172]), .B0_t (THETA_n179), .Z0_t (StateFromRhoPi[48]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U354 ( .A0_t (StateOut[164]), .B0_t (THETA_n179), .Z0_t (StateFromRhoPi[31]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U353 ( .A0_t (THETA_n178), .B0_t (THETA_n177), .Z0_t (THETA_n179) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U352 ( .A0_t (StateOut[75]), .B0_t (THETA_n176), .Z0_t (StateFromRhoPi[197]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U351 ( .A0_t (StateOut[67]), .B0_t (THETA_n176), .Z0_t (StateFromRhoPi[128]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U350 ( .A0_t (StateOut[59]), .B0_t (THETA_n176), .Z0_t (StateFromRhoPi[109]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U349 ( .A0_t (StateOut[51]), .B0_t (THETA_n176), .Z0_t (StateFromRhoPi[47]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U348 ( .A0_t (StateOut[43]), .B0_t (THETA_n176), .Z0_t (StateFromRhoPi[20]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U347 ( .A0_t (THETA_n175), .B0_t (THETA_n177), .Z0_t (THETA_n176) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U346 ( .A0_t (OutData[3]), .B0_t (THETA_n174), .Z0_t (THETA_n177) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U345 ( .A0_t (THETA_n173), .B0_t (THETA_n172), .Z0_t (THETA_n174) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U344 ( .A0_t (StateOut[11]), .B0_t (StateOut[19]), .Z0_t (THETA_n172) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U343 ( .A0_t (StateOut[35]), .B0_t (StateOut[27]), .Z0_t (THETA_n173) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U342 ( .A0_t (StateOut[193]), .B0_t (THETA_n171), .Z0_t (StateFromRhoPi[167]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U341 ( .A0_t (StateOut[185]), .B0_t (THETA_n171), .Z0_t (StateFromRhoPi[137]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U340 ( .A0_t (StateOut[177]), .B0_t (THETA_n171), .Z0_t (StateFromRhoPi[112]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U339 ( .A0_t (StateOut[169]), .B0_t (THETA_n171), .Z0_t (StateFromRhoPi[53]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U338 ( .A0_t (StateOut[161]), .B0_t (THETA_n171), .Z0_t (StateFromRhoPi[28]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U337 ( .A0_t (THETA_n170), .B0_t (THETA_n169), .Z0_t (THETA_n171) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U336 ( .A0_t (StateOut[72]), .B0_t (THETA_n168), .Z0_t (StateFromRhoPi[194]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U335 ( .A0_t (StateOut[64]), .B0_t (THETA_n168), .Z0_t (StateFromRhoPi[133]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U334 ( .A0_t (StateOut[56]), .B0_t (THETA_n168), .Z0_t (StateFromRhoPi[106]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U333 ( .A0_t (StateOut[48]), .B0_t (THETA_n168), .Z0_t (StateFromRhoPi[44]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U332 ( .A0_t (StateOut[40]), .B0_t (THETA_n168), .Z0_t (StateFromRhoPi[17]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U331 ( .A0_t (THETA_n167), .B0_t (THETA_n169), .Z0_t (THETA_n168) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U330 ( .A0_t (OutData[0]), .B0_t (THETA_n166), .Z0_t (THETA_n169) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U329 ( .A0_t (THETA_n165), .B0_t (THETA_n164), .Z0_t (THETA_n166) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U328 ( .A0_t (StateOut[8]), .B0_t (StateOut[16]), .Z0_t (THETA_n164) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U327 ( .A0_t (StateOut[32]), .B0_t (StateOut[24]), .Z0_t (THETA_n165) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U326 ( .A0_t (StateOut[154]), .B0_t (THETA_n163), .Z0_t (StateFromRhoPi[186]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U325 ( .A0_t (StateOut[146]), .B0_t (THETA_n163), .Z0_t (StateFromRhoPi[127]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U324 ( .A0_t (StateOut[138]), .B0_t (THETA_n163), .Z0_t (StateFromRhoPi[99]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U323 ( .A0_t (StateOut[130]), .B0_t (THETA_n163), .Z0_t (StateFromRhoPi[73]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U322 ( .A0_t (StateOut[122]), .B0_t (THETA_n163), .Z0_t (StateFromRhoPi[14]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U321 ( .A0_t (THETA_n162), .B0_t (THETA_n175), .Z0_t (THETA_n163) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U320 ( .A0_t (StateOut[82]), .B0_t (THETA_n161), .Z0_t (THETA_n175) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U319 ( .A0_t (THETA_n160), .B0_t (THETA_n159), .Z0_t (THETA_n161) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U318 ( .A0_t (StateOut[90]), .B0_t (StateOut[98]), .Z0_t (THETA_n159) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U317 ( .A0_t (StateOut[114]), .B0_t (StateOut[106]), .Z0_t (THETA_n160) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U316 ( .A0_t (StateOut[33]), .B0_t (THETA_n158), .Z0_t (StateFromRhoPi[179]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U315 ( .A0_t (StateOut[25]), .B0_t (THETA_n158), .Z0_t (StateFromRhoPi[154]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U314 ( .A0_t (StateOut[17]), .B0_t (THETA_n158), .Z0_t (StateFromRhoPi[92]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U313 ( .A0_t (StateOut[9]), .B0_t (THETA_n158), .Z0_t (StateFromRhoPi[69]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U312 ( .A0_t (OutData[1]), .B0_t (THETA_n158), .Z0_t (StateFromRhoPi[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U311 ( .A0_t (THETA_n191), .B0_t (THETA_n162), .Z0_t (THETA_n158) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U310 ( .A0_t (StateOut[177]), .B0_t (THETA_n157), .Z0_t (THETA_n162) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U309 ( .A0_t (THETA_n156), .B0_t (THETA_n155), .Z0_t (THETA_n157) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U308 ( .A0_t (StateOut[169]), .B0_t (StateOut[161]), .Z0_t (THETA_n155) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U307 ( .A0_t (StateOut[185]), .B0_t (StateOut[193]), .Z0_t (THETA_n156) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U306 ( .A0_t (StateOut[64]), .B0_t (THETA_n154), .Z0_t (THETA_n191) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U305 ( .A0_t (THETA_n153), .B0_t (THETA_n152), .Z0_t (THETA_n154) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U304 ( .A0_t (StateOut[48]), .B0_t (StateOut[40]), .Z0_t (THETA_n152) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U303 ( .A0_t (StateOut[72]), .B0_t (StateOut[56]), .Z0_t (THETA_n153) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U302 ( .A0_t (StateOut[114]), .B0_t (THETA_n151), .Z0_t (StateFromRhoPi[175]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U301 ( .A0_t (StateOut[106]), .B0_t (THETA_n151), .Z0_t (StateFromRhoPi[145]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U300 ( .A0_t (StateOut[98]), .B0_t (THETA_n151), .Z0_t (StateFromRhoPi[85]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U299 ( .A0_t (StateOut[90]), .B0_t (THETA_n151), .Z0_t (StateFromRhoPi[56]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U298 ( .A0_t (StateOut[82]), .B0_t (THETA_n151), .Z0_t (StateFromRhoPi[32]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U297 ( .A0_t (THETA_n150), .B0_t (THETA_n170), .Z0_t (THETA_n151) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U296 ( .A0_t (StateOut[121]), .B0_t (THETA_n149), .Z0_t (THETA_n170) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U295 ( .A0_t (THETA_n148), .B0_t (THETA_n147), .Z0_t (THETA_n149) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U294 ( .A0_t (StateOut[129]), .B0_t (StateOut[137]), .Z0_t (THETA_n147) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U293 ( .A0_t (StateOut[153]), .B0_t (StateOut[145]), .Z0_t (THETA_n148) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U292 ( .A0_t (StateOut[153]), .B0_t (THETA_n146), .Z0_t (StateFromRhoPi[185]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U291 ( .A0_t (StateOut[145]), .B0_t (THETA_n146), .Z0_t (StateFromRhoPi[126]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U290 ( .A0_t (StateOut[137]), .B0_t (THETA_n146), .Z0_t (StateFromRhoPi[98]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U289 ( .A0_t (StateOut[129]), .B0_t (THETA_n146), .Z0_t (StateFromRhoPi[72]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U288 ( .A0_t (StateOut[121]), .B0_t (THETA_n146), .Z0_t (StateFromRhoPi[13]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U287 ( .A0_t (THETA_n145), .B0_t (THETA_n144), .Z0_t (THETA_n146) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U286 ( .A0_t (StateOut[74]), .B0_t (THETA_n143), .Z0_t (StateFromRhoPi[196]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U285 ( .A0_t (StateOut[66]), .B0_t (THETA_n143), .Z0_t (StateFromRhoPi[135]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U284 ( .A0_t (StateOut[58]), .B0_t (THETA_n143), .Z0_t (StateFromRhoPi[108]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U283 ( .A0_t (StateOut[50]), .B0_t (THETA_n143), .Z0_t (StateFromRhoPi[46]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U282 ( .A0_t (StateOut[42]), .B0_t (THETA_n143), .Z0_t (StateFromRhoPi[19]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U281 ( .A0_t (THETA_n142), .B0_t (THETA_n144), .Z0_t (THETA_n143) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U280 ( .A0_t (StateOut[81]), .B0_t (THETA_n141), .Z0_t (THETA_n144) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U279 ( .A0_t (THETA_n140), .B0_t (THETA_n139), .Z0_t (THETA_n141) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U278 ( .A0_t (StateOut[89]), .B0_t (StateOut[97]), .Z0_t (THETA_n139) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U277 ( .A0_t (StateOut[113]), .B0_t (StateOut[105]), .Z0_t (THETA_n140) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U276 ( .A0_t (StateOut[32]), .B0_t (THETA_n138), .Z0_t (StateFromRhoPi[178]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U275 ( .A0_t (StateOut[24]), .B0_t (THETA_n138), .Z0_t (StateFromRhoPi[153]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U274 ( .A0_t (StateOut[16]), .B0_t (THETA_n138), .Z0_t (StateFromRhoPi[91]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U273 ( .A0_t (StateOut[8]), .B0_t (THETA_n138), .Z0_t (StateFromRhoPi[68]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U272 ( .A0_t (OutData[0]), .B0_t (THETA_n138), .Z0_t (StateFromRhoPi[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U271 ( .A0_t (THETA_n183), .B0_t (THETA_n145), .Z0_t (THETA_n138) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U270 ( .A0_t (StateOut[160]), .B0_t (THETA_n137), .Z0_t (THETA_n145) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U269 ( .A0_t (THETA_n136), .B0_t (THETA_n135), .Z0_t (THETA_n137) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U268 ( .A0_t (StateOut[168]), .B0_t (StateOut[176]), .Z0_t (THETA_n135) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U267 ( .A0_t (StateOut[192]), .B0_t (StateOut[184]), .Z0_t (THETA_n136) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U266 ( .A0_t (StateOut[47]), .B0_t (THETA_n134), .Z0_t (THETA_n183) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U265 ( .A0_t (THETA_n133), .B0_t (THETA_n132), .Z0_t (THETA_n134) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U264 ( .A0_t (StateOut[55]), .B0_t (StateOut[63]), .Z0_t (THETA_n132) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U263 ( .A0_t (StateOut[79]), .B0_t (StateOut[71]), .Z0_t (THETA_n133) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U262 ( .A0_t (StateOut[192]), .B0_t (THETA_n131), .Z0_t (StateFromRhoPi[166]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U261 ( .A0_t (StateOut[184]), .B0_t (THETA_n131), .Z0_t (StateFromRhoPi[136]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U260 ( .A0_t (StateOut[176]), .B0_t (THETA_n131), .Z0_t (StateFromRhoPi[119]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U259 ( .A0_t (StateOut[168]), .B0_t (THETA_n131), .Z0_t (StateFromRhoPi[52]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U258 ( .A0_t (StateOut[160]), .B0_t (THETA_n131), .Z0_t (StateFromRhoPi[27]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U257 ( .A0_t (THETA_n130), .B0_t (THETA_n129), .Z0_t (THETA_n131) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U256 ( .A0_t (StateOut[79]), .B0_t (THETA_n128), .Z0_t (StateFromRhoPi[193]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U255 ( .A0_t (StateOut[71]), .B0_t (THETA_n128), .Z0_t (StateFromRhoPi[132]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U254 ( .A0_t (StateOut[63]), .B0_t (THETA_n128), .Z0_t (StateFromRhoPi[105]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U253 ( .A0_t (StateOut[55]), .B0_t (THETA_n128), .Z0_t (StateFromRhoPi[43]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U252 ( .A0_t (StateOut[47]), .B0_t (THETA_n128), .Z0_t (StateFromRhoPi[16]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U251 ( .A0_t (THETA_n127), .B0_t (THETA_n129), .Z0_t (THETA_n128) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U250 ( .A0_t (OutData[7]), .B0_t (THETA_n126), .Z0_t (THETA_n129) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U249 ( .A0_t (THETA_n125), .B0_t (THETA_n124), .Z0_t (THETA_n126) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U248 ( .A0_t (StateOut[15]), .B0_t (StateOut[23]), .Z0_t (THETA_n124) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U247 ( .A0_t (StateOut[39]), .B0_t (StateOut[31]), .Z0_t (THETA_n125) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U246 ( .A0_t (StateOut[117]), .B0_t (THETA_n123), .Z0_t (StateFromRhoPi[170]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U245 ( .A0_t (StateOut[109]), .B0_t (THETA_n123), .Z0_t (StateFromRhoPi[148]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U244 ( .A0_t (StateOut[101]), .B0_t (THETA_n123), .Z0_t (StateFromRhoPi[80]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U243 ( .A0_t (StateOut[93]), .B0_t (THETA_n123), .Z0_t (StateFromRhoPi[59]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U242 ( .A0_t (StateOut[85]), .B0_t (THETA_n123), .Z0_t (StateFromRhoPi[35]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U241 ( .A0_t (THETA_n122), .B0_t (THETA_n178), .Z0_t (THETA_n123) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U240 ( .A0_t (StateOut[124]), .B0_t (THETA_n121), .Z0_t (THETA_n178) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U239 ( .A0_t (THETA_n120), .B0_t (THETA_n119), .Z0_t (THETA_n121) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U238 ( .A0_t (StateOut[132]), .B0_t (StateOut[140]), .Z0_t (THETA_n119) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U237 ( .A0_t (StateOut[156]), .B0_t (StateOut[148]), .Z0_t (THETA_n120) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U236 ( .A0_t (StateOut[152]), .B0_t (THETA_n118), .Z0_t (StateFromRhoPi[184]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U235 ( .A0_t (StateOut[144]), .B0_t (THETA_n118), .Z0_t (StateFromRhoPi[125]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U234 ( .A0_t (StateOut[136]), .B0_t (THETA_n118), .Z0_t (StateFromRhoPi[97]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U233 ( .A0_t (StateOut[128]), .B0_t (THETA_n118), .Z0_t (StateFromRhoPi[79]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U232 ( .A0_t (StateOut[120]), .B0_t (THETA_n118), .Z0_t (StateFromRhoPi[12]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U231 ( .A0_t (THETA_n117), .B0_t (THETA_n116), .Z0_t (THETA_n118) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U230 ( .A0_t (StateOut[73]), .B0_t (THETA_n115), .Z0_t (StateFromRhoPi[195]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U229 ( .A0_t (StateOut[65]), .B0_t (THETA_n115), .Z0_t (StateFromRhoPi[134]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U228 ( .A0_t (StateOut[57]), .B0_t (THETA_n115), .Z0_t (StateFromRhoPi[107]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U227 ( .A0_t (StateOut[49]), .B0_t (THETA_n115), .Z0_t (StateFromRhoPi[45]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U226 ( .A0_t (StateOut[41]), .B0_t (THETA_n115), .Z0_t (StateFromRhoPi[18]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U225 ( .A0_t (THETA_n114), .B0_t (THETA_n116), .Z0_t (THETA_n115) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U224 ( .A0_t (StateOut[96]), .B0_t (THETA_n113), .Z0_t (THETA_n116) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U223 ( .A0_t (THETA_n112), .B0_t (THETA_n111), .Z0_t (THETA_n113) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U222 ( .A0_t (StateOut[88]), .B0_t (StateOut[80]), .Z0_t (THETA_n111) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U221 ( .A0_t (StateOut[104]), .B0_t (StateOut[112]), .Z0_t (THETA_n112) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U220 ( .A0_t (StateOut[113]), .B0_t (THETA_n110), .Z0_t (StateFromRhoPi[174]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U219 ( .A0_t (StateOut[105]), .B0_t (THETA_n110), .Z0_t (StateFromRhoPi[144]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U218 ( .A0_t (StateOut[97]), .B0_t (THETA_n110), .Z0_t (StateFromRhoPi[84]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U217 ( .A0_t (StateOut[89]), .B0_t (THETA_n110), .Z0_t (StateFromRhoPi[63]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U216 ( .A0_t (StateOut[81]), .B0_t (THETA_n110), .Z0_t (StateFromRhoPi[39]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U215 ( .A0_t (THETA_n109), .B0_t (THETA_n130), .Z0_t (THETA_n110) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U214 ( .A0_t (StateOut[144]), .B0_t (THETA_n108), .Z0_t (THETA_n130) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U213 ( .A0_t (THETA_n107), .B0_t (THETA_n106), .Z0_t (THETA_n108) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U212 ( .A0_t (StateOut[128]), .B0_t (StateOut[120]), .Z0_t (THETA_n106) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U211 ( .A0_t (StateOut[152]), .B0_t (StateOut[136]), .Z0_t (THETA_n107) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U210 ( .A0_t (StateOut[34]), .B0_t (THETA_n105), .Z0_t (StateFromRhoPi[180]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U209 ( .A0_t (StateOut[26]), .B0_t (THETA_n105), .Z0_t (StateFromRhoPi[155]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U208 ( .A0_t (StateOut[18]), .B0_t (THETA_n105), .Z0_t (StateFromRhoPi[93]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U207 ( .A0_t (StateOut[10]), .B0_t (THETA_n105), .Z0_t (StateFromRhoPi[70]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U206 ( .A0_t (OutData[2]), .B0_t (THETA_n105), .Z0_t (StateFromRhoPi[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U205 ( .A0_t (THETA_n104), .B0_t (THETA_n109), .Z0_t (THETA_n105) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U204 ( .A0_t (StateOut[57]), .B0_t (THETA_n103), .Z0_t (THETA_n109) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U203 ( .A0_t (THETA_n102), .B0_t (THETA_n101), .Z0_t (THETA_n103) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U202 ( .A0_t (StateOut[49]), .B0_t (StateOut[41]), .Z0_t (THETA_n101) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U201 ( .A0_t (StateOut[65]), .B0_t (StateOut[73]), .Z0_t (THETA_n102) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U200 ( .A0_t (StateOut[39]), .B0_t (THETA_n100), .Z0_t (StateFromRhoPi[177]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U199 ( .A0_t (StateOut[31]), .B0_t (THETA_n100), .Z0_t (StateFromRhoPi[152]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U198 ( .A0_t (StateOut[23]), .B0_t (THETA_n100), .Z0_t (StateFromRhoPi[90]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U197 ( .A0_t (StateOut[15]), .B0_t (THETA_n100), .Z0_t (StateFromRhoPi[67]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U196 ( .A0_t (OutData[7]), .B0_t (THETA_n100), .Z0_t (StateFromRhoPi[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U195 ( .A0_t (THETA_n99), .B0_t (THETA_n117), .Z0_t (THETA_n100) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U194 ( .A0_t (StateOut[183]), .B0_t (THETA_n98), .Z0_t (THETA_n117) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U193 ( .A0_t (THETA_n97), .B0_t (THETA_n96), .Z0_t (THETA_n98) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U192 ( .A0_t (StateOut[175]), .B0_t (StateOut[167]), .Z0_t (THETA_n96) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U191 ( .A0_t (StateOut[191]), .B0_t (StateOut[199]), .Z0_t (THETA_n97) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U190 ( .A0_t (StateOut[118]), .B0_t (THETA_n95), .Z0_t (StateFromRhoPi[171]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U189 ( .A0_t (StateOut[110]), .B0_t (THETA_n95), .Z0_t (StateFromRhoPi[149]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U188 ( .A0_t (StateOut[102]), .B0_t (THETA_n95), .Z0_t (StateFromRhoPi[81]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U187 ( .A0_t (StateOut[94]), .B0_t (THETA_n95), .Z0_t (StateFromRhoPi[60]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U186 ( .A0_t (StateOut[86]), .B0_t (THETA_n95), .Z0_t (StateFromRhoPi[36]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U185 ( .A0_t (THETA_n94), .B0_t (THETA_n99), .Z0_t (THETA_n95) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U184 ( .A0_t (StateOut[62]), .B0_t (THETA_n93), .Z0_t (THETA_n99) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U183 ( .A0_t (THETA_n92), .B0_t (THETA_n91), .Z0_t (THETA_n93) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U182 ( .A0_t (StateOut[54]), .B0_t (StateOut[46]), .Z0_t (THETA_n91) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U181 ( .A0_t (StateOut[70]), .B0_t (StateOut[78]), .Z0_t (THETA_n92) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U180 ( .A0_t (StateOut[159]), .B0_t (THETA_n90), .Z0_t (StateFromRhoPi[191]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U179 ( .A0_t (StateOut[151]), .B0_t (THETA_n90), .Z0_t (StateFromRhoPi[124]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U178 ( .A0_t (StateOut[143]), .B0_t (THETA_n90), .Z0_t (StateFromRhoPi[96]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U177 ( .A0_t (StateOut[135]), .B0_t (THETA_n90), .Z0_t (StateFromRhoPi[78]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U176 ( .A0_t (StateOut[127]), .B0_t (THETA_n90), .Z0_t (StateFromRhoPi[11]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U175 ( .A0_t (THETA_n89), .B0_t (THETA_n167), .Z0_t (THETA_n90) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U174 ( .A0_t (StateOut[103]), .B0_t (THETA_n88), .Z0_t (THETA_n167) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U173 ( .A0_t (THETA_n87), .B0_t (THETA_n86), .Z0_t (THETA_n88) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U172 ( .A0_t (StateOut[95]), .B0_t (StateOut[87]), .Z0_t (THETA_n86) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U171 ( .A0_t (StateOut[111]), .B0_t (StateOut[119]), .Z0_t (THETA_n87) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U170 ( .A0_t (StateOut[38]), .B0_t (THETA_n85), .Z0_t (StateFromRhoPi[176]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U169 ( .A0_t (StateOut[30]), .B0_t (THETA_n85), .Z0_t (StateFromRhoPi[159]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U168 ( .A0_t (StateOut[22]), .B0_t (THETA_n85), .Z0_t (StateFromRhoPi[89]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U167 ( .A0_t (StateOut[14]), .B0_t (THETA_n85), .Z0_t (StateFromRhoPi[66]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U166 ( .A0_t (OutData[6]), .B0_t (THETA_n85), .Z0_t (StateFromRhoPi[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U165 ( .A0_t (THETA_n122), .B0_t (THETA_n89), .Z0_t (THETA_n85) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U164 ( .A0_t (StateOut[182]), .B0_t (THETA_n84), .Z0_t (THETA_n89) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U163 ( .A0_t (THETA_n83), .B0_t (THETA_n82), .Z0_t (THETA_n84) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U162 ( .A0_t (StateOut[174]), .B0_t (StateOut[166]), .Z0_t (THETA_n82) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U161 ( .A0_t (StateOut[190]), .B0_t (StateOut[198]), .Z0_t (THETA_n83) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U160 ( .A0_t (StateOut[45]), .B0_t (THETA_n81), .Z0_t (THETA_n122) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U159 ( .A0_t (THETA_n80), .B0_t (THETA_n79), .Z0_t (THETA_n81) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U158 ( .A0_t (StateOut[53]), .B0_t (StateOut[61]), .Z0_t (THETA_n79) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U157 ( .A0_t (StateOut[77]), .B0_t (StateOut[69]), .Z0_t (THETA_n80) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U156 ( .A0_t (StateOut[195]), .B0_t (THETA_n78), .Z0_t (StateFromRhoPi[161]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U155 ( .A0_t (StateOut[187]), .B0_t (THETA_n78), .Z0_t (StateFromRhoPi[139]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U154 ( .A0_t (StateOut[179]), .B0_t (THETA_n78), .Z0_t (StateFromRhoPi[114]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U153 ( .A0_t (StateOut[171]), .B0_t (THETA_n78), .Z0_t (StateFromRhoPi[55]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U152 ( .A0_t (StateOut[163]), .B0_t (THETA_n78), .Z0_t (StateFromRhoPi[30]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U151 ( .A0_t (THETA_n77), .B0_t (THETA_n142), .Z0_t (THETA_n78) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U150 ( .A0_t (StateOut[26]), .B0_t (THETA_n76), .Z0_t (THETA_n142) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U149 ( .A0_t (THETA_n75), .B0_t (THETA_n74), .Z0_t (THETA_n76) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U148 ( .A0_t (StateOut[10]), .B0_t (OutData[2]), .Z0_t (THETA_n74) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U147 ( .A0_t (StateOut[34]), .B0_t (StateOut[18]), .Z0_t (THETA_n75) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U146 ( .A0_t (StateOut[197]), .B0_t (THETA_n73), .Z0_t (StateFromRhoPi[163]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U145 ( .A0_t (StateOut[189]), .B0_t (THETA_n73), .Z0_t (StateFromRhoPi[141]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U144 ( .A0_t (StateOut[181]), .B0_t (THETA_n73), .Z0_t (StateFromRhoPi[116]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U143 ( .A0_t (StateOut[173]), .B0_t (THETA_n73), .Z0_t (StateFromRhoPi[49]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U142 ( .A0_t (StateOut[165]), .B0_t (THETA_n73), .Z0_t (StateFromRhoPi[24]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U141 ( .A0_t (THETA_n72), .B0_t (THETA_n94), .Z0_t (THETA_n73) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U140 ( .A0_t (StateOut[125]), .B0_t (THETA_n71), .Z0_t (THETA_n94) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U139 ( .A0_t (THETA_n70), .B0_t (THETA_n69), .Z0_t (THETA_n71) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U138 ( .A0_t (StateOut[133]), .B0_t (StateOut[141]), .Z0_t (THETA_n69) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U137 ( .A0_t (StateOut[157]), .B0_t (StateOut[149]), .Z0_t (THETA_n70) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U136 ( .A0_t (StateOut[76]), .B0_t (THETA_n68), .Z0_t (StateFromRhoPi[198]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U135 ( .A0_t (StateOut[68]), .B0_t (THETA_n68), .Z0_t (StateFromRhoPi[129]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U134 ( .A0_t (StateOut[60]), .B0_t (THETA_n68), .Z0_t (StateFromRhoPi[110]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U133 ( .A0_t (StateOut[52]), .B0_t (THETA_n68), .Z0_t (StateFromRhoPi[40]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U132 ( .A0_t (StateOut[44]), .B0_t (THETA_n68), .Z0_t (StateFromRhoPi[21]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U131 ( .A0_t (THETA_n67), .B0_t (THETA_n72), .Z0_t (THETA_n68) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U130 ( .A0_t (OutData[4]), .B0_t (THETA_n66), .Z0_t (THETA_n72) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U129 ( .A0_t (THETA_n65), .B0_t (THETA_n64), .Z0_t (THETA_n66) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U128 ( .A0_t (StateOut[12]), .B0_t (StateOut[20]), .Z0_t (THETA_n64) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U127 ( .A0_t (StateOut[36]), .B0_t (StateOut[28]), .Z0_t (THETA_n65) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U126 ( .A0_t (StateOut[116]), .B0_t (THETA_n63), .Z0_t (StateFromRhoPi[169]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U125 ( .A0_t (StateOut[108]), .B0_t (THETA_n63), .Z0_t (StateFromRhoPi[147]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U124 ( .A0_t (StateOut[100]), .B0_t (THETA_n63), .Z0_t (StateFromRhoPi[87]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U123 ( .A0_t (StateOut[92]), .B0_t (THETA_n63), .Z0_t (StateFromRhoPi[58]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U122 ( .A0_t (StateOut[84]), .B0_t (THETA_n63), .Z0_t (StateFromRhoPi[34]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U121 ( .A0_t (THETA_n62), .B0_t (THETA_n77), .Z0_t (THETA_n63) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U120 ( .A0_t (StateOut[123]), .B0_t (THETA_n61), .Z0_t (THETA_n77) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U119 ( .A0_t (THETA_n60), .B0_t (THETA_n59), .Z0_t (THETA_n61) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U118 ( .A0_t (StateOut[131]), .B0_t (StateOut[139]), .Z0_t (THETA_n59) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U117 ( .A0_t (StateOut[155]), .B0_t (StateOut[147]), .Z0_t (THETA_n60) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U116 ( .A0_t (StateOut[37]), .B0_t (THETA_n58), .Z0_t (StateFromRhoPi[183]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U115 ( .A0_t (StateOut[29]), .B0_t (THETA_n58), .Z0_t (StateFromRhoPi[158]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U114 ( .A0_t (StateOut[21]), .B0_t (THETA_n58), .Z0_t (StateFromRhoPi[88]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U113 ( .A0_t (StateOut[13]), .B0_t (THETA_n58), .Z0_t (StateFromRhoPi[65]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U112 ( .A0_t (OutData[5]), .B0_t (THETA_n58), .Z0_t (StateFromRhoPi[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U111 ( .A0_t (THETA_n57), .B0_t (THETA_n62), .Z0_t (THETA_n58) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U110 ( .A0_t (StateOut[60]), .B0_t (THETA_n56), .Z0_t (THETA_n62) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U109 ( .A0_t (THETA_n55), .B0_t (THETA_n54), .Z0_t (THETA_n56) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U108 ( .A0_t (StateOut[52]), .B0_t (StateOut[44]), .Z0_t (THETA_n54) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U107 ( .A0_t (StateOut[68]), .B0_t (StateOut[76]), .Z0_t (THETA_n55) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U106 ( .A0_t (StateOut[115]), .B0_t (THETA_n53), .Z0_t (StateFromRhoPi[168]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U105 ( .A0_t (StateOut[107]), .B0_t (THETA_n53), .Z0_t (StateFromRhoPi[146]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U104 ( .A0_t (StateOut[99]), .B0_t (THETA_n53), .Z0_t (StateFromRhoPi[86]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U103 ( .A0_t (StateOut[91]), .B0_t (THETA_n53), .Z0_t (StateFromRhoPi[57]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U102 ( .A0_t (StateOut[83]), .B0_t (THETA_n53), .Z0_t (StateFromRhoPi[33]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U101 ( .A0_t (THETA_n52), .B0_t (THETA_n51), .Z0_t (THETA_n53) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U100 ( .A0_t (StateOut[36]), .B0_t (THETA_n50), .Z0_t (StateFromRhoPi[182]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U99 ( .A0_t (StateOut[28]), .B0_t (THETA_n50), .Z0_t (StateFromRhoPi[157]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U98 ( .A0_t (StateOut[20]), .B0_t (THETA_n50), .Z0_t (StateFromRhoPi[95]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U97 ( .A0_t (StateOut[12]), .B0_t (THETA_n50), .Z0_t (StateFromRhoPi[64]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U96 ( .A0_t (OutData[4]), .B0_t (THETA_n50), .Z0_t (StateFromRhoPi[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U95 ( .A0_t (THETA_n49), .B0_t (THETA_n51), .Z0_t (THETA_n50) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U94 ( .A0_t (StateOut[59]), .B0_t (THETA_n48), .Z0_t (THETA_n51) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U93 ( .A0_t (THETA_n47), .B0_t (THETA_n46), .Z0_t (THETA_n48) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U92 ( .A0_t (StateOut[51]), .B0_t (StateOut[43]), .Z0_t (THETA_n46) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U91 ( .A0_t (StateOut[67]), .B0_t (StateOut[75]), .Z0_t (THETA_n47) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U90 ( .A0_t (StateOut[77]), .B0_t (THETA_n45), .Z0_t (StateFromRhoPi[199]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U89 ( .A0_t (StateOut[69]), .B0_t (THETA_n45), .Z0_t (StateFromRhoPi[130]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U88 ( .A0_t (StateOut[61]), .B0_t (THETA_n45), .Z0_t (StateFromRhoPi[111]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U87 ( .A0_t (StateOut[53]), .B0_t (THETA_n45), .Z0_t (StateFromRhoPi[41]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U86 ( .A0_t (StateOut[45]), .B0_t (THETA_n45), .Z0_t (StateFromRhoPi[22]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U85 ( .A0_t (THETA_n44), .B0_t (THETA_n186), .Z0_t (THETA_n45) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U84 ( .A0_t (StateOut[29]), .B0_t (THETA_n43), .Z0_t (THETA_n186) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U83 ( .A0_t (THETA_n42), .B0_t (THETA_n41), .Z0_t (THETA_n43) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U82 ( .A0_t (StateOut[13]), .B0_t (OutData[5]), .Z0_t (THETA_n41) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U81 ( .A0_t (StateOut[37]), .B0_t (StateOut[21]), .Z0_t (THETA_n42) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U80 ( .A0_t (StateOut[35]), .B0_t (THETA_n40), .Z0_t (StateFromRhoPi[181]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U79 ( .A0_t (StateOut[27]), .B0_t (THETA_n40), .Z0_t (StateFromRhoPi[156]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U78 ( .A0_t (StateOut[19]), .B0_t (THETA_n40), .Z0_t (StateFromRhoPi[94]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U77 ( .A0_t (StateOut[11]), .B0_t (THETA_n40), .Z0_t (StateFromRhoPi[71]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U76 ( .A0_t (OutData[3]), .B0_t (THETA_n40), .Z0_t (StateFromRhoPi[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U75 ( .A0_t (THETA_n39), .B0_t (THETA_n150), .Z0_t (THETA_n40) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U74 ( .A0_t (StateOut[66]), .B0_t (THETA_n38), .Z0_t (THETA_n150) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U73 ( .A0_t (THETA_n37), .B0_t (THETA_n36), .Z0_t (THETA_n38) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U72 ( .A0_t (StateOut[50]), .B0_t (StateOut[42]), .Z0_t (THETA_n36) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U71 ( .A0_t (StateOut[74]), .B0_t (StateOut[58]), .Z0_t (THETA_n37) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U70 ( .A0_t (StateOut[158]), .B0_t (THETA_n35), .Z0_t (StateFromRhoPi[190]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U69 ( .A0_t (StateOut[150]), .B0_t (THETA_n35), .Z0_t (StateFromRhoPi[123]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U68 ( .A0_t (StateOut[142]), .B0_t (THETA_n35), .Z0_t (StateFromRhoPi[103]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U67 ( .A0_t (StateOut[134]), .B0_t (THETA_n35), .Z0_t (StateFromRhoPi[77]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U66 ( .A0_t (StateOut[126]), .B0_t (THETA_n35), .Z0_t (StateFromRhoPi[10]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U65 ( .A0_t (THETA_n127), .B0_t (THETA_n57), .Z0_t (THETA_n35) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U64 ( .A0_t (StateOut[181]), .B0_t (THETA_n34), .Z0_t (THETA_n57) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U63 ( .A0_t (THETA_n33), .B0_t (THETA_n32), .Z0_t (THETA_n34) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U62 ( .A0_t (StateOut[173]), .B0_t (StateOut[165]), .Z0_t (THETA_n32) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U61 ( .A0_t (StateOut[189]), .B0_t (StateOut[197]), .Z0_t (THETA_n33) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U60 ( .A0_t (StateOut[110]), .B0_t (THETA_n31), .Z0_t (THETA_n127) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U59 ( .A0_t (THETA_n30), .B0_t (THETA_n29), .Z0_t (THETA_n31) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U58 ( .A0_t (StateOut[94]), .B0_t (StateOut[86]), .Z0_t (THETA_n29) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U57 ( .A0_t (StateOut[118]), .B0_t (StateOut[102]), .Z0_t (THETA_n30) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U56 ( .A0_t (StateOut[157]), .B0_t (THETA_n28), .Z0_t (StateFromRhoPi[189]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U55 ( .A0_t (StateOut[149]), .B0_t (THETA_n28), .Z0_t (StateFromRhoPi[122]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U54 ( .A0_t (StateOut[141]), .B0_t (THETA_n28), .Z0_t (StateFromRhoPi[102]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U53 ( .A0_t (StateOut[133]), .B0_t (THETA_n28), .Z0_t (StateFromRhoPi[76]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U52 ( .A0_t (StateOut[125]), .B0_t (THETA_n28), .Z0_t (StateFromRhoPi[9]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U51 ( .A0_t (THETA_n196), .B0_t (THETA_n49), .Z0_t (THETA_n28) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U50 ( .A0_t (StateOut[180]), .B0_t (THETA_n27), .Z0_t (THETA_n49) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U49 ( .A0_t (THETA_n26), .B0_t (THETA_n25), .Z0_t (THETA_n27) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U48 ( .A0_t (StateOut[172]), .B0_t (StateOut[164]), .Z0_t (THETA_n25) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U47 ( .A0_t (StateOut[188]), .B0_t (StateOut[196]), .Z0_t (THETA_n26) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U46 ( .A0_t (StateOut[109]), .B0_t (THETA_n24), .Z0_t (THETA_n196) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U45 ( .A0_t (THETA_n23), .B0_t (THETA_n22), .Z0_t (THETA_n24) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U44 ( .A0_t (StateOut[93]), .B0_t (StateOut[85]), .Z0_t (THETA_n22) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U43 ( .A0_t (StateOut[117]), .B0_t (StateOut[101]), .Z0_t (THETA_n23) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U42 ( .A0_t (StateOut[194]), .B0_t (THETA_n21), .Z0_t (StateFromRhoPi[160]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U41 ( .A0_t (StateOut[186]), .B0_t (THETA_n21), .Z0_t (StateFromRhoPi[138]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U40 ( .A0_t (StateOut[178]), .B0_t (THETA_n21), .Z0_t (StateFromRhoPi[113]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U39 ( .A0_t (StateOut[170]), .B0_t (THETA_n21), .Z0_t (StateFromRhoPi[54]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U38 ( .A0_t (StateOut[162]), .B0_t (THETA_n21), .Z0_t (StateFromRhoPi[29]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U37 ( .A0_t (THETA_n114), .B0_t (THETA_n52), .Z0_t (THETA_n21) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U36 ( .A0_t (StateOut[138]), .B0_t (THETA_n20), .Z0_t (THETA_n52) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U35 ( .A0_t (THETA_n19), .B0_t (THETA_n18), .Z0_t (THETA_n20) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U34 ( .A0_t (StateOut[130]), .B0_t (StateOut[122]), .Z0_t (THETA_n18) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U33 ( .A0_t (StateOut[146]), .B0_t (StateOut[154]), .Z0_t (THETA_n19) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U32 ( .A0_t (StateOut[17]), .B0_t (THETA_n17), .Z0_t (THETA_n114) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U31 ( .A0_t (THETA_n16), .B0_t (THETA_n15), .Z0_t (THETA_n17) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U30 ( .A0_t (StateOut[9]), .B0_t (OutData[1]), .Z0_t (THETA_n15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U29 ( .A0_t (StateOut[25]), .B0_t (StateOut[33]), .Z0_t (THETA_n16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U28 ( .A0_t (StateOut[156]), .B0_t (THETA_n14), .Z0_t (StateFromRhoPi[188]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U27 ( .A0_t (StateOut[148]), .B0_t (THETA_n14), .Z0_t (StateFromRhoPi[121]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U26 ( .A0_t (StateOut[140]), .B0_t (THETA_n14), .Z0_t (StateFromRhoPi[101]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U25 ( .A0_t (StateOut[132]), .B0_t (THETA_n14), .Z0_t (StateFromRhoPi[75]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U24 ( .A0_t (StateOut[124]), .B0_t (THETA_n14), .Z0_t (StateFromRhoPi[8]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U23 ( .A0_t (THETA_n44), .B0_t (THETA_n39), .Z0_t (THETA_n14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U22 ( .A0_t (StateOut[179]), .B0_t (THETA_n13), .Z0_t (THETA_n39) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U21 ( .A0_t (THETA_n12), .B0_t (THETA_n11), .Z0_t (THETA_n13) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U20 ( .A0_t (StateOut[171]), .B0_t (StateOut[163]), .Z0_t (THETA_n11) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U19 ( .A0_t (StateOut[187]), .B0_t (StateOut[195]), .Z0_t (THETA_n12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U18 ( .A0_t (StateOut[100]), .B0_t (THETA_n10), .Z0_t (THETA_n44) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U17 ( .A0_t (THETA_n9), .B0_t (THETA_n8), .Z0_t (THETA_n10) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U16 ( .A0_t (StateOut[92]), .B0_t (StateOut[84]), .Z0_t (THETA_n8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U15 ( .A0_t (StateOut[108]), .B0_t (StateOut[116]), .Z0_t (THETA_n9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U14 ( .A0_t (StateOut[155]), .B0_t (THETA_n7), .Z0_t (StateFromRhoPi[187]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U13 ( .A0_t (StateOut[147]), .B0_t (THETA_n7), .Z0_t (StateFromRhoPi[120]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U12 ( .A0_t (StateOut[139]), .B0_t (THETA_n7), .Z0_t (StateFromRhoPi[100]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U11 ( .A0_t (StateOut[131]), .B0_t (THETA_n7), .Z0_t (StateFromRhoPi[74]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U10 ( .A0_t (StateOut[123]), .B0_t (THETA_n7), .Z0_t (StateFromRhoPi[15]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U9 ( .A0_t (THETA_n104), .B0_t (THETA_n67), .Z0_t (THETA_n7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U8 ( .A0_t (StateOut[107]), .B0_t (THETA_n6), .Z0_t (THETA_n67) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U7 ( .A0_t (THETA_n5), .B0_t (THETA_n4), .Z0_t (THETA_n6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U6 ( .A0_t (StateOut[91]), .B0_t (StateOut[83]), .Z0_t (THETA_n4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U5 ( .A0_t (StateOut[115]), .B0_t (StateOut[99]), .Z0_t (THETA_n5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U4 ( .A0_t (StateOut[186]), .B0_t (THETA_n3), .Z0_t (THETA_n104) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U3 ( .A0_t (THETA_n2), .B0_t (THETA_n1), .Z0_t (THETA_n3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) THETA_U2 ( .A0_t (StateOut[170]), .B0_t (StateOut[162]), .Z0_t (THETA_n1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) THETA_U1 ( .A0_t (StateOut[194]), .B0_t (StateOut[178]), .Z0_t (THETA_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_U4 ( .A0_t (CHI_ChiOut[0]), .B0_t (IotaRC[0]), .Z0_t (StateFromChi[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_U3 ( .A0_t (CHI_ChiOut[1]), .B0_t (IotaRC[1]), .Z0_t (StateFromChi[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_U2 ( .A0_t (CHI_ChiOut_7), .B0_t (IotaRC_7), .Z0_t (StateFromChi[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_U1 ( .A0_t (CHI_ChiOut_3), .B0_t (IotaRC_3), .Z0_t (StateFromChi[3]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[40]), .B0_t (StateFromRhoPi[80]), .Z0_t (CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_and_xor_inst_a_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_and_xor_inst_a_nxy), .B0_t (StateFromRhoPi[0]), .Z0_t (CHI_ChiOut[0]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[80]), .B0_t (StateFromRhoPi[120]), .Z0_t (CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_and_xor_inst_b_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_and_xor_inst_b_nxy), .B0_t (StateFromRhoPi[40]), .Z0_t (StateFromChi[40]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[120]), .B0_t (StateFromRhoPi[160]), .Z0_t (CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_and_xor_inst_c_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_and_xor_inst_c_nxy), .B0_t (StateFromRhoPi[80]), .Z0_t (StateFromChi[80]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[160]), .B0_t (StateFromRhoPi[0]), .Z0_t (CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_and_xor_inst_d_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_and_xor_inst_d_nxy), .B0_t (StateFromRhoPi[120]), .Z0_t (StateFromChi[120]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[0]), .B0_t (StateFromRhoPi[40]), .Z0_t (CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_and_xor_inst_e_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_0__GEN_ROWS_0__sbox_and_xor_inst_e_nxy), .B0_t (StateFromRhoPi[160]), .Z0_t (StateFromChi[160]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[48]), .B0_t (StateFromRhoPi[88]), .Z0_t (CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_and_xor_inst_a_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_and_xor_inst_a_nxy), .B0_t (StateFromRhoPi[8]), .Z0_t (StateFromChi[8]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[88]), .B0_t (StateFromRhoPi[128]), .Z0_t (CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_and_xor_inst_b_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_and_xor_inst_b_nxy), .B0_t (StateFromRhoPi[48]), .Z0_t (StateFromChi[48]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[128]), .B0_t (StateFromRhoPi[168]), .Z0_t (CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_and_xor_inst_c_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_and_xor_inst_c_nxy), .B0_t (StateFromRhoPi[88]), .Z0_t (StateFromChi[88]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[168]), .B0_t (StateFromRhoPi[8]), .Z0_t (CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_and_xor_inst_d_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_and_xor_inst_d_nxy), .B0_t (StateFromRhoPi[128]), .Z0_t (StateFromChi[128]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[8]), .B0_t (StateFromRhoPi[48]), .Z0_t (CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_and_xor_inst_e_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_0__GEN_ROWS_1__sbox_and_xor_inst_e_nxy), .B0_t (StateFromRhoPi[168]), .Z0_t (StateFromChi[168]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[56]), .B0_t (StateFromRhoPi[96]), .Z0_t (CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_and_xor_inst_a_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_and_xor_inst_a_nxy), .B0_t (StateFromRhoPi[16]), .Z0_t (StateFromChi[16]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[96]), .B0_t (StateFromRhoPi[136]), .Z0_t (CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_and_xor_inst_b_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_and_xor_inst_b_nxy), .B0_t (StateFromRhoPi[56]), .Z0_t (StateFromChi[56]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[136]), .B0_t (StateFromRhoPi[176]), .Z0_t (CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_and_xor_inst_c_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_and_xor_inst_c_nxy), .B0_t (StateFromRhoPi[96]), .Z0_t (StateFromChi[96]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[176]), .B0_t (StateFromRhoPi[16]), .Z0_t (CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_and_xor_inst_d_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_and_xor_inst_d_nxy), .B0_t (StateFromRhoPi[136]), .Z0_t (StateFromChi[136]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[16]), .B0_t (StateFromRhoPi[56]), .Z0_t (CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_and_xor_inst_e_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_0__GEN_ROWS_2__sbox_and_xor_inst_e_nxy), .B0_t (StateFromRhoPi[176]), .Z0_t (StateFromChi[176]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[64]), .B0_t (StateFromRhoPi[104]), .Z0_t (CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_and_xor_inst_a_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_and_xor_inst_a_nxy), .B0_t (StateFromRhoPi[24]), .Z0_t (StateFromChi[24]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[104]), .B0_t (StateFromRhoPi[144]), .Z0_t (CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_and_xor_inst_b_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_and_xor_inst_b_nxy), .B0_t (StateFromRhoPi[64]), .Z0_t (StateFromChi[64]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[144]), .B0_t (StateFromRhoPi[184]), .Z0_t (CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_and_xor_inst_c_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_and_xor_inst_c_nxy), .B0_t (StateFromRhoPi[104]), .Z0_t (StateFromChi[104]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[184]), .B0_t (StateFromRhoPi[24]), .Z0_t (CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_and_xor_inst_d_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_and_xor_inst_d_nxy), .B0_t (StateFromRhoPi[144]), .Z0_t (StateFromChi[144]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[24]), .B0_t (StateFromRhoPi[64]), .Z0_t (CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_and_xor_inst_e_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_0__GEN_ROWS_3__sbox_and_xor_inst_e_nxy), .B0_t (StateFromRhoPi[184]), .Z0_t (StateFromChi[184]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[72]), .B0_t (StateFromRhoPi[112]), .Z0_t (CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_and_xor_inst_a_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_and_xor_inst_a_nxy), .B0_t (StateFromRhoPi[32]), .Z0_t (StateFromChi[32]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[112]), .B0_t (StateFromRhoPi[152]), .Z0_t (CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_and_xor_inst_b_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_and_xor_inst_b_nxy), .B0_t (StateFromRhoPi[72]), .Z0_t (StateFromChi[72]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[152]), .B0_t (StateFromRhoPi[192]), .Z0_t (CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_and_xor_inst_c_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_and_xor_inst_c_nxy), .B0_t (StateFromRhoPi[112]), .Z0_t (StateFromChi[112]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[192]), .B0_t (StateFromRhoPi[32]), .Z0_t (CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_and_xor_inst_d_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_and_xor_inst_d_nxy), .B0_t (StateFromRhoPi[152]), .Z0_t (StateFromChi[152]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[32]), .B0_t (StateFromRhoPi[72]), .Z0_t (CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_and_xor_inst_e_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_0__GEN_ROWS_4__sbox_and_xor_inst_e_nxy), .B0_t (StateFromRhoPi[192]), .Z0_t (StateFromChi[192]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_0__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[41]), .B0_t (StateFromRhoPi[81]), .Z0_t (CHI_GEN_SLICES_1__GEN_ROWS_0__sbox_and_xor_inst_a_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_0__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_1__GEN_ROWS_0__sbox_and_xor_inst_a_nxy), .B0_t (StateFromRhoPi[1]), .Z0_t (CHI_ChiOut[1]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_0__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[81]), .B0_t (StateFromRhoPi[121]), .Z0_t (CHI_GEN_SLICES_1__GEN_ROWS_0__sbox_and_xor_inst_b_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_0__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_1__GEN_ROWS_0__sbox_and_xor_inst_b_nxy), .B0_t (StateFromRhoPi[41]), .Z0_t (StateFromChi[41]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_0__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[121]), .B0_t (StateFromRhoPi[161]), .Z0_t (CHI_GEN_SLICES_1__GEN_ROWS_0__sbox_and_xor_inst_c_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_0__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_1__GEN_ROWS_0__sbox_and_xor_inst_c_nxy), .B0_t (StateFromRhoPi[81]), .Z0_t (StateFromChi[81]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_0__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[161]), .B0_t (StateFromRhoPi[1]), .Z0_t (CHI_GEN_SLICES_1__GEN_ROWS_0__sbox_and_xor_inst_d_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_0__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_1__GEN_ROWS_0__sbox_and_xor_inst_d_nxy), .B0_t (StateFromRhoPi[121]), .Z0_t (StateFromChi[121]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_0__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[1]), .B0_t (StateFromRhoPi[41]), .Z0_t (CHI_GEN_SLICES_1__GEN_ROWS_0__sbox_and_xor_inst_e_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_0__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_1__GEN_ROWS_0__sbox_and_xor_inst_e_nxy), .B0_t (StateFromRhoPi[161]), .Z0_t (StateFromChi[161]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_1__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[49]), .B0_t (StateFromRhoPi[89]), .Z0_t (CHI_GEN_SLICES_1__GEN_ROWS_1__sbox_and_xor_inst_a_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_1__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_1__GEN_ROWS_1__sbox_and_xor_inst_a_nxy), .B0_t (StateFromRhoPi[9]), .Z0_t (StateFromChi[9]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_1__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[89]), .B0_t (StateFromRhoPi[129]), .Z0_t (CHI_GEN_SLICES_1__GEN_ROWS_1__sbox_and_xor_inst_b_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_1__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_1__GEN_ROWS_1__sbox_and_xor_inst_b_nxy), .B0_t (StateFromRhoPi[49]), .Z0_t (StateFromChi[49]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_1__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[129]), .B0_t (StateFromRhoPi[169]), .Z0_t (CHI_GEN_SLICES_1__GEN_ROWS_1__sbox_and_xor_inst_c_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_1__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_1__GEN_ROWS_1__sbox_and_xor_inst_c_nxy), .B0_t (StateFromRhoPi[89]), .Z0_t (StateFromChi[89]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_1__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[169]), .B0_t (StateFromRhoPi[9]), .Z0_t (CHI_GEN_SLICES_1__GEN_ROWS_1__sbox_and_xor_inst_d_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_1__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_1__GEN_ROWS_1__sbox_and_xor_inst_d_nxy), .B0_t (StateFromRhoPi[129]), .Z0_t (StateFromChi[129]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_1__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[9]), .B0_t (StateFromRhoPi[49]), .Z0_t (CHI_GEN_SLICES_1__GEN_ROWS_1__sbox_and_xor_inst_e_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_1__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_1__GEN_ROWS_1__sbox_and_xor_inst_e_nxy), .B0_t (StateFromRhoPi[169]), .Z0_t (StateFromChi[169]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_2__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[57]), .B0_t (StateFromRhoPi[97]), .Z0_t (CHI_GEN_SLICES_1__GEN_ROWS_2__sbox_and_xor_inst_a_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_2__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_1__GEN_ROWS_2__sbox_and_xor_inst_a_nxy), .B0_t (StateFromRhoPi[17]), .Z0_t (StateFromChi[17]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_2__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[97]), .B0_t (StateFromRhoPi[137]), .Z0_t (CHI_GEN_SLICES_1__GEN_ROWS_2__sbox_and_xor_inst_b_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_2__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_1__GEN_ROWS_2__sbox_and_xor_inst_b_nxy), .B0_t (StateFromRhoPi[57]), .Z0_t (StateFromChi[57]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_2__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[137]), .B0_t (StateFromRhoPi[177]), .Z0_t (CHI_GEN_SLICES_1__GEN_ROWS_2__sbox_and_xor_inst_c_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_2__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_1__GEN_ROWS_2__sbox_and_xor_inst_c_nxy), .B0_t (StateFromRhoPi[97]), .Z0_t (StateFromChi[97]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_2__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[177]), .B0_t (StateFromRhoPi[17]), .Z0_t (CHI_GEN_SLICES_1__GEN_ROWS_2__sbox_and_xor_inst_d_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_2__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_1__GEN_ROWS_2__sbox_and_xor_inst_d_nxy), .B0_t (StateFromRhoPi[137]), .Z0_t (StateFromChi[137]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_2__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[17]), .B0_t (StateFromRhoPi[57]), .Z0_t (CHI_GEN_SLICES_1__GEN_ROWS_2__sbox_and_xor_inst_e_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_2__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_1__GEN_ROWS_2__sbox_and_xor_inst_e_nxy), .B0_t (StateFromRhoPi[177]), .Z0_t (StateFromChi[177]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_3__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[65]), .B0_t (StateFromRhoPi[105]), .Z0_t (CHI_GEN_SLICES_1__GEN_ROWS_3__sbox_and_xor_inst_a_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_3__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_1__GEN_ROWS_3__sbox_and_xor_inst_a_nxy), .B0_t (StateFromRhoPi[25]), .Z0_t (StateFromChi[25]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_3__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[105]), .B0_t (StateFromRhoPi[145]), .Z0_t (CHI_GEN_SLICES_1__GEN_ROWS_3__sbox_and_xor_inst_b_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_3__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_1__GEN_ROWS_3__sbox_and_xor_inst_b_nxy), .B0_t (StateFromRhoPi[65]), .Z0_t (StateFromChi[65]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_3__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[145]), .B0_t (StateFromRhoPi[185]), .Z0_t (CHI_GEN_SLICES_1__GEN_ROWS_3__sbox_and_xor_inst_c_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_3__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_1__GEN_ROWS_3__sbox_and_xor_inst_c_nxy), .B0_t (StateFromRhoPi[105]), .Z0_t (StateFromChi[105]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_3__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[185]), .B0_t (StateFromRhoPi[25]), .Z0_t (CHI_GEN_SLICES_1__GEN_ROWS_3__sbox_and_xor_inst_d_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_3__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_1__GEN_ROWS_3__sbox_and_xor_inst_d_nxy), .B0_t (StateFromRhoPi[145]), .Z0_t (StateFromChi[145]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_3__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[25]), .B0_t (StateFromRhoPi[65]), .Z0_t (CHI_GEN_SLICES_1__GEN_ROWS_3__sbox_and_xor_inst_e_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_3__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_1__GEN_ROWS_3__sbox_and_xor_inst_e_nxy), .B0_t (StateFromRhoPi[185]), .Z0_t (StateFromChi[185]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_4__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[73]), .B0_t (StateFromRhoPi[113]), .Z0_t (CHI_GEN_SLICES_1__GEN_ROWS_4__sbox_and_xor_inst_a_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_4__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_1__GEN_ROWS_4__sbox_and_xor_inst_a_nxy), .B0_t (StateFromRhoPi[33]), .Z0_t (StateFromChi[33]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_4__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[113]), .B0_t (StateFromRhoPi[153]), .Z0_t (CHI_GEN_SLICES_1__GEN_ROWS_4__sbox_and_xor_inst_b_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_4__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_1__GEN_ROWS_4__sbox_and_xor_inst_b_nxy), .B0_t (StateFromRhoPi[73]), .Z0_t (StateFromChi[73]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_4__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[153]), .B0_t (StateFromRhoPi[193]), .Z0_t (CHI_GEN_SLICES_1__GEN_ROWS_4__sbox_and_xor_inst_c_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_4__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_1__GEN_ROWS_4__sbox_and_xor_inst_c_nxy), .B0_t (StateFromRhoPi[113]), .Z0_t (StateFromChi[113]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_4__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[193]), .B0_t (StateFromRhoPi[33]), .Z0_t (CHI_GEN_SLICES_1__GEN_ROWS_4__sbox_and_xor_inst_d_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_4__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_1__GEN_ROWS_4__sbox_and_xor_inst_d_nxy), .B0_t (StateFromRhoPi[153]), .Z0_t (StateFromChi[153]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_4__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[33]), .B0_t (StateFromRhoPi[73]), .Z0_t (CHI_GEN_SLICES_1__GEN_ROWS_4__sbox_and_xor_inst_e_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_1__GEN_ROWS_4__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_1__GEN_ROWS_4__sbox_and_xor_inst_e_nxy), .B0_t (StateFromRhoPi[193]), .Z0_t (StateFromChi[193]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_0__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[42]), .B0_t (StateFromRhoPi[82]), .Z0_t (CHI_GEN_SLICES_2__GEN_ROWS_0__sbox_and_xor_inst_a_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_0__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_2__GEN_ROWS_0__sbox_and_xor_inst_a_nxy), .B0_t (StateFromRhoPi[2]), .Z0_t (StateFromChi[2]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_0__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[82]), .B0_t (StateFromRhoPi[122]), .Z0_t (CHI_GEN_SLICES_2__GEN_ROWS_0__sbox_and_xor_inst_b_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_0__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_2__GEN_ROWS_0__sbox_and_xor_inst_b_nxy), .B0_t (StateFromRhoPi[42]), .Z0_t (StateFromChi[42]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_0__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[122]), .B0_t (StateFromRhoPi[162]), .Z0_t (CHI_GEN_SLICES_2__GEN_ROWS_0__sbox_and_xor_inst_c_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_0__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_2__GEN_ROWS_0__sbox_and_xor_inst_c_nxy), .B0_t (StateFromRhoPi[82]), .Z0_t (StateFromChi[82]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_0__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[162]), .B0_t (StateFromRhoPi[2]), .Z0_t (CHI_GEN_SLICES_2__GEN_ROWS_0__sbox_and_xor_inst_d_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_0__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_2__GEN_ROWS_0__sbox_and_xor_inst_d_nxy), .B0_t (StateFromRhoPi[122]), .Z0_t (StateFromChi[122]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_0__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[2]), .B0_t (StateFromRhoPi[42]), .Z0_t (CHI_GEN_SLICES_2__GEN_ROWS_0__sbox_and_xor_inst_e_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_0__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_2__GEN_ROWS_0__sbox_and_xor_inst_e_nxy), .B0_t (StateFromRhoPi[162]), .Z0_t (StateFromChi[162]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_1__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[50]), .B0_t (StateFromRhoPi[90]), .Z0_t (CHI_GEN_SLICES_2__GEN_ROWS_1__sbox_and_xor_inst_a_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_1__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_2__GEN_ROWS_1__sbox_and_xor_inst_a_nxy), .B0_t (StateFromRhoPi[10]), .Z0_t (StateFromChi[10]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_1__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[90]), .B0_t (StateFromRhoPi[130]), .Z0_t (CHI_GEN_SLICES_2__GEN_ROWS_1__sbox_and_xor_inst_b_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_1__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_2__GEN_ROWS_1__sbox_and_xor_inst_b_nxy), .B0_t (StateFromRhoPi[50]), .Z0_t (StateFromChi[50]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_1__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[130]), .B0_t (StateFromRhoPi[170]), .Z0_t (CHI_GEN_SLICES_2__GEN_ROWS_1__sbox_and_xor_inst_c_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_1__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_2__GEN_ROWS_1__sbox_and_xor_inst_c_nxy), .B0_t (StateFromRhoPi[90]), .Z0_t (StateFromChi[90]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_1__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[170]), .B0_t (StateFromRhoPi[10]), .Z0_t (CHI_GEN_SLICES_2__GEN_ROWS_1__sbox_and_xor_inst_d_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_1__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_2__GEN_ROWS_1__sbox_and_xor_inst_d_nxy), .B0_t (StateFromRhoPi[130]), .Z0_t (StateFromChi[130]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_1__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[10]), .B0_t (StateFromRhoPi[50]), .Z0_t (CHI_GEN_SLICES_2__GEN_ROWS_1__sbox_and_xor_inst_e_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_1__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_2__GEN_ROWS_1__sbox_and_xor_inst_e_nxy), .B0_t (StateFromRhoPi[170]), .Z0_t (StateFromChi[170]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_2__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[58]), .B0_t (StateFromRhoPi[98]), .Z0_t (CHI_GEN_SLICES_2__GEN_ROWS_2__sbox_and_xor_inst_a_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_2__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_2__GEN_ROWS_2__sbox_and_xor_inst_a_nxy), .B0_t (StateFromRhoPi[18]), .Z0_t (StateFromChi[18]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_2__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[98]), .B0_t (StateFromRhoPi[138]), .Z0_t (CHI_GEN_SLICES_2__GEN_ROWS_2__sbox_and_xor_inst_b_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_2__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_2__GEN_ROWS_2__sbox_and_xor_inst_b_nxy), .B0_t (StateFromRhoPi[58]), .Z0_t (StateFromChi[58]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_2__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[138]), .B0_t (StateFromRhoPi[178]), .Z0_t (CHI_GEN_SLICES_2__GEN_ROWS_2__sbox_and_xor_inst_c_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_2__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_2__GEN_ROWS_2__sbox_and_xor_inst_c_nxy), .B0_t (StateFromRhoPi[98]), .Z0_t (StateFromChi[98]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_2__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[178]), .B0_t (StateFromRhoPi[18]), .Z0_t (CHI_GEN_SLICES_2__GEN_ROWS_2__sbox_and_xor_inst_d_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_2__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_2__GEN_ROWS_2__sbox_and_xor_inst_d_nxy), .B0_t (StateFromRhoPi[138]), .Z0_t (StateFromChi[138]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_2__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[18]), .B0_t (StateFromRhoPi[58]), .Z0_t (CHI_GEN_SLICES_2__GEN_ROWS_2__sbox_and_xor_inst_e_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_2__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_2__GEN_ROWS_2__sbox_and_xor_inst_e_nxy), .B0_t (StateFromRhoPi[178]), .Z0_t (StateFromChi[178]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_3__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[66]), .B0_t (StateFromRhoPi[106]), .Z0_t (CHI_GEN_SLICES_2__GEN_ROWS_3__sbox_and_xor_inst_a_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_3__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_2__GEN_ROWS_3__sbox_and_xor_inst_a_nxy), .B0_t (StateFromRhoPi[26]), .Z0_t (StateFromChi[26]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_3__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[106]), .B0_t (StateFromRhoPi[146]), .Z0_t (CHI_GEN_SLICES_2__GEN_ROWS_3__sbox_and_xor_inst_b_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_3__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_2__GEN_ROWS_3__sbox_and_xor_inst_b_nxy), .B0_t (StateFromRhoPi[66]), .Z0_t (StateFromChi[66]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_3__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[146]), .B0_t (StateFromRhoPi[186]), .Z0_t (CHI_GEN_SLICES_2__GEN_ROWS_3__sbox_and_xor_inst_c_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_3__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_2__GEN_ROWS_3__sbox_and_xor_inst_c_nxy), .B0_t (StateFromRhoPi[106]), .Z0_t (StateFromChi[106]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_3__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[186]), .B0_t (StateFromRhoPi[26]), .Z0_t (CHI_GEN_SLICES_2__GEN_ROWS_3__sbox_and_xor_inst_d_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_3__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_2__GEN_ROWS_3__sbox_and_xor_inst_d_nxy), .B0_t (StateFromRhoPi[146]), .Z0_t (StateFromChi[146]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_3__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[26]), .B0_t (StateFromRhoPi[66]), .Z0_t (CHI_GEN_SLICES_2__GEN_ROWS_3__sbox_and_xor_inst_e_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_3__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_2__GEN_ROWS_3__sbox_and_xor_inst_e_nxy), .B0_t (StateFromRhoPi[186]), .Z0_t (StateFromChi[186]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_4__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[74]), .B0_t (StateFromRhoPi[114]), .Z0_t (CHI_GEN_SLICES_2__GEN_ROWS_4__sbox_and_xor_inst_a_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_4__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_2__GEN_ROWS_4__sbox_and_xor_inst_a_nxy), .B0_t (StateFromRhoPi[34]), .Z0_t (StateFromChi[34]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_4__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[114]), .B0_t (StateFromRhoPi[154]), .Z0_t (CHI_GEN_SLICES_2__GEN_ROWS_4__sbox_and_xor_inst_b_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_4__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_2__GEN_ROWS_4__sbox_and_xor_inst_b_nxy), .B0_t (StateFromRhoPi[74]), .Z0_t (StateFromChi[74]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_4__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[154]), .B0_t (StateFromRhoPi[194]), .Z0_t (CHI_GEN_SLICES_2__GEN_ROWS_4__sbox_and_xor_inst_c_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_4__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_2__GEN_ROWS_4__sbox_and_xor_inst_c_nxy), .B0_t (StateFromRhoPi[114]), .Z0_t (StateFromChi[114]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_4__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[194]), .B0_t (StateFromRhoPi[34]), .Z0_t (CHI_GEN_SLICES_2__GEN_ROWS_4__sbox_and_xor_inst_d_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_4__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_2__GEN_ROWS_4__sbox_and_xor_inst_d_nxy), .B0_t (StateFromRhoPi[154]), .Z0_t (StateFromChi[154]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_4__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[34]), .B0_t (StateFromRhoPi[74]), .Z0_t (CHI_GEN_SLICES_2__GEN_ROWS_4__sbox_and_xor_inst_e_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_2__GEN_ROWS_4__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_2__GEN_ROWS_4__sbox_and_xor_inst_e_nxy), .B0_t (StateFromRhoPi[194]), .Z0_t (StateFromChi[194]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_0__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[43]), .B0_t (StateFromRhoPi[83]), .Z0_t (CHI_GEN_SLICES_3__GEN_ROWS_0__sbox_and_xor_inst_a_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_0__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_3__GEN_ROWS_0__sbox_and_xor_inst_a_nxy), .B0_t (StateFromRhoPi[3]), .Z0_t (CHI_ChiOut_3) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_0__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[83]), .B0_t (StateFromRhoPi[123]), .Z0_t (CHI_GEN_SLICES_3__GEN_ROWS_0__sbox_and_xor_inst_b_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_0__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_3__GEN_ROWS_0__sbox_and_xor_inst_b_nxy), .B0_t (StateFromRhoPi[43]), .Z0_t (StateFromChi[43]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_0__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[123]), .B0_t (StateFromRhoPi[163]), .Z0_t (CHI_GEN_SLICES_3__GEN_ROWS_0__sbox_and_xor_inst_c_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_0__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_3__GEN_ROWS_0__sbox_and_xor_inst_c_nxy), .B0_t (StateFromRhoPi[83]), .Z0_t (StateFromChi[83]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_0__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[163]), .B0_t (StateFromRhoPi[3]), .Z0_t (CHI_GEN_SLICES_3__GEN_ROWS_0__sbox_and_xor_inst_d_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_0__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_3__GEN_ROWS_0__sbox_and_xor_inst_d_nxy), .B0_t (StateFromRhoPi[123]), .Z0_t (StateFromChi[123]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_0__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[3]), .B0_t (StateFromRhoPi[43]), .Z0_t (CHI_GEN_SLICES_3__GEN_ROWS_0__sbox_and_xor_inst_e_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_0__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_3__GEN_ROWS_0__sbox_and_xor_inst_e_nxy), .B0_t (StateFromRhoPi[163]), .Z0_t (StateFromChi[163]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_1__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[51]), .B0_t (StateFromRhoPi[91]), .Z0_t (CHI_GEN_SLICES_3__GEN_ROWS_1__sbox_and_xor_inst_a_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_1__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_3__GEN_ROWS_1__sbox_and_xor_inst_a_nxy), .B0_t (StateFromRhoPi[11]), .Z0_t (StateFromChi[11]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_1__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[91]), .B0_t (StateFromRhoPi[131]), .Z0_t (CHI_GEN_SLICES_3__GEN_ROWS_1__sbox_and_xor_inst_b_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_1__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_3__GEN_ROWS_1__sbox_and_xor_inst_b_nxy), .B0_t (StateFromRhoPi[51]), .Z0_t (StateFromChi[51]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_1__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[131]), .B0_t (StateFromRhoPi[171]), .Z0_t (CHI_GEN_SLICES_3__GEN_ROWS_1__sbox_and_xor_inst_c_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_1__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_3__GEN_ROWS_1__sbox_and_xor_inst_c_nxy), .B0_t (StateFromRhoPi[91]), .Z0_t (StateFromChi[91]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_1__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[171]), .B0_t (StateFromRhoPi[11]), .Z0_t (CHI_GEN_SLICES_3__GEN_ROWS_1__sbox_and_xor_inst_d_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_1__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_3__GEN_ROWS_1__sbox_and_xor_inst_d_nxy), .B0_t (StateFromRhoPi[131]), .Z0_t (StateFromChi[131]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_1__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[11]), .B0_t (StateFromRhoPi[51]), .Z0_t (CHI_GEN_SLICES_3__GEN_ROWS_1__sbox_and_xor_inst_e_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_1__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_3__GEN_ROWS_1__sbox_and_xor_inst_e_nxy), .B0_t (StateFromRhoPi[171]), .Z0_t (StateFromChi[171]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_2__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[59]), .B0_t (StateFromRhoPi[99]), .Z0_t (CHI_GEN_SLICES_3__GEN_ROWS_2__sbox_and_xor_inst_a_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_2__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_3__GEN_ROWS_2__sbox_and_xor_inst_a_nxy), .B0_t (StateFromRhoPi[19]), .Z0_t (StateFromChi[19]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_2__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[99]), .B0_t (StateFromRhoPi[139]), .Z0_t (CHI_GEN_SLICES_3__GEN_ROWS_2__sbox_and_xor_inst_b_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_2__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_3__GEN_ROWS_2__sbox_and_xor_inst_b_nxy), .B0_t (StateFromRhoPi[59]), .Z0_t (StateFromChi[59]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_2__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[139]), .B0_t (StateFromRhoPi[179]), .Z0_t (CHI_GEN_SLICES_3__GEN_ROWS_2__sbox_and_xor_inst_c_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_2__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_3__GEN_ROWS_2__sbox_and_xor_inst_c_nxy), .B0_t (StateFromRhoPi[99]), .Z0_t (StateFromChi[99]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_2__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[179]), .B0_t (StateFromRhoPi[19]), .Z0_t (CHI_GEN_SLICES_3__GEN_ROWS_2__sbox_and_xor_inst_d_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_2__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_3__GEN_ROWS_2__sbox_and_xor_inst_d_nxy), .B0_t (StateFromRhoPi[139]), .Z0_t (StateFromChi[139]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_2__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[19]), .B0_t (StateFromRhoPi[59]), .Z0_t (CHI_GEN_SLICES_3__GEN_ROWS_2__sbox_and_xor_inst_e_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_2__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_3__GEN_ROWS_2__sbox_and_xor_inst_e_nxy), .B0_t (StateFromRhoPi[179]), .Z0_t (StateFromChi[179]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_3__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[67]), .B0_t (StateFromRhoPi[107]), .Z0_t (CHI_GEN_SLICES_3__GEN_ROWS_3__sbox_and_xor_inst_a_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_3__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_3__GEN_ROWS_3__sbox_and_xor_inst_a_nxy), .B0_t (StateFromRhoPi[27]), .Z0_t (StateFromChi[27]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_3__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[107]), .B0_t (StateFromRhoPi[147]), .Z0_t (CHI_GEN_SLICES_3__GEN_ROWS_3__sbox_and_xor_inst_b_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_3__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_3__GEN_ROWS_3__sbox_and_xor_inst_b_nxy), .B0_t (StateFromRhoPi[67]), .Z0_t (StateFromChi[67]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_3__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[147]), .B0_t (StateFromRhoPi[187]), .Z0_t (CHI_GEN_SLICES_3__GEN_ROWS_3__sbox_and_xor_inst_c_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_3__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_3__GEN_ROWS_3__sbox_and_xor_inst_c_nxy), .B0_t (StateFromRhoPi[107]), .Z0_t (StateFromChi[107]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_3__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[187]), .B0_t (StateFromRhoPi[27]), .Z0_t (CHI_GEN_SLICES_3__GEN_ROWS_3__sbox_and_xor_inst_d_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_3__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_3__GEN_ROWS_3__sbox_and_xor_inst_d_nxy), .B0_t (StateFromRhoPi[147]), .Z0_t (StateFromChi[147]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_3__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[27]), .B0_t (StateFromRhoPi[67]), .Z0_t (CHI_GEN_SLICES_3__GEN_ROWS_3__sbox_and_xor_inst_e_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_3__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_3__GEN_ROWS_3__sbox_and_xor_inst_e_nxy), .B0_t (StateFromRhoPi[187]), .Z0_t (StateFromChi[187]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_4__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[75]), .B0_t (StateFromRhoPi[115]), .Z0_t (CHI_GEN_SLICES_3__GEN_ROWS_4__sbox_and_xor_inst_a_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_4__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_3__GEN_ROWS_4__sbox_and_xor_inst_a_nxy), .B0_t (StateFromRhoPi[35]), .Z0_t (StateFromChi[35]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_4__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[115]), .B0_t (StateFromRhoPi[155]), .Z0_t (CHI_GEN_SLICES_3__GEN_ROWS_4__sbox_and_xor_inst_b_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_4__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_3__GEN_ROWS_4__sbox_and_xor_inst_b_nxy), .B0_t (StateFromRhoPi[75]), .Z0_t (StateFromChi[75]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_4__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[155]), .B0_t (StateFromRhoPi[195]), .Z0_t (CHI_GEN_SLICES_3__GEN_ROWS_4__sbox_and_xor_inst_c_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_4__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_3__GEN_ROWS_4__sbox_and_xor_inst_c_nxy), .B0_t (StateFromRhoPi[115]), .Z0_t (StateFromChi[115]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_4__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[195]), .B0_t (StateFromRhoPi[35]), .Z0_t (CHI_GEN_SLICES_3__GEN_ROWS_4__sbox_and_xor_inst_d_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_4__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_3__GEN_ROWS_4__sbox_and_xor_inst_d_nxy), .B0_t (StateFromRhoPi[155]), .Z0_t (StateFromChi[155]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_4__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[35]), .B0_t (StateFromRhoPi[75]), .Z0_t (CHI_GEN_SLICES_3__GEN_ROWS_4__sbox_and_xor_inst_e_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_3__GEN_ROWS_4__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_3__GEN_ROWS_4__sbox_and_xor_inst_e_nxy), .B0_t (StateFromRhoPi[195]), .Z0_t (StateFromChi[195]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_0__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[44]), .B0_t (StateFromRhoPi[84]), .Z0_t (CHI_GEN_SLICES_4__GEN_ROWS_0__sbox_and_xor_inst_a_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_0__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_4__GEN_ROWS_0__sbox_and_xor_inst_a_nxy), .B0_t (StateFromRhoPi[4]), .Z0_t (StateFromChi[4]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_0__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[84]), .B0_t (StateFromRhoPi[124]), .Z0_t (CHI_GEN_SLICES_4__GEN_ROWS_0__sbox_and_xor_inst_b_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_0__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_4__GEN_ROWS_0__sbox_and_xor_inst_b_nxy), .B0_t (StateFromRhoPi[44]), .Z0_t (StateFromChi[44]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_0__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[124]), .B0_t (StateFromRhoPi[164]), .Z0_t (CHI_GEN_SLICES_4__GEN_ROWS_0__sbox_and_xor_inst_c_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_0__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_4__GEN_ROWS_0__sbox_and_xor_inst_c_nxy), .B0_t (StateFromRhoPi[84]), .Z0_t (StateFromChi[84]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_0__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[164]), .B0_t (StateFromRhoPi[4]), .Z0_t (CHI_GEN_SLICES_4__GEN_ROWS_0__sbox_and_xor_inst_d_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_0__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_4__GEN_ROWS_0__sbox_and_xor_inst_d_nxy), .B0_t (StateFromRhoPi[124]), .Z0_t (StateFromChi[124]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_0__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[4]), .B0_t (StateFromRhoPi[44]), .Z0_t (CHI_GEN_SLICES_4__GEN_ROWS_0__sbox_and_xor_inst_e_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_0__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_4__GEN_ROWS_0__sbox_and_xor_inst_e_nxy), .B0_t (StateFromRhoPi[164]), .Z0_t (StateFromChi[164]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_1__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[52]), .B0_t (StateFromRhoPi[92]), .Z0_t (CHI_GEN_SLICES_4__GEN_ROWS_1__sbox_and_xor_inst_a_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_1__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_4__GEN_ROWS_1__sbox_and_xor_inst_a_nxy), .B0_t (StateFromRhoPi[12]), .Z0_t (StateFromChi[12]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_1__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[92]), .B0_t (StateFromRhoPi[132]), .Z0_t (CHI_GEN_SLICES_4__GEN_ROWS_1__sbox_and_xor_inst_b_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_1__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_4__GEN_ROWS_1__sbox_and_xor_inst_b_nxy), .B0_t (StateFromRhoPi[52]), .Z0_t (StateFromChi[52]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_1__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[132]), .B0_t (StateFromRhoPi[172]), .Z0_t (CHI_GEN_SLICES_4__GEN_ROWS_1__sbox_and_xor_inst_c_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_1__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_4__GEN_ROWS_1__sbox_and_xor_inst_c_nxy), .B0_t (StateFromRhoPi[92]), .Z0_t (StateFromChi[92]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_1__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[172]), .B0_t (StateFromRhoPi[12]), .Z0_t (CHI_GEN_SLICES_4__GEN_ROWS_1__sbox_and_xor_inst_d_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_1__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_4__GEN_ROWS_1__sbox_and_xor_inst_d_nxy), .B0_t (StateFromRhoPi[132]), .Z0_t (StateFromChi[132]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_1__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[12]), .B0_t (StateFromRhoPi[52]), .Z0_t (CHI_GEN_SLICES_4__GEN_ROWS_1__sbox_and_xor_inst_e_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_1__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_4__GEN_ROWS_1__sbox_and_xor_inst_e_nxy), .B0_t (StateFromRhoPi[172]), .Z0_t (StateFromChi[172]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_2__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[60]), .B0_t (StateFromRhoPi[100]), .Z0_t (CHI_GEN_SLICES_4__GEN_ROWS_2__sbox_and_xor_inst_a_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_2__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_4__GEN_ROWS_2__sbox_and_xor_inst_a_nxy), .B0_t (StateFromRhoPi[20]), .Z0_t (StateFromChi[20]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_2__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[100]), .B0_t (StateFromRhoPi[140]), .Z0_t (CHI_GEN_SLICES_4__GEN_ROWS_2__sbox_and_xor_inst_b_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_2__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_4__GEN_ROWS_2__sbox_and_xor_inst_b_nxy), .B0_t (StateFromRhoPi[60]), .Z0_t (StateFromChi[60]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_2__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[140]), .B0_t (StateFromRhoPi[180]), .Z0_t (CHI_GEN_SLICES_4__GEN_ROWS_2__sbox_and_xor_inst_c_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_2__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_4__GEN_ROWS_2__sbox_and_xor_inst_c_nxy), .B0_t (StateFromRhoPi[100]), .Z0_t (StateFromChi[100]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_2__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[180]), .B0_t (StateFromRhoPi[20]), .Z0_t (CHI_GEN_SLICES_4__GEN_ROWS_2__sbox_and_xor_inst_d_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_2__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_4__GEN_ROWS_2__sbox_and_xor_inst_d_nxy), .B0_t (StateFromRhoPi[140]), .Z0_t (StateFromChi[140]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_2__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[20]), .B0_t (StateFromRhoPi[60]), .Z0_t (CHI_GEN_SLICES_4__GEN_ROWS_2__sbox_and_xor_inst_e_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_2__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_4__GEN_ROWS_2__sbox_and_xor_inst_e_nxy), .B0_t (StateFromRhoPi[180]), .Z0_t (StateFromChi[180]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_3__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[68]), .B0_t (StateFromRhoPi[108]), .Z0_t (CHI_GEN_SLICES_4__GEN_ROWS_3__sbox_and_xor_inst_a_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_3__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_4__GEN_ROWS_3__sbox_and_xor_inst_a_nxy), .B0_t (StateFromRhoPi[28]), .Z0_t (StateFromChi[28]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_3__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[108]), .B0_t (StateFromRhoPi[148]), .Z0_t (CHI_GEN_SLICES_4__GEN_ROWS_3__sbox_and_xor_inst_b_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_3__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_4__GEN_ROWS_3__sbox_and_xor_inst_b_nxy), .B0_t (StateFromRhoPi[68]), .Z0_t (StateFromChi[68]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_3__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[148]), .B0_t (StateFromRhoPi[188]), .Z0_t (CHI_GEN_SLICES_4__GEN_ROWS_3__sbox_and_xor_inst_c_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_3__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_4__GEN_ROWS_3__sbox_and_xor_inst_c_nxy), .B0_t (StateFromRhoPi[108]), .Z0_t (StateFromChi[108]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_3__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[188]), .B0_t (StateFromRhoPi[28]), .Z0_t (CHI_GEN_SLICES_4__GEN_ROWS_3__sbox_and_xor_inst_d_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_3__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_4__GEN_ROWS_3__sbox_and_xor_inst_d_nxy), .B0_t (StateFromRhoPi[148]), .Z0_t (StateFromChi[148]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_3__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[28]), .B0_t (StateFromRhoPi[68]), .Z0_t (CHI_GEN_SLICES_4__GEN_ROWS_3__sbox_and_xor_inst_e_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_3__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_4__GEN_ROWS_3__sbox_and_xor_inst_e_nxy), .B0_t (StateFromRhoPi[188]), .Z0_t (StateFromChi[188]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_4__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[76]), .B0_t (StateFromRhoPi[116]), .Z0_t (CHI_GEN_SLICES_4__GEN_ROWS_4__sbox_and_xor_inst_a_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_4__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_4__GEN_ROWS_4__sbox_and_xor_inst_a_nxy), .B0_t (StateFromRhoPi[36]), .Z0_t (StateFromChi[36]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_4__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[116]), .B0_t (StateFromRhoPi[156]), .Z0_t (CHI_GEN_SLICES_4__GEN_ROWS_4__sbox_and_xor_inst_b_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_4__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_4__GEN_ROWS_4__sbox_and_xor_inst_b_nxy), .B0_t (StateFromRhoPi[76]), .Z0_t (StateFromChi[76]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_4__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[156]), .B0_t (StateFromRhoPi[196]), .Z0_t (CHI_GEN_SLICES_4__GEN_ROWS_4__sbox_and_xor_inst_c_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_4__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_4__GEN_ROWS_4__sbox_and_xor_inst_c_nxy), .B0_t (StateFromRhoPi[116]), .Z0_t (StateFromChi[116]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_4__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[196]), .B0_t (StateFromRhoPi[36]), .Z0_t (CHI_GEN_SLICES_4__GEN_ROWS_4__sbox_and_xor_inst_d_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_4__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_4__GEN_ROWS_4__sbox_and_xor_inst_d_nxy), .B0_t (StateFromRhoPi[156]), .Z0_t (StateFromChi[156]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_4__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[36]), .B0_t (StateFromRhoPi[76]), .Z0_t (CHI_GEN_SLICES_4__GEN_ROWS_4__sbox_and_xor_inst_e_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_4__GEN_ROWS_4__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_4__GEN_ROWS_4__sbox_and_xor_inst_e_nxy), .B0_t (StateFromRhoPi[196]), .Z0_t (StateFromChi[196]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_0__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[45]), .B0_t (StateFromRhoPi[85]), .Z0_t (CHI_GEN_SLICES_5__GEN_ROWS_0__sbox_and_xor_inst_a_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_0__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_5__GEN_ROWS_0__sbox_and_xor_inst_a_nxy), .B0_t (StateFromRhoPi[5]), .Z0_t (StateFromChi[5]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_0__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[85]), .B0_t (StateFromRhoPi[125]), .Z0_t (CHI_GEN_SLICES_5__GEN_ROWS_0__sbox_and_xor_inst_b_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_0__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_5__GEN_ROWS_0__sbox_and_xor_inst_b_nxy), .B0_t (StateFromRhoPi[45]), .Z0_t (StateFromChi[45]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_0__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[125]), .B0_t (StateFromRhoPi[165]), .Z0_t (CHI_GEN_SLICES_5__GEN_ROWS_0__sbox_and_xor_inst_c_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_0__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_5__GEN_ROWS_0__sbox_and_xor_inst_c_nxy), .B0_t (StateFromRhoPi[85]), .Z0_t (StateFromChi[85]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_0__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[165]), .B0_t (StateFromRhoPi[5]), .Z0_t (CHI_GEN_SLICES_5__GEN_ROWS_0__sbox_and_xor_inst_d_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_0__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_5__GEN_ROWS_0__sbox_and_xor_inst_d_nxy), .B0_t (StateFromRhoPi[125]), .Z0_t (StateFromChi[125]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_0__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[5]), .B0_t (StateFromRhoPi[45]), .Z0_t (CHI_GEN_SLICES_5__GEN_ROWS_0__sbox_and_xor_inst_e_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_0__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_5__GEN_ROWS_0__sbox_and_xor_inst_e_nxy), .B0_t (StateFromRhoPi[165]), .Z0_t (StateFromChi[165]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_1__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[53]), .B0_t (StateFromRhoPi[93]), .Z0_t (CHI_GEN_SLICES_5__GEN_ROWS_1__sbox_and_xor_inst_a_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_1__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_5__GEN_ROWS_1__sbox_and_xor_inst_a_nxy), .B0_t (StateFromRhoPi[13]), .Z0_t (StateFromChi[13]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_1__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[93]), .B0_t (StateFromRhoPi[133]), .Z0_t (CHI_GEN_SLICES_5__GEN_ROWS_1__sbox_and_xor_inst_b_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_1__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_5__GEN_ROWS_1__sbox_and_xor_inst_b_nxy), .B0_t (StateFromRhoPi[53]), .Z0_t (StateFromChi[53]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_1__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[133]), .B0_t (StateFromRhoPi[173]), .Z0_t (CHI_GEN_SLICES_5__GEN_ROWS_1__sbox_and_xor_inst_c_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_1__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_5__GEN_ROWS_1__sbox_and_xor_inst_c_nxy), .B0_t (StateFromRhoPi[93]), .Z0_t (StateFromChi[93]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_1__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[173]), .B0_t (StateFromRhoPi[13]), .Z0_t (CHI_GEN_SLICES_5__GEN_ROWS_1__sbox_and_xor_inst_d_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_1__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_5__GEN_ROWS_1__sbox_and_xor_inst_d_nxy), .B0_t (StateFromRhoPi[133]), .Z0_t (StateFromChi[133]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_1__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[13]), .B0_t (StateFromRhoPi[53]), .Z0_t (CHI_GEN_SLICES_5__GEN_ROWS_1__sbox_and_xor_inst_e_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_1__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_5__GEN_ROWS_1__sbox_and_xor_inst_e_nxy), .B0_t (StateFromRhoPi[173]), .Z0_t (StateFromChi[173]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_2__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[61]), .B0_t (StateFromRhoPi[101]), .Z0_t (CHI_GEN_SLICES_5__GEN_ROWS_2__sbox_and_xor_inst_a_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_2__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_5__GEN_ROWS_2__sbox_and_xor_inst_a_nxy), .B0_t (StateFromRhoPi[21]), .Z0_t (StateFromChi[21]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_2__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[101]), .B0_t (StateFromRhoPi[141]), .Z0_t (CHI_GEN_SLICES_5__GEN_ROWS_2__sbox_and_xor_inst_b_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_2__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_5__GEN_ROWS_2__sbox_and_xor_inst_b_nxy), .B0_t (StateFromRhoPi[61]), .Z0_t (StateFromChi[61]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_2__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[141]), .B0_t (StateFromRhoPi[181]), .Z0_t (CHI_GEN_SLICES_5__GEN_ROWS_2__sbox_and_xor_inst_c_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_2__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_5__GEN_ROWS_2__sbox_and_xor_inst_c_nxy), .B0_t (StateFromRhoPi[101]), .Z0_t (StateFromChi[101]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_2__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[181]), .B0_t (StateFromRhoPi[21]), .Z0_t (CHI_GEN_SLICES_5__GEN_ROWS_2__sbox_and_xor_inst_d_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_2__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_5__GEN_ROWS_2__sbox_and_xor_inst_d_nxy), .B0_t (StateFromRhoPi[141]), .Z0_t (StateFromChi[141]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_2__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[21]), .B0_t (StateFromRhoPi[61]), .Z0_t (CHI_GEN_SLICES_5__GEN_ROWS_2__sbox_and_xor_inst_e_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_2__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_5__GEN_ROWS_2__sbox_and_xor_inst_e_nxy), .B0_t (StateFromRhoPi[181]), .Z0_t (StateFromChi[181]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_3__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[69]), .B0_t (StateFromRhoPi[109]), .Z0_t (CHI_GEN_SLICES_5__GEN_ROWS_3__sbox_and_xor_inst_a_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_3__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_5__GEN_ROWS_3__sbox_and_xor_inst_a_nxy), .B0_t (StateFromRhoPi[29]), .Z0_t (StateFromChi[29]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_3__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[109]), .B0_t (StateFromRhoPi[149]), .Z0_t (CHI_GEN_SLICES_5__GEN_ROWS_3__sbox_and_xor_inst_b_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_3__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_5__GEN_ROWS_3__sbox_and_xor_inst_b_nxy), .B0_t (StateFromRhoPi[69]), .Z0_t (StateFromChi[69]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_3__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[149]), .B0_t (StateFromRhoPi[189]), .Z0_t (CHI_GEN_SLICES_5__GEN_ROWS_3__sbox_and_xor_inst_c_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_3__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_5__GEN_ROWS_3__sbox_and_xor_inst_c_nxy), .B0_t (StateFromRhoPi[109]), .Z0_t (StateFromChi[109]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_3__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[189]), .B0_t (StateFromRhoPi[29]), .Z0_t (CHI_GEN_SLICES_5__GEN_ROWS_3__sbox_and_xor_inst_d_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_3__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_5__GEN_ROWS_3__sbox_and_xor_inst_d_nxy), .B0_t (StateFromRhoPi[149]), .Z0_t (StateFromChi[149]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_3__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[29]), .B0_t (StateFromRhoPi[69]), .Z0_t (CHI_GEN_SLICES_5__GEN_ROWS_3__sbox_and_xor_inst_e_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_3__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_5__GEN_ROWS_3__sbox_and_xor_inst_e_nxy), .B0_t (StateFromRhoPi[189]), .Z0_t (StateFromChi[189]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_4__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[77]), .B0_t (StateFromRhoPi[117]), .Z0_t (CHI_GEN_SLICES_5__GEN_ROWS_4__sbox_and_xor_inst_a_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_4__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_5__GEN_ROWS_4__sbox_and_xor_inst_a_nxy), .B0_t (StateFromRhoPi[37]), .Z0_t (StateFromChi[37]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_4__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[117]), .B0_t (StateFromRhoPi[157]), .Z0_t (CHI_GEN_SLICES_5__GEN_ROWS_4__sbox_and_xor_inst_b_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_4__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_5__GEN_ROWS_4__sbox_and_xor_inst_b_nxy), .B0_t (StateFromRhoPi[77]), .Z0_t (StateFromChi[77]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_4__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[157]), .B0_t (StateFromRhoPi[197]), .Z0_t (CHI_GEN_SLICES_5__GEN_ROWS_4__sbox_and_xor_inst_c_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_4__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_5__GEN_ROWS_4__sbox_and_xor_inst_c_nxy), .B0_t (StateFromRhoPi[117]), .Z0_t (StateFromChi[117]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_4__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[197]), .B0_t (StateFromRhoPi[37]), .Z0_t (CHI_GEN_SLICES_5__GEN_ROWS_4__sbox_and_xor_inst_d_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_4__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_5__GEN_ROWS_4__sbox_and_xor_inst_d_nxy), .B0_t (StateFromRhoPi[157]), .Z0_t (StateFromChi[157]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_4__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[37]), .B0_t (StateFromRhoPi[77]), .Z0_t (CHI_GEN_SLICES_5__GEN_ROWS_4__sbox_and_xor_inst_e_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_5__GEN_ROWS_4__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_5__GEN_ROWS_4__sbox_and_xor_inst_e_nxy), .B0_t (StateFromRhoPi[197]), .Z0_t (StateFromChi[197]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_0__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[46]), .B0_t (StateFromRhoPi[86]), .Z0_t (CHI_GEN_SLICES_6__GEN_ROWS_0__sbox_and_xor_inst_a_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_0__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_6__GEN_ROWS_0__sbox_and_xor_inst_a_nxy), .B0_t (StateFromRhoPi[6]), .Z0_t (StateFromChi[6]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_0__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[86]), .B0_t (StateFromRhoPi[126]), .Z0_t (CHI_GEN_SLICES_6__GEN_ROWS_0__sbox_and_xor_inst_b_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_0__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_6__GEN_ROWS_0__sbox_and_xor_inst_b_nxy), .B0_t (StateFromRhoPi[46]), .Z0_t (StateFromChi[46]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_0__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[126]), .B0_t (StateFromRhoPi[166]), .Z0_t (CHI_GEN_SLICES_6__GEN_ROWS_0__sbox_and_xor_inst_c_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_0__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_6__GEN_ROWS_0__sbox_and_xor_inst_c_nxy), .B0_t (StateFromRhoPi[86]), .Z0_t (StateFromChi[86]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_0__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[166]), .B0_t (StateFromRhoPi[6]), .Z0_t (CHI_GEN_SLICES_6__GEN_ROWS_0__sbox_and_xor_inst_d_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_0__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_6__GEN_ROWS_0__sbox_and_xor_inst_d_nxy), .B0_t (StateFromRhoPi[126]), .Z0_t (StateFromChi[126]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_0__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[6]), .B0_t (StateFromRhoPi[46]), .Z0_t (CHI_GEN_SLICES_6__GEN_ROWS_0__sbox_and_xor_inst_e_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_0__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_6__GEN_ROWS_0__sbox_and_xor_inst_e_nxy), .B0_t (StateFromRhoPi[166]), .Z0_t (StateFromChi[166]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_1__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[54]), .B0_t (StateFromRhoPi[94]), .Z0_t (CHI_GEN_SLICES_6__GEN_ROWS_1__sbox_and_xor_inst_a_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_1__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_6__GEN_ROWS_1__sbox_and_xor_inst_a_nxy), .B0_t (StateFromRhoPi[14]), .Z0_t (StateFromChi[14]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_1__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[94]), .B0_t (StateFromRhoPi[134]), .Z0_t (CHI_GEN_SLICES_6__GEN_ROWS_1__sbox_and_xor_inst_b_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_1__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_6__GEN_ROWS_1__sbox_and_xor_inst_b_nxy), .B0_t (StateFromRhoPi[54]), .Z0_t (StateFromChi[54]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_1__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[134]), .B0_t (StateFromRhoPi[174]), .Z0_t (CHI_GEN_SLICES_6__GEN_ROWS_1__sbox_and_xor_inst_c_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_1__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_6__GEN_ROWS_1__sbox_and_xor_inst_c_nxy), .B0_t (StateFromRhoPi[94]), .Z0_t (StateFromChi[94]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_1__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[174]), .B0_t (StateFromRhoPi[14]), .Z0_t (CHI_GEN_SLICES_6__GEN_ROWS_1__sbox_and_xor_inst_d_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_1__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_6__GEN_ROWS_1__sbox_and_xor_inst_d_nxy), .B0_t (StateFromRhoPi[134]), .Z0_t (StateFromChi[134]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_1__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[14]), .B0_t (StateFromRhoPi[54]), .Z0_t (CHI_GEN_SLICES_6__GEN_ROWS_1__sbox_and_xor_inst_e_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_1__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_6__GEN_ROWS_1__sbox_and_xor_inst_e_nxy), .B0_t (StateFromRhoPi[174]), .Z0_t (StateFromChi[174]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_2__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[62]), .B0_t (StateFromRhoPi[102]), .Z0_t (CHI_GEN_SLICES_6__GEN_ROWS_2__sbox_and_xor_inst_a_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_2__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_6__GEN_ROWS_2__sbox_and_xor_inst_a_nxy), .B0_t (StateFromRhoPi[22]), .Z0_t (StateFromChi[22]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_2__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[102]), .B0_t (StateFromRhoPi[142]), .Z0_t (CHI_GEN_SLICES_6__GEN_ROWS_2__sbox_and_xor_inst_b_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_2__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_6__GEN_ROWS_2__sbox_and_xor_inst_b_nxy), .B0_t (StateFromRhoPi[62]), .Z0_t (StateFromChi[62]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_2__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[142]), .B0_t (StateFromRhoPi[182]), .Z0_t (CHI_GEN_SLICES_6__GEN_ROWS_2__sbox_and_xor_inst_c_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_2__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_6__GEN_ROWS_2__sbox_and_xor_inst_c_nxy), .B0_t (StateFromRhoPi[102]), .Z0_t (StateFromChi[102]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_2__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[182]), .B0_t (StateFromRhoPi[22]), .Z0_t (CHI_GEN_SLICES_6__GEN_ROWS_2__sbox_and_xor_inst_d_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_2__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_6__GEN_ROWS_2__sbox_and_xor_inst_d_nxy), .B0_t (StateFromRhoPi[142]), .Z0_t (StateFromChi[142]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_2__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[22]), .B0_t (StateFromRhoPi[62]), .Z0_t (CHI_GEN_SLICES_6__GEN_ROWS_2__sbox_and_xor_inst_e_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_2__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_6__GEN_ROWS_2__sbox_and_xor_inst_e_nxy), .B0_t (StateFromRhoPi[182]), .Z0_t (StateFromChi[182]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_3__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[70]), .B0_t (StateFromRhoPi[110]), .Z0_t (CHI_GEN_SLICES_6__GEN_ROWS_3__sbox_and_xor_inst_a_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_3__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_6__GEN_ROWS_3__sbox_and_xor_inst_a_nxy), .B0_t (StateFromRhoPi[30]), .Z0_t (StateFromChi[30]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_3__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[110]), .B0_t (StateFromRhoPi[150]), .Z0_t (CHI_GEN_SLICES_6__GEN_ROWS_3__sbox_and_xor_inst_b_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_3__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_6__GEN_ROWS_3__sbox_and_xor_inst_b_nxy), .B0_t (StateFromRhoPi[70]), .Z0_t (StateFromChi[70]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_3__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[150]), .B0_t (StateFromRhoPi[190]), .Z0_t (CHI_GEN_SLICES_6__GEN_ROWS_3__sbox_and_xor_inst_c_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_3__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_6__GEN_ROWS_3__sbox_and_xor_inst_c_nxy), .B0_t (StateFromRhoPi[110]), .Z0_t (StateFromChi[110]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_3__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[190]), .B0_t (StateFromRhoPi[30]), .Z0_t (CHI_GEN_SLICES_6__GEN_ROWS_3__sbox_and_xor_inst_d_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_3__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_6__GEN_ROWS_3__sbox_and_xor_inst_d_nxy), .B0_t (StateFromRhoPi[150]), .Z0_t (StateFromChi[150]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_3__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[30]), .B0_t (StateFromRhoPi[70]), .Z0_t (CHI_GEN_SLICES_6__GEN_ROWS_3__sbox_and_xor_inst_e_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_3__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_6__GEN_ROWS_3__sbox_and_xor_inst_e_nxy), .B0_t (StateFromRhoPi[190]), .Z0_t (StateFromChi[190]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_4__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[78]), .B0_t (StateFromRhoPi[118]), .Z0_t (CHI_GEN_SLICES_6__GEN_ROWS_4__sbox_and_xor_inst_a_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_4__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_6__GEN_ROWS_4__sbox_and_xor_inst_a_nxy), .B0_t (StateFromRhoPi[38]), .Z0_t (StateFromChi[38]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_4__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[118]), .B0_t (StateFromRhoPi[158]), .Z0_t (CHI_GEN_SLICES_6__GEN_ROWS_4__sbox_and_xor_inst_b_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_4__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_6__GEN_ROWS_4__sbox_and_xor_inst_b_nxy), .B0_t (StateFromRhoPi[78]), .Z0_t (StateFromChi[78]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_4__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[158]), .B0_t (StateFromRhoPi[198]), .Z0_t (CHI_GEN_SLICES_6__GEN_ROWS_4__sbox_and_xor_inst_c_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_4__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_6__GEN_ROWS_4__sbox_and_xor_inst_c_nxy), .B0_t (StateFromRhoPi[118]), .Z0_t (StateFromChi[118]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_4__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[198]), .B0_t (StateFromRhoPi[38]), .Z0_t (CHI_GEN_SLICES_6__GEN_ROWS_4__sbox_and_xor_inst_d_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_4__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_6__GEN_ROWS_4__sbox_and_xor_inst_d_nxy), .B0_t (StateFromRhoPi[158]), .Z0_t (StateFromChi[158]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_4__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[38]), .B0_t (StateFromRhoPi[78]), .Z0_t (CHI_GEN_SLICES_6__GEN_ROWS_4__sbox_and_xor_inst_e_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_6__GEN_ROWS_4__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_6__GEN_ROWS_4__sbox_and_xor_inst_e_nxy), .B0_t (StateFromRhoPi[198]), .Z0_t (StateFromChi[198]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_0__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[47]), .B0_t (StateFromRhoPi[87]), .Z0_t (CHI_GEN_SLICES_7__GEN_ROWS_0__sbox_and_xor_inst_a_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_0__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_7__GEN_ROWS_0__sbox_and_xor_inst_a_nxy), .B0_t (StateFromRhoPi[7]), .Z0_t (CHI_ChiOut_7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_0__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[87]), .B0_t (StateFromRhoPi[127]), .Z0_t (CHI_GEN_SLICES_7__GEN_ROWS_0__sbox_and_xor_inst_b_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_0__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_7__GEN_ROWS_0__sbox_and_xor_inst_b_nxy), .B0_t (StateFromRhoPi[47]), .Z0_t (StateFromChi[47]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_0__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[127]), .B0_t (StateFromRhoPi[167]), .Z0_t (CHI_GEN_SLICES_7__GEN_ROWS_0__sbox_and_xor_inst_c_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_0__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_7__GEN_ROWS_0__sbox_and_xor_inst_c_nxy), .B0_t (StateFromRhoPi[87]), .Z0_t (StateFromChi[87]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_0__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[167]), .B0_t (StateFromRhoPi[7]), .Z0_t (CHI_GEN_SLICES_7__GEN_ROWS_0__sbox_and_xor_inst_d_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_0__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_7__GEN_ROWS_0__sbox_and_xor_inst_d_nxy), .B0_t (StateFromRhoPi[127]), .Z0_t (StateFromChi[127]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_0__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[7]), .B0_t (StateFromRhoPi[47]), .Z0_t (CHI_GEN_SLICES_7__GEN_ROWS_0__sbox_and_xor_inst_e_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_0__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_7__GEN_ROWS_0__sbox_and_xor_inst_e_nxy), .B0_t (StateFromRhoPi[167]), .Z0_t (StateFromChi[167]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_1__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[55]), .B0_t (StateFromRhoPi[95]), .Z0_t (CHI_GEN_SLICES_7__GEN_ROWS_1__sbox_and_xor_inst_a_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_1__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_7__GEN_ROWS_1__sbox_and_xor_inst_a_nxy), .B0_t (StateFromRhoPi[15]), .Z0_t (StateFromChi[15]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_1__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[95]), .B0_t (StateFromRhoPi[135]), .Z0_t (CHI_GEN_SLICES_7__GEN_ROWS_1__sbox_and_xor_inst_b_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_1__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_7__GEN_ROWS_1__sbox_and_xor_inst_b_nxy), .B0_t (StateFromRhoPi[55]), .Z0_t (StateFromChi[55]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_1__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[135]), .B0_t (StateFromRhoPi[175]), .Z0_t (CHI_GEN_SLICES_7__GEN_ROWS_1__sbox_and_xor_inst_c_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_1__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_7__GEN_ROWS_1__sbox_and_xor_inst_c_nxy), .B0_t (StateFromRhoPi[95]), .Z0_t (StateFromChi[95]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_1__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[175]), .B0_t (StateFromRhoPi[15]), .Z0_t (CHI_GEN_SLICES_7__GEN_ROWS_1__sbox_and_xor_inst_d_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_1__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_7__GEN_ROWS_1__sbox_and_xor_inst_d_nxy), .B0_t (StateFromRhoPi[135]), .Z0_t (StateFromChi[135]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_1__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[15]), .B0_t (StateFromRhoPi[55]), .Z0_t (CHI_GEN_SLICES_7__GEN_ROWS_1__sbox_and_xor_inst_e_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_1__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_7__GEN_ROWS_1__sbox_and_xor_inst_e_nxy), .B0_t (StateFromRhoPi[175]), .Z0_t (StateFromChi[175]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_2__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[63]), .B0_t (StateFromRhoPi[103]), .Z0_t (CHI_GEN_SLICES_7__GEN_ROWS_2__sbox_and_xor_inst_a_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_2__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_7__GEN_ROWS_2__sbox_and_xor_inst_a_nxy), .B0_t (StateFromRhoPi[23]), .Z0_t (StateFromChi[23]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_2__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[103]), .B0_t (StateFromRhoPi[143]), .Z0_t (CHI_GEN_SLICES_7__GEN_ROWS_2__sbox_and_xor_inst_b_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_2__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_7__GEN_ROWS_2__sbox_and_xor_inst_b_nxy), .B0_t (StateFromRhoPi[63]), .Z0_t (StateFromChi[63]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_2__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[143]), .B0_t (StateFromRhoPi[183]), .Z0_t (CHI_GEN_SLICES_7__GEN_ROWS_2__sbox_and_xor_inst_c_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_2__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_7__GEN_ROWS_2__sbox_and_xor_inst_c_nxy), .B0_t (StateFromRhoPi[103]), .Z0_t (StateFromChi[103]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_2__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[183]), .B0_t (StateFromRhoPi[23]), .Z0_t (CHI_GEN_SLICES_7__GEN_ROWS_2__sbox_and_xor_inst_d_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_2__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_7__GEN_ROWS_2__sbox_and_xor_inst_d_nxy), .B0_t (StateFromRhoPi[143]), .Z0_t (StateFromChi[143]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_2__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[23]), .B0_t (StateFromRhoPi[63]), .Z0_t (CHI_GEN_SLICES_7__GEN_ROWS_2__sbox_and_xor_inst_e_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_2__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_7__GEN_ROWS_2__sbox_and_xor_inst_e_nxy), .B0_t (StateFromRhoPi[183]), .Z0_t (StateFromChi[183]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_3__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[71]), .B0_t (StateFromRhoPi[111]), .Z0_t (CHI_GEN_SLICES_7__GEN_ROWS_3__sbox_and_xor_inst_a_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_3__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_7__GEN_ROWS_3__sbox_and_xor_inst_a_nxy), .B0_t (StateFromRhoPi[31]), .Z0_t (StateFromChi[31]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_3__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[111]), .B0_t (StateFromRhoPi[151]), .Z0_t (CHI_GEN_SLICES_7__GEN_ROWS_3__sbox_and_xor_inst_b_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_3__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_7__GEN_ROWS_3__sbox_and_xor_inst_b_nxy), .B0_t (StateFromRhoPi[71]), .Z0_t (StateFromChi[71]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_3__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[151]), .B0_t (StateFromRhoPi[191]), .Z0_t (CHI_GEN_SLICES_7__GEN_ROWS_3__sbox_and_xor_inst_c_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_3__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_7__GEN_ROWS_3__sbox_and_xor_inst_c_nxy), .B0_t (StateFromRhoPi[111]), .Z0_t (StateFromChi[111]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_3__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[191]), .B0_t (StateFromRhoPi[31]), .Z0_t (CHI_GEN_SLICES_7__GEN_ROWS_3__sbox_and_xor_inst_d_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_3__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_7__GEN_ROWS_3__sbox_and_xor_inst_d_nxy), .B0_t (StateFromRhoPi[151]), .Z0_t (StateFromChi[151]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_3__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[31]), .B0_t (StateFromRhoPi[71]), .Z0_t (CHI_GEN_SLICES_7__GEN_ROWS_3__sbox_and_xor_inst_e_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_3__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_7__GEN_ROWS_3__sbox_and_xor_inst_e_nxy), .B0_t (StateFromRhoPi[191]), .Z0_t (StateFromChi[191]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_4__sbox_and_xor_inst_a_instA_U1 ( .A0_t (StateFromRhoPi[79]), .B0_t (StateFromRhoPi[119]), .Z0_t (CHI_GEN_SLICES_7__GEN_ROWS_4__sbox_and_xor_inst_a_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_4__sbox_and_xor_inst_a_instX_U1 ( .A0_t (CHI_GEN_SLICES_7__GEN_ROWS_4__sbox_and_xor_inst_a_nxy), .B0_t (StateFromRhoPi[39]), .Z0_t (StateFromChi[39]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_4__sbox_and_xor_inst_b_instA_U1 ( .A0_t (StateFromRhoPi[119]), .B0_t (StateFromRhoPi[159]), .Z0_t (CHI_GEN_SLICES_7__GEN_ROWS_4__sbox_and_xor_inst_b_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_4__sbox_and_xor_inst_b_instX_U1 ( .A0_t (CHI_GEN_SLICES_7__GEN_ROWS_4__sbox_and_xor_inst_b_nxy), .B0_t (StateFromRhoPi[79]), .Z0_t (StateFromChi[79]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_4__sbox_and_xor_inst_c_instA_U1 ( .A0_t (StateFromRhoPi[159]), .B0_t (StateFromRhoPi[199]), .Z0_t (CHI_GEN_SLICES_7__GEN_ROWS_4__sbox_and_xor_inst_c_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_4__sbox_and_xor_inst_c_instX_U1 ( .A0_t (CHI_GEN_SLICES_7__GEN_ROWS_4__sbox_and_xor_inst_c_nxy), .B0_t (StateFromRhoPi[119]), .Z0_t (StateFromChi[119]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_4__sbox_and_xor_inst_d_instA_U1 ( .A0_t (StateFromRhoPi[199]), .B0_t (StateFromRhoPi[39]), .Z0_t (CHI_GEN_SLICES_7__GEN_ROWS_4__sbox_and_xor_inst_d_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_4__sbox_and_xor_inst_d_instX_U1 ( .A0_t (CHI_GEN_SLICES_7__GEN_ROWS_4__sbox_and_xor_inst_d_nxy), .B0_t (StateFromRhoPi[159]), .Z0_t (StateFromChi[159]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_4__sbox_and_xor_inst_e_instA_U1 ( .A0_t (StateFromRhoPi[39]), .B0_t (StateFromRhoPi[79]), .Z0_t (CHI_GEN_SLICES_7__GEN_ROWS_4__sbox_and_xor_inst_e_nxy) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) CHI_GEN_SLICES_7__GEN_ROWS_4__sbox_and_xor_inst_e_instX_U1 ( .A0_t (CHI_GEN_SLICES_7__GEN_ROWS_4__sbox_and_xor_inst_e_nxy), .B0_t (StateFromRhoPi[199]), .Z0_t (StateFromChi[199]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b1), .NL(1'b1)) KECCAK_CONTROL_U42 ( .A0_t (KECCAK_CONTROL_n47), .B0_t (Reset), .Z0_t (KECCAK_CONTROL_CtrlStatexDP[0]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_U41 ( .A0_t (KECCAK_CONTROL_n45), .B0_t (KECCAK_CONTROL_CtrlStatexDP[0]), .Z0_t (KECCAK_CONTROL_n47) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_U40 ( .A0_t (KECCAK_CONTROL_CtrlStatexDP_reg_1__Q), .B0_t (KECCAK_CONTROL_CtrlStatexDP[2]), .Z0_t (KECCAK_CONTROL_n45) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) KECCAK_CONTROL_U39 ( .A0_t (Reset), .B0_t (KECCAK_CONTROL_n44), .Z0_t (KECCAK_CONTROL_RoundCountxDP[4]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b0)) KECCAK_CONTROL_U38 ( .A0_t (KECCAK_CONTROL_RoundCountxDP[4]), .B0_t (KECCAK_CONTROL_n43), .Z0_t (KECCAK_CONTROL_n44) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) KECCAK_CONTROL_U37 ( .A0_t (KECCAK_CONTROL_RoundCountxDP[4]), .B0_t (KECCAK_CONTROL_n34), .Z0_t (KECCAK_CONTROL_RoundCountLastxDP_reg_Q) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_U36 ( .A0_t (Reset), .B0_t (KECCAK_CONTROL_n33), .Z0_t (KECCAK_CONTROL_n34) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_U35 ( .A0_t (KECCAK_CONTROL_n32), .B0_t (KECCAK_CONTROL_RoundCountxDP[1]), .Z0_t (KECCAK_CONTROL_n33) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_U34 ( .A0_t (KECCAK_CONTROL_RoundCountxDP[0]), .B0_t (KECCAK_CONTROL_n30), .Z0_t (KECCAK_CONTROL_n32) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) KECCAK_CONTROL_U33 ( .A0_t (Reset), .B0_t (KECCAK_CONTROL_n29), .Z0_t (KECCAK_CONTROL_CtrlStatexDP[2]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_U32 ( .A0_t (KECCAK_CONTROL_CtrlStatexDP[2]), .B0_t (KECCAK_CONTROL_n28), .Z0_t (KECCAK_CONTROL_n29) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_U31 ( .A0_t (KECCAK_CONTROL_n27), .B0_t (KECCAK_CONTROL_RoundCountLastxDP_reg_Q), .Z0_t (KECCAK_CONTROL_n28) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_U30 ( .A0_t (KECCAK_CONTROL_CtrlStatexDP[0]), .B0_t (KECCAK_CONTROL_CtrlStatexDP_reg_1__Q), .Z0_t (KECCAK_CONTROL_n27) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) KECCAK_CONTROL_U29 ( .A0_t (Reset), .B0_t (KECCAK_CONTROL_n25), .Z0_t (KECCAK_CONTROL_RoundCountxDP[2]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b0)) KECCAK_CONTROL_U28 ( .A0_t (KECCAK_CONTROL_RoundCountxDP[2]), .B0_t (KECCAK_CONTROL_n23), .Z0_t (KECCAK_CONTROL_n25) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) KECCAK_CONTROL_U27 ( .A0_t (Reset), .B0_t (KECCAK_CONTROL_n22), .Z0_t (KECCAK_CONTROL_CtrlStatexDP_reg_1__Q) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_U26 ( .A0_t (KECCAK_CONTROL_n21), .B0_t (KECCAK_CONTROL_n20), .Z0_t (KECCAK_CONTROL_n22) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_U25 ( .A0_t (KECCAK_CONTROL_CtrlStatexDP[2]), .B0_t (KECCAK_CONTROL_CtrlStatexDP[0]), .Z0_t (KECCAK_CONTROL_n20) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_U24 ( .A0_t (KECCAK_CONTROL_CtrlStatexDP_reg_1__Q), .B0_t (KECCAK_CONTROL_n19), .Z0_t (KECCAK_CONTROL_n21) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_U23 ( .A0_t (KECCAK_CONTROL_CtrlStatexDP[2]), .B0_t (KECCAK_CONTROL_RoundCountLastxDP_reg_Q), .Z0_t (KECCAK_CONTROL_n19) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) KECCAK_CONTROL_U22 ( .A0_t (Reset), .B0_t (KECCAK_CONTROL_n18), .Z0_t (KECCAK_CONTROL_RoundCountxDP[1]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) KECCAK_CONTROL_U21 ( .A0_t (KECCAK_CONTROL_n17), .B0_t (KECCAK_CONTROL_RoundCountxDP[1]), .Z0_t (KECCAK_CONTROL_n18) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) KECCAK_CONTROL_U20 ( .A0_t (KECCAK_CONTROL_n16), .B0_t (KECCAK_CONTROL_n15), .Z0_t (KECCAK_CONTROL_RoundCountxDP[3]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_U19 ( .A0_t (KECCAK_CONTROL_RoundCountxDP[3]), .B0_t (KECCAK_CONTROL_n14), .Z0_t (KECCAK_CONTROL_n15) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_U18 ( .A0_t (KECCAK_CONTROL_RoundCountxDP[2]), .B0_t (KECCAK_CONTROL_n23), .Z0_t (KECCAK_CONTROL_n14) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_U16 ( .A0_t (Reset), .B0_t (KECCAK_CONTROL_n43), .Z0_t (KECCAK_CONTROL_n16) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_U15 ( .A0_t (KECCAK_CONTROL_n30), .B0_t (KECCAK_CONTROL_n23), .Z0_t (KECCAK_CONTROL_n43) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_U14 ( .A0_t (KECCAK_CONTROL_n17), .B0_t (KECCAK_CONTROL_RoundCountxDP[1]), .Z0_t (KECCAK_CONTROL_n23) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_U12 ( .A0_t (KECCAK_CONTROL_n13), .B0_t (KECCAK_CONTROL_RoundCountxDP[0]), .Z0_t (KECCAK_CONTROL_n17) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_U11 ( .A0_t (KECCAK_CONTROL_RoundCountxDP[3]), .B0_t (KECCAK_CONTROL_RoundCountxDP[2]), .Z0_t (KECCAK_CONTROL_n30) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) KECCAK_CONTROL_U9 ( .A0_t (Reset), .B0_t (KECCAK_CONTROL_n11), .Z0_t (KECCAK_CONTROL_RoundCountxDP[0]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b0)) KECCAK_CONTROL_U8 ( .A0_t (KECCAK_CONTROL_RoundCountxDP[0]), .B0_t (KECCAK_CONTROL_n13), .Z0_t (KECCAK_CONTROL_n11) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_U7 ( .A0_t (KECCAK_CONTROL_n10), .B0_t (KECCAK_CONTROL_CtrlStatexDP[2]), .Z0_t (KECCAK_CONTROL_n13) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b0)) KECCAK_CONTROL_U5 ( .A0_t (KECCAK_CONTROL_CtrlStatexDP[0]), .B0_t (KECCAK_CONTROL_CtrlStatexDP_reg_1__Q), .Z0_t (KECCAK_CONTROL_n10) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_U2 ( .A0_t (KECCAK_CONTROL_CtrlStatexDP[2]), .B0_t (KECCAK_CONTROL_n8), .Z0_t (Ready) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_U1 ( .A0_t (KECCAK_CONTROL_CtrlStatexDP_reg_1__Q), .B0_t (KECCAK_CONTROL_CtrlStatexDP[0]), .Z0_t (KECCAK_CONTROL_n8) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_RC_GEN_U35 ( .A0_t (KECCAK_CONTROL_RC_GEN_n3), .B0_t (KECCAK_CONTROL_RC_GEN_n28), .Z0_t (KECCAK_CONTROL_RC_GEN_n24) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_RC_GEN_U34 ( .A0_t (KECCAK_CONTROL_RC_GEN_n27), .B0_t (KECCAK_CONTROL_RC_GEN_n26), .Z0_t (KECCAK_CONTROL_RC_GEN_n28) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_RC_GEN_U33 ( .A0_t (KECCAK_CONTROL_RoundCountxDP[4]), .B0_t (KECCAK_CONTROL_RC_GEN_n25), .Z0_t (IotaRC_3) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_RC_GEN_U31 ( .A0_t (KECCAK_CONTROL_RC_GEN_n22), .B0_t (KECCAK_CONTROL_RC_GEN_n19), .Z0_t (KECCAK_CONTROL_RC_GEN_n25) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_RC_GEN_U30 ( .A0_t (KECCAK_CONTROL_RoundCountxDP[0]), .B0_t (KECCAK_CONTROL_RC_GEN_n18), .Z0_t (KECCAK_CONTROL_RC_GEN_n19) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_RC_GEN_U29 ( .A0_t (KECCAK_CONTROL_RoundCountxDP[3]), .B0_t (KECCAK_CONTROL_RC_GEN_n17), .Z0_t (KECCAK_CONTROL_RC_GEN_n18) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_RC_GEN_U27 ( .A0_t (KECCAK_CONTROL_RC_GEN_n27), .B0_t (KECCAK_CONTROL_RC_GEN_n15), .Z0_t (KECCAK_CONTROL_RC_GEN_n17) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_RC_GEN_U24 ( .A0_t (KECCAK_CONTROL_RC_GEN_n14), .B0_t (KECCAK_CONTROL_RC_GEN_n13), .Z0_t (KECCAK_CONTROL_RC_GEN_n22) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_RC_GEN_U23 ( .A0_t (KECCAK_CONTROL_RoundCountxDP[3]), .B0_t (KECCAK_CONTROL_RC_GEN_n27), .Z0_t (KECCAK_CONTROL_RC_GEN_n13) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_RC_GEN_U22 ( .A0_t (KECCAK_CONTROL_RoundCountxDP[2]), .B0_t (KECCAK_CONTROL_RoundCountxDP[1]), .Z0_t (KECCAK_CONTROL_RC_GEN_n27) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_RC_GEN_U21 ( .A0_t (KECCAK_CONTROL_RoundCountxDP[2]), .B0_t (KECCAK_CONTROL_RC_GEN_n12), .Z0_t (KECCAK_CONTROL_RC_GEN_n14) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_RC_GEN_U20 ( .A0_t (KECCAK_CONTROL_RC_GEN_n11), .B0_t (KECCAK_CONTROL_RoundCountxDP[0]), .Z0_t (KECCAK_CONTROL_RC_GEN_n12) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_RC_GEN_U18 ( .A0_t (KECCAK_CONTROL_RoundCountxDP[0]), .B0_t (KECCAK_CONTROL_RC_GEN_n9), .Z0_t (KECCAK_CONTROL_RC_GEN_n30) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_RC_GEN_U17 ( .A0_t (KECCAK_CONTROL_RC_GEN_n9), .B0_t (KECCAK_CONTROL_RC_GEN_n8), .Z0_t (KECCAK_CONTROL_RC_GEN_n20) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_RC_GEN_U16 ( .A0_t (KECCAK_CONTROL_RC_GEN_n3), .B0_t (KECCAK_CONTROL_RoundCountxDP[4]), .Z0_t (KECCAK_CONTROL_RC_GEN_n8) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_RC_GEN_U15 ( .A0_t (KECCAK_CONTROL_RC_GEN_n15), .B0_t (KECCAK_CONTROL_RoundCountxDP[3]), .Z0_t (KECCAK_CONTROL_RC_GEN_n9) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_RC_GEN_U14 ( .A0_t (KECCAK_CONTROL_RoundCountxDP[4]), .B0_t (KECCAK_CONTROL_RC_GEN_n6), .Z0_t (IotaRC[0]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_RC_GEN_U13 ( .A0_t (KECCAK_CONTROL_RoundCountxDP[2]), .B0_t (KECCAK_CONTROL_RC_GEN_n5), .Z0_t (KECCAK_CONTROL_RC_GEN_n6) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_RC_GEN_U12 ( .A0_t (KECCAK_CONTROL_RC_GEN_n4), .B0_t (KECCAK_CONTROL_RoundCountxDP[0]), .Z0_t (KECCAK_CONTROL_RC_GEN_n5) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_RC_GEN_U11 ( .A0_t (KECCAK_CONTROL_RC_GEN_n11), .B0_t (KECCAK_CONTROL_RC_GEN_n3), .Z0_t (KECCAK_CONTROL_RC_GEN_n4) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_RC_GEN_U9 ( .A0_t (KECCAK_CONTROL_RoundCountxDP[4]), .B0_t (KECCAK_CONTROL_RC_GEN_n2), .Z0_t (KECCAK_CONTROL_RC_GEN_n21) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_RC_GEN_U8 ( .A0_t (KECCAK_CONTROL_RC_GEN_n26), .B0_t (KECCAK_CONTROL_RC_GEN_n3), .Z0_t (KECCAK_CONTROL_RC_GEN_n2) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_RC_GEN_U7 ( .A0_t (KECCAK_CONTROL_RoundCountxDP[3]), .B0_t (KECCAK_CONTROL_RoundCountxDP[1]), .Z0_t (KECCAK_CONTROL_RC_GEN_n3) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_RC_GEN_U6 ( .A0_t (KECCAK_CONTROL_RoundCountxDP[2]), .B0_t (KECCAK_CONTROL_RC_GEN_n11), .Z0_t (KECCAK_CONTROL_RC_GEN_n26) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_RC_GEN_U5 ( .A0_t (KECCAK_CONTROL_RoundCountxDP[1]), .B0_t (KECCAK_CONTROL_RoundCountxDP[3]), .Z0_t (KECCAK_CONTROL_RC_GEN_n11) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) KECCAK_CONTROL_RC_GEN_U2 ( .A0_t (KECCAK_CONTROL_RC_GEN_n15), .B0_t (KECCAK_CONTROL_RoundCountxDP[3]), .Z0_t (KECCAK_CONTROL_RC_GEN_n23) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_RC_GEN_U1 ( .A0_t (KECCAK_CONTROL_RoundCountxDP[2]), .B0_t (KECCAK_CONTROL_RoundCountxDP[1]), .Z0_t (KECCAK_CONTROL_RC_GEN_n15) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) KECCAK_CONTROL_RC_GEN_U25_XOR1_U1 ( .A0_t (KECCAK_CONTROL_RC_GEN_n21), .B0_t (KECCAK_CONTROL_RC_GEN_n20), .Z0_t (KECCAK_CONTROL_RC_GEN_U25_X) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_RC_GEN_U25_AND1_U1 ( .A0_t (KECCAK_CONTROL_RoundCountxDP[0]), .B0_t (KECCAK_CONTROL_RC_GEN_U25_X), .Z0_t (KECCAK_CONTROL_RC_GEN_U25_Y) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) KECCAK_CONTROL_RC_GEN_U25_XOR2_U1 ( .A0_t (KECCAK_CONTROL_RC_GEN_U25_Y), .B0_t (KECCAK_CONTROL_RC_GEN_n21), .Z0_t (IotaRC_7) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) KECCAK_CONTROL_RC_GEN_U28_XOR1_U1 ( .A0_t (KECCAK_CONTROL_RC_GEN_n24), .B0_t (KECCAK_CONTROL_RC_GEN_n23), .Z0_t (KECCAK_CONTROL_RC_GEN_U28_X) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_RC_GEN_U28_AND1_U1 ( .A0_t (KECCAK_CONTROL_RoundCountxDP[0]), .B0_t (KECCAK_CONTROL_RC_GEN_U28_X), .Z0_t (KECCAK_CONTROL_RC_GEN_U28_Y) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) KECCAK_CONTROL_RC_GEN_U28_XOR2_U1 ( .A0_t (KECCAK_CONTROL_RC_GEN_U28_Y), .B0_t (KECCAK_CONTROL_RC_GEN_n24), .Z0_t (KECCAK_CONTROL_RC_GEN_n31) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) KECCAK_CONTROL_RC_GEN_U32_XOR1_U1 ( .A0_t (KECCAK_CONTROL_RC_GEN_n31), .B0_t (KECCAK_CONTROL_RC_GEN_n30), .Z0_t (KECCAK_CONTROL_RC_GEN_U32_X) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) KECCAK_CONTROL_RC_GEN_U32_AND1_U1 ( .A0_t (KECCAK_CONTROL_RoundCountxDP[4]), .B0_t (KECCAK_CONTROL_RC_GEN_U32_X), .Z0_t (KECCAK_CONTROL_RC_GEN_U32_Y) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) KECCAK_CONTROL_RC_GEN_U32_XOR2_U1 ( .A0_t (KECCAK_CONTROL_RC_GEN_U32_Y), .B0_t (KECCAK_CONTROL_RC_GEN_n31), .Z0_t (IotaRC[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U810_XOR1_U1 ( .A0_t (StateOut[11]), .B0_t (StateFromChi[3]), .Z0_t (U810_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U810_AND1_U1 ( .A0_t (n9), .B0_t (U810_X), .Z0_t (U810_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U810_XOR2_U1 ( .A0_t (U810_Y), .B0_t (StateOut[11]), .Z0_t (OutData[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U812_XOR1_U1 ( .A0_t (StateOut[15]), .B0_t (StateFromChi[7]), .Z0_t (U812_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U812_AND1_U1 ( .A0_t (n9), .B0_t (U812_X), .Z0_t (U812_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U812_XOR2_U1 ( .A0_t (U812_Y), .B0_t (StateOut[15]), .Z0_t (OutData[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U814_XOR1_U1 ( .A0_t (StateOut[8]), .B0_t (StateFromChi[0]), .Z0_t (U814_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U814_AND1_U1 ( .A0_t (n9), .B0_t (U814_X), .Z0_t (U814_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U814_XOR2_U1 ( .A0_t (U814_Y), .B0_t (StateOut[8]), .Z0_t (OutData[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U816_XOR1_U1 ( .A0_t (StateOut[9]), .B0_t (StateFromChi[1]), .Z0_t (U816_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U816_AND1_U1 ( .A0_t (n9), .B0_t (U816_X), .Z0_t (U816_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U816_XOR2_U1 ( .A0_t (U816_Y), .B0_t (StateOut[9]), .Z0_t (OutData[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U817_XOR1_U1 ( .A0_t (StateOut[47]), .B0_t (StateFromChi[39]), .Z0_t (U817_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U817_AND1_U1 ( .A0_t (n9), .B0_t (U817_X), .Z0_t (U817_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U817_XOR2_U1 ( .A0_t (U817_Y), .B0_t (StateOut[47]), .Z0_t (StateOut[39]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U818_XOR1_U1 ( .A0_t (StateOut[71]), .B0_t (StateFromChi[63]), .Z0_t (U818_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U818_AND1_U1 ( .A0_t (n9), .B0_t (U818_X), .Z0_t (U818_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U818_XOR2_U1 ( .A0_t (U818_Y), .B0_t (StateOut[71]), .Z0_t (StateOut[63]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U820_XOR1_U1 ( .A0_t (StateOut[95]), .B0_t (StateFromChi[87]), .Z0_t (U820_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U820_AND1_U1 ( .A0_t (n9), .B0_t (U820_X), .Z0_t (U820_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U820_XOR2_U1 ( .A0_t (U820_Y), .B0_t (StateOut[95]), .Z0_t (StateOut[87]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U821_XOR1_U1 ( .A0_t (StateOut[127]), .B0_t (StateFromChi[119]), .Z0_t (U821_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U821_AND1_U1 ( .A0_t (n9), .B0_t (U821_X), .Z0_t (U821_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U821_XOR2_U1 ( .A0_t (U821_Y), .B0_t (StateOut[127]), .Z0_t (StateOut[119]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U822_XOR1_U1 ( .A0_t (StateOut[151]), .B0_t (StateFromChi[143]), .Z0_t (U822_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U822_AND1_U1 ( .A0_t (n9), .B0_t (U822_X), .Z0_t (U822_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U822_XOR2_U1 ( .A0_t (U822_Y), .B0_t (StateOut[151]), .Z0_t (StateOut[143]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U823_XOR1_U1 ( .A0_t (StateOut[159]), .B0_t (StateFromChi[151]), .Z0_t (U823_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U823_AND1_U1 ( .A0_t (n9), .B0_t (U823_X), .Z0_t (U823_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U823_XOR2_U1 ( .A0_t (U823_Y), .B0_t (StateOut[159]), .Z0_t (StateOut[151]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U824_XOR1_U1 ( .A0_t (StateOut[175]), .B0_t (StateFromChi[167]), .Z0_t (U824_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U824_AND1_U1 ( .A0_t (n9), .B0_t (U824_X), .Z0_t (U824_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U824_XOR2_U1 ( .A0_t (U824_Y), .B0_t (StateOut[175]), .Z0_t (StateOut[167]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U825_XOR1_U1 ( .A0_t (StateOut[46]), .B0_t (StateFromChi[38]), .Z0_t (U825_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U825_AND1_U1 ( .A0_t (n9), .B0_t (U825_X), .Z0_t (U825_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U825_XOR2_U1 ( .A0_t (U825_Y), .B0_t (StateOut[46]), .Z0_t (StateOut[38]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U827_XOR1_U1 ( .A0_t (StateOut[70]), .B0_t (StateFromChi[62]), .Z0_t (U827_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U827_AND1_U1 ( .A0_t (n9), .B0_t (U827_X), .Z0_t (U827_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U827_XOR2_U1 ( .A0_t (U827_Y), .B0_t (StateOut[70]), .Z0_t (StateOut[62]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U828_XOR1_U1 ( .A0_t (StateOut[126]), .B0_t (StateFromChi[118]), .Z0_t (U828_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U828_AND1_U1 ( .A0_t (n9), .B0_t (U828_X), .Z0_t (U828_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U828_XOR2_U1 ( .A0_t (U828_Y), .B0_t (StateOut[126]), .Z0_t (StateOut[118]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U830_XOR1_U1 ( .A0_t (StateOut[150]), .B0_t (StateFromChi[142]), .Z0_t (U830_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U830_AND1_U1 ( .A0_t (n9), .B0_t (U830_X), .Z0_t (U830_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U830_XOR2_U1 ( .A0_t (U830_Y), .B0_t (StateOut[150]), .Z0_t (StateOut[142]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U831_XOR1_U1 ( .A0_t (StateOut[158]), .B0_t (StateFromChi[150]), .Z0_t (U831_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U831_AND1_U1 ( .A0_t (n9), .B0_t (U831_X), .Z0_t (U831_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U831_XOR2_U1 ( .A0_t (U831_Y), .B0_t (StateOut[158]), .Z0_t (StateOut[150]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U832_XOR1_U1 ( .A0_t (StateOut[174]), .B0_t (StateFromChi[166]), .Z0_t (U832_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U832_AND1_U1 ( .A0_t (n9), .B0_t (U832_X), .Z0_t (U832_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U832_XOR2_U1 ( .A0_t (U832_Y), .B0_t (StateOut[174]), .Z0_t (StateOut[166]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U833_XOR1_U1 ( .A0_t (StateOut[182]), .B0_t (StateFromChi[174]), .Z0_t (U833_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U833_AND1_U1 ( .A0_t (n9), .B0_t (U833_X), .Z0_t (U833_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U833_XOR2_U1 ( .A0_t (U833_Y), .B0_t (StateOut[182]), .Z0_t (StateOut[174]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U834_XOR1_U1 ( .A0_t (StateOut[45]), .B0_t (StateFromChi[37]), .Z0_t (U834_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U834_AND1_U1 ( .A0_t (n9), .B0_t (U834_X), .Z0_t (U834_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U834_XOR2_U1 ( .A0_t (U834_Y), .B0_t (StateOut[45]), .Z0_t (StateOut[37]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U835_XOR1_U1 ( .A0_t (StateOut[61]), .B0_t (StateFromChi[53]), .Z0_t (U835_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U835_AND1_U1 ( .A0_t (n9), .B0_t (U835_X), .Z0_t (U835_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U835_XOR2_U1 ( .A0_t (U835_Y), .B0_t (StateOut[61]), .Z0_t (StateOut[53]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U836_XOR1_U1 ( .A0_t (StateOut[69]), .B0_t (StateFromChi[61]), .Z0_t (U836_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U836_AND1_U1 ( .A0_t (n9), .B0_t (U836_X), .Z0_t (U836_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U836_XOR2_U1 ( .A0_t (U836_Y), .B0_t (StateOut[69]), .Z0_t (StateOut[61]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U837_XOR1_U1 ( .A0_t (StateOut[77]), .B0_t (StateFromChi[69]), .Z0_t (U837_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U837_AND1_U1 ( .A0_t (n9), .B0_t (U837_X), .Z0_t (U837_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U837_XOR2_U1 ( .A0_t (U837_Y), .B0_t (StateOut[77]), .Z0_t (StateOut[69]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U838_XOR1_U1 ( .A0_t (StateOut[125]), .B0_t (StateFromChi[117]), .Z0_t (U838_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U838_AND1_U1 ( .A0_t (n9), .B0_t (U838_X), .Z0_t (U838_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U838_XOR2_U1 ( .A0_t (U838_Y), .B0_t (StateOut[125]), .Z0_t (StateOut[117]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U839_XOR1_U1 ( .A0_t (StateOut[149]), .B0_t (StateFromChi[141]), .Z0_t (U839_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U839_AND1_U1 ( .A0_t (n9), .B0_t (U839_X), .Z0_t (U839_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U839_XOR2_U1 ( .A0_t (U839_Y), .B0_t (StateOut[149]), .Z0_t (StateOut[141]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U841_XOR1_U1 ( .A0_t (StateOut[157]), .B0_t (StateFromChi[149]), .Z0_t (U841_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U841_AND1_U1 ( .A0_t (n9), .B0_t (U841_X), .Z0_t (U841_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U841_XOR2_U1 ( .A0_t (U841_Y), .B0_t (StateOut[157]), .Z0_t (StateOut[149]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U842_XOR1_U1 ( .A0_t (StateOut[173]), .B0_t (StateFromChi[165]), .Z0_t (U842_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U842_AND1_U1 ( .A0_t (n9), .B0_t (U842_X), .Z0_t (U842_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U842_XOR2_U1 ( .A0_t (U842_Y), .B0_t (StateOut[173]), .Z0_t (StateOut[165]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U843_XOR1_U1 ( .A0_t (StateOut[181]), .B0_t (StateFromChi[173]), .Z0_t (U843_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U843_AND1_U1 ( .A0_t (n9), .B0_t (U843_X), .Z0_t (U843_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U843_XOR2_U1 ( .A0_t (U843_Y), .B0_t (StateOut[181]), .Z0_t (StateOut[173]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U844_XOR1_U1 ( .A0_t (StateOut[36]), .B0_t (StateFromChi[28]), .Z0_t (U844_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U844_AND1_U1 ( .A0_t (n9), .B0_t (U844_X), .Z0_t (U844_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U844_XOR2_U1 ( .A0_t (U844_Y), .B0_t (StateOut[36]), .Z0_t (StateOut[28]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U845_XOR1_U1 ( .A0_t (StateOut[44]), .B0_t (StateFromChi[36]), .Z0_t (U845_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U845_AND1_U1 ( .A0_t (n9), .B0_t (U845_X), .Z0_t (U845_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U845_XOR2_U1 ( .A0_t (U845_Y), .B0_t (StateOut[44]), .Z0_t (StateOut[36]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U846_XOR1_U1 ( .A0_t (StateOut[60]), .B0_t (StateFromChi[52]), .Z0_t (U846_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U846_AND1_U1 ( .A0_t (n9), .B0_t (U846_X), .Z0_t (U846_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U846_XOR2_U1 ( .A0_t (U846_Y), .B0_t (StateOut[60]), .Z0_t (StateOut[52]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U847_XOR1_U1 ( .A0_t (StateOut[68]), .B0_t (StateFromChi[60]), .Z0_t (U847_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U847_AND1_U1 ( .A0_t (n9), .B0_t (U847_X), .Z0_t (U847_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U847_XOR2_U1 ( .A0_t (U847_Y), .B0_t (StateOut[68]), .Z0_t (StateOut[60]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U848_XOR1_U1 ( .A0_t (StateOut[92]), .B0_t (StateFromChi[84]), .Z0_t (U848_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U848_AND1_U1 ( .A0_t (n9), .B0_t (U848_X), .Z0_t (U848_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U848_XOR2_U1 ( .A0_t (U848_Y), .B0_t (StateOut[92]), .Z0_t (StateOut[84]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U849_XOR1_U1 ( .A0_t (StateOut[100]), .B0_t (StateFromChi[92]), .Z0_t (U849_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U849_AND1_U1 ( .A0_t (n9), .B0_t (U849_X), .Z0_t (U849_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U849_XOR2_U1 ( .A0_t (U849_Y), .B0_t (StateOut[100]), .Z0_t (StateOut[92]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U850_XOR1_U1 ( .A0_t (StateOut[124]), .B0_t (StateFromChi[116]), .Z0_t (U850_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U850_AND1_U1 ( .A0_t (n9), .B0_t (U850_X), .Z0_t (U850_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U850_XOR2_U1 ( .A0_t (U850_Y), .B0_t (StateOut[124]), .Z0_t (StateOut[116]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U851_XOR1_U1 ( .A0_t (StateOut[172]), .B0_t (StateFromChi[164]), .Z0_t (U851_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U851_AND1_U1 ( .A0_t (n9), .B0_t (U851_X), .Z0_t (U851_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U851_XOR2_U1 ( .A0_t (U851_Y), .B0_t (StateOut[172]), .Z0_t (StateOut[164]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U852_XOR1_U1 ( .A0_t (StateOut[180]), .B0_t (StateFromChi[172]), .Z0_t (U852_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U852_AND1_U1 ( .A0_t (n9), .B0_t (U852_X), .Z0_t (U852_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U852_XOR2_U1 ( .A0_t (U852_Y), .B0_t (StateOut[180]), .Z0_t (StateOut[172]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U853_XOR1_U1 ( .A0_t (StateOut[35]), .B0_t (StateFromChi[27]), .Z0_t (U853_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U853_AND1_U1 ( .A0_t (n9), .B0_t (U853_X), .Z0_t (U853_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U853_XOR2_U1 ( .A0_t (U853_Y), .B0_t (StateOut[35]), .Z0_t (StateOut[27]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U854_XOR1_U1 ( .A0_t (StateOut[59]), .B0_t (StateFromChi[51]), .Z0_t (U854_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U854_AND1_U1 ( .A0_t (n9), .B0_t (U854_X), .Z0_t (U854_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U854_XOR2_U1 ( .A0_t (U854_Y), .B0_t (StateOut[59]), .Z0_t (StateOut[51]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U855_XOR1_U1 ( .A0_t (StateOut[91]), .B0_t (StateFromChi[83]), .Z0_t (U855_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U855_AND1_U1 ( .A0_t (n9), .B0_t (U855_X), .Z0_t (U855_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U855_XOR2_U1 ( .A0_t (U855_Y), .B0_t (StateOut[91]), .Z0_t (StateOut[83]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U856_XOR1_U1 ( .A0_t (StateOut[155]), .B0_t (StateFromChi[147]), .Z0_t (U856_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U856_AND1_U1 ( .A0_t (n9), .B0_t (U856_X), .Z0_t (U856_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U856_XOR2_U1 ( .A0_t (U856_Y), .B0_t (StateOut[155]), .Z0_t (StateOut[147]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U857_XOR1_U1 ( .A0_t (StateOut[171]), .B0_t (StateFromChi[163]), .Z0_t (U857_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U857_AND1_U1 ( .A0_t (n9), .B0_t (U857_X), .Z0_t (U857_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U857_XOR2_U1 ( .A0_t (U857_Y), .B0_t (StateOut[171]), .Z0_t (StateOut[163]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U858_XOR1_U1 ( .A0_t (StateOut[179]), .B0_t (StateFromChi[171]), .Z0_t (U858_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U858_AND1_U1 ( .A0_t (n9), .B0_t (U858_X), .Z0_t (U858_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U858_XOR2_U1 ( .A0_t (U858_Y), .B0_t (StateOut[179]), .Z0_t (StateOut[171]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U859_XOR1_U1 ( .A0_t (StateOut[187]), .B0_t (StateFromChi[179]), .Z0_t (U859_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U859_AND1_U1 ( .A0_t (n9), .B0_t (U859_X), .Z0_t (U859_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U859_XOR2_U1 ( .A0_t (U859_Y), .B0_t (StateOut[187]), .Z0_t (StateOut[179]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U860_XOR1_U1 ( .A0_t (StateOut[34]), .B0_t (StateFromChi[26]), .Z0_t (U860_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U860_AND1_U1 ( .A0_t (n9), .B0_t (U860_X), .Z0_t (U860_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U860_XOR2_U1 ( .A0_t (U860_Y), .B0_t (StateOut[34]), .Z0_t (StateOut[26]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U861_XOR1_U1 ( .A0_t (StateOut[42]), .B0_t (StateFromChi[34]), .Z0_t (U861_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U861_AND1_U1 ( .A0_t (n9), .B0_t (U861_X), .Z0_t (U861_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U861_XOR2_U1 ( .A0_t (U861_Y), .B0_t (StateOut[42]), .Z0_t (StateOut[34]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U862_XOR1_U1 ( .A0_t (StateOut[58]), .B0_t (StateFromChi[50]), .Z0_t (U862_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U862_AND1_U1 ( .A0_t (n9), .B0_t (U862_X), .Z0_t (U862_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U862_XOR2_U1 ( .A0_t (U862_Y), .B0_t (StateOut[58]), .Z0_t (StateOut[50]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U863_XOR1_U1 ( .A0_t (StateOut[66]), .B0_t (StateFromChi[58]), .Z0_t (U863_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U863_AND1_U1 ( .A0_t (n9), .B0_t (U863_X), .Z0_t (U863_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U863_XOR2_U1 ( .A0_t (U863_Y), .B0_t (StateOut[66]), .Z0_t (StateOut[58]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U864_XOR1_U1 ( .A0_t (StateOut[90]), .B0_t (StateFromChi[82]), .Z0_t (U864_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U864_AND1_U1 ( .A0_t (n9), .B0_t (U864_X), .Z0_t (U864_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U864_XOR2_U1 ( .A0_t (U864_Y), .B0_t (StateOut[90]), .Z0_t (StateOut[82]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U865_XOR1_U1 ( .A0_t (StateOut[162]), .B0_t (StateFromChi[154]), .Z0_t (U865_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U865_AND1_U1 ( .A0_t (n9), .B0_t (U865_X), .Z0_t (U865_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U865_XOR2_U1 ( .A0_t (U865_Y), .B0_t (StateOut[162]), .Z0_t (StateOut[154]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U866_XOR1_U1 ( .A0_t (StateOut[33]), .B0_t (StateFromChi[25]), .Z0_t (U866_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U866_AND1_U1 ( .A0_t (n9), .B0_t (U866_X), .Z0_t (U866_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U866_XOR2_U1 ( .A0_t (U866_Y), .B0_t (StateOut[33]), .Z0_t (StateOut[25]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U867_XOR1_U1 ( .A0_t (StateOut[57]), .B0_t (StateFromChi[49]), .Z0_t (U867_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U867_AND1_U1 ( .A0_t (n9), .B0_t (U867_X), .Z0_t (U867_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U867_XOR2_U1 ( .A0_t (U867_Y), .B0_t (StateOut[57]), .Z0_t (StateOut[49]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U868_XOR1_U1 ( .A0_t (StateOut[89]), .B0_t (StateFromChi[81]), .Z0_t (U868_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U868_AND1_U1 ( .A0_t (n9), .B0_t (U868_X), .Z0_t (U868_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U868_XOR2_U1 ( .A0_t (U868_Y), .B0_t (StateOut[89]), .Z0_t (StateOut[81]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U869_XOR1_U1 ( .A0_t (StateOut[145]), .B0_t (StateFromChi[137]), .Z0_t (U869_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U869_AND1_U1 ( .A0_t (n9), .B0_t (U869_X), .Z0_t (U869_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U869_XOR2_U1 ( .A0_t (U869_Y), .B0_t (StateOut[145]), .Z0_t (StateOut[137]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U870_XOR1_U1 ( .A0_t (StateOut[177]), .B0_t (StateFromChi[169]), .Z0_t (U870_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U870_AND1_U1 ( .A0_t (n9), .B0_t (U870_X), .Z0_t (U870_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U870_XOR2_U1 ( .A0_t (U870_Y), .B0_t (StateOut[177]), .Z0_t (StateOut[169]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U871_XOR1_U1 ( .A0_t (StateOut[32]), .B0_t (StateFromChi[24]), .Z0_t (U871_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U871_AND1_U1 ( .A0_t (n9), .B0_t (U871_X), .Z0_t (U871_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U871_XOR2_U1 ( .A0_t (U871_Y), .B0_t (StateOut[32]), .Z0_t (StateOut[24]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U872_XOR1_U1 ( .A0_t (StateOut[120]), .B0_t (StateFromChi[112]), .Z0_t (U872_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U872_AND1_U1 ( .A0_t (n9), .B0_t (U872_X), .Z0_t (U872_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U872_XOR2_U1 ( .A0_t (U872_Y), .B0_t (StateOut[120]), .Z0_t (StateOut[112]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U873_XOR1_U1 ( .A0_t (StateOut[144]), .B0_t (StateFromChi[136]), .Z0_t (U873_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U873_AND1_U1 ( .A0_t (n9), .B0_t (U873_X), .Z0_t (U873_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U873_XOR2_U1 ( .A0_t (U873_Y), .B0_t (StateOut[144]), .Z0_t (StateOut[136]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U874_XOR1_U1 ( .A0_t (StateOut[152]), .B0_t (StateFromChi[144]), .Z0_t (U874_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U874_AND1_U1 ( .A0_t (n9), .B0_t (U874_X), .Z0_t (U874_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U874_XOR2_U1 ( .A0_t (U874_Y), .B0_t (StateOut[152]), .Z0_t (StateOut[144]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U875_XOR1_U1 ( .A0_t (StateOut[31]), .B0_t (StateFromChi[23]), .Z0_t (U875_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U875_AND1_U1 ( .A0_t (n9), .B0_t (U875_X), .Z0_t (U875_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U875_XOR2_U1 ( .A0_t (U875_Y), .B0_t (StateOut[31]), .Z0_t (StateOut[23]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U876_XOR1_U1 ( .A0_t (StateOut[39]), .B0_t (StateFromChi[31]), .Z0_t (U876_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U876_AND1_U1 ( .A0_t (n9), .B0_t (U876_X), .Z0_t (U876_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U876_XOR2_U1 ( .A0_t (U876_Y), .B0_t (StateOut[39]), .Z0_t (StateOut[31]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U877_XOR1_U1 ( .A0_t (StateOut[63]), .B0_t (StateFromChi[55]), .Z0_t (U877_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U877_AND1_U1 ( .A0_t (n9), .B0_t (U877_X), .Z0_t (U877_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U877_XOR2_U1 ( .A0_t (U877_Y), .B0_t (StateOut[63]), .Z0_t (StateOut[55]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U878_XOR1_U1 ( .A0_t (StateOut[119]), .B0_t (StateFromChi[111]), .Z0_t (U878_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U878_AND1_U1 ( .A0_t (n9), .B0_t (U878_X), .Z0_t (U878_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U878_XOR2_U1 ( .A0_t (U878_Y), .B0_t (StateOut[119]), .Z0_t (StateOut[111]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U879_XOR1_U1 ( .A0_t (StateOut[183]), .B0_t (StateFromChi[175]), .Z0_t (U879_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U879_AND1_U1 ( .A0_t (n9), .B0_t (U879_X), .Z0_t (U879_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U879_XOR2_U1 ( .A0_t (U879_Y), .B0_t (StateOut[183]), .Z0_t (StateOut[175]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U880_XOR1_U1 ( .A0_t (InData[7]), .B0_t (StateFromChi[199]), .Z0_t (U880_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U880_AND1_U1 ( .A0_t (n9), .B0_t (U880_X), .Z0_t (U880_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U880_XOR2_U1 ( .A0_t (U880_Y), .B0_t (InData[7]), .Z0_t (StateOut[199]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U881_XOR1_U1 ( .A0_t (StateOut[30]), .B0_t (StateFromChi[22]), .Z0_t (U881_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U881_AND1_U1 ( .A0_t (n9), .B0_t (U881_X), .Z0_t (U881_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U881_XOR2_U1 ( .A0_t (U881_Y), .B0_t (StateOut[30]), .Z0_t (StateOut[22]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U882_XOR1_U1 ( .A0_t (StateOut[38]), .B0_t (StateFromChi[30]), .Z0_t (U882_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U882_AND1_U1 ( .A0_t (n9), .B0_t (U882_X), .Z0_t (U882_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U882_XOR2_U1 ( .A0_t (U882_Y), .B0_t (StateOut[38]), .Z0_t (StateOut[30]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U883_XOR1_U1 ( .A0_t (StateOut[62]), .B0_t (StateFromChi[54]), .Z0_t (U883_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U883_AND1_U1 ( .A0_t (n9), .B0_t (U883_X), .Z0_t (U883_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U883_XOR2_U1 ( .A0_t (U883_Y), .B0_t (StateOut[62]), .Z0_t (StateOut[54]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U884_XOR1_U1 ( .A0_t (StateOut[94]), .B0_t (StateFromChi[86]), .Z0_t (U884_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U884_AND1_U1 ( .A0_t (n9), .B0_t (U884_X), .Z0_t (U884_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U884_XOR2_U1 ( .A0_t (U884_Y), .B0_t (StateOut[94]), .Z0_t (StateOut[86]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U885_XOR1_U1 ( .A0_t (StateOut[118]), .B0_t (StateFromChi[110]), .Z0_t (U885_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U885_AND1_U1 ( .A0_t (n9), .B0_t (U885_X), .Z0_t (U885_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U885_XOR2_U1 ( .A0_t (U885_Y), .B0_t (StateOut[118]), .Z0_t (StateOut[110]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U886_XOR1_U1 ( .A0_t (InData[6]), .B0_t (StateFromChi[198]), .Z0_t (U886_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U886_AND1_U1 ( .A0_t (n9), .B0_t (U886_X), .Z0_t (U886_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U886_XOR2_U1 ( .A0_t (U886_Y), .B0_t (InData[6]), .Z0_t (StateOut[198]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U887_XOR1_U1 ( .A0_t (StateOut[29]), .B0_t (StateFromChi[21]), .Z0_t (U887_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U887_AND1_U1 ( .A0_t (n9), .B0_t (U887_X), .Z0_t (U887_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U887_XOR2_U1 ( .A0_t (U887_Y), .B0_t (StateOut[29]), .Z0_t (StateOut[21]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U888_XOR1_U1 ( .A0_t (StateOut[37]), .B0_t (StateFromChi[29]), .Z0_t (U888_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U888_AND1_U1 ( .A0_t (n9), .B0_t (U888_X), .Z0_t (U888_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U888_XOR2_U1 ( .A0_t (U888_Y), .B0_t (StateOut[37]), .Z0_t (StateOut[29]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U889_XOR1_U1 ( .A0_t (StateOut[93]), .B0_t (StateFromChi[85]), .Z0_t (U889_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U889_AND1_U1 ( .A0_t (n9), .B0_t (U889_X), .Z0_t (U889_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U889_XOR2_U1 ( .A0_t (U889_Y), .B0_t (StateOut[93]), .Z0_t (StateOut[85]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U890_XOR1_U1 ( .A0_t (StateOut[141]), .B0_t (StateFromChi[133]), .Z0_t (U890_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U890_AND1_U1 ( .A0_t (n9), .B0_t (U890_X), .Z0_t (U890_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U890_XOR2_U1 ( .A0_t (U890_Y), .B0_t (StateOut[141]), .Z0_t (StateOut[133]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U891_XOR1_U1 ( .A0_t (StateOut[52]), .B0_t (StateFromChi[44]), .Z0_t (U891_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U891_AND1_U1 ( .A0_t (n9), .B0_t (U891_X), .Z0_t (U891_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U891_XOR2_U1 ( .A0_t (U891_Y), .B0_t (StateOut[52]), .Z0_t (StateOut[44]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U892_XOR1_U1 ( .A0_t (StateOut[76]), .B0_t (StateFromChi[68]), .Z0_t (U892_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U892_AND1_U1 ( .A0_t (n9), .B0_t (U892_X), .Z0_t (U892_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U892_XOR2_U1 ( .A0_t (U892_Y), .B0_t (StateOut[76]), .Z0_t (StateOut[68]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U893_XOR1_U1 ( .A0_t (StateOut[140]), .B0_t (StateFromChi[132]), .Z0_t (U893_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U893_AND1_U1 ( .A0_t (n9), .B0_t (U893_X), .Z0_t (U893_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U893_XOR2_U1 ( .A0_t (U893_Y), .B0_t (StateOut[140]), .Z0_t (StateOut[132]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U894_XOR1_U1 ( .A0_t (StateOut[148]), .B0_t (StateFromChi[140]), .Z0_t (U894_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U894_AND1_U1 ( .A0_t (n9), .B0_t (U894_X), .Z0_t (U894_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U894_XOR2_U1 ( .A0_t (U894_Y), .B0_t (StateOut[148]), .Z0_t (StateOut[140]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U895_XOR1_U1 ( .A0_t (StateOut[156]), .B0_t (StateFromChi[148]), .Z0_t (U895_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U895_AND1_U1 ( .A0_t (n9), .B0_t (U895_X), .Z0_t (U895_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U895_XOR2_U1 ( .A0_t (U895_Y), .B0_t (StateOut[156]), .Z0_t (StateOut[148]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U896_XOR1_U1 ( .A0_t (StateOut[43]), .B0_t (StateFromChi[35]), .Z0_t (U896_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U896_AND1_U1 ( .A0_t (n9), .B0_t (U896_X), .Z0_t (U896_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U896_XOR2_U1 ( .A0_t (U896_Y), .B0_t (StateOut[43]), .Z0_t (StateOut[35]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U897_XOR1_U1 ( .A0_t (StateOut[51]), .B0_t (StateFromChi[43]), .Z0_t (U897_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U897_AND1_U1 ( .A0_t (n9), .B0_t (U897_X), .Z0_t (U897_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U897_XOR2_U1 ( .A0_t (U897_Y), .B0_t (StateOut[51]), .Z0_t (StateOut[43]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U898_XOR1_U1 ( .A0_t (StateOut[67]), .B0_t (StateFromChi[59]), .Z0_t (U898_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U898_AND1_U1 ( .A0_t (n9), .B0_t (U898_X), .Z0_t (U898_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U898_XOR2_U1 ( .A0_t (U898_Y), .B0_t (StateOut[67]), .Z0_t (StateOut[59]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U899_XOR1_U1 ( .A0_t (StateOut[75]), .B0_t (StateFromChi[67]), .Z0_t (U899_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U899_AND1_U1 ( .A0_t (n9), .B0_t (U899_X), .Z0_t (U899_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U899_XOR2_U1 ( .A0_t (U899_Y), .B0_t (StateOut[75]), .Z0_t (StateOut[67]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U900_XOR1_U1 ( .A0_t (StateOut[99]), .B0_t (StateFromChi[91]), .Z0_t (U900_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U900_AND1_U1 ( .A0_t (n9), .B0_t (U900_X), .Z0_t (U900_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U900_XOR2_U1 ( .A0_t (U900_Y), .B0_t (StateOut[99]), .Z0_t (StateOut[91]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U901_XOR1_U1 ( .A0_t (StateOut[123]), .B0_t (StateFromChi[115]), .Z0_t (U901_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U901_AND1_U1 ( .A0_t (n9), .B0_t (U901_X), .Z0_t (U901_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U901_XOR2_U1 ( .A0_t (U901_Y), .B0_t (StateOut[123]), .Z0_t (StateOut[115]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U902_XOR1_U1 ( .A0_t (StateOut[139]), .B0_t (StateFromChi[131]), .Z0_t (U902_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U902_AND1_U1 ( .A0_t (n9), .B0_t (U902_X), .Z0_t (U902_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U902_XOR2_U1 ( .A0_t (U902_Y), .B0_t (StateOut[139]), .Z0_t (StateOut[131]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U903_XOR1_U1 ( .A0_t (StateOut[147]), .B0_t (StateFromChi[139]), .Z0_t (U903_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U903_AND1_U1 ( .A0_t (n9), .B0_t (U903_X), .Z0_t (U903_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U903_XOR2_U1 ( .A0_t (U903_Y), .B0_t (StateOut[147]), .Z0_t (StateOut[139]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U904_XOR1_U1 ( .A0_t (StateOut[50]), .B0_t (StateFromChi[42]), .Z0_t (U904_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U904_AND1_U1 ( .A0_t (n9), .B0_t (U904_X), .Z0_t (U904_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U904_XOR2_U1 ( .A0_t (U904_Y), .B0_t (StateOut[50]), .Z0_t (StateOut[42]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U905_XOR1_U1 ( .A0_t (StateOut[98]), .B0_t (StateFromChi[90]), .Z0_t (U905_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U905_AND1_U1 ( .A0_t (n9), .B0_t (U905_X), .Z0_t (U905_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U905_XOR2_U1 ( .A0_t (U905_Y), .B0_t (StateOut[98]), .Z0_t (StateOut[90]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U906_XOR1_U1 ( .A0_t (StateOut[114]), .B0_t (StateFromChi[106]), .Z0_t (U906_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U906_AND1_U1 ( .A0_t (n9), .B0_t (U906_X), .Z0_t (U906_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U906_XOR2_U1 ( .A0_t (U906_Y), .B0_t (StateOut[114]), .Z0_t (StateOut[106]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U907_XOR1_U1 ( .A0_t (StateOut[122]), .B0_t (StateFromChi[114]), .Z0_t (U907_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U907_AND1_U1 ( .A0_t (n9), .B0_t (U907_X), .Z0_t (U907_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U907_XOR2_U1 ( .A0_t (U907_Y), .B0_t (StateOut[122]), .Z0_t (StateOut[114]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U908_XOR1_U1 ( .A0_t (StateOut[138]), .B0_t (StateFromChi[130]), .Z0_t (U908_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U908_AND1_U1 ( .A0_t (n9), .B0_t (U908_X), .Z0_t (U908_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U908_XOR2_U1 ( .A0_t (U908_Y), .B0_t (StateOut[138]), .Z0_t (StateOut[130]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U909_XOR1_U1 ( .A0_t (StateOut[146]), .B0_t (StateFromChi[138]), .Z0_t (U909_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U909_AND1_U1 ( .A0_t (n9), .B0_t (U909_X), .Z0_t (U909_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U909_XOR2_U1 ( .A0_t (U909_Y), .B0_t (StateOut[146]), .Z0_t (StateOut[138]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U910_XOR1_U1 ( .A0_t (StateOut[154]), .B0_t (StateFromChi[146]), .Z0_t (U910_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U910_AND1_U1 ( .A0_t (n9), .B0_t (U910_X), .Z0_t (U910_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U910_XOR2_U1 ( .A0_t (U910_Y), .B0_t (StateOut[154]), .Z0_t (StateOut[146]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U911_XOR1_U1 ( .A0_t (StateOut[170]), .B0_t (StateFromChi[162]), .Z0_t (U911_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U911_AND1_U1 ( .A0_t (n9), .B0_t (U911_X), .Z0_t (U911_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U911_XOR2_U1 ( .A0_t (U911_Y), .B0_t (StateOut[170]), .Z0_t (StateOut[162]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U912_XOR1_U1 ( .A0_t (StateOut[178]), .B0_t (StateFromChi[170]), .Z0_t (U912_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U912_AND1_U1 ( .A0_t (n9), .B0_t (U912_X), .Z0_t (U912_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U912_XOR2_U1 ( .A0_t (U912_Y), .B0_t (StateOut[178]), .Z0_t (StateOut[170]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U913_XOR1_U1 ( .A0_t (StateOut[186]), .B0_t (StateFromChi[178]), .Z0_t (U913_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U913_AND1_U1 ( .A0_t (n9), .B0_t (U913_X), .Z0_t (U913_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U913_XOR2_U1 ( .A0_t (U913_Y), .B0_t (StateOut[186]), .Z0_t (StateOut[178]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U914_XOR1_U1 ( .A0_t (InData[2]), .B0_t (StateFromChi[194]), .Z0_t (U914_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U914_AND1_U1 ( .A0_t (n9), .B0_t (U914_X), .Z0_t (U914_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U914_XOR2_U1 ( .A0_t (U914_Y), .B0_t (InData[2]), .Z0_t (StateOut[194]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U915_XOR1_U1 ( .A0_t (StateOut[25]), .B0_t (StateFromChi[17]), .Z0_t (U915_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U915_AND1_U1 ( .A0_t (n9), .B0_t (U915_X), .Z0_t (U915_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U915_XOR2_U1 ( .A0_t (U915_Y), .B0_t (StateOut[25]), .Z0_t (StateOut[17]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U916_XOR1_U1 ( .A0_t (StateOut[41]), .B0_t (StateFromChi[33]), .Z0_t (U916_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U916_AND1_U1 ( .A0_t (n9), .B0_t (U916_X), .Z0_t (U916_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U916_XOR2_U1 ( .A0_t (U916_Y), .B0_t (StateOut[41]), .Z0_t (StateOut[33]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U917_XOR1_U1 ( .A0_t (StateOut[49]), .B0_t (StateFromChi[41]), .Z0_t (U917_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U917_AND1_U1 ( .A0_t (n9), .B0_t (U917_X), .Z0_t (U917_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U917_XOR2_U1 ( .A0_t (U917_Y), .B0_t (StateOut[49]), .Z0_t (StateOut[41]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U918_XOR1_U1 ( .A0_t (StateOut[65]), .B0_t (StateFromChi[57]), .Z0_t (U918_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U918_AND1_U1 ( .A0_t (n9), .B0_t (U918_X), .Z0_t (U918_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U918_XOR2_U1 ( .A0_t (U918_Y), .B0_t (StateOut[65]), .Z0_t (StateOut[57]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U919_XOR1_U1 ( .A0_t (StateOut[113]), .B0_t (StateFromChi[105]), .Z0_t (U919_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U919_AND1_U1 ( .A0_t (n9), .B0_t (U919_X), .Z0_t (U919_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U919_XOR2_U1 ( .A0_t (U919_Y), .B0_t (StateOut[113]), .Z0_t (StateOut[105]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U920_XOR1_U1 ( .A0_t (StateOut[121]), .B0_t (StateFromChi[113]), .Z0_t (U920_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U920_AND1_U1 ( .A0_t (n9), .B0_t (U920_X), .Z0_t (U920_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U920_XOR2_U1 ( .A0_t (U920_Y), .B0_t (StateOut[121]), .Z0_t (StateOut[113]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U921_XOR1_U1 ( .A0_t (StateOut[137]), .B0_t (StateFromChi[129]), .Z0_t (U921_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U921_AND1_U1 ( .A0_t (n9), .B0_t (U921_X), .Z0_t (U921_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U921_XOR2_U1 ( .A0_t (U921_Y), .B0_t (StateOut[137]), .Z0_t (StateOut[129]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U922_XOR1_U1 ( .A0_t (StateOut[153]), .B0_t (StateFromChi[145]), .Z0_t (U922_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U922_AND1_U1 ( .A0_t (n9), .B0_t (U922_X), .Z0_t (U922_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U922_XOR2_U1 ( .A0_t (U922_Y), .B0_t (StateOut[153]), .Z0_t (StateOut[145]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U923_XOR1_U1 ( .A0_t (StateOut[161]), .B0_t (StateFromChi[153]), .Z0_t (U923_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U923_AND1_U1 ( .A0_t (n9), .B0_t (U923_X), .Z0_t (U923_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U923_XOR2_U1 ( .A0_t (U923_Y), .B0_t (StateOut[161]), .Z0_t (StateOut[153]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U924_XOR1_U1 ( .A0_t (StateOut[169]), .B0_t (StateFromChi[161]), .Z0_t (U924_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U924_AND1_U1 ( .A0_t (n9), .B0_t (U924_X), .Z0_t (U924_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U924_XOR2_U1 ( .A0_t (U924_Y), .B0_t (StateOut[169]), .Z0_t (StateOut[161]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U925_XOR1_U1 ( .A0_t (StateOut[185]), .B0_t (StateFromChi[177]), .Z0_t (U925_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U925_AND1_U1 ( .A0_t (n9), .B0_t (U925_X), .Z0_t (U925_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U925_XOR2_U1 ( .A0_t (U925_Y), .B0_t (StateOut[185]), .Z0_t (StateOut[177]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U926_XOR1_U1 ( .A0_t (InData[1]), .B0_t (StateFromChi[193]), .Z0_t (U926_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U926_AND1_U1 ( .A0_t (n9), .B0_t (U926_X), .Z0_t (U926_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U926_XOR2_U1 ( .A0_t (U926_Y), .B0_t (InData[1]), .Z0_t (StateOut[193]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U927_XOR1_U1 ( .A0_t (StateOut[24]), .B0_t (StateFromChi[16]), .Z0_t (U927_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U927_AND1_U1 ( .A0_t (n9), .B0_t (U927_X), .Z0_t (U927_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U927_XOR2_U1 ( .A0_t (U927_Y), .B0_t (StateOut[24]), .Z0_t (StateOut[16]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U928_XOR1_U1 ( .A0_t (StateOut[40]), .B0_t (StateFromChi[32]), .Z0_t (U928_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U928_AND1_U1 ( .A0_t (n9), .B0_t (U928_X), .Z0_t (U928_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U928_XOR2_U1 ( .A0_t (U928_Y), .B0_t (StateOut[40]), .Z0_t (StateOut[32]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U929_XOR1_U1 ( .A0_t (StateOut[48]), .B0_t (StateFromChi[40]), .Z0_t (U929_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U929_AND1_U1 ( .A0_t (n9), .B0_t (U929_X), .Z0_t (U929_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U929_XOR2_U1 ( .A0_t (U929_Y), .B0_t (StateOut[48]), .Z0_t (StateOut[40]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U930_XOR1_U1 ( .A0_t (StateOut[56]), .B0_t (StateFromChi[48]), .Z0_t (U930_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U930_AND1_U1 ( .A0_t (n9), .B0_t (U930_X), .Z0_t (U930_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U930_XOR2_U1 ( .A0_t (U930_Y), .B0_t (StateOut[56]), .Z0_t (StateOut[48]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U931_XOR1_U1 ( .A0_t (StateOut[64]), .B0_t (StateFromChi[56]), .Z0_t (U931_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U931_AND1_U1 ( .A0_t (n9), .B0_t (U931_X), .Z0_t (U931_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U931_XOR2_U1 ( .A0_t (U931_Y), .B0_t (StateOut[64]), .Z0_t (StateOut[56]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U932_XOR1_U1 ( .A0_t (StateOut[88]), .B0_t (StateFromChi[80]), .Z0_t (U932_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U932_AND1_U1 ( .A0_t (n9), .B0_t (U932_X), .Z0_t (U932_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U932_XOR2_U1 ( .A0_t (U932_Y), .B0_t (StateOut[88]), .Z0_t (StateOut[80]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U933_XOR1_U1 ( .A0_t (StateOut[112]), .B0_t (StateFromChi[104]), .Z0_t (U933_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U933_AND1_U1 ( .A0_t (n9), .B0_t (U933_X), .Z0_t (U933_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U933_XOR2_U1 ( .A0_t (U933_Y), .B0_t (StateOut[112]), .Z0_t (StateOut[104]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U934_XOR1_U1 ( .A0_t (StateOut[160]), .B0_t (StateFromChi[152]), .Z0_t (U934_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U934_AND1_U1 ( .A0_t (n9), .B0_t (U934_X), .Z0_t (U934_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U934_XOR2_U1 ( .A0_t (U934_Y), .B0_t (StateOut[160]), .Z0_t (StateOut[152]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U935_XOR1_U1 ( .A0_t (StateOut[168]), .B0_t (StateFromChi[160]), .Z0_t (U935_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U935_AND1_U1 ( .A0_t (n9), .B0_t (U935_X), .Z0_t (U935_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U935_XOR2_U1 ( .A0_t (U935_Y), .B0_t (StateOut[168]), .Z0_t (StateOut[160]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U936_XOR1_U1 ( .A0_t (StateOut[176]), .B0_t (StateFromChi[168]), .Z0_t (U936_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U936_AND1_U1 ( .A0_t (n9), .B0_t (U936_X), .Z0_t (U936_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U936_XOR2_U1 ( .A0_t (U936_Y), .B0_t (StateOut[176]), .Z0_t (StateOut[168]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U937_XOR1_U1 ( .A0_t (InData[0]), .B0_t (StateFromChi[192]), .Z0_t (U937_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U937_AND1_U1 ( .A0_t (n9), .B0_t (U937_X), .Z0_t (U937_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U937_XOR2_U1 ( .A0_t (U937_Y), .B0_t (InData[0]), .Z0_t (StateOut[192]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U938_XOR1_U1 ( .A0_t (StateOut[23]), .B0_t (StateFromChi[15]), .Z0_t (U938_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U938_AND1_U1 ( .A0_t (n9), .B0_t (U938_X), .Z0_t (U938_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U938_XOR2_U1 ( .A0_t (U938_Y), .B0_t (StateOut[23]), .Z0_t (StateOut[15]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U939_XOR1_U1 ( .A0_t (StateOut[55]), .B0_t (StateFromChi[47]), .Z0_t (U939_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U939_AND1_U1 ( .A0_t (n9), .B0_t (U939_X), .Z0_t (U939_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U939_XOR2_U1 ( .A0_t (U939_Y), .B0_t (StateOut[55]), .Z0_t (StateOut[47]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U940_XOR1_U1 ( .A0_t (StateOut[79]), .B0_t (StateFromChi[71]), .Z0_t (U940_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U940_AND1_U1 ( .A0_t (n9), .B0_t (U940_X), .Z0_t (U940_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U940_XOR2_U1 ( .A0_t (U940_Y), .B0_t (StateOut[79]), .Z0_t (StateOut[71]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U941_XOR1_U1 ( .A0_t (StateOut[87]), .B0_t (StateFromChi[79]), .Z0_t (U941_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U941_AND1_U1 ( .A0_t (n9), .B0_t (U941_X), .Z0_t (U941_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U941_XOR2_U1 ( .A0_t (U941_Y), .B0_t (StateOut[87]), .Z0_t (StateOut[79]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U942_XOR1_U1 ( .A0_t (StateOut[103]), .B0_t (StateFromChi[95]), .Z0_t (U942_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U942_AND1_U1 ( .A0_t (n9), .B0_t (U942_X), .Z0_t (U942_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U942_XOR2_U1 ( .A0_t (U942_Y), .B0_t (StateOut[103]), .Z0_t (StateOut[95]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U943_XOR1_U1 ( .A0_t (StateOut[111]), .B0_t (StateFromChi[103]), .Z0_t (U943_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U943_AND1_U1 ( .A0_t (n9), .B0_t (U943_X), .Z0_t (U943_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U943_XOR2_U1 ( .A0_t (U943_Y), .B0_t (StateOut[111]), .Z0_t (StateOut[103]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U944_XOR1_U1 ( .A0_t (StateOut[135]), .B0_t (StateFromChi[127]), .Z0_t (U944_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U944_AND1_U1 ( .A0_t (n9), .B0_t (U944_X), .Z0_t (U944_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U944_XOR2_U1 ( .A0_t (U944_Y), .B0_t (StateOut[135]), .Z0_t (StateOut[127]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U945_XOR1_U1 ( .A0_t (StateOut[143]), .B0_t (StateFromChi[135]), .Z0_t (U945_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U945_AND1_U1 ( .A0_t (n9), .B0_t (U945_X), .Z0_t (U945_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U945_XOR2_U1 ( .A0_t (U945_Y), .B0_t (StateOut[143]), .Z0_t (StateOut[135]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U946_XOR1_U1 ( .A0_t (StateOut[167]), .B0_t (StateFromChi[159]), .Z0_t (U946_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U946_AND1_U1 ( .A0_t (n9), .B0_t (U946_X), .Z0_t (U946_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U946_XOR2_U1 ( .A0_t (U946_Y), .B0_t (StateOut[167]), .Z0_t (StateOut[159]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U947_XOR1_U1 ( .A0_t (StateOut[191]), .B0_t (StateFromChi[183]), .Z0_t (U947_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U947_AND1_U1 ( .A0_t (n9), .B0_t (U947_X), .Z0_t (U947_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U947_XOR2_U1 ( .A0_t (U947_Y), .B0_t (StateOut[191]), .Z0_t (StateOut[183]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U948_XOR1_U1 ( .A0_t (StateOut[199]), .B0_t (StateFromChi[191]), .Z0_t (U948_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U948_AND1_U1 ( .A0_t (n9), .B0_t (U948_X), .Z0_t (U948_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U948_XOR2_U1 ( .A0_t (U948_Y), .B0_t (StateOut[199]), .Z0_t (StateOut[191]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U949_XOR1_U1 ( .A0_t (StateOut[22]), .B0_t (StateFromChi[14]), .Z0_t (U949_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U949_AND1_U1 ( .A0_t (n9), .B0_t (U949_X), .Z0_t (U949_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U949_XOR2_U1 ( .A0_t (U949_Y), .B0_t (StateOut[22]), .Z0_t (StateOut[14]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U950_XOR1_U1 ( .A0_t (StateOut[54]), .B0_t (StateFromChi[46]), .Z0_t (U950_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U950_AND1_U1 ( .A0_t (n9), .B0_t (U950_X), .Z0_t (U950_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U950_XOR2_U1 ( .A0_t (U950_Y), .B0_t (StateOut[54]), .Z0_t (StateOut[46]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U951_XOR1_U1 ( .A0_t (StateOut[78]), .B0_t (StateFromChi[70]), .Z0_t (U951_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U951_AND1_U1 ( .A0_t (n9), .B0_t (U951_X), .Z0_t (U951_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U951_XOR2_U1 ( .A0_t (U951_Y), .B0_t (StateOut[78]), .Z0_t (StateOut[70]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U952_XOR1_U1 ( .A0_t (StateOut[86]), .B0_t (StateFromChi[78]), .Z0_t (U952_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U952_AND1_U1 ( .A0_t (n9), .B0_t (U952_X), .Z0_t (U952_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U952_XOR2_U1 ( .A0_t (U952_Y), .B0_t (StateOut[86]), .Z0_t (StateOut[78]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U953_XOR1_U1 ( .A0_t (StateOut[102]), .B0_t (StateFromChi[94]), .Z0_t (U953_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U953_AND1_U1 ( .A0_t (n9), .B0_t (U953_X), .Z0_t (U953_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U953_XOR2_U1 ( .A0_t (U953_Y), .B0_t (StateOut[102]), .Z0_t (StateOut[94]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U954_XOR1_U1 ( .A0_t (StateOut[110]), .B0_t (StateFromChi[102]), .Z0_t (U954_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U954_AND1_U1 ( .A0_t (n9), .B0_t (U954_X), .Z0_t (U954_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U954_XOR2_U1 ( .A0_t (U954_Y), .B0_t (StateOut[110]), .Z0_t (StateOut[102]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U955_XOR1_U1 ( .A0_t (StateOut[134]), .B0_t (StateFromChi[126]), .Z0_t (U955_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U955_AND1_U1 ( .A0_t (n9), .B0_t (U955_X), .Z0_t (U955_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U955_XOR2_U1 ( .A0_t (U955_Y), .B0_t (StateOut[134]), .Z0_t (StateOut[126]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U956_XOR1_U1 ( .A0_t (StateOut[142]), .B0_t (StateFromChi[134]), .Z0_t (U956_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U956_AND1_U1 ( .A0_t (n9), .B0_t (U956_X), .Z0_t (U956_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U956_XOR2_U1 ( .A0_t (U956_Y), .B0_t (StateOut[142]), .Z0_t (StateOut[134]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U957_XOR1_U1 ( .A0_t (StateOut[166]), .B0_t (StateFromChi[158]), .Z0_t (U957_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U957_AND1_U1 ( .A0_t (n9), .B0_t (U957_X), .Z0_t (U957_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U957_XOR2_U1 ( .A0_t (U957_Y), .B0_t (StateOut[166]), .Z0_t (StateOut[158]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U958_XOR1_U1 ( .A0_t (StateOut[190]), .B0_t (StateFromChi[182]), .Z0_t (U958_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U958_AND1_U1 ( .A0_t (n9), .B0_t (U958_X), .Z0_t (U958_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U958_XOR2_U1 ( .A0_t (U958_Y), .B0_t (StateOut[190]), .Z0_t (StateOut[182]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U959_XOR1_U1 ( .A0_t (StateOut[198]), .B0_t (StateFromChi[190]), .Z0_t (U959_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U959_AND1_U1 ( .A0_t (n9), .B0_t (U959_X), .Z0_t (U959_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U959_XOR2_U1 ( .A0_t (U959_Y), .B0_t (StateOut[198]), .Z0_t (StateOut[190]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U960_XOR1_U1 ( .A0_t (StateOut[21]), .B0_t (StateFromChi[13]), .Z0_t (U960_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U960_AND1_U1 ( .A0_t (n9), .B0_t (U960_X), .Z0_t (U960_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U960_XOR2_U1 ( .A0_t (U960_Y), .B0_t (StateOut[21]), .Z0_t (StateOut[13]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U961_XOR1_U1 ( .A0_t (StateOut[53]), .B0_t (StateFromChi[45]), .Z0_t (U961_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U961_AND1_U1 ( .A0_t (n9), .B0_t (U961_X), .Z0_t (U961_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U961_XOR2_U1 ( .A0_t (U961_Y), .B0_t (StateOut[53]), .Z0_t (StateOut[45]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U962_XOR1_U1 ( .A0_t (StateOut[85]), .B0_t (StateFromChi[77]), .Z0_t (U962_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U962_AND1_U1 ( .A0_t (n9), .B0_t (U962_X), .Z0_t (U962_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U962_XOR2_U1 ( .A0_t (U962_Y), .B0_t (StateOut[85]), .Z0_t (StateOut[77]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U963_XOR1_U1 ( .A0_t (StateOut[101]), .B0_t (StateFromChi[93]), .Z0_t (U963_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U963_AND1_U1 ( .A0_t (n9), .B0_t (U963_X), .Z0_t (U963_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U963_XOR2_U1 ( .A0_t (U963_Y), .B0_t (StateOut[101]), .Z0_t (StateOut[93]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U964_XOR1_U1 ( .A0_t (StateOut[109]), .B0_t (StateFromChi[101]), .Z0_t (U964_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U964_AND1_U1 ( .A0_t (n9), .B0_t (U964_X), .Z0_t (U964_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U964_XOR2_U1 ( .A0_t (U964_Y), .B0_t (StateOut[109]), .Z0_t (StateOut[101]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U965_XOR1_U1 ( .A0_t (StateOut[117]), .B0_t (StateFromChi[109]), .Z0_t (U965_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U965_AND1_U1 ( .A0_t (n9), .B0_t (U965_X), .Z0_t (U965_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U965_XOR2_U1 ( .A0_t (U965_Y), .B0_t (StateOut[117]), .Z0_t (StateOut[109]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U966_XOR1_U1 ( .A0_t (StateOut[133]), .B0_t (StateFromChi[125]), .Z0_t (U966_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U966_AND1_U1 ( .A0_t (n9), .B0_t (U966_X), .Z0_t (U966_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U966_XOR2_U1 ( .A0_t (U966_Y), .B0_t (StateOut[133]), .Z0_t (StateOut[125]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U967_XOR1_U1 ( .A0_t (StateOut[165]), .B0_t (StateFromChi[157]), .Z0_t (U967_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U967_AND1_U1 ( .A0_t (n9), .B0_t (U967_X), .Z0_t (U967_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U967_XOR2_U1 ( .A0_t (U967_Y), .B0_t (StateOut[165]), .Z0_t (StateOut[157]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U968_XOR1_U1 ( .A0_t (StateOut[189]), .B0_t (StateFromChi[181]), .Z0_t (U968_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U968_AND1_U1 ( .A0_t (n9), .B0_t (U968_X), .Z0_t (U968_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U968_XOR2_U1 ( .A0_t (U968_Y), .B0_t (StateOut[189]), .Z0_t (StateOut[181]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U969_XOR1_U1 ( .A0_t (StateOut[197]), .B0_t (StateFromChi[189]), .Z0_t (U969_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U969_AND1_U1 ( .A0_t (n9), .B0_t (U969_X), .Z0_t (U969_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U969_XOR2_U1 ( .A0_t (U969_Y), .B0_t (StateOut[197]), .Z0_t (StateOut[189]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U970_XOR1_U1 ( .A0_t (InData[5]), .B0_t (StateFromChi[197]), .Z0_t (U970_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U970_AND1_U1 ( .A0_t (n9), .B0_t (U970_X), .Z0_t (U970_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U970_XOR2_U1 ( .A0_t (U970_Y), .B0_t (InData[5]), .Z0_t (StateOut[197]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U971_XOR1_U1 ( .A0_t (StateOut[20]), .B0_t (StateFromChi[12]), .Z0_t (U971_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U971_AND1_U1 ( .A0_t (n9), .B0_t (U971_X), .Z0_t (U971_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U971_XOR2_U1 ( .A0_t (U971_Y), .B0_t (StateOut[20]), .Z0_t (StateOut[12]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U972_XOR1_U1 ( .A0_t (StateOut[28]), .B0_t (StateFromChi[20]), .Z0_t (U972_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U972_AND1_U1 ( .A0_t (n9), .B0_t (U972_X), .Z0_t (U972_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U972_XOR2_U1 ( .A0_t (U972_Y), .B0_t (StateOut[28]), .Z0_t (StateOut[20]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U973_XOR1_U1 ( .A0_t (StateOut[84]), .B0_t (StateFromChi[76]), .Z0_t (U973_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U973_AND1_U1 ( .A0_t (n9), .B0_t (U973_X), .Z0_t (U973_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U973_XOR2_U1 ( .A0_t (U973_Y), .B0_t (StateOut[84]), .Z0_t (StateOut[76]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U974_XOR1_U1 ( .A0_t (StateOut[108]), .B0_t (StateFromChi[100]), .Z0_t (U974_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U974_AND1_U1 ( .A0_t (n9), .B0_t (U974_X), .Z0_t (U974_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U974_XOR2_U1 ( .A0_t (U974_Y), .B0_t (StateOut[108]), .Z0_t (StateOut[100]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U975_XOR1_U1 ( .A0_t (StateOut[116]), .B0_t (StateFromChi[108]), .Z0_t (U975_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U975_AND1_U1 ( .A0_t (n9), .B0_t (U975_X), .Z0_t (U975_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U975_XOR2_U1 ( .A0_t (U975_Y), .B0_t (StateOut[116]), .Z0_t (StateOut[108]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U976_XOR1_U1 ( .A0_t (StateOut[132]), .B0_t (StateFromChi[124]), .Z0_t (U976_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U976_AND1_U1 ( .A0_t (n9), .B0_t (U976_X), .Z0_t (U976_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U976_XOR2_U1 ( .A0_t (U976_Y), .B0_t (StateOut[132]), .Z0_t (StateOut[124]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U977_XOR1_U1 ( .A0_t (StateOut[164]), .B0_t (StateFromChi[156]), .Z0_t (U977_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U977_AND1_U1 ( .A0_t (n9), .B0_t (U977_X), .Z0_t (U977_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U977_XOR2_U1 ( .A0_t (U977_Y), .B0_t (StateOut[164]), .Z0_t (StateOut[156]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U978_XOR1_U1 ( .A0_t (StateOut[188]), .B0_t (StateFromChi[180]), .Z0_t (U978_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U978_AND1_U1 ( .A0_t (n9), .B0_t (U978_X), .Z0_t (U978_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U978_XOR2_U1 ( .A0_t (U978_Y), .B0_t (StateOut[188]), .Z0_t (StateOut[180]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U979_XOR1_U1 ( .A0_t (StateOut[196]), .B0_t (StateFromChi[188]), .Z0_t (U979_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U979_AND1_U1 ( .A0_t (n9), .B0_t (U979_X), .Z0_t (U979_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U979_XOR2_U1 ( .A0_t (U979_Y), .B0_t (StateOut[196]), .Z0_t (StateOut[188]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U980_XOR1_U1 ( .A0_t (InData[4]), .B0_t (StateFromChi[196]), .Z0_t (U980_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U980_AND1_U1 ( .A0_t (n9), .B0_t (U980_X), .Z0_t (U980_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U980_XOR2_U1 ( .A0_t (U980_Y), .B0_t (InData[4]), .Z0_t (StateOut[196]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U981_XOR1_U1 ( .A0_t (StateOut[19]), .B0_t (StateFromChi[11]), .Z0_t (U981_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U981_AND1_U1 ( .A0_t (n9), .B0_t (U981_X), .Z0_t (U981_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U981_XOR2_U1 ( .A0_t (U981_Y), .B0_t (StateOut[19]), .Z0_t (StateOut[11]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U982_XOR1_U1 ( .A0_t (StateOut[27]), .B0_t (StateFromChi[19]), .Z0_t (U982_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U982_AND1_U1 ( .A0_t (n9), .B0_t (U982_X), .Z0_t (U982_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U982_XOR2_U1 ( .A0_t (U982_Y), .B0_t (StateOut[27]), .Z0_t (StateOut[19]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U983_XOR1_U1 ( .A0_t (StateOut[83]), .B0_t (StateFromChi[75]), .Z0_t (U983_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U983_AND1_U1 ( .A0_t (n9), .B0_t (U983_X), .Z0_t (U983_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U983_XOR2_U1 ( .A0_t (U983_Y), .B0_t (StateOut[83]), .Z0_t (StateOut[75]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U984_XOR1_U1 ( .A0_t (StateOut[107]), .B0_t (StateFromChi[99]), .Z0_t (U984_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U984_AND1_U1 ( .A0_t (n9), .B0_t (U984_X), .Z0_t (U984_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U984_XOR2_U1 ( .A0_t (U984_Y), .B0_t (StateOut[107]), .Z0_t (StateOut[99]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U985_XOR1_U1 ( .A0_t (StateOut[115]), .B0_t (StateFromChi[107]), .Z0_t (U985_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U985_AND1_U1 ( .A0_t (n9), .B0_t (U985_X), .Z0_t (U985_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U985_XOR2_U1 ( .A0_t (U985_Y), .B0_t (StateOut[115]), .Z0_t (StateOut[107]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U986_XOR1_U1 ( .A0_t (StateOut[131]), .B0_t (StateFromChi[123]), .Z0_t (U986_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U986_AND1_U1 ( .A0_t (n9), .B0_t (U986_X), .Z0_t (U986_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U986_XOR2_U1 ( .A0_t (U986_Y), .B0_t (StateOut[131]), .Z0_t (StateOut[123]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U987_XOR1_U1 ( .A0_t (StateOut[163]), .B0_t (StateFromChi[155]), .Z0_t (U987_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U987_AND1_U1 ( .A0_t (n9), .B0_t (U987_X), .Z0_t (U987_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U987_XOR2_U1 ( .A0_t (U987_Y), .B0_t (StateOut[163]), .Z0_t (StateOut[155]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U988_XOR1_U1 ( .A0_t (StateOut[195]), .B0_t (StateFromChi[187]), .Z0_t (U988_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U988_AND1_U1 ( .A0_t (n9), .B0_t (U988_X), .Z0_t (U988_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U988_XOR2_U1 ( .A0_t (U988_Y), .B0_t (StateOut[195]), .Z0_t (StateOut[187]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U989_XOR1_U1 ( .A0_t (InData[3]), .B0_t (StateFromChi[195]), .Z0_t (U989_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U989_AND1_U1 ( .A0_t (n9), .B0_t (U989_X), .Z0_t (U989_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U989_XOR2_U1 ( .A0_t (U989_Y), .B0_t (InData[3]), .Z0_t (StateOut[195]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U990_XOR1_U1 ( .A0_t (StateOut[18]), .B0_t (StateFromChi[10]), .Z0_t (U990_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U990_AND1_U1 ( .A0_t (n9), .B0_t (U990_X), .Z0_t (U990_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U990_XOR2_U1 ( .A0_t (U990_Y), .B0_t (StateOut[18]), .Z0_t (StateOut[10]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U991_XOR1_U1 ( .A0_t (StateOut[26]), .B0_t (StateFromChi[18]), .Z0_t (U991_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U991_AND1_U1 ( .A0_t (n9), .B0_t (U991_X), .Z0_t (U991_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U991_XOR2_U1 ( .A0_t (U991_Y), .B0_t (StateOut[26]), .Z0_t (StateOut[18]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U992_XOR1_U1 ( .A0_t (StateOut[74]), .B0_t (StateFromChi[66]), .Z0_t (U992_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U992_AND1_U1 ( .A0_t (n9), .B0_t (U992_X), .Z0_t (U992_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U992_XOR2_U1 ( .A0_t (U992_Y), .B0_t (StateOut[74]), .Z0_t (StateOut[66]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U993_XOR1_U1 ( .A0_t (StateOut[82]), .B0_t (StateFromChi[74]), .Z0_t (U993_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U993_AND1_U1 ( .A0_t (n9), .B0_t (U993_X), .Z0_t (U993_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U993_XOR2_U1 ( .A0_t (U993_Y), .B0_t (StateOut[82]), .Z0_t (StateOut[74]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U994_XOR1_U1 ( .A0_t (StateOut[106]), .B0_t (StateFromChi[98]), .Z0_t (U994_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U994_AND1_U1 ( .A0_t (n9), .B0_t (U994_X), .Z0_t (U994_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U994_XOR2_U1 ( .A0_t (U994_Y), .B0_t (StateOut[106]), .Z0_t (StateOut[98]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U995_XOR1_U1 ( .A0_t (StateOut[130]), .B0_t (StateFromChi[122]), .Z0_t (U995_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U995_AND1_U1 ( .A0_t (n9), .B0_t (U995_X), .Z0_t (U995_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U995_XOR2_U1 ( .A0_t (U995_Y), .B0_t (StateOut[130]), .Z0_t (StateOut[122]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U996_XOR1_U1 ( .A0_t (StateOut[194]), .B0_t (StateFromChi[186]), .Z0_t (U996_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U996_AND1_U1 ( .A0_t (n9), .B0_t (U996_X), .Z0_t (U996_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U996_XOR2_U1 ( .A0_t (U996_Y), .B0_t (StateOut[194]), .Z0_t (StateOut[186]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U997_XOR1_U1 ( .A0_t (StateOut[17]), .B0_t (StateFromChi[9]), .Z0_t (U997_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U997_AND1_U1 ( .A0_t (n9), .B0_t (U997_X), .Z0_t (U997_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U997_XOR2_U1 ( .A0_t (U997_Y), .B0_t (StateOut[17]), .Z0_t (StateOut[9]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U998_XOR1_U1 ( .A0_t (StateOut[73]), .B0_t (StateFromChi[65]), .Z0_t (U998_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U998_AND1_U1 ( .A0_t (n9), .B0_t (U998_X), .Z0_t (U998_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U998_XOR2_U1 ( .A0_t (U998_Y), .B0_t (StateOut[73]), .Z0_t (StateOut[65]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U999_XOR1_U1 ( .A0_t (StateOut[81]), .B0_t (StateFromChi[73]), .Z0_t (U999_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U999_AND1_U1 ( .A0_t (n9), .B0_t (U999_X), .Z0_t (U999_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U999_XOR2_U1 ( .A0_t (U999_Y), .B0_t (StateOut[81]), .Z0_t (StateOut[73]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1000_XOR1_U1 ( .A0_t (StateOut[97]), .B0_t (StateFromChi[89]), .Z0_t (U1000_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1000_AND1_U1 ( .A0_t (n9), .B0_t (U1000_X), .Z0_t (U1000_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U1000_XOR2_U1 ( .A0_t (U1000_Y), .B0_t (StateOut[97]), .Z0_t (StateOut[89]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1001_XOR1_U1 ( .A0_t (StateOut[105]), .B0_t (StateFromChi[97]), .Z0_t (U1001_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1001_AND1_U1 ( .A0_t (n9), .B0_t (U1001_X), .Z0_t (U1001_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U1001_XOR2_U1 ( .A0_t (U1001_Y), .B0_t (StateOut[105]), .Z0_t (StateOut[97]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1002_XOR1_U1 ( .A0_t (StateOut[129]), .B0_t (StateFromChi[121]), .Z0_t (U1002_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1002_AND1_U1 ( .A0_t (n9), .B0_t (U1002_X), .Z0_t (U1002_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U1002_XOR2_U1 ( .A0_t (U1002_Y), .B0_t (StateOut[129]), .Z0_t (StateOut[121]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1003_XOR1_U1 ( .A0_t (StateOut[193]), .B0_t (StateFromChi[185]), .Z0_t (U1003_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1003_AND1_U1 ( .A0_t (n9), .B0_t (U1003_X), .Z0_t (U1003_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U1003_XOR2_U1 ( .A0_t (U1003_Y), .B0_t (StateOut[193]), .Z0_t (StateOut[185]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1004_XOR1_U1 ( .A0_t (StateOut[16]), .B0_t (StateFromChi[8]), .Z0_t (U1004_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1004_AND1_U1 ( .A0_t (n9), .B0_t (U1004_X), .Z0_t (U1004_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U1004_XOR2_U1 ( .A0_t (U1004_Y), .B0_t (StateOut[16]), .Z0_t (StateOut[8]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1005_XOR1_U1 ( .A0_t (StateOut[72]), .B0_t (StateFromChi[64]), .Z0_t (U1005_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1005_AND1_U1 ( .A0_t (n9), .B0_t (U1005_X), .Z0_t (U1005_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U1005_XOR2_U1 ( .A0_t (U1005_Y), .B0_t (StateOut[72]), .Z0_t (StateOut[64]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1006_XOR1_U1 ( .A0_t (StateOut[80]), .B0_t (StateFromChi[72]), .Z0_t (U1006_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1006_AND1_U1 ( .A0_t (n9), .B0_t (U1006_X), .Z0_t (U1006_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U1006_XOR2_U1 ( .A0_t (U1006_Y), .B0_t (StateOut[80]), .Z0_t (StateOut[72]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1007_XOR1_U1 ( .A0_t (StateOut[96]), .B0_t (StateFromChi[88]), .Z0_t (U1007_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1007_AND1_U1 ( .A0_t (n9), .B0_t (U1007_X), .Z0_t (U1007_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U1007_XOR2_U1 ( .A0_t (U1007_Y), .B0_t (StateOut[96]), .Z0_t (StateOut[88]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1008_XOR1_U1 ( .A0_t (StateOut[104]), .B0_t (StateFromChi[96]), .Z0_t (U1008_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1008_AND1_U1 ( .A0_t (n9), .B0_t (U1008_X), .Z0_t (U1008_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U1008_XOR2_U1 ( .A0_t (U1008_Y), .B0_t (StateOut[104]), .Z0_t (StateOut[96]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1009_XOR1_U1 ( .A0_t (StateOut[128]), .B0_t (StateFromChi[120]), .Z0_t (U1009_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1009_AND1_U1 ( .A0_t (n9), .B0_t (U1009_X), .Z0_t (U1009_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U1009_XOR2_U1 ( .A0_t (U1009_Y), .B0_t (StateOut[128]), .Z0_t (StateOut[120]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1010_XOR1_U1 ( .A0_t (StateOut[136]), .B0_t (StateFromChi[128]), .Z0_t (U1010_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1010_AND1_U1 ( .A0_t (n9), .B0_t (U1010_X), .Z0_t (U1010_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U1010_XOR2_U1 ( .A0_t (U1010_Y), .B0_t (StateOut[136]), .Z0_t (StateOut[128]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1011_XOR1_U1 ( .A0_t (StateOut[184]), .B0_t (StateFromChi[176]), .Z0_t (U1011_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1011_AND1_U1 ( .A0_t (n9), .B0_t (U1011_X), .Z0_t (U1011_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U1011_XOR2_U1 ( .A0_t (U1011_Y), .B0_t (StateOut[184]), .Z0_t (StateOut[176]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1012_XOR1_U1 ( .A0_t (StateOut[192]), .B0_t (StateFromChi[184]), .Z0_t (U1012_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1012_AND1_U1 ( .A0_t (n9), .B0_t (U1012_X), .Z0_t (U1012_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U1012_XOR2_U1 ( .A0_t (U1012_Y), .B0_t (StateOut[192]), .Z0_t (StateOut[184]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1013_XOR1_U1 ( .A0_t (StateOut[14]), .B0_t (StateFromChi[6]), .Z0_t (U1013_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1013_AND1_U1 ( .A0_t (n9), .B0_t (U1013_X), .Z0_t (U1013_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U1013_XOR2_U1 ( .A0_t (U1013_Y), .B0_t (StateOut[14]), .Z0_t (OutData[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1014_XOR1_U1 ( .A0_t (StateOut[13]), .B0_t (StateFromChi[5]), .Z0_t (U1014_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1014_AND1_U1 ( .A0_t (n9), .B0_t (U1014_X), .Z0_t (U1014_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U1014_XOR2_U1 ( .A0_t (U1014_Y), .B0_t (StateOut[13]), .Z0_t (OutData[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1015_XOR1_U1 ( .A0_t (StateOut[12]), .B0_t (StateFromChi[4]), .Z0_t (U1015_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1015_AND1_U1 ( .A0_t (n9), .B0_t (U1015_X), .Z0_t (U1015_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U1015_XOR2_U1 ( .A0_t (U1015_Y), .B0_t (StateOut[12]), .Z0_t (OutData[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1016_XOR1_U1 ( .A0_t (StateOut[10]), .B0_t (StateFromChi[2]), .Z0_t (U1016_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U1016_AND1_U1 ( .A0_t (n9), .B0_t (U1016_X), .Z0_t (U1016_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) U1016_XOR2_U1 ( .A0_t (U1016_Y), .B0_t (StateOut[10]), .Z0_t (OutData[2]) ) ;

    /* register cells */
endmodule
